magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< pwell >>
rect -76 -26 452 226
<< mvnmos >>
rect 0 0 160 200
rect 216 0 376 200
<< mvndiff >>
rect -50 0 0 200
rect 160 182 216 200
rect 160 148 171 182
rect 205 148 216 182
rect 160 114 216 148
rect 160 80 171 114
rect 205 80 216 114
rect 160 46 216 80
rect 160 12 171 46
rect 205 12 216 46
rect 160 0 216 12
rect 376 0 426 200
<< mvndiffc >>
rect 171 148 205 182
rect 171 80 205 114
rect 171 12 205 46
<< poly >>
rect 0 200 160 226
rect 216 200 376 226
rect 0 -26 160 0
rect 216 -26 376 0
<< locali >>
rect 171 182 205 198
rect 171 114 205 148
rect 171 46 205 80
rect 171 -4 205 12
<< metal1 >>
rect -51 -16 -5 186
rect 381 -16 427 186
use hvDFL1sd2_CDNS_52468879185133  hvDFL1sd2_CDNS_52468879185133_0
timestamp 1704896540
transform 1 0 160 0 1 0
box 0 0 1 1
use hvDFM1sd_CDNS_52468879185147  hvDFM1sd_CDNS_52468879185147_0
timestamp 1704896540
transform -1 0 0 0 1 0
box -26 -26 79 226
use hvDFM1sd_CDNS_52468879185147  hvDFM1sd_CDNS_52468879185147_1
timestamp 1704896540
transform 1 0 376 0 1 0
box -26 -26 79 226
<< labels >>
flabel comment s -28 85 -28 85 0 FreeSans 300 0 0 0 S
flabel comment s 188 97 188 97 0 FreeSans 300 0 0 0 D
flabel comment s 404 85 404 85 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 85981374
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85979984
<< end >>
