magic
tech sky130A
timestamp 1704896540
<< properties >>
string GDS_END 78412332
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 78411564
<< end >>
