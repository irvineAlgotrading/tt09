magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -77 1179 1723 1285
rect -77 925 77 1179
rect 1569 925 1723 1179
<< pwell >>
rect -67 341 359 427
rect 273 43 359 341
rect 1262 341 1713 427
rect 1262 43 1348 341
rect 273 -43 1348 43
<< psubdiff >>
rect -41 367 -17 401
rect 17 367 65 401
rect 99 367 135 401
rect 169 367 205 401
rect 239 377 333 401
rect 239 367 299 377
rect 299 296 333 343
rect 299 215 333 262
rect 299 134 333 181
rect 1288 367 1312 401
rect 1346 367 1391 401
rect 1425 367 1469 401
rect 1503 367 1547 401
rect 1581 367 1629 401
rect 1663 367 1687 401
rect 1288 284 1322 367
rect 1288 203 1322 250
rect 299 17 333 100
rect 1288 122 1322 169
rect 1288 41 1322 88
rect 299 -17 323 17
rect 357 -17 396 17
rect 430 -17 468 17
rect 502 -17 540 17
rect 574 -17 612 17
rect 646 -17 684 17
rect 718 -17 756 17
rect 790 -17 828 17
rect 862 -17 900 17
rect 934 -17 972 17
rect 1006 -17 1044 17
rect 1078 -17 1116 17
rect 1150 -17 1188 17
rect 1222 7 1288 17
rect 1222 -17 1322 7
<< nsubdiff >>
rect -41 1215 -17 1249
rect 17 1215 75 1249
rect 109 1215 145 1249
rect 179 1215 215 1249
rect 249 1215 285 1249
rect 319 1215 355 1249
rect 389 1215 425 1249
rect 459 1215 495 1249
rect 529 1215 565 1249
rect 599 1215 635 1249
rect 669 1215 705 1249
rect 739 1215 775 1249
rect 809 1215 845 1249
rect 879 1215 915 1249
rect 949 1215 985 1249
rect 1019 1215 1054 1249
rect 1088 1215 1123 1249
rect 1157 1215 1192 1249
rect 1226 1215 1261 1249
rect 1295 1215 1330 1249
rect 1364 1215 1399 1249
rect 1433 1215 1468 1249
rect 1502 1215 1537 1249
rect 1571 1215 1629 1249
rect 1663 1215 1687 1249
<< psubdiffcont >>
rect -17 367 17 401
rect 65 367 99 401
rect 135 367 169 401
rect 205 367 239 401
rect 299 343 333 377
rect 299 262 333 296
rect 299 181 333 215
rect 299 100 333 134
rect 1312 367 1346 401
rect 1391 367 1425 401
rect 1469 367 1503 401
rect 1547 367 1581 401
rect 1629 367 1663 401
rect 1288 250 1322 284
rect 1288 169 1322 203
rect 1288 88 1322 122
rect 323 -17 357 17
rect 396 -17 430 17
rect 468 -17 502 17
rect 540 -17 574 17
rect 612 -17 646 17
rect 684 -17 718 17
rect 756 -17 790 17
rect 828 -17 862 17
rect 900 -17 934 17
rect 972 -17 1006 17
rect 1044 -17 1078 17
rect 1116 -17 1150 17
rect 1188 -17 1222 17
rect 1288 7 1322 41
<< nsubdiffcont >>
rect -17 1215 17 1249
rect 75 1215 109 1249
rect 145 1215 179 1249
rect 215 1215 249 1249
rect 285 1215 319 1249
rect 355 1215 389 1249
rect 425 1215 459 1249
rect 495 1215 529 1249
rect 565 1215 599 1249
rect 635 1215 669 1249
rect 705 1215 739 1249
rect 775 1215 809 1249
rect 845 1215 879 1249
rect 915 1215 949 1249
rect 985 1215 1019 1249
rect 1054 1215 1088 1249
rect 1123 1215 1157 1249
rect 1192 1215 1226 1249
rect 1261 1215 1295 1249
rect 1330 1215 1364 1249
rect 1399 1215 1433 1249
rect 1468 1215 1502 1249
rect 1537 1215 1571 1249
rect 1629 1215 1663 1249
<< poly >>
rect 28 929 228 936
rect 284 929 484 936
rect 28 883 484 929
rect 540 883 740 935
rect 28 867 740 883
rect 28 833 323 867
rect 357 833 391 867
rect 425 833 459 867
rect 493 833 527 867
rect 561 833 595 867
rect 629 833 663 867
rect 697 833 740 867
rect 28 817 740 833
rect 906 883 1106 936
rect 1418 935 1618 936
rect 1162 883 1618 935
rect 906 867 1618 883
rect 906 833 1017 867
rect 1051 833 1085 867
rect 1119 833 1153 867
rect 1187 833 1221 867
rect 1255 833 1289 867
rect 1323 833 1618 867
rect 906 817 1618 833
rect 28 767 228 817
rect 1418 767 1618 817
rect 578 101 712 123
rect 578 67 594 101
rect 628 67 662 101
rect 696 67 712 101
rect 578 51 712 67
rect 930 101 1064 124
rect 930 67 946 101
rect 980 67 1014 101
rect 1048 67 1064 101
rect 930 51 1064 67
<< polycont >>
rect 323 833 357 867
rect 391 833 425 867
rect 459 833 493 867
rect 527 833 561 867
rect 595 833 629 867
rect 663 833 697 867
rect 1017 833 1051 867
rect 1085 833 1119 867
rect 1153 833 1187 867
rect 1221 833 1255 867
rect 1289 833 1323 867
rect 594 67 628 101
rect 662 67 696 101
rect 946 67 980 101
rect 1014 67 1048 101
<< locali >>
rect -33 1215 -17 1249
rect 17 1215 75 1249
rect 109 1215 145 1249
rect 179 1215 215 1249
rect 249 1215 285 1249
rect 319 1215 355 1249
rect 389 1215 425 1249
rect 459 1215 495 1249
rect 529 1215 565 1249
rect 599 1215 635 1249
rect 669 1215 705 1249
rect 739 1215 775 1249
rect 809 1215 845 1249
rect 879 1215 915 1249
rect 949 1215 985 1249
rect 1019 1215 1054 1249
rect 1088 1215 1123 1249
rect 1157 1215 1192 1249
rect 1226 1215 1261 1249
rect 1295 1215 1330 1249
rect 1364 1215 1399 1249
rect 1433 1215 1468 1249
rect 1502 1215 1537 1249
rect 1571 1215 1629 1249
rect 1663 1215 1679 1249
rect -17 1019 17 1057
rect 495 1019 529 1057
rect -17 947 17 985
rect 239 739 273 1008
rect 495 947 529 985
rect 1117 1019 1151 1057
rect 307 833 323 867
rect 357 833 391 867
rect 425 833 459 867
rect 493 833 527 867
rect 573 833 595 867
rect 645 833 663 867
rect 697 833 713 867
rect 751 793 785 983
rect 861 867 895 963
rect 1117 947 1151 985
rect 1629 1019 1663 1057
rect 859 833 897 867
rect 1001 833 1005 867
rect 1051 833 1077 867
rect 1119 833 1153 867
rect 1187 833 1221 867
rect 1255 833 1289 867
rect 1323 833 1339 867
rect 749 759 787 793
rect 751 753 785 759
rect 861 741 895 833
rect 1373 739 1407 963
rect 1629 947 1663 985
rect -17 541 17 579
rect -17 469 17 507
rect 495 541 529 579
rect 495 469 529 507
rect 1117 541 1151 579
rect 1117 469 1151 507
rect 1629 541 1663 579
rect 1629 469 1663 507
rect -33 367 -17 401
rect 17 367 65 401
rect 99 367 135 401
rect 169 367 205 401
rect 239 377 333 401
rect 239 367 299 377
rect 299 296 333 343
rect 299 215 333 262
rect 299 134 333 181
rect 1288 367 1312 401
rect 1346 367 1391 401
rect 1425 367 1469 401
rect 1503 367 1547 401
rect 1581 367 1629 401
rect 1663 367 1679 401
rect 1288 284 1322 367
rect 1288 203 1322 250
rect 1288 122 1322 169
rect 299 17 333 100
rect 594 101 696 117
rect 628 67 662 101
rect 594 51 696 67
rect 946 101 1048 117
rect 980 67 1014 101
rect 946 51 1048 67
rect 1288 41 1322 88
rect 299 -17 323 17
rect 357 -17 396 17
rect 430 -17 468 17
rect 502 -17 540 17
rect 574 -17 612 17
rect 646 -17 684 17
rect 718 -17 756 17
rect 790 -17 828 17
rect 862 -17 900 17
rect 934 -17 972 17
rect 1006 -17 1044 17
rect 1078 -17 1116 17
rect 1150 -17 1188 17
rect 1222 7 1288 17
rect 1222 -17 1322 7
<< viali >>
rect -17 1057 17 1091
rect -17 985 17 1019
rect 495 1057 529 1091
rect -17 913 17 947
rect 495 985 529 1019
rect 1117 1057 1151 1091
rect 1117 985 1151 1019
rect 495 913 529 947
rect 539 833 561 867
rect 561 833 573 867
rect 611 833 629 867
rect 629 833 645 867
rect 1629 1057 1663 1091
rect 1629 985 1663 1019
rect 1117 913 1151 947
rect 825 833 859 867
rect 897 833 931 867
rect 1005 833 1017 867
rect 1017 833 1039 867
rect 1077 833 1085 867
rect 1085 833 1111 867
rect 715 759 749 793
rect 787 759 821 793
rect 1629 913 1663 947
rect -17 579 17 613
rect -17 507 17 541
rect -17 435 17 469
rect 495 579 529 613
rect 495 507 529 541
rect 495 435 529 469
rect 1117 579 1151 613
rect 1117 507 1151 541
rect 1117 435 1151 469
rect 1629 579 1663 613
rect 1629 507 1663 541
rect 1629 435 1663 469
<< metal1 >>
rect -61 1091 1707 1103
rect -61 1057 -17 1091
rect 17 1057 495 1091
rect 529 1057 1117 1091
rect 1151 1057 1629 1091
rect 1663 1057 1707 1091
rect -61 1019 1707 1057
rect -61 985 -17 1019
rect 17 985 495 1019
rect 529 985 1117 1019
rect 1151 985 1629 1019
rect 1663 985 1707 1019
rect -61 947 1707 985
rect -61 913 -17 947
rect 17 913 495 947
rect 529 913 1117 947
rect 1151 913 1629 947
rect 1663 913 1707 947
rect -61 901 1707 913
rect 527 867 943 873
rect 527 833 539 867
rect 573 833 611 867
rect 645 833 825 867
rect 859 833 897 867
rect 931 833 943 867
rect 527 827 943 833
rect 993 867 1123 873
rect 993 833 1005 867
rect 1039 833 1077 867
rect 1111 833 1123 867
rect 993 827 1123 833
tri 965 799 993 827 se
rect 993 799 1032 827
tri 1032 799 1060 827 nw
rect 703 793 986 799
rect 703 759 715 793
rect 749 759 787 793
rect 821 759 986 793
rect 703 753 986 759
tri 986 753 1032 799 nw
rect -61 613 1712 625
rect -61 579 -17 613
rect 17 579 495 613
rect 529 579 1117 613
rect 1151 579 1629 613
rect 1663 579 1712 613
rect -61 541 1712 579
rect -61 507 -17 541
rect 17 507 495 541
rect 529 507 1117 541
rect 1151 507 1629 541
rect 1663 507 1712 541
rect -61 469 1712 507
rect -61 435 -17 469
rect 17 435 495 469
rect 529 435 1117 469
rect 1151 435 1629 469
rect 1663 435 1712 469
rect -61 423 1712 435
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1704896540
transform -1 0 821 0 1 759
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1704896540
transform -1 0 931 0 -1 867
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1704896540
transform 1 0 1005 0 -1 867
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1704896540
transform 1 0 539 0 -1 867
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1704896540
transform 0 -1 529 -1 0 1091
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_1
timestamp 1704896540
transform 0 -1 1151 -1 0 613
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_2
timestamp 1704896540
transform 0 -1 1151 -1 0 1091
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_3
timestamp 1704896540
transform 0 -1 529 -1 0 613
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_4
timestamp 1704896540
transform 0 1 1629 -1 0 613
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_5
timestamp 1704896540
transform 0 1 1629 -1 0 1091
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_6
timestamp 1704896540
transform 0 1 -17 -1 0 613
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_7
timestamp 1704896540
transform 0 1 -17 -1 0 1091
box 0 0 1 1
use nfet_CDNS_524688791851172  nfet_CDNS_524688791851172_0
timestamp 1704896540
transform -1 0 1618 0 1 541
box -79 -26 279 226
use nfet_CDNS_524688791851172  nfet_CDNS_524688791851172_1
timestamp 1704896540
transform 1 0 28 0 1 541
box -79 -26 279 226
use nfet_CDNS_524688791851173  nfet_CDNS_524688791851173_0
timestamp 1704896540
transform -1 0 1106 0 -1 749
box -79 -26 279 626
use nfet_CDNS_524688791851173  nfet_CDNS_524688791851173_1
timestamp 1704896540
transform 1 0 540 0 -1 749
box -79 -26 279 626
use pfet_CDNS_524688791851170  pfet_CDNS_524688791851170_0
timestamp 1704896540
transform -1 0 1106 0 -1 1161
box -89 -36 289 236
use pfet_CDNS_524688791851170  pfet_CDNS_524688791851170_1
timestamp 1704896540
transform 1 0 540 0 -1 1161
box -89 -36 289 236
use pfet_CDNS_524688791851171  pfet_CDNS_524688791851171_0
timestamp 1704896540
transform 1 0 28 0 -1 1161
box -89 -36 545 236
use pfet_CDNS_524688791851171  pfet_CDNS_524688791851171_1
timestamp 1704896540
transform 1 0 1162 0 -1 1161
box -89 -36 545 236
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_0
timestamp 1704896540
transform -1 0 712 0 1 51
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_1
timestamp 1704896540
transform -1 0 1064 0 1 51
box 0 0 1 1
use PYL1_CDNS_52468879185289  PYL1_CDNS_52468879185289_0
timestamp 1704896540
transform 0 -1 1339 1 0 817
box 0 0 1 1
use PYL1_CDNS_52468879185327  PYL1_CDNS_52468879185327_0
timestamp 1704896540
transform 0 -1 713 1 0 817
box 0 0 1 1
<< properties >>
string GDS_END 85524846
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85517018
string path 0.375 30.800 40.775 30.800 
<< end >>
