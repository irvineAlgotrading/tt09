magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -66 377 738 897
<< pwell >>
rect 4 43 668 299
rect -26 -43 698 43
<< mvnmos >>
rect 87 189 187 273
rect 313 123 413 273
rect 485 123 585 273
<< mvpmos >>
rect 137 443 237 593
rect 313 443 413 743
rect 485 443 585 743
<< mvndiff >>
rect 30 248 87 273
rect 30 214 42 248
rect 76 214 87 248
rect 30 189 87 214
rect 187 265 313 273
rect 187 248 268 265
rect 187 214 198 248
rect 232 231 268 248
rect 302 231 313 265
rect 232 214 313 231
rect 187 189 313 214
rect 256 165 313 189
rect 256 131 268 165
rect 302 131 313 165
rect 256 123 313 131
rect 413 123 485 273
rect 585 265 642 273
rect 585 231 596 265
rect 630 231 642 265
rect 585 165 642 231
rect 585 131 596 165
rect 630 131 642 165
rect 585 123 642 131
<< mvpdiff >>
rect 256 735 313 743
rect 256 701 268 735
rect 302 701 313 735
rect 256 654 313 701
rect 256 620 268 654
rect 302 620 313 654
rect 256 593 313 620
rect 80 585 137 593
rect 80 551 92 585
rect 126 551 137 585
rect 80 485 137 551
rect 80 451 92 485
rect 126 451 137 485
rect 80 443 137 451
rect 237 571 313 593
rect 237 537 268 571
rect 302 537 313 571
rect 237 490 313 537
rect 237 456 268 490
rect 302 456 313 490
rect 237 443 313 456
rect 413 443 485 743
rect 585 735 642 743
rect 585 701 596 735
rect 630 701 642 735
rect 585 652 642 701
rect 585 618 596 652
rect 630 618 642 652
rect 585 568 642 618
rect 585 534 596 568
rect 630 534 642 568
rect 585 485 642 534
rect 585 451 596 485
rect 630 451 642 485
rect 585 443 642 451
<< mvndiffc >>
rect 42 214 76 248
rect 198 214 232 248
rect 268 231 302 265
rect 268 131 302 165
rect 596 231 630 265
rect 596 131 630 165
<< mvpdiffc >>
rect 268 701 302 735
rect 268 620 302 654
rect 92 551 126 585
rect 92 451 126 485
rect 268 537 302 571
rect 268 456 302 490
rect 596 701 630 735
rect 596 618 630 652
rect 596 534 630 568
rect 596 451 630 485
<< mvpsubdiff >>
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 672 831
<< mvpsubdiffcont >>
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
<< poly >>
rect 313 743 413 769
rect 485 743 585 769
rect 137 593 237 619
rect 137 417 237 443
rect 313 421 413 443
rect 87 349 237 417
rect 87 315 119 349
rect 153 315 187 349
rect 221 315 237 349
rect 279 395 413 421
rect 279 361 295 395
rect 329 361 363 395
rect 397 361 413 395
rect 485 391 585 443
rect 279 341 413 361
rect 455 375 589 391
rect 455 341 471 375
rect 505 341 539 375
rect 573 341 589 375
rect 455 325 589 341
rect 87 299 237 315
rect 87 273 187 299
rect 313 273 413 299
rect 485 273 585 325
rect 87 101 187 189
rect 313 101 413 123
rect 87 28 413 101
rect 485 97 585 123
<< polycont >>
rect 119 315 153 349
rect 187 315 221 349
rect 295 361 329 395
rect 363 361 397 395
rect 471 341 505 375
rect 539 341 573 375
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 672 831
rect 166 735 560 751
rect 200 701 238 735
rect 302 701 310 735
rect 344 701 382 735
rect 416 701 454 735
rect 488 701 526 735
rect 166 654 560 701
rect 166 620 268 654
rect 302 620 560 654
rect 35 585 130 601
rect 35 551 92 585
rect 126 551 130 585
rect 35 485 130 551
rect 35 451 92 485
rect 126 451 130 485
rect 166 571 560 620
rect 166 537 268 571
rect 302 542 560 571
rect 596 735 647 751
rect 630 701 647 735
rect 596 652 647 701
rect 630 618 647 652
rect 596 568 647 618
rect 302 537 455 542
rect 166 490 455 537
rect 630 534 647 568
rect 166 456 268 490
rect 302 456 455 490
rect 35 420 130 451
rect 35 395 413 420
rect 35 386 295 395
rect 35 267 69 386
rect 329 361 363 395
rect 397 361 413 395
rect 489 391 562 508
rect 596 485 647 534
rect 630 451 647 485
rect 596 425 647 451
rect 103 349 261 350
rect 103 315 119 349
rect 153 315 187 349
rect 221 315 261 349
rect 295 345 413 361
rect 455 375 573 391
rect 455 341 471 375
rect 505 341 539 375
rect 455 325 573 341
rect 103 301 261 315
rect 35 248 76 267
rect 35 214 42 248
rect 35 181 76 214
rect 110 265 455 267
rect 110 248 268 265
rect 110 214 198 248
rect 232 231 268 248
rect 302 231 455 265
rect 489 232 562 325
rect 607 291 647 425
rect 596 265 647 291
rect 232 214 455 231
rect 110 198 455 214
rect 630 231 647 265
rect 110 165 560 198
rect 110 147 268 165
rect 94 131 268 147
rect 302 131 560 165
rect 94 113 560 131
rect 596 165 647 231
rect 630 131 647 165
rect 596 115 647 131
rect 128 79 166 113
rect 200 79 238 113
rect 272 79 310 113
rect 344 79 382 113
rect 416 79 454 113
rect 488 79 526 113
rect 94 73 560 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 166 701 200 735
rect 238 701 268 735
rect 268 701 272 735
rect 310 701 344 735
rect 382 701 416 735
rect 454 701 488 735
rect 526 701 560 735
rect 94 79 128 113
rect 166 79 200 113
rect 238 79 272 113
rect 310 79 344 113
rect 382 79 416 113
rect 454 79 488 113
rect 526 79 560 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 831 672 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 672 831
rect 0 791 672 797
rect 0 735 672 763
rect 0 701 166 735
rect 200 701 238 735
rect 272 701 310 735
rect 344 701 382 735
rect 416 701 454 735
rect 488 701 526 735
rect 560 701 672 735
rect 0 689 672 701
rect 0 113 672 125
rect 0 79 94 113
rect 128 79 166 113
rect 200 79 238 113
rect 272 79 310 113
rect 344 79 382 113
rect 416 79 454 113
rect 488 79 526 113
rect 560 79 672 113
rect 0 51 672 79
rect 0 17 672 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -23 672 -17
<< labels >>
rlabel comment s 0 0 0 0 4 einvp_1
flabel metal1 s 0 51 672 125 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel metal1 s 0 0 672 23 0 FreeSans 340 0 0 0 VNB
port 4 nsew ground bidirectional
flabel metal1 s 0 689 672 763 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 791 672 814 0 FreeSans 340 0 0 0 VPB
port 5 nsew power bidirectional
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 TE
port 2 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 TE
port 2 nsew signal input
flabel locali s 607 168 641 202 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 607 464 641 498 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 607 538 641 572 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 607 612 641 646 0 FreeSans 340 0 0 0 Z
port 7 nsew signal output
flabel locali s 511 242 545 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 511 464 545 498 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 672 814
string GDS_END 1239596
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 1230040
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
<< end >>
