magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -89 -36 245 236
<< pmos >>
rect 0 0 50 200
rect 106 0 156 200
<< pdiff >>
rect -50 0 0 200
rect 50 182 106 200
rect 50 148 61 182
rect 95 148 106 182
rect 50 114 106 148
rect 50 80 61 114
rect 95 80 106 114
rect 50 46 106 80
rect 50 12 61 46
rect 95 12 106 46
rect 50 0 106 12
rect 156 182 209 200
rect 156 148 167 182
rect 201 148 209 182
rect 156 114 209 148
rect 156 80 167 114
rect 201 80 209 114
rect 156 46 209 80
rect 156 12 167 46
rect 201 12 209 46
rect 156 0 209 12
<< pdiffc >>
rect 61 148 95 182
rect 61 80 95 114
rect 61 12 95 46
rect 167 148 201 182
rect 167 80 201 114
rect 167 12 201 46
<< poly >>
rect 0 200 50 226
rect 106 200 156 226
rect 0 -26 50 0
rect 106 -26 156 0
<< locali >>
rect 61 182 95 198
rect 61 114 95 148
rect 61 46 95 80
rect 61 -4 95 12
rect 167 182 201 198
rect 167 114 201 148
rect 167 46 201 80
rect 167 -4 201 12
<< metal1 >>
rect -51 -16 -5 186
use DFL1sd2_CDNS_52468879185419  DFL1sd2_CDNS_52468879185419_0
timestamp 1704896540
transform 1 0 50 0 1 0
box 0 0 1 1
use DFL1sd_CDNS_5246887918529  DFL1sd_CDNS_5246887918529_0
timestamp 1704896540
transform 1 0 156 0 1 0
box 0 0 1 1
use DFM1sd_CDNS_524688791851377  DFM1sd_CDNS_524688791851377_0
timestamp 1704896540
transform -1 0 0 0 1 0
box -36 -36 89 236
<< labels >>
flabel comment s -28 85 -28 85 0 FreeSans 300 0 0 0 S
flabel comment s 78 97 78 97 0 FreeSans 300 0 0 0 D
flabel comment s 184 97 184 97 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 85950364
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85948978
<< end >>
