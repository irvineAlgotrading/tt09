magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -66 377 160 1251
rect 560 403 1054 863
rect 1454 493 2178 1251
rect 1960 377 2178 493
<< pwell >>
rect -26 1585 2138 1671
rect 668 1195 1394 1585
rect 1850 1345 2108 1585
rect 1174 317 1900 433
rect 600 43 1900 317
rect -26 -43 2138 43
<< locali >>
rect 0 1611 2112 1645
rect 0 797 160 831
rect 499 306 561 440
rect 2024 881 2090 1525
rect 1743 797 2112 831
rect 0 -17 2112 17
<< obsli1 >>
rect 660 1543 1402 1577
rect 660 1217 778 1543
rect 842 1199 908 1509
rect 972 1233 1090 1543
rect 1154 1199 1220 1509
rect 1284 1233 1402 1543
rect 1842 1367 1960 1549
rect 842 1133 1586 1199
rect 618 1033 1132 1099
rect 618 399 684 1033
rect 718 671 956 805
rect 1520 787 1586 1133
rect 1727 1107 1793 1311
rect 1643 1041 1793 1107
rect 1475 721 1609 787
rect 748 465 866 671
rect 1520 625 1586 687
rect 1643 625 1709 1041
rect 1842 960 1960 1189
rect 1758 881 1960 960
rect 930 495 996 623
rect 1520 559 1709 625
rect 1788 559 1906 741
rect 1643 495 1709 559
rect 930 433 1314 495
rect 1066 429 1314 433
rect 1348 429 1726 495
rect 618 349 969 399
rect 618 137 684 349
rect 1066 295 1132 429
rect 748 85 866 295
rect 930 229 1132 295
rect 930 137 996 229
rect 1166 85 1284 395
rect 1348 119 1414 429
rect 1478 85 1596 395
rect 1660 119 1726 429
rect 1790 85 1908 395
rect 748 51 1908 85
<< metal1 >>
rect 0 1605 2112 1651
rect 0 1503 2112 1577
rect 0 865 2112 939
rect 0 791 2112 837
rect 0 689 2112 763
rect 14 604 2098 661
rect 0 51 2112 125
rect 0 -23 2112 23
<< labels >>
rlabel locali s 499 306 561 440 6 A
port 1 nsew signal input
rlabel metal1 s 14 604 2098 661 6 LOWHVPWR
port 2 nsew power bidirectional
rlabel nwell s 560 403 1054 863 6 LOWHVPWR
port 2 nsew power bidirectional
rlabel metal1 s 0 1503 2112 1577 6 VGND
port 3 nsew ground bidirectional
rlabel metal1 s 0 51 2112 125 6 VGND
port 3 nsew ground bidirectional
rlabel metal1 s 0 -23 2112 23 8 VNB
port 4 nsew ground bidirectional
rlabel pwell s -26 -43 2138 43 8 VNB
port 4 nsew ground bidirectional
rlabel pwell s 600 43 1900 317 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 1174 317 1900 433 6 VNB
port 4 nsew ground bidirectional
rlabel metal1 s 0 1605 2112 1651 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 1850 1345 2108 1585 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 668 1195 1394 1585 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s -26 1585 2138 1671 6 VNB
port 4 nsew ground bidirectional
rlabel locali s 0 1611 2112 1645 6 VNB
port 4 nsew ground bidirectional
rlabel locali s 0 -17 2112 17 8 VNB
port 4 nsew ground bidirectional
rlabel metal1 s 0 791 2112 837 6 VPB
port 5 nsew power bidirectional
rlabel nwell s 1960 377 2178 493 6 VPB
port 5 nsew power bidirectional
rlabel nwell s 1454 493 2178 1251 6 VPB
port 5 nsew power bidirectional
rlabel nwell s -66 377 160 1251 6 VPB
port 5 nsew power bidirectional
rlabel locali s 1743 797 2112 831 6 VPB
port 5 nsew power bidirectional
rlabel locali s 0 797 160 831 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 865 2112 939 6 VPWR
port 6 nsew power bidirectional
rlabel metal1 s 0 689 2112 763 6 VPWR
port 6 nsew power bidirectional
rlabel locali s 2024 881 2090 1525 6 X
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2112 1628
string LEFclass CORE
string LEFsite unithvdbl
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 167916
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 146448
<< end >>
