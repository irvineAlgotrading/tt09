magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< pwell >>
rect -68 -26 1748 92
<< ndiff >>
rect -42 50 0 66
rect -42 16 -34 50
rect -42 0 0 16
rect 1680 50 1722 66
rect 1714 16 1722 50
rect 1680 0 1722 16
<< ndiffc >>
rect -34 16 0 50
rect 1680 16 1714 50
<< ndiffres >>
rect 0 0 1680 66
<< locali >>
rect -34 50 0 66
rect -34 0 0 16
rect 1680 50 1714 66
rect 1680 0 1714 16
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_0
timestamp 1704896540
transform -1 0 8 0 1 4
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_1
timestamp 1704896540
transform 1 0 1672 0 1 4
box 0 0 1 1
<< properties >>
string GDS_END 86217574
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86217072
<< end >>
