magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -119 -66 975 266
<< mvpmos >>
rect 0 0 400 200
rect 456 0 856 200
<< mvpdiff >>
rect -53 182 0 200
rect -53 148 -45 182
rect -11 148 0 182
rect -53 114 0 148
rect -53 80 -45 114
rect -11 80 0 114
rect -53 46 0 80
rect -53 12 -45 46
rect -11 12 0 46
rect -53 0 0 12
rect 400 182 456 200
rect 400 148 411 182
rect 445 148 456 182
rect 400 114 456 148
rect 400 80 411 114
rect 445 80 456 114
rect 400 46 456 80
rect 400 12 411 46
rect 445 12 456 46
rect 400 0 456 12
rect 856 182 909 200
rect 856 148 867 182
rect 901 148 909 182
rect 856 114 909 148
rect 856 80 867 114
rect 901 80 909 114
rect 856 46 909 80
rect 856 12 867 46
rect 901 12 909 46
rect 856 0 909 12
<< mvpdiffc >>
rect -45 148 -11 182
rect -45 80 -11 114
rect -45 12 -11 46
rect 411 148 445 182
rect 411 80 445 114
rect 411 12 445 46
rect 867 148 901 182
rect 867 80 901 114
rect 867 12 901 46
<< poly >>
rect 0 200 400 232
rect 456 200 856 232
rect 0 -32 400 0
rect 456 -32 856 0
<< locali >>
rect -45 182 -11 198
rect -45 114 -11 148
rect -45 46 -11 80
rect -45 -4 -11 12
rect 411 182 445 198
rect 411 114 445 148
rect 411 46 445 80
rect 411 -4 445 12
rect 867 182 901 198
rect 867 114 901 148
rect 867 46 901 80
rect 867 -4 901 12
use DFL1sd2_CDNS_52468879185419  DFL1sd2_CDNS_52468879185419_0
timestamp 1704896540
transform 1 0 400 0 1 0
box 0 0 1 1
use DFL1sd_CDNS_5246887918529  DFL1sd_CDNS_5246887918529_0
timestamp 1704896540
transform -1 0 0 0 1 0
box 0 0 1 1
use DFL1sd_CDNS_5246887918529  DFL1sd_CDNS_5246887918529_1
timestamp 1704896540
transform 1 0 856 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s -28 97 -28 97 0 FreeSans 300 0 0 0 S
flabel comment s 428 97 428 97 0 FreeSans 300 0 0 0 D
flabel comment s 884 97 884 97 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 6682394
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 6680882
<< end >>
