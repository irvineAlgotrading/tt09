magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -119 -66 1311 266
<< mvpmos >>
rect 0 0 100 200
rect 156 0 256 200
rect 312 0 412 200
rect 468 0 568 200
rect 624 0 724 200
rect 780 0 880 200
rect 936 0 1036 200
rect 1092 0 1192 200
<< mvpdiff >>
rect -53 182 0 200
rect -53 148 -45 182
rect -11 148 0 182
rect -53 114 0 148
rect -53 80 -45 114
rect -11 80 0 114
rect -53 46 0 80
rect -53 12 -45 46
rect -11 12 0 46
rect -53 0 0 12
rect 100 182 156 200
rect 100 148 111 182
rect 145 148 156 182
rect 100 114 156 148
rect 100 80 111 114
rect 145 80 156 114
rect 100 46 156 80
rect 100 12 111 46
rect 145 12 156 46
rect 100 0 156 12
rect 256 182 312 200
rect 256 148 267 182
rect 301 148 312 182
rect 256 114 312 148
rect 256 80 267 114
rect 301 80 312 114
rect 256 46 312 80
rect 256 12 267 46
rect 301 12 312 46
rect 256 0 312 12
rect 412 182 468 200
rect 412 148 423 182
rect 457 148 468 182
rect 412 114 468 148
rect 412 80 423 114
rect 457 80 468 114
rect 412 46 468 80
rect 412 12 423 46
rect 457 12 468 46
rect 412 0 468 12
rect 568 182 624 200
rect 568 148 579 182
rect 613 148 624 182
rect 568 114 624 148
rect 568 80 579 114
rect 613 80 624 114
rect 568 46 624 80
rect 568 12 579 46
rect 613 12 624 46
rect 568 0 624 12
rect 724 182 780 200
rect 724 148 735 182
rect 769 148 780 182
rect 724 114 780 148
rect 724 80 735 114
rect 769 80 780 114
rect 724 46 780 80
rect 724 12 735 46
rect 769 12 780 46
rect 724 0 780 12
rect 880 182 936 200
rect 880 148 891 182
rect 925 148 936 182
rect 880 114 936 148
rect 880 80 891 114
rect 925 80 936 114
rect 880 46 936 80
rect 880 12 891 46
rect 925 12 936 46
rect 880 0 936 12
rect 1036 182 1092 200
rect 1036 148 1047 182
rect 1081 148 1092 182
rect 1036 114 1092 148
rect 1036 80 1047 114
rect 1081 80 1092 114
rect 1036 46 1092 80
rect 1036 12 1047 46
rect 1081 12 1092 46
rect 1036 0 1092 12
rect 1192 182 1245 200
rect 1192 148 1203 182
rect 1237 148 1245 182
rect 1192 114 1245 148
rect 1192 80 1203 114
rect 1237 80 1245 114
rect 1192 46 1245 80
rect 1192 12 1203 46
rect 1237 12 1245 46
rect 1192 0 1245 12
<< mvpdiffc >>
rect -45 148 -11 182
rect -45 80 -11 114
rect -45 12 -11 46
rect 111 148 145 182
rect 111 80 145 114
rect 111 12 145 46
rect 267 148 301 182
rect 267 80 301 114
rect 267 12 301 46
rect 423 148 457 182
rect 423 80 457 114
rect 423 12 457 46
rect 579 148 613 182
rect 579 80 613 114
rect 579 12 613 46
rect 735 148 769 182
rect 735 80 769 114
rect 735 12 769 46
rect 891 148 925 182
rect 891 80 925 114
rect 891 12 925 46
rect 1047 148 1081 182
rect 1047 80 1081 114
rect 1047 12 1081 46
rect 1203 148 1237 182
rect 1203 80 1237 114
rect 1203 12 1237 46
<< poly >>
rect 0 200 100 252
rect 156 200 256 252
rect 312 200 412 252
rect 468 200 568 252
rect 624 200 724 252
rect 780 200 880 252
rect 936 200 1036 252
rect 1092 200 1192 252
rect 0 -52 100 0
rect 156 -52 256 0
rect 312 -52 412 0
rect 468 -52 568 0
rect 624 -52 724 0
rect 780 -52 880 0
rect 936 -52 1036 0
rect 1092 -52 1192 0
<< locali >>
rect -45 182 -11 198
rect -45 114 -11 148
rect -45 46 -11 80
rect -45 -4 -11 12
rect 111 182 145 198
rect 111 114 145 148
rect 111 46 145 80
rect 111 -4 145 12
rect 267 182 301 198
rect 267 114 301 148
rect 267 46 301 80
rect 267 -4 301 12
rect 423 182 457 198
rect 423 114 457 148
rect 423 46 457 80
rect 423 -4 457 12
rect 579 182 613 198
rect 579 114 613 148
rect 579 46 613 80
rect 579 -4 613 12
rect 735 182 769 198
rect 735 114 769 148
rect 735 46 769 80
rect 735 -4 769 12
rect 891 182 925 198
rect 891 114 925 148
rect 891 46 925 80
rect 891 -4 925 12
rect 1047 182 1081 198
rect 1047 114 1081 148
rect 1047 46 1081 80
rect 1047 -4 1081 12
rect 1203 182 1237 198
rect 1203 114 1237 148
rect 1203 46 1237 80
rect 1203 -4 1237 12
use DFL1sd_CDNS_5246887918529  DFL1sd_CDNS_5246887918529_0
timestamp 1704896540
transform 1 0 1192 0 1 0
box 0 0 1 1
use hvDFL1sd2_CDNS_52468879185110  hvDFL1sd2_CDNS_52468879185110_0
timestamp 1704896540
transform 1 0 1036 0 1 0
box 0 0 1 1
use hvDFL1sd2_CDNS_52468879185110  hvDFL1sd2_CDNS_52468879185110_1
timestamp 1704896540
transform 1 0 880 0 1 0
box 0 0 1 1
use hvDFL1sd2_CDNS_52468879185110  hvDFL1sd2_CDNS_52468879185110_2
timestamp 1704896540
transform 1 0 724 0 1 0
box 0 0 1 1
use hvDFL1sd2_CDNS_52468879185110  hvDFL1sd2_CDNS_52468879185110_3
timestamp 1704896540
transform 1 0 568 0 1 0
box 0 0 1 1
use hvDFL1sd2_CDNS_52468879185110  hvDFL1sd2_CDNS_52468879185110_4
timestamp 1704896540
transform 1 0 412 0 1 0
box 0 0 1 1
use hvDFL1sd2_CDNS_52468879185110  hvDFL1sd2_CDNS_52468879185110_5
timestamp 1704896540
transform 1 0 256 0 1 0
box 0 0 1 1
use hvDFL1sd2_CDNS_52468879185110  hvDFL1sd2_CDNS_52468879185110_6
timestamp 1704896540
transform 1 0 100 0 1 0
box 0 0 1 1
use hvDFL1sd_CDNS_5246887918589  hvDFL1sd_CDNS_5246887918589_0
timestamp 1704896540
transform -1 0 0 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s -28 97 -28 97 0 FreeSans 300 0 0 0 S
flabel comment s 128 97 128 97 0 FreeSans 300 0 0 0 D
flabel comment s 284 97 284 97 0 FreeSans 300 0 0 0 S
flabel comment s 440 97 440 97 0 FreeSans 300 0 0 0 D
flabel comment s 596 97 596 97 0 FreeSans 300 0 0 0 S
flabel comment s 752 97 752 97 0 FreeSans 300 0 0 0 D
flabel comment s 908 97 908 97 0 FreeSans 300 0 0 0 S
flabel comment s 1064 97 1064 97 0 FreeSans 300 0 0 0 D
flabel comment s 1220 97 1220 97 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 80249060
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 80244544
<< end >>
