magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 1 21 643 203
rect 30 -17 64 21
<< locali >>
rect 106 51 155 493
rect 289 202 371 323
rect 481 280 522 397
rect 405 205 522 280
rect 573 199 625 290
<< obsli1 >>
rect 0 527 644 561
rect 18 327 69 527
rect 21 17 69 177
rect 189 437 359 527
rect 393 401 445 493
rect 221 357 445 401
rect 221 266 255 357
rect 189 168 255 266
rect 559 330 624 527
rect 189 127 359 168
rect 189 17 255 93
rect 293 51 359 127
rect 393 127 624 165
rect 393 93 435 127
rect 569 99 624 127
rect 469 17 535 93
rect 0 -17 644 17
<< metal1 >>
rect 0 496 644 592
rect 0 -48 644 48
<< labels >>
rlabel locali s 573 199 625 290 6 A1
port 1 nsew signal input
rlabel locali s 405 205 522 280 6 A2
port 2 nsew signal input
rlabel locali s 481 280 522 397 6 A2
port 2 nsew signal input
rlabel locali s 289 202 371 323 6 B1
port 3 nsew signal input
rlabel metal1 s 0 -48 644 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 21 643 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 682 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 644 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 106 51 155 493 6 X
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 644 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1271234
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1265726
<< end >>
