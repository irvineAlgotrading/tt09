magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< metal2 >>
rect 0 785 136 794
rect 0 0 136 9
<< via2 >>
rect 0 9 136 785
<< metal3 >>
rect -5 785 141 790
rect -5 9 0 785
rect 136 9 141 785
rect -5 4 141 9
<< properties >>
string GDS_END 85412056
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85410644
<< end >>
