magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect 13240 3885 14184 4064
rect 13240 3337 14621 3885
rect 12841 3307 14621 3337
rect 12462 3128 14621 3307
rect 12462 3079 14126 3128
rect 13240 2414 14126 3079
rect 8777 912 8943 1644
<< pwell >>
rect 10107 2074 10193 2186
rect 11043 2074 11129 2186
<< mvpsubdiff >>
rect 10133 2100 10167 2160
rect 11069 2100 11103 2160
<< mvnsubdiff >>
rect 12528 3210 13058 3241
rect 12528 3176 12552 3210
rect 12586 3176 12627 3210
rect 12661 3176 12702 3210
rect 12736 3176 12777 3210
rect 12811 3176 12852 3210
rect 12886 3176 12926 3210
rect 12960 3176 13000 3210
rect 13034 3176 13058 3210
rect 12528 3145 13058 3176
rect 8843 1554 8877 1578
rect 8843 1480 8877 1520
rect 8843 1406 8877 1446
rect 8843 1332 8877 1372
rect 8843 1258 8877 1298
rect 8843 1184 8877 1224
rect 8843 1110 8877 1150
rect 8843 1036 8877 1076
rect 8843 978 8877 1002
<< mvnsubdiffcont >>
rect 12552 3176 12586 3210
rect 12627 3176 12661 3210
rect 12702 3176 12736 3210
rect 12777 3176 12811 3210
rect 12852 3176 12886 3210
rect 12926 3176 12960 3210
rect 13000 3176 13034 3210
rect 8843 1520 8877 1554
rect 8843 1446 8877 1480
rect 8843 1372 8877 1406
rect 8843 1298 8877 1332
rect 8843 1224 8877 1258
rect 8843 1150 8877 1184
rect 8843 1076 8877 1110
rect 8843 1002 8877 1036
<< poly >>
rect 14345 3531 14479 3547
rect 14345 3497 14361 3531
rect 14395 3497 14429 3531
rect 14463 3497 14479 3531
rect 14345 3481 14479 3497
rect 13809 3299 14065 3315
rect 13809 3265 13825 3299
rect 13859 3265 13920 3299
rect 13954 3265 14015 3299
rect 14049 3265 14065 3299
rect 13809 3249 14065 3265
rect 13359 3161 14007 3177
rect 13359 3127 13375 3161
rect 13409 3127 13447 3161
rect 13481 3127 13519 3161
rect 13553 3127 13592 3161
rect 13626 3127 13665 3161
rect 13699 3127 13738 3161
rect 13772 3127 13811 3161
rect 13845 3127 13884 3161
rect 13918 3127 13957 3161
rect 13991 3127 14007 3161
rect 13359 3111 14007 3127
rect 14267 3136 14387 3169
rect 14267 3102 14305 3136
rect 14339 3102 14387 3136
rect 14267 3068 14387 3102
rect 14267 3034 14305 3068
rect 14339 3034 14387 3068
rect 14267 3001 14387 3034
rect 14443 3136 14563 3169
rect 14443 3102 14491 3136
rect 14525 3102 14563 3136
rect 14443 3068 14563 3102
rect 14443 3034 14491 3068
rect 14525 3034 14563 3068
rect 14443 3001 14563 3034
rect 13112 2924 13188 2940
rect 13112 2890 13138 2924
rect 13172 2890 13188 2924
rect 13112 2848 13188 2890
rect 13112 2814 13138 2848
rect 13172 2814 13188 2848
rect 13112 2771 13188 2814
rect 13112 2737 13138 2771
rect 13172 2737 13188 2771
rect 13112 2694 13188 2737
rect 13112 2660 13138 2694
rect 13172 2660 13188 2694
rect 13112 2644 13188 2660
rect 14267 2671 14401 2687
rect 14267 2637 14283 2671
rect 14317 2637 14351 2671
rect 14385 2637 14401 2671
rect 14267 2621 14401 2637
rect 13112 2572 13188 2588
rect 13112 2538 13138 2572
rect 13172 2538 13188 2572
rect 13112 2492 13188 2538
rect 14315 2546 14449 2562
rect 14315 2512 14331 2546
rect 14365 2512 14399 2546
rect 14433 2512 14449 2546
rect 14315 2496 14449 2512
rect 13112 2488 13138 2492
rect 13122 2458 13138 2488
rect 13172 2458 13188 2492
rect 13122 2442 13188 2458
rect 10294 2126 10414 2134
rect 10470 2126 10590 2134
rect 10646 2126 10766 2134
rect 10822 2126 10942 2134
rect 9018 1728 9138 1814
rect 9018 1694 9061 1728
rect 9095 1694 9138 1728
rect 9018 1660 9138 1694
rect 9018 1626 9061 1660
rect 9095 1626 9138 1660
rect 9018 1604 9138 1626
rect 9194 1728 9314 1814
rect 9194 1694 9237 1728
rect 9271 1694 9314 1728
rect 9194 1660 9314 1694
rect 9194 1626 9237 1660
rect 9271 1626 9314 1660
rect 9194 1604 9314 1626
rect 9398 1728 9518 1814
rect 9398 1694 9414 1728
rect 9448 1694 9518 1728
rect 9398 1660 9518 1694
rect 9398 1626 9414 1660
rect 9448 1626 9518 1660
rect 9398 1604 9518 1626
rect 9865 220 9921 292
<< polycont >>
rect 14361 3497 14395 3531
rect 14429 3497 14463 3531
rect 13825 3265 13859 3299
rect 13920 3265 13954 3299
rect 14015 3265 14049 3299
rect 13375 3127 13409 3161
rect 13447 3127 13481 3161
rect 13519 3127 13553 3161
rect 13592 3127 13626 3161
rect 13665 3127 13699 3161
rect 13738 3127 13772 3161
rect 13811 3127 13845 3161
rect 13884 3127 13918 3161
rect 13957 3127 13991 3161
rect 14305 3102 14339 3136
rect 14305 3034 14339 3068
rect 14491 3102 14525 3136
rect 14491 3034 14525 3068
rect 13138 2890 13172 2924
rect 13138 2814 13172 2848
rect 13138 2737 13172 2771
rect 13138 2660 13172 2694
rect 14283 2637 14317 2671
rect 14351 2637 14385 2671
rect 13138 2538 13172 2572
rect 14331 2512 14365 2546
rect 14399 2512 14433 2546
rect 13138 2458 13172 2492
rect 9061 1694 9095 1728
rect 9061 1626 9095 1660
rect 9237 1694 9271 1728
rect 9237 1626 9271 1660
rect 9414 1694 9448 1728
rect 9414 1626 9448 1660
<< locali >>
rect 14304 4029 14697 4047
rect 14304 3995 14315 4029
rect 14349 3995 14417 4029
rect 14451 3995 14697 4029
rect 10043 3692 10173 3906
rect 10043 3658 10055 3692
rect 10089 3658 10127 3692
rect 10161 3658 10173 3692
rect 10300 3538 10371 3906
rect 13764 3765 13798 3826
rect 13764 3671 13798 3731
rect 14076 3765 14110 3826
rect 13764 3577 13798 3637
rect 13920 3577 13954 3638
rect 14076 3671 14110 3731
rect 14076 3577 14110 3637
rect 10334 3504 10372 3538
rect 13920 3483 13954 3543
rect 13920 3389 13954 3449
rect 12528 3210 13058 3303
rect 13809 3265 13825 3299
rect 13859 3265 13886 3299
rect 13954 3265 14015 3299
rect 14053 3265 14065 3299
rect 12528 3176 12552 3210
rect 12586 3176 12627 3210
rect 12661 3176 12702 3210
rect 12736 3176 12777 3210
rect 12811 3176 12852 3210
rect 12886 3176 12926 3210
rect 12960 3176 13000 3210
rect 13034 3176 13058 3210
rect 12528 3149 13058 3176
rect 13359 3159 13375 3161
rect 12528 3115 12651 3149
rect 12685 3115 12723 3149
rect 12757 3115 13058 3149
rect 13135 3127 13375 3159
rect 13409 3127 13447 3161
rect 13481 3127 13519 3161
rect 13553 3127 13592 3161
rect 13626 3127 13665 3161
rect 13699 3127 13738 3161
rect 13772 3127 13811 3161
rect 13845 3127 13884 3161
rect 13918 3157 13957 3161
rect 13991 3157 14007 3161
rect 13923 3127 13957 3157
rect 13135 3123 13889 3127
rect 13923 3123 13961 3127
rect 13995 3123 14007 3157
rect 13135 3119 14007 3123
rect 14146 3152 14186 3989
rect 14304 3976 14697 3995
rect 14315 3695 14349 3733
rect 14516 3596 14554 3630
rect 14379 3531 14417 3537
rect 14395 3503 14417 3531
rect 14345 3497 14361 3503
rect 14395 3497 14429 3503
rect 14463 3497 14479 3531
rect 14222 3384 14256 3423
rect 14222 3311 14256 3350
rect 14573 3242 14607 3345
rect 14644 3152 14697 3976
rect 14146 3136 14339 3152
rect 12539 2945 12577 2979
rect 12611 2945 12650 2979
rect 12684 2945 12723 2979
rect 13135 2924 13175 3119
rect 14146 3102 14305 3136
rect 14146 3068 14339 3102
rect 13135 2890 13138 2924
rect 13172 2890 13175 2924
rect 13135 2848 13175 2890
rect 13314 2987 13348 3031
rect 13314 2909 13348 2953
rect 13666 2987 13700 3031
rect 13666 2909 13700 2953
rect 14018 2987 14052 3031
rect 14146 3034 14305 3068
rect 14146 3018 14339 3034
rect 14491 3136 14697 3152
rect 14525 3102 14697 3136
rect 14491 3068 14697 3102
rect 14525 3034 14697 3068
rect 14491 3018 14697 3034
rect 14018 2909 14052 2953
rect 14222 2911 14256 2949
rect 13135 2814 13138 2848
rect 13172 2814 13175 2848
rect 14383 2831 14447 2975
rect 12854 2776 12924 2810
rect 12958 2776 13028 2810
rect 13135 2771 13175 2814
rect 13135 2737 13138 2771
rect 13172 2737 13175 2771
rect 13135 2694 13175 2737
rect 14222 2754 14256 2792
rect 14383 2797 14400 2831
rect 14434 2797 14447 2831
rect 14383 2759 14447 2797
rect 14383 2725 14400 2759
rect 14434 2725 14447 2759
rect 14383 2713 14447 2725
rect 13135 2660 13138 2694
rect 13172 2660 13175 2694
rect 13135 2644 13175 2660
rect 12539 2599 12577 2633
rect 12611 2599 12650 2633
rect 12684 2599 12723 2633
rect 13491 2614 13525 2664
rect 13138 2572 13172 2588
rect 13138 2499 13172 2537
rect 13491 2529 13525 2580
rect 14614 2671 14697 3018
rect 13843 2614 13877 2664
rect 14267 2637 14283 2671
rect 14317 2637 14351 2671
rect 14385 2637 14697 2671
rect 14267 2622 14697 2637
rect 13843 2529 13877 2580
rect 14192 2548 14230 2582
rect 12844 2443 12882 2477
rect 12916 2443 12955 2477
rect 12989 2443 13028 2477
rect 13138 2442 13172 2458
rect 14158 2474 14264 2548
rect 14314 2546 14713 2579
rect 14314 2512 14331 2546
rect 14365 2512 14399 2546
rect 14433 2512 14713 2546
rect 14158 2368 14330 2474
rect 14452 2390 14486 2428
rect 14647 2353 14713 2512
rect 14647 2319 14669 2353
rect 14703 2319 14713 2353
rect 14647 2281 14713 2319
rect 14647 2247 14669 2281
rect 14703 2247 14713 2281
rect 14647 2235 14713 2247
rect 10133 2120 10167 2158
rect 11069 2120 11103 2158
rect 8959 1990 8993 2028
rect 9339 1990 9373 2028
rect 9149 1800 9183 1834
rect 8959 1766 9464 1800
rect 8843 1554 8877 1578
rect 8959 1553 8993 1766
rect 9398 1728 9464 1766
rect 9529 1738 9563 1836
rect 9045 1694 9061 1728
rect 9095 1694 9111 1728
rect 9045 1660 9111 1694
rect 9045 1656 9061 1660
rect 9095 1656 9111 1660
rect 9221 1694 9237 1728
rect 9271 1694 9287 1728
rect 9221 1660 9287 1694
rect 9221 1656 9237 1660
rect 9095 1626 9099 1656
rect 9061 1622 9099 1626
rect 9234 1626 9237 1656
rect 9271 1656 9287 1660
rect 9398 1694 9414 1728
rect 9448 1694 9464 1728
rect 9548 1704 9586 1738
rect 9398 1660 9464 1694
rect 9271 1626 9272 1656
rect 9234 1622 9272 1626
rect 9398 1626 9414 1660
rect 9448 1626 9464 1660
rect 9529 1556 9563 1704
rect 8843 1480 8877 1520
rect 8843 1406 8877 1446
rect 8993 1390 9031 1424
rect 8843 1332 8877 1372
rect 8843 1258 8877 1298
rect 8843 1184 8877 1224
rect 8843 1110 8877 1150
rect 8843 1051 8877 1076
rect 8843 979 8877 1002
rect 9339 979 9373 1017
rect 9758 725 9796 759
rect 9830 725 9842 759
rect 6410 267 6448 301
rect 9760 270 9842 725
rect 9865 236 9922 270
<< viali >>
rect 14315 3995 14349 4029
rect 14417 3995 14451 4029
rect 10055 3658 10089 3692
rect 10127 3658 10161 3692
rect 13764 3826 13798 3860
rect 13764 3731 13798 3765
rect 14076 3826 14110 3860
rect 14076 3731 14110 3765
rect 13764 3637 13798 3671
rect 13764 3543 13798 3577
rect 13920 3638 13954 3672
rect 13920 3543 13954 3577
rect 14076 3637 14110 3671
rect 14076 3543 14110 3577
rect 10300 3504 10334 3538
rect 10372 3504 10406 3538
rect 13920 3449 13954 3483
rect 13920 3355 13954 3389
rect 13886 3265 13920 3299
rect 14019 3265 14049 3299
rect 14049 3265 14053 3299
rect 12651 3115 12685 3149
rect 12723 3115 12757 3149
rect 13889 3127 13918 3157
rect 13918 3127 13923 3157
rect 13961 3127 13991 3157
rect 13991 3127 13995 3157
rect 13889 3123 13923 3127
rect 13961 3123 13995 3127
rect 14315 3733 14349 3767
rect 14315 3661 14349 3695
rect 14482 3596 14516 3630
rect 14554 3596 14588 3630
rect 14345 3531 14379 3537
rect 14417 3531 14451 3537
rect 14345 3503 14361 3531
rect 14361 3503 14379 3531
rect 14417 3503 14429 3531
rect 14429 3503 14451 3531
rect 14222 3423 14256 3457
rect 14222 3350 14256 3384
rect 14222 3277 14256 3311
rect 14573 3345 14607 3379
rect 14573 3208 14607 3242
rect 12505 2945 12539 2979
rect 12577 2945 12611 2979
rect 12650 2945 12684 2979
rect 12723 2945 12757 2979
rect 13314 3031 13348 3065
rect 13314 2953 13348 2987
rect 13314 2875 13348 2909
rect 13666 3031 13700 3065
rect 13666 2953 13700 2987
rect 13666 2875 13700 2909
rect 14018 3031 14052 3065
rect 14018 2953 14052 2987
rect 14018 2875 14052 2909
rect 14222 2949 14256 2983
rect 14222 2877 14256 2911
rect 12820 2776 12854 2810
rect 12924 2776 12958 2810
rect 13028 2776 13062 2810
rect 14222 2792 14256 2826
rect 14222 2720 14256 2754
rect 14400 2797 14434 2831
rect 14400 2725 14434 2759
rect 13491 2664 13525 2698
rect 12505 2599 12539 2633
rect 12577 2599 12611 2633
rect 12650 2599 12684 2633
rect 12723 2599 12757 2633
rect 13138 2538 13172 2571
rect 13138 2537 13172 2538
rect 13138 2492 13172 2499
rect 13491 2580 13525 2614
rect 13491 2495 13525 2529
rect 13843 2664 13877 2698
rect 13843 2580 13877 2614
rect 13843 2495 13877 2529
rect 14158 2548 14192 2582
rect 14230 2548 14264 2582
rect 12810 2443 12844 2477
rect 12882 2443 12916 2477
rect 12955 2443 12989 2477
rect 13028 2443 13062 2477
rect 13138 2465 13172 2492
rect 14452 2428 14486 2462
rect 14452 2356 14486 2390
rect 14669 2319 14703 2353
rect 14669 2247 14703 2281
rect 10133 2158 10167 2192
rect 10133 2086 10167 2120
rect 11069 2158 11103 2192
rect 11069 2086 11103 2120
rect 8959 2028 8993 2062
rect 8959 1956 8993 1990
rect 9339 2028 9373 2062
rect 9339 1956 9373 1990
rect 9027 1622 9061 1656
rect 9099 1622 9133 1656
rect 9200 1622 9234 1656
rect 9514 1704 9548 1738
rect 9586 1704 9620 1738
rect 9272 1622 9306 1656
rect 8959 1390 8993 1424
rect 9031 1390 9065 1424
rect 8843 1036 8877 1051
rect 8843 1017 8877 1036
rect 8843 945 8877 979
rect 9339 1017 9373 1051
rect 9339 945 9373 979
rect 9724 725 9758 759
rect 9796 725 9830 759
rect 6376 267 6410 301
rect 6448 267 6482 301
<< metal1 >>
rect 8847 4441 8877 4493
rect 8929 4441 8941 4493
rect 8993 4441 14375 4493
tri 14247 4413 14275 4441 ne
rect 14275 4413 14375 4441
rect 6994 4407 11490 4413
rect 7046 4361 11490 4407
rect 11491 4362 11492 4412
rect 11528 4362 11529 4412
rect 11530 4361 11618 4413
rect 11670 4361 11682 4413
rect 11734 4361 13607 4413
rect 13659 4361 13671 4413
rect 13723 4361 13729 4413
tri 14275 4385 14303 4413 ne
rect 6994 4342 7046 4355
rect 6994 4284 7046 4290
rect 8676 4327 11490 4333
rect 11492 4332 11528 4333
rect 8728 4281 11490 4327
rect 11491 4282 11529 4332
rect 11492 4281 11528 4282
rect 11530 4281 11618 4333
rect 11670 4281 11682 4333
rect 11734 4281 11791 4333
rect 11792 4282 11793 4332
rect 11829 4282 11830 4332
rect 11831 4281 11850 4333
rect 11902 4281 11914 4333
rect 11966 4289 12303 4333
tri 12303 4289 12347 4333 sw
rect 11966 4281 12347 4289
rect 8676 4263 8728 4275
tri 12270 4249 12302 4281 ne
rect 8676 4205 8728 4211
tri 12282 4092 12302 4112 se
rect 12302 4092 12347 4281
tri 11814 4089 11817 4092 se
tri 12281 4091 12282 4092 se
rect 12282 4091 12347 4092
tri 11947 4089 11949 4091 sw
tri 12279 4089 12281 4091 se
rect 12281 4089 12347 4091
tri 12277 4087 12279 4089 se
rect 12279 4087 12347 4089
tri 12347 4087 12399 4139 sw
rect 13601 4087 13607 4093
tri 11814 4040 11817 4043 ne
tri 11947 4041 11949 4043 nw
rect 13120 4041 13607 4087
rect 13659 4041 13671 4093
rect 13723 4041 13729 4093
rect 14303 4053 14375 4413
rect 14303 4029 14463 4053
rect 14303 3995 14315 4029
rect 14349 3995 14417 4029
rect 14451 3995 14463 4029
rect 8210 3959 8999 3987
rect 14303 3971 14463 3995
rect 151 3866 14355 3872
rect 151 3814 11699 3866
rect 11751 3814 12671 3866
rect 12723 3814 13701 3866
rect 13753 3860 13789 3866
rect 13841 3860 14355 3866
rect 13753 3826 13764 3860
rect 13841 3826 14076 3860
rect 14110 3826 14355 3860
rect 13753 3814 13789 3826
rect 13841 3814 14355 3826
rect 151 3784 14355 3814
rect 151 3732 11699 3784
rect 11751 3732 12671 3784
rect 12723 3732 13701 3784
rect 13753 3765 13789 3784
rect 13841 3767 14355 3784
rect 13841 3765 14315 3767
rect 13753 3732 13764 3765
rect 13841 3732 14076 3765
rect 151 3731 13764 3732
rect 13798 3731 14076 3732
rect 14110 3733 14315 3765
rect 14349 3733 14355 3767
rect 14110 3731 14355 3733
rect 151 3726 14355 3731
tri 13688 3698 13716 3726 ne
rect 13716 3698 13843 3726
rect 9735 3692 10173 3698
tri 13716 3695 13719 3698 ne
rect 13719 3695 13843 3698
tri 13843 3695 13874 3726 nw
tri 14000 3695 14031 3726 ne
rect 14031 3695 14355 3726
rect 9787 3658 10055 3692
rect 10089 3658 10127 3692
rect 10161 3658 10173 3692
tri 13719 3672 13742 3695 ne
rect 13742 3672 13820 3695
tri 13820 3672 13843 3695 nw
tri 14031 3684 14042 3695 ne
rect 14042 3684 14315 3695
rect 13914 3672 13960 3684
tri 13742 3671 13743 3672 ne
rect 13743 3671 13804 3672
rect 9787 3652 10173 3658
tri 13743 3656 13758 3671 ne
rect 9787 3640 9797 3652
rect 9735 3637 9797 3640
tri 9797 3637 9812 3652 nw
rect 13758 3637 13764 3671
rect 13798 3637 13804 3671
tri 13804 3656 13820 3672 nw
rect 9735 3630 9790 3637
tri 9790 3630 9797 3637 nw
rect 9735 3628 9787 3630
tri 9787 3627 9790 3630 nw
rect 9735 3570 9787 3576
rect 13758 3577 13804 3637
rect 9980 3498 9986 3550
rect 10038 3498 10050 3550
rect 10102 3538 10468 3550
rect 10102 3504 10300 3538
rect 10334 3504 10372 3538
rect 10406 3504 10468 3538
rect 13758 3543 13764 3577
rect 13798 3543 13804 3577
rect 13758 3531 13804 3543
rect 13914 3638 13920 3672
rect 13954 3638 13960 3672
tri 14042 3671 14055 3684 ne
rect 14055 3671 14315 3684
tri 14055 3656 14070 3671 ne
rect 13914 3577 13960 3638
rect 13914 3543 13920 3577
rect 13954 3543 13960 3577
rect 10102 3498 10468 3504
rect 13914 3503 13960 3543
rect 14070 3637 14076 3671
rect 14110 3661 14315 3671
rect 14349 3661 14355 3695
tri 14355 3693 14388 3726 nw
rect 14110 3649 14355 3661
rect 14110 3637 14133 3649
rect 14070 3630 14133 3637
tri 14133 3630 14152 3649 nw
tri 14187 3630 14206 3649 ne
rect 14206 3630 14282 3649
tri 14282 3630 14301 3649 nw
rect 14470 3630 14735 3636
rect 14070 3577 14116 3630
tri 14116 3613 14133 3630 nw
tri 14206 3620 14216 3630 ne
rect 14070 3543 14076 3577
rect 14110 3543 14116 3577
rect 14070 3531 14116 3543
tri 13960 3503 13981 3524 sw
rect 13521 3457 13558 3489
rect 13914 3483 13981 3503
rect 13914 3449 13920 3483
rect 13954 3457 13981 3483
tri 13981 3457 14027 3503 sw
rect 14216 3457 14262 3630
tri 14262 3610 14282 3630 nw
rect 14470 3596 14482 3630
rect 14516 3596 14554 3630
rect 14588 3596 14735 3630
rect 14470 3590 14735 3596
tri 14658 3559 14689 3590 ne
rect 13954 3454 14027 3457
tri 14027 3454 14030 3457 sw
rect 13954 3449 14178 3454
rect 13914 3448 14178 3449
tri 7522 3355 7537 3370 se
rect 7537 3355 8947 3370
tri 7517 3350 7522 3355 se
rect 7522 3350 8947 3355
tri 7512 3345 7517 3350 se
rect 7517 3345 8947 3350
rect 13113 3346 13119 3398
rect 13171 3346 13183 3398
rect 13235 3346 13241 3398
rect 13914 3396 14126 3448
rect 13914 3389 14178 3396
rect 13914 3355 13920 3389
rect 13954 3384 14178 3389
rect 13954 3355 14126 3384
tri 7478 3311 7512 3345 se
rect 7512 3318 8947 3345
rect 13914 3343 14126 3355
tri 14109 3326 14126 3343 ne
rect 14126 3326 14178 3332
rect 14216 3423 14222 3457
rect 14256 3423 14262 3457
rect 14216 3384 14262 3423
rect 14216 3350 14222 3384
rect 14256 3350 14262 3384
rect 7512 3311 7540 3318
tri 7540 3311 7547 3318 nw
tri 8922 3311 8929 3318 ne
rect 8929 3311 8947 3318
tri 7475 3308 7478 3311 se
rect 7478 3308 7537 3311
tri 7537 3308 7540 3311 nw
tri 8929 3308 8932 3311 ne
rect 8932 3308 8947 3311
tri 7466 3299 7475 3308 se
rect 7475 3299 7528 3308
tri 7528 3299 7537 3308 nw
tri 8932 3299 8941 3308 ne
rect 8941 3299 8947 3308
rect 14216 3311 14262 3350
tri 7461 3294 7466 3299 se
rect 7466 3294 7523 3299
tri 7523 3294 7528 3299 nw
tri 8941 3294 8946 3299 ne
rect 8946 3294 8947 3299
rect 13874 3299 13969 3305
rect 14021 3299 14033 3305
rect 6856 3242 6862 3294
rect 6914 3242 6926 3294
rect 6978 3265 7494 3294
tri 7494 3265 7523 3294 nw
tri 8946 3293 8947 3294 ne
rect 6978 3242 7471 3265
tri 7471 3242 7494 3265 nw
rect 13206 3246 13212 3298
rect 13264 3246 13276 3298
rect 13328 3246 13334 3298
rect 13874 3265 13886 3299
rect 13920 3265 13969 3299
rect 13874 3253 13969 3265
rect 14021 3253 14033 3265
rect 14085 3253 14091 3305
rect 14216 3277 14222 3311
rect 14256 3277 14262 3311
rect 14216 3265 14262 3277
rect 14333 3537 14463 3543
rect 14333 3503 14345 3537
rect 14379 3503 14417 3537
rect 14451 3503 14463 3537
rect 14333 3497 14463 3503
tri 14328 3265 14333 3270 se
rect 14333 3265 14361 3497
tri 14361 3447 14411 3497 nw
tri 14316 3253 14328 3265 se
rect 14328 3253 14361 3265
tri 14309 3246 14316 3253 se
rect 14316 3246 14361 3253
tri 14305 3242 14309 3246 se
rect 14309 3242 14361 3246
rect 151 3048 11231 3214
rect 11862 3190 11868 3242
rect 11920 3190 11932 3242
rect 11984 3218 11990 3242
tri 11990 3218 12014 3242 sw
tri 14285 3222 14305 3242 se
rect 14305 3222 14361 3242
tri 13782 3218 13786 3222 se
rect 13786 3218 14361 3222
rect 11984 3194 14361 3218
rect 14567 3379 14614 3391
rect 14567 3345 14573 3379
rect 14607 3345 14614 3379
rect 14567 3242 14614 3345
rect 14567 3208 14573 3242
rect 14607 3208 14614 3242
rect 11984 3190 13814 3194
tri 13814 3190 13818 3194 nw
rect 12639 3107 12645 3159
rect 12697 3107 12711 3159
rect 12763 3107 12769 3159
rect 13877 3157 14007 3163
rect 13877 3123 13889 3157
rect 13923 3123 13961 3157
rect 13995 3145 14007 3157
tri 14007 3145 14025 3163 sw
rect 13995 3123 14209 3145
rect 13877 3108 14209 3123
tri 14181 3107 14182 3108 ne
rect 14182 3107 14209 3108
tri 14182 3106 14183 3107 ne
rect 14183 3106 14209 3107
tri 11806 3100 11812 3106 ne
tri 11940 3100 11946 3106 nw
tri 14183 3100 14189 3106 ne
rect 14189 3100 14209 3106
tri 14189 3080 14209 3100 ne
tri 14209 3092 14262 3145 sw
rect 14209 3080 14262 3092
tri 14209 3077 14212 3080 ne
rect 14212 3077 14262 3080
rect 151 3031 1021 3048
tri 1021 3031 1038 3048 nw
tri 1152 3031 1169 3048 ne
rect 1169 3031 11231 3048
rect 151 3012 1002 3031
tri 1002 3012 1021 3031 nw
tri 1169 3012 1188 3031 ne
rect 1188 3012 11231 3031
rect 13306 3071 14061 3077
tri 14212 3073 14216 3077 ne
rect 13306 3065 13701 3071
rect 13306 3031 13314 3065
rect 13348 3031 13666 3065
rect 13700 3031 13701 3065
rect 13306 3019 13701 3031
rect 13753 3019 13789 3071
rect 13841 3065 14061 3071
rect 13841 3031 14018 3065
rect 14052 3031 14061 3065
rect 13841 3019 14061 3031
tri 9701 2987 9726 3012 ne
rect 9726 2987 9778 3012
tri 9778 2987 9803 3012 nw
rect 13306 2997 14061 3019
rect 13306 2987 13701 2997
rect 9727 2985 9777 2986
rect 9726 2949 9778 2985
rect 9727 2948 9777 2949
rect 9726 2911 9778 2947
rect 12493 2979 12769 2985
rect 12493 2945 12505 2979
rect 12539 2945 12577 2979
rect 12611 2945 12650 2979
rect 12684 2945 12723 2979
rect 12757 2953 12769 2979
tri 12769 2953 12770 2954 sw
rect 13306 2953 13314 2987
rect 13348 2953 13666 2987
rect 13700 2953 13701 2987
rect 12757 2949 12770 2953
tri 12770 2949 12774 2953 sw
rect 12757 2945 12774 2949
tri 9778 2911 9796 2929 sw
tri 11977 2911 11995 2929 ne
rect 11995 2911 12010 2929
rect 9726 2909 9796 2911
tri 9796 2909 9798 2911 sw
tri 11995 2909 11997 2911 ne
rect 11997 2909 12010 2911
rect 9726 2904 9798 2909
tri 9798 2904 9803 2909 sw
tri 11997 2904 12002 2909 ne
rect 12002 2904 12010 2909
rect 9726 2852 9910 2904
rect 9962 2852 9974 2904
rect 10026 2852 10032 2904
tri 12002 2896 12010 2904 ne
rect 12493 2924 12774 2945
tri 12774 2924 12799 2949 sw
rect 13306 2945 13701 2953
rect 13753 2945 13789 2997
rect 13841 2987 14061 2997
rect 13841 2953 14018 2987
rect 14052 2953 14061 2987
rect 13841 2945 14061 2953
rect 12493 2911 13189 2924
tri 13189 2911 13202 2924 sw
rect 13306 2922 14061 2945
rect 12493 2909 13202 2911
tri 13202 2909 13204 2911 sw
rect 13306 2909 13701 2922
rect 12493 2875 13204 2909
tri 13204 2875 13238 2909 sw
rect 13306 2875 13314 2909
rect 13348 2875 13666 2909
rect 13700 2875 13701 2909
rect 12493 2850 13238 2875
rect 12493 2831 12779 2850
tri 12779 2831 12798 2850 nw
tri 13168 2831 13187 2850 ne
rect 13187 2834 13238 2850
tri 13238 2834 13279 2875 sw
rect 13306 2870 13701 2875
rect 13753 2870 13789 2922
rect 13841 2909 14061 2922
rect 13841 2875 14018 2909
rect 14052 2875 14061 2909
rect 13841 2870 14061 2875
rect 13306 2863 14061 2870
rect 14216 2983 14262 3077
tri 14559 2993 14567 3001 se
rect 14567 2993 14614 3208
rect 14216 2949 14222 2983
rect 14256 2964 14262 2983
tri 14262 2964 14291 2993 sw
tri 14530 2964 14559 2993 se
rect 14559 2964 14614 2993
rect 14256 2949 14614 2964
rect 14216 2911 14614 2949
rect 14216 2877 14222 2911
rect 14256 2904 14614 2911
rect 14256 2877 14263 2904
rect 14216 2865 14263 2877
tri 14263 2865 14302 2904 nw
rect 13187 2831 14087 2834
rect 12493 2826 12774 2831
tri 12774 2826 12779 2831 nw
tri 13187 2829 13189 2831 ne
rect 13189 2829 14087 2831
tri 13189 2826 13192 2829 ne
rect 13192 2826 14087 2829
tri 11809 2800 11812 2803 se
tri 11940 2800 11943 2803 sw
tri 11809 2751 11812 2754 ne
tri 11940 2751 11943 2754 nw
tri 11985 2720 12010 2745 se
tri 11963 2698 11985 2720 se
rect 11985 2698 12010 2720
tri 11953 2688 11963 2698 se
rect 11963 2688 12010 2698
tri 12263 2720 12288 2745 sw
tri 12468 2720 12493 2745 se
rect 12493 2720 12769 2826
tri 12769 2821 12774 2826 nw
tri 13192 2821 13197 2826 ne
rect 13197 2821 14087 2826
tri 13197 2816 13202 2821 ne
rect 13202 2816 14087 2821
rect 12263 2698 12288 2720
tri 12288 2698 12310 2720 sw
tri 12446 2698 12468 2720 se
rect 12468 2698 12769 2720
rect 12263 2688 12310 2698
tri 12310 2688 12320 2698 sw
tri 12436 2688 12446 2698 se
rect 12446 2688 12769 2698
rect 151 2664 9751 2688
tri 9751 2664 9775 2688 sw
tri 9983 2664 10007 2688 se
rect 10007 2664 12769 2688
rect 151 2643 9775 2664
tri 9775 2643 9796 2664 sw
tri 9962 2643 9983 2664 se
rect 9983 2643 12769 2664
rect 151 2633 12769 2643
rect 151 2599 12505 2633
rect 12539 2599 12577 2633
rect 12611 2599 12650 2633
rect 12684 2599 12723 2633
rect 12757 2599 12769 2633
rect 12808 2810 13155 2816
rect 12808 2776 12820 2810
rect 12854 2776 12924 2810
rect 12958 2776 13028 2810
rect 13062 2776 13155 2810
tri 13202 2792 13226 2816 ne
rect 13226 2792 14087 2816
rect 12808 2740 13155 2776
tri 13226 2771 13247 2792 ne
rect 13247 2771 14087 2792
rect 14216 2826 14262 2865
tri 14262 2864 14263 2865 nw
rect 14216 2792 14222 2826
rect 14256 2792 14262 2826
tri 14087 2771 14090 2774 sw
tri 14005 2759 14017 2771 ne
rect 14017 2759 14090 2771
tri 14090 2759 14102 2771 sw
tri 14017 2754 14022 2759 ne
rect 14022 2754 14102 2759
tri 14102 2754 14107 2759 sw
rect 14216 2754 14262 2792
tri 14022 2750 14026 2754 ne
rect 14026 2750 14107 2754
tri 14107 2750 14111 2754 sw
tri 13155 2740 13165 2750 sw
tri 14026 2740 14036 2750 ne
rect 14036 2740 14111 2750
rect 12808 2734 13165 2740
rect 12808 2682 13113 2734
tri 13165 2720 13185 2740 sw
tri 14036 2720 14056 2740 ne
rect 14056 2720 14111 2740
tri 14111 2720 14141 2750 sw
rect 14216 2720 14222 2754
rect 14256 2720 14262 2754
rect 14394 2831 14440 2843
rect 14394 2797 14400 2831
rect 14434 2797 14440 2831
rect 14394 2759 14440 2797
rect 14394 2725 14400 2759
rect 14434 2725 14440 2759
rect 13165 2710 13185 2720
tri 13185 2710 13195 2720 sw
tri 14056 2711 14065 2720 ne
rect 14065 2711 14141 2720
tri 13478 2710 13479 2711 se
rect 13479 2710 13883 2711
rect 13165 2698 13883 2710
rect 13165 2682 13491 2698
rect 12808 2670 13491 2682
rect 12808 2618 13113 2670
rect 13165 2664 13491 2670
rect 13525 2664 13843 2698
rect 13877 2664 13883 2698
tri 14065 2690 14086 2711 ne
rect 14086 2690 14141 2711
tri 14086 2665 14111 2690 ne
rect 14111 2665 14141 2690
tri 14141 2665 14196 2720 sw
rect 14216 2708 14262 2720
tri 14381 2708 14394 2721 se
rect 14394 2708 14440 2725
tri 14338 2665 14381 2708 se
rect 14381 2673 14440 2708
rect 14381 2665 14432 2673
tri 14432 2665 14440 2673 nw
rect 13165 2618 13883 2664
tri 14111 2632 14144 2665 ne
rect 12808 2614 13883 2618
rect 12808 2612 13491 2614
rect 151 2502 12769 2599
tri 13439 2583 13468 2612 ne
rect 13468 2583 13491 2612
rect 13132 2571 13178 2583
tri 13468 2580 13471 2583 ne
rect 13471 2580 13491 2583
rect 13525 2580 13843 2614
rect 13877 2580 13883 2614
tri 13471 2572 13479 2580 ne
rect 13132 2537 13138 2571
rect 13172 2537 13178 2571
rect 151 2486 11407 2502
rect 12105 2499 12118 2502
tri 12118 2499 12121 2502 nw
rect 13132 2499 13178 2537
tri 12105 2486 12118 2499 nw
rect 12798 2477 13074 2483
tri 11809 2448 11812 2451 se
tri 11940 2448 11943 2451 sw
rect 12798 2443 12810 2477
rect 12844 2443 12882 2477
rect 12916 2443 12955 2477
rect 12989 2443 13028 2477
rect 13062 2443 13074 2477
tri 11809 2399 11812 2402 ne
tri 11940 2399 11943 2402 nw
rect 12798 2392 13074 2443
rect 13132 2465 13138 2499
rect 13172 2465 13178 2499
rect 13479 2529 13883 2580
rect 14144 2582 14305 2665
rect 13479 2495 13491 2529
rect 13525 2495 13843 2529
rect 13877 2495 13883 2529
rect 13132 2462 13178 2465
tri 13178 2462 13205 2489 sw
rect 13479 2483 13883 2495
rect 14039 2547 14091 2553
rect 14144 2548 14158 2582
rect 14192 2548 14230 2582
rect 14264 2548 14305 2582
rect 14144 2538 14305 2548
tri 14305 2538 14432 2665 nw
tri 14037 2483 14039 2485 se
rect 14039 2483 14091 2495
tri 14667 2485 14689 2507 se
rect 14689 2485 14735 3590
tri 14016 2462 14037 2483 se
rect 14037 2462 14039 2483
rect 13132 2455 13205 2462
tri 13205 2455 13212 2462 sw
tri 14009 2455 14016 2462 se
rect 14016 2455 14039 2462
rect 13132 2431 14039 2455
tri 14091 2462 14114 2485 sw
tri 14659 2477 14667 2485 se
rect 14667 2477 14735 2485
tri 14449 2474 14452 2477 se
rect 14452 2474 14735 2477
tri 14434 2462 14446 2474 se
rect 14446 2462 14735 2474
rect 14091 2455 14114 2462
tri 14114 2455 14121 2462 sw
tri 14427 2455 14434 2462 se
rect 14434 2455 14452 2462
rect 14091 2431 14452 2455
rect 13132 2428 14452 2431
rect 14486 2431 14735 2462
rect 14486 2428 14492 2431
rect 13132 2423 14492 2428
tri 14413 2422 14414 2423 ne
rect 14414 2422 14492 2423
tri 13074 2392 13104 2422 sw
tri 14414 2392 14444 2422 ne
rect 14444 2392 14492 2422
tri 14492 2401 14522 2431 nw
rect 12798 2340 13168 2392
rect 13220 2340 13232 2392
rect 13284 2340 14040 2392
rect 14092 2340 14104 2392
rect 14156 2340 14162 2392
tri 14444 2390 14446 2392 ne
rect 14446 2390 14492 2392
rect 14446 2356 14452 2390
rect 14486 2356 14492 2390
rect 14446 2344 14492 2356
rect 14659 2353 14711 2365
rect 14659 2319 14669 2353
rect 14703 2319 14711 2353
rect 14659 2281 14711 2319
rect 14659 2247 14669 2281
rect 14703 2247 14711 2281
rect 151 2192 11407 2204
rect 151 2158 10133 2192
rect 10167 2158 11069 2192
rect 11103 2158 11407 2192
rect 151 2120 11407 2158
rect 151 2086 10133 2120
rect 10167 2086 11069 2120
rect 11103 2086 11407 2120
rect 151 2074 11407 2086
tri 8928 2062 8940 2074 ne
rect 8940 2062 9379 2074
tri 8940 2049 8953 2062 ne
rect 8953 2028 8959 2062
rect 8993 2028 9339 2062
rect 9373 2028 9379 2062
tri 9379 2049 9404 2074 nw
rect 8953 1990 9379 2028
rect 8953 1956 8959 1990
rect 8993 1956 9339 1990
rect 9373 1956 9379 1990
rect 8953 1944 9379 1956
rect 9436 1994 9577 2046
rect 9579 2045 9615 2046
rect 9578 1995 9616 2045
rect 9579 1994 9615 1995
rect 9617 1994 9665 2046
rect 9717 1994 9729 2046
rect 9781 1994 9787 2046
tri 9787 1994 9797 2004 sw
rect 9904 1994 9910 2046
rect 9962 1994 9974 2046
rect 10026 1994 10032 2046
rect 6711 1871 6862 1923
rect 6914 1871 6926 1923
rect 6978 1871 7443 1923
tri 9411 1890 9436 1915 se
rect 9436 1890 9488 1994
tri 9488 1969 9513 1994 nw
tri 9723 1969 9748 1994 ne
rect 9748 1969 9797 1994
tri 9748 1920 9797 1969 ne
tri 9797 1926 9865 1994 sw
tri 9955 1969 9980 1994 ne
rect 9980 1969 10032 1994
rect 9981 1967 10031 1968
tri 14643 1931 14659 1947 se
rect 14659 1931 14711 2247
rect 9981 1930 10031 1931
tri 14642 1930 14643 1931 se
rect 14643 1930 14711 1931
tri 14641 1929 14642 1930 se
rect 14642 1929 14711 1930
tri 9977 1926 9980 1929 se
rect 9980 1926 10032 1929
rect 9797 1920 9865 1926
tri 9797 1915 9802 1920 ne
rect 9802 1915 9865 1920
tri 9488 1890 9513 1915 sw
tri 9802 1890 9827 1915 ne
rect 9827 1904 9865 1915
tri 9865 1904 9887 1926 sw
tri 9955 1904 9977 1926 se
rect 9977 1904 10032 1926
rect 9827 1890 10032 1904
rect 7058 1822 7161 1843
tri 7161 1822 7182 1843 sw
rect 8779 1838 8785 1890
rect 8837 1838 8849 1890
rect 8901 1838 9514 1890
rect 9516 1889 9552 1890
rect 9515 1839 9553 1889
rect 9516 1838 9552 1839
rect 9554 1838 9665 1890
rect 9717 1838 9729 1890
rect 9781 1838 9787 1890
tri 9827 1852 9865 1890 ne
rect 9865 1852 10032 1890
tri 14594 1882 14641 1929 se
rect 14641 1925 14711 1929
rect 14641 1882 14668 1925
tri 14668 1882 14711 1925 nw
tri 14572 1860 14594 1882 se
tri 9955 1838 9969 1852 ne
rect 9969 1838 10032 1852
tri 9555 1822 9571 1838 ne
rect 9571 1822 9632 1838
rect 7058 1791 7182 1822
tri 7139 1748 7182 1791 ne
tri 7182 1748 7256 1822 sw
tri 9571 1813 9580 1822 ne
rect 9580 1813 9632 1822
tri 9632 1813 9657 1838 nw
tri 9969 1827 9980 1838 ne
rect 9581 1811 9631 1812
rect 9581 1774 9631 1775
tri 9555 1748 9580 1773 se
rect 9580 1748 9632 1773
tri 9632 1748 9657 1773 sw
tri 9955 1748 9980 1773 se
rect 9980 1748 10032 1838
rect 11586 1808 11592 1860
rect 11644 1808 11656 1860
rect 11708 1808 14594 1860
tri 14594 1808 14668 1882 nw
tri 7182 1738 7192 1748 ne
rect 7192 1738 9712 1748
tri 7192 1704 7226 1738 ne
rect 7226 1704 9514 1738
rect 9548 1704 9586 1738
rect 9620 1704 9712 1738
tri 7226 1696 7234 1704 ne
rect 7234 1696 9712 1704
rect 9713 1697 9714 1747
rect 9750 1697 9751 1747
rect 9752 1696 10032 1748
rect 8871 1616 8877 1668
rect 8929 1616 8941 1668
rect 8993 1656 9145 1668
rect 8993 1622 9027 1656
rect 9061 1622 9099 1656
rect 9133 1622 9145 1656
rect 8993 1616 9145 1622
rect 9188 1656 9318 1662
rect 9188 1622 9200 1656
rect 9234 1622 9272 1656
rect 9306 1622 9318 1656
rect 9188 1616 9318 1622
rect 151 1458 11407 1588
tri 8710 1424 8716 1430 se
rect 8716 1424 9077 1430
tri 8676 1390 8710 1424 se
rect 8710 1390 8959 1424
rect 8993 1390 9031 1424
rect 9065 1390 9077 1424
tri 8653 1367 8676 1390 se
rect 8676 1384 9077 1390
rect 8676 1367 8716 1384
tri 8716 1367 8733 1384 nw
tri 8642 1356 8653 1367 se
tri 7786 1340 7802 1356 se
rect 7802 1340 8653 1356
rect 6407 1288 6413 1340
rect 6465 1288 6477 1340
rect 6529 1311 7406 1340
tri 7406 1311 7435 1340 sw
tri 7757 1311 7786 1340 se
rect 7786 1311 8653 1340
rect 6529 1288 7435 1311
tri 7384 1237 7435 1288 ne
tri 7435 1237 7509 1311 sw
tri 7740 1294 7757 1311 se
rect 7757 1304 8653 1311
tri 8653 1304 8716 1367 nw
rect 7757 1294 7802 1304
tri 7802 1294 7812 1304 nw
tri 8713 1294 8720 1301 se
rect 8720 1294 9346 1301
tri 7683 1237 7740 1294 se
rect 7740 1237 7745 1294
tri 7745 1237 7802 1294 nw
tri 8661 1242 8713 1294 se
rect 8713 1249 9346 1294
rect 8713 1242 8735 1249
tri 8735 1242 8742 1249 nw
tri 7435 1185 7487 1237 ne
rect 7487 1185 7693 1237
tri 7693 1185 7745 1237 nw
rect 7805 1190 7811 1242
rect 7863 1190 7875 1242
rect 7927 1190 8683 1242
tri 8683 1190 8735 1242 nw
rect 8779 1091 8785 1143
rect 8837 1091 8849 1143
rect 8901 1091 8907 1143
rect 151 1051 11407 1063
rect 151 1017 8843 1051
rect 8877 1017 9339 1051
rect 9373 1017 11407 1051
rect 151 979 11407 1017
rect 151 945 8843 979
rect 8877 945 9339 979
rect 9373 945 11407 979
rect 151 861 11407 945
rect 8947 787 8999 833
rect 8960 728 8971 739
rect 9659 719 9665 771
rect 9717 759 9729 771
rect 9781 759 9842 771
rect 9717 725 9724 759
rect 9781 725 9796 759
rect 9830 725 9842 759
rect 9717 719 9729 725
rect 9781 719 9842 725
rect 7805 621 7811 673
rect 7863 621 7875 673
rect 7927 621 7933 673
rect 56 409 11312 537
rect 11367 409 11407 537
rect 56 335 9588 409
tri 9588 375 9622 409 nw
rect 11186 375 11204 409
tri 11204 375 11238 409 nw
tri 11186 357 11204 375 nw
rect 6364 301 6413 307
rect 6465 301 6477 307
rect 6364 267 6376 301
rect 6410 267 6413 301
rect 6364 255 6413 267
rect 6465 255 6477 267
rect 6529 255 6535 307
rect 6756 276 6771 290
rect 7012 255 8710 307
rect 6875 38 6881 90
rect 6933 38 6945 90
rect 6997 38 7003 90
<< rmetal1 >>
rect 11490 4412 11492 4413
rect 11490 4362 11491 4412
rect 11490 4361 11492 4362
rect 11528 4412 11530 4413
rect 11529 4362 11530 4412
rect 11528 4361 11530 4362
rect 11490 4332 11492 4333
rect 11528 4332 11530 4333
rect 11490 4282 11491 4332
rect 11529 4282 11530 4332
rect 11490 4281 11492 4282
rect 11528 4281 11530 4282
rect 11791 4332 11793 4333
rect 11791 4282 11792 4332
rect 11791 4281 11793 4282
rect 11829 4332 11831 4333
rect 11830 4282 11831 4332
rect 11829 4281 11831 4282
rect 9726 2986 9778 2987
rect 9726 2985 9727 2986
rect 9777 2985 9778 2986
rect 9726 2948 9727 2949
rect 9777 2948 9778 2949
rect 9726 2947 9778 2948
rect 9577 2045 9579 2046
rect 9615 2045 9617 2046
rect 9577 1995 9578 2045
rect 9616 1995 9617 2045
rect 9577 1994 9579 1995
rect 9615 1994 9617 1995
rect 9980 1968 10032 1969
rect 9980 1967 9981 1968
rect 10031 1967 10032 1968
rect 9980 1930 9981 1931
rect 10031 1930 10032 1931
rect 9980 1929 10032 1930
rect 9514 1889 9516 1890
rect 9552 1889 9554 1890
rect 9514 1839 9515 1889
rect 9553 1839 9554 1889
rect 9514 1838 9516 1839
rect 9552 1838 9554 1839
rect 9580 1812 9632 1813
rect 9580 1811 9581 1812
rect 9631 1811 9632 1812
rect 9580 1774 9581 1775
rect 9631 1774 9632 1775
rect 9580 1773 9632 1774
rect 9712 1747 9714 1748
rect 9712 1697 9713 1747
rect 9712 1696 9714 1697
rect 9750 1747 9752 1748
rect 9751 1697 9752 1747
rect 9750 1696 9752 1697
<< via1 >>
rect 8877 4441 8929 4493
rect 8941 4441 8993 4493
rect 6994 4355 7046 4407
rect 11618 4361 11670 4413
rect 11682 4361 11734 4413
rect 13607 4361 13659 4413
rect 13671 4361 13723 4413
rect 6994 4290 7046 4342
rect 8676 4275 8728 4327
rect 11618 4281 11670 4333
rect 11682 4281 11734 4333
rect 11850 4281 11902 4333
rect 11914 4281 11966 4333
rect 8676 4211 8728 4263
rect 13607 4041 13659 4093
rect 13671 4041 13723 4093
rect 11699 3814 11751 3866
rect 12671 3814 12723 3866
rect 13701 3814 13753 3866
rect 13789 3860 13841 3866
rect 13789 3826 13798 3860
rect 13798 3826 13841 3860
rect 13789 3814 13841 3826
rect 11699 3732 11751 3784
rect 12671 3732 12723 3784
rect 13701 3732 13753 3784
rect 13789 3765 13841 3784
rect 13789 3732 13798 3765
rect 13798 3732 13841 3765
rect 9735 3640 9787 3692
rect 9735 3576 9787 3628
rect 9986 3498 10038 3550
rect 10050 3498 10102 3550
rect 13119 3346 13171 3398
rect 13183 3346 13235 3398
rect 14126 3396 14178 3448
rect 14126 3332 14178 3384
rect 13969 3299 14021 3305
rect 14033 3299 14085 3305
rect 6862 3242 6914 3294
rect 6926 3242 6978 3294
rect 13212 3246 13264 3298
rect 13276 3246 13328 3298
rect 13969 3265 14019 3299
rect 14019 3265 14021 3299
rect 14033 3265 14053 3299
rect 14053 3265 14085 3299
rect 13969 3253 14021 3265
rect 14033 3253 14085 3265
rect 11868 3190 11920 3242
rect 11932 3190 11984 3242
rect 12645 3149 12697 3159
rect 12645 3115 12651 3149
rect 12651 3115 12685 3149
rect 12685 3115 12697 3149
rect 12645 3107 12697 3115
rect 12711 3149 12763 3159
rect 12711 3115 12723 3149
rect 12723 3115 12757 3149
rect 12757 3115 12763 3149
rect 12711 3107 12763 3115
rect 13701 3019 13753 3071
rect 13789 3019 13841 3071
rect 9910 2852 9962 2904
rect 9974 2852 10026 2904
rect 13701 2945 13753 2997
rect 13789 2945 13841 2997
rect 13701 2870 13753 2922
rect 13789 2870 13841 2922
rect 13113 2682 13165 2734
rect 13113 2618 13165 2670
rect 14039 2495 14091 2547
rect 14039 2431 14091 2483
rect 13168 2340 13220 2392
rect 13232 2340 13284 2392
rect 14040 2340 14092 2392
rect 14104 2340 14156 2392
rect 9665 1994 9717 2046
rect 9729 1994 9781 2046
rect 9910 1994 9962 2046
rect 9974 1994 10026 2046
rect 6862 1871 6914 1923
rect 6926 1871 6978 1923
rect 8785 1838 8837 1890
rect 8849 1838 8901 1890
rect 9665 1838 9717 1890
rect 9729 1838 9781 1890
rect 11592 1808 11644 1860
rect 11656 1808 11708 1860
rect 8877 1616 8929 1668
rect 8941 1616 8993 1668
rect 6413 1288 6465 1340
rect 6477 1288 6529 1340
rect 7811 1190 7863 1242
rect 7875 1190 7927 1242
rect 8785 1091 8837 1143
rect 8849 1091 8901 1143
rect 9665 719 9717 771
rect 9729 759 9781 771
rect 9729 725 9758 759
rect 9758 725 9781 759
rect 9729 719 9781 725
rect 7811 621 7863 673
rect 7875 621 7927 673
rect 6413 301 6465 307
rect 6477 301 6529 307
rect 6413 267 6448 301
rect 6448 267 6465 301
rect 6477 267 6482 301
rect 6482 267 6529 301
rect 6413 255 6465 267
rect 6477 255 6529 267
rect 6881 38 6933 90
rect 6945 38 6997 90
<< metal2 >>
rect 8871 4441 8877 4493
rect 8929 4441 8941 4493
rect 8993 4441 8999 4493
tri 8915 4413 8943 4441 ne
rect 8943 4413 8999 4441
rect 6994 4407 7046 4413
tri 8943 4409 8947 4413 ne
rect 6994 4342 7046 4355
tri 6977 3550 6994 3567 se
rect 6994 3550 7046 4290
tri 6925 3498 6977 3550 se
rect 6977 3545 7046 3550
rect 6977 3498 6999 3545
tri 6999 3498 7046 3545 nw
rect 8676 4327 8728 4333
rect 8676 4263 8728 4275
tri 6920 3493 6925 3498 se
rect 6925 3493 6994 3498
tri 6994 3493 6999 3498 nw
tri 6875 3448 6920 3493 se
rect 6920 3448 6949 3493
tri 6949 3448 6994 3493 nw
tri 6846 3419 6875 3448 se
rect 6875 3419 6920 3448
tri 6920 3419 6949 3448 nw
rect 8676 3419 8728 4211
tri 8914 4041 8947 4074 se
rect 8947 4041 8999 4413
rect 11612 4361 11618 4413
rect 11670 4361 11682 4413
rect 11734 4361 11740 4413
rect 11612 4333 11740 4361
rect 13601 4361 13607 4413
rect 13659 4361 13671 4413
rect 13723 4361 13729 4413
rect 11612 4281 11618 4333
rect 11670 4281 11682 4333
rect 11734 4281 11740 4333
tri 11812 4281 11844 4313 se
rect 11844 4281 11850 4333
rect 11902 4281 11914 4333
rect 11966 4281 11972 4333
tri 11784 4253 11812 4281 se
rect 11812 4253 11972 4281
tri 8910 4037 8914 4041 se
rect 8914 4037 8999 4041
rect 11675 4198 11972 4253
rect 11675 4093 11727 4198
tri 11727 4162 11763 4198 nw
rect 11676 4091 11726 4092
rect 11675 4055 11727 4091
rect 11676 4054 11726 4055
rect 11675 3872 11727 4053
rect 13601 4093 13729 4361
rect 13601 4041 13607 4093
rect 13659 4041 13671 4093
rect 13723 4041 13729 4093
tri 11817 4017 11840 4040 ne
rect 11907 4017 11924 4040
tri 11924 4017 11947 4040 nw
tri 11907 4000 11924 4017 nw
tri 11727 3872 11775 3920 sw
rect 11675 3866 11775 3872
rect 11675 3814 11699 3866
rect 11751 3814 11775 3866
rect 11675 3784 11775 3814
rect 11675 3732 11699 3784
rect 11751 3732 11775 3784
rect 11675 3726 11775 3732
rect 12639 3866 12747 3872
rect 12639 3814 12671 3866
rect 12723 3814 12747 3866
rect 12639 3784 12747 3814
rect 12639 3732 12671 3784
rect 12723 3732 12747 3784
rect 9735 3692 9787 3698
rect 9735 3628 9787 3640
tri 6825 3398 6846 3419 se
rect 6846 3398 6899 3419
tri 6899 3398 6920 3419 nw
tri 8676 3398 8697 3419 ne
rect 8697 3412 8728 3419
tri 8728 3412 8757 3441 sw
rect 8697 3398 8757 3412
tri 8757 3398 8771 3412 sw
tri 6773 3346 6825 3398 se
rect 6825 3346 6847 3398
tri 6847 3346 6899 3398 nw
tri 8697 3367 8728 3398 ne
rect 8728 3367 8771 3398
tri 8728 3346 8749 3367 ne
rect 8749 3346 8771 3367
tri 8771 3346 8823 3398 sw
tri 6772 3345 6773 3346 se
rect 6773 3345 6846 3346
tri 6846 3345 6847 3346 nw
tri 8749 3345 8750 3346 ne
rect 8750 3345 8823 3346
tri 6766 3339 6772 3345 se
rect 6772 3339 6833 3345
rect 6766 3332 6833 3339
tri 6833 3332 6846 3345 nw
tri 8750 3338 8757 3345 ne
rect 8757 3338 8823 3345
tri 8823 3338 8831 3346 sw
tri 8757 3332 8763 3338 ne
rect 8763 3332 8831 3338
rect 6766 1843 6818 3332
tri 6818 3317 6833 3332 nw
tri 8763 3317 8778 3332 ne
rect 8778 3317 8831 3332
tri 8778 3316 8779 3317 ne
rect 6856 3242 6862 3294
rect 6914 3242 6926 3294
rect 6978 3242 6984 3294
rect 6856 1923 6908 3242
tri 6908 3217 6933 3242 nw
tri 6908 1923 6933 1948 sw
rect 6856 1871 6862 1923
rect 6914 1871 6926 1923
rect 6978 1871 6984 1923
rect 8779 1890 8831 3317
rect 6766 1791 6875 1843
rect 8779 1838 8785 1890
rect 8837 1838 8849 1890
rect 8901 1838 8907 1890
rect 6407 1288 6413 1340
rect 6465 1288 6477 1340
rect 6529 1288 6535 1340
rect 6407 307 6478 1288
tri 6478 1263 6503 1288 nw
rect 7805 1190 7811 1242
rect 7863 1190 7875 1242
rect 7927 1190 7933 1242
rect 7805 673 7872 1190
tri 7872 1165 7897 1190 nw
rect 8779 1143 8843 1838
tri 8843 1813 8868 1838 nw
tri 8922 1668 8947 1693 se
rect 8947 1668 8999 3242
tri 9710 2046 9735 2071 se
rect 9735 2046 9787 3576
rect 9980 3498 9986 3550
rect 10038 3498 10050 3550
rect 10102 3498 10108 3550
rect 9815 2932 9873 2984
tri 9973 2922 9980 2929 se
rect 9980 2922 10032 3498
tri 10032 3473 10057 3498 nw
tri 11714 3246 11737 3269 sw
rect 11714 3242 11737 3246
tri 11737 3242 11741 3246 sw
tri 9955 2904 9973 2922 se
rect 9973 2904 10032 2922
rect 9904 2852 9910 2904
rect 9962 2852 9974 2904
rect 10026 2852 10032 2904
tri 9955 2827 9980 2852 ne
tri 9955 2046 9980 2071 se
rect 9980 2046 10032 2852
rect 9659 1994 9665 2046
rect 9717 1994 9729 2046
rect 9781 1994 9787 2046
rect 9904 1994 9910 2046
rect 9962 1994 9974 2046
rect 10026 1994 10032 2046
rect 11586 3190 11868 3242
rect 11920 3190 11932 3242
rect 11984 3190 11990 3242
rect 8871 1616 8877 1668
rect 8929 1616 8941 1668
rect 8993 1616 8999 1668
tri 8922 1591 8947 1616 ne
rect 8947 1221 8999 1616
rect 9659 1838 9665 1890
rect 9717 1838 9729 1890
rect 9781 1838 9787 1890
rect 9346 1249 9393 1301
tri 8843 1143 8868 1168 sw
rect 8779 1091 8785 1143
rect 8837 1091 8849 1143
rect 8901 1091 8907 1143
rect 9659 771 9787 1838
rect 9659 719 9665 771
rect 9717 719 9729 771
rect 9781 719 9787 771
rect 11586 1860 11714 3190
tri 11714 3162 11742 3190 nw
rect 12639 3159 12747 3732
rect 13700 3866 13841 3872
rect 13700 3814 13701 3866
rect 13753 3814 13789 3866
rect 13700 3784 13841 3814
rect 13700 3732 13701 3784
rect 13753 3732 13789 3784
rect 13113 3346 13119 3398
rect 13171 3346 13183 3398
rect 13235 3346 13241 3398
rect 13113 3332 13186 3346
tri 13186 3332 13200 3346 nw
rect 12639 3107 12645 3159
rect 12697 3107 12711 3159
rect 12763 3107 12769 3159
rect 13113 2734 13165 3332
tri 13165 3311 13186 3332 nw
rect 13113 2670 13165 2682
rect 13113 2612 13165 2618
rect 13206 3246 13212 3298
rect 13264 3246 13276 3298
rect 13328 3246 13334 3298
tri 13174 2392 13206 2424 se
rect 13206 2392 13258 3246
tri 13258 3210 13294 3246 nw
rect 13700 3071 13841 3732
rect 14126 3448 14178 3454
rect 14126 3384 14178 3396
rect 14126 3326 14178 3332
rect 13963 3253 13969 3305
rect 14021 3253 14033 3305
rect 14085 3253 14091 3305
tri 14004 3218 14039 3253 ne
rect 13700 3019 13701 3071
rect 13753 3019 13789 3071
rect 13700 2997 13841 3019
rect 13700 2945 13701 2997
rect 13753 2945 13789 2997
rect 13700 2922 13841 2945
rect 13700 2870 13701 2922
rect 13753 2870 13789 2922
rect 13700 2864 13841 2870
rect 14039 2547 14091 3253
rect 14039 2483 14091 2495
rect 14039 2425 14091 2431
tri 13258 2392 13290 2424 sw
rect 14126 2392 14162 3326
rect 13162 2340 13168 2392
rect 13220 2340 13232 2392
rect 13284 2340 13290 2392
rect 14034 2340 14040 2392
rect 14092 2340 14104 2392
rect 14156 2340 14162 2392
rect 11586 1808 11592 1860
rect 11644 1808 11656 1860
rect 11708 1808 11714 1860
tri 7872 673 7897 698 sw
rect 7805 621 7811 673
rect 7863 621 7875 673
rect 7927 621 7933 673
tri 6478 307 6503 332 sw
rect 6407 255 6413 307
rect 6465 255 6477 307
rect 6529 255 6535 307
tri 6841 221 6875 255 ne
rect 6875 90 6927 275
rect 11586 255 11714 1808
tri 6927 90 6961 124 sw
rect 6875 38 6881 90
rect 6933 38 6945 90
rect 6997 38 7003 90
<< rmetal2 >>
rect 11675 4092 11727 4093
rect 11675 4091 11676 4092
rect 11726 4091 11727 4092
rect 11675 4054 11676 4055
rect 11726 4054 11727 4055
rect 11675 4053 11727 4054
use hvnTran_CDNS_52468879185363  hvnTran_CDNS_52468879185363_0
timestamp 1704896540
transform 1 0 9398 0 1 1838
box -93 -26 199 226
use hvnTran_CDNS_52468879185364  hvnTran_CDNS_52468879185364_0
timestamp 1704896540
transform 1 0 9018 0 1 1838
box -93 -26 389 226
use hvpTran_CDNS_52468879185361  hvpTran_CDNS_52468879185361_0
timestamp 1704896540
transform -1 0 9314 0 -1 1578
box -133 -66 236 666
use hvpTran_CDNS_52468879185361  hvpTran_CDNS_52468879185361_1
timestamp 1704896540
transform 1 0 9018 0 -1 1578
box -133 -66 236 666
use hvpTran_CDNS_52468879185362  hvpTran_CDNS_52468879185362_0
timestamp 1704896540
transform 1 0 9398 0 -1 1578
box -133 -66 239 666
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1704896540
transform 0 -1 9373 -1 0 1051
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1704896540
transform 0 -1 8877 -1 0 1051
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1704896540
transform -1 0 9830 0 1 725
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1704896540
transform 0 1 9339 1 0 1956
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_4
timestamp 1704896540
transform 0 1 8959 1 0 1956
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_5
timestamp 1704896540
transform 0 -1 10167 1 0 2086
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_6
timestamp 1704896540
transform 0 -1 11103 1 0 2086
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_7
timestamp 1704896540
transform 1 0 9200 0 -1 1656
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_8
timestamp 1704896540
transform 1 0 9027 0 -1 1656
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_9
timestamp 1704896540
transform 1 0 8959 0 -1 1424
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_10
timestamp 1704896540
transform 1 0 9514 0 -1 1738
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_11
timestamp 1704896540
transform 1 0 10055 0 1 3658
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_12
timestamp 1704896540
transform 1 0 10300 0 1 3504
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_13
timestamp 1704896540
transform 1 0 6376 0 1 267
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1704896540
transform 0 -1 9787 -1 0 3698
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_1
timestamp 1704896540
transform -1 0 7933 0 1 621
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_2
timestamp 1704896540
transform -1 0 7933 0 1 1190
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_3
timestamp 1704896540
transform -1 0 8999 0 1 1616
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_4
timestamp 1704896540
transform -1 0 10032 0 1 1994
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_5
timestamp 1704896540
transform -1 0 10032 0 1 2852
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_6
timestamp 1704896540
transform 1 0 9659 0 1 1838
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_7
timestamp 1704896540
transform 1 0 6856 0 1 3242
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_8
timestamp 1704896540
transform 1 0 6856 0 1 1871
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_9
timestamp 1704896540
transform 1 0 9659 0 1 719
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_10
timestamp 1704896540
transform 1 0 8779 0 1 1838
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_11
timestamp 1704896540
transform 1 0 8779 0 1 1091
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_12
timestamp 1704896540
transform 1 0 6407 0 1 1288
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_13
timestamp 1704896540
transform 1 0 6407 0 1 255
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_14
timestamp 1704896540
transform 1 0 9980 0 1 3498
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_15
timestamp 1704896540
transform 1 0 9659 0 1 1994
box 0 0 1 1
use nfet_CDNS_524688791851409  nfet_CDNS_524688791851409_0
timestamp 1704896540
transform 1 0 14267 0 1 2713
box -79 -26 199 110
use nfet_CDNS_524688791851409  nfet_CDNS_524688791851409_1
timestamp 1704896540
transform 1 0 14267 0 1 2891
box -79 -26 199 110
use nfet_CDNS_524688791851410  nfet_CDNS_524688791851410_0
timestamp 1704896540
transform -1 0 14441 0 -1 2470
box -79 -26 179 110
use nfet_CDNS_524688791851411  nfet_CDNS_524688791851411_0
timestamp 1704896540
transform 0 1 12486 -1 0 2588
box -79 -26 179 626
use nfet_CDNS_524688791851412  nfet_CDNS_524688791851412_0
timestamp 1704896540
transform 0 1 12486 -1 0 2940
box -79 -26 375 626
use pfet_CDNS_52468879185663  pfet_CDNS_52468879185663_0
timestamp 1704896540
transform 1 0 14267 0 1 3194
box -119 -66 415 266
use pfet_CDNS_524688791851413  pfet_CDNS_524688791851413_0
timestamp 1704896540
transform -1 0 14007 0 -1 3079
box -119 -66 767 666
use pfet_CDNS_524688791851414  pfet_CDNS_524688791851414_0
timestamp 1704896540
transform 1 0 14360 0 1 3579
box -119 -66 219 266
use pfet_CDNS_524688791851415  pfet_CDNS_524688791851415_0
timestamp 1704896540
transform 1 0 13809 0 1 3347
box -119 -66 375 666
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_0
timestamp 1704896540
transform 0 1 9398 1 0 1610
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_1
timestamp 1704896540
transform 0 1 9221 1 0 1610
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_2
timestamp 1704896540
transform 0 1 9045 1 0 1610
box 0 0 1 1
use sky130_fd_io__sio_com_pdpredrvr_pbias  sky130_fd_io__sio_com_pdpredrvr_pbias_0
timestamp 1704896540
transform -1 0 20219 0 1 -2765
box 11364 2974 20068 5671
use sky130_fd_io__sio_com_pdpredrvr_strong_nr2  sky130_fd_io__sio_com_pdpredrvr_strong_nr2_0
timestamp 1704896540
transform -1 0 11407 0 1 2124
box -307 10 3426 1950
use sky130_fd_io__sio_com_pdpredrvr_strong_nr2_a  sky130_fd_io__sio_com_pdpredrvr_strong_nr2_a_0
timestamp 1704896540
transform -1 0 11186 0 -1 2126
box -528 0 2606 1910
use sky130_fd_io__sio_com_pdpredrvr_strong_nr2_i2c  sky130_fd_io__sio_com_pdpredrvr_strong_nr2_i2c_0
timestamp 1704896540
transform 1 0 11139 0 1 2297
box 112 77 2613 1798
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851254  sky130_fd_io__sio_tk_em1o_CDNS_524688791851254_0
timestamp 1704896540
transform 0 -1 10032 -1 0 2021
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851254  sky130_fd_io__sio_tk_em1o_CDNS_524688791851254_1
timestamp 1704896540
transform 0 1 9580 1 0 1721
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851254  sky130_fd_io__sio_tk_em1o_CDNS_524688791851254_2
timestamp 1704896540
transform 1 0 11438 0 -1 4413
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851254  sky130_fd_io__sio_tk_em1o_CDNS_524688791851254_3
timestamp 1704896540
transform 1 0 9660 0 1 1696
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851254  sky130_fd_io__sio_tk_em1o_CDNS_524688791851254_4
timestamp 1704896540
transform 1 0 11739 0 1 4281
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851255  sky130_fd_io__sio_tk_em1s_CDNS_524688791851255_0
timestamp 1704896540
transform 0 -1 9778 -1 0 3039
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851255  sky130_fd_io__sio_tk_em1s_CDNS_524688791851255_1
timestamp 1704896540
transform -1 0 9669 0 1 1994
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851255  sky130_fd_io__sio_tk_em1s_CDNS_524688791851255_2
timestamp 1704896540
transform -1 0 11582 0 1 4281
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851255  sky130_fd_io__sio_tk_em1s_CDNS_524688791851255_3
timestamp 1704896540
transform -1 0 9606 0 -1 1890
box 0 0 1 1
use sky130_fd_io__sio_tk_em2s_CDNS_524688791851404  sky130_fd_io__sio_tk_em2s_CDNS_524688791851404_0
timestamp 1704896540
transform 0 1 11675 -1 0 4145
box 0 0 1 1
<< labels >>
flabel comment s 13246 2670 13246 2670 0 FreeSans 200 0 0 0 i2c_mode_enable_h_n
flabel comment s 14324 3086 14324 3086 0 FreeSans 200 0 0 0 i2c_mode_h_n
flabel comment s 6484 1312 6484 1312 0 FreeSans 300 0 0 0 en_fast_h
flabel comment s 8461 1341 8461 1341 0 FreeSans 300 0 0 0 en_fast_h
flabel comment s 9614 1726 9614 1726 0 FreeSans 300 0 0 0 en_fast_h_n
flabel comment s 7048 1826 7048 1826 0 FreeSans 300 0 0 0 en_fast_h_n
flabel comment s 8849 1882 8849 1882 0 FreeSans 300 0 0 0 pbias
flabel comment s 10358 3923 10358 3923 0 FreeSans 100 0 0 0 li_jumper_ok
flabel comment s 10107 1682 10107 1682 0 FreeSans 300 0 0 0 pbias
flabel comment s 9992 2350 9992 2350 0 FreeSans 300 90 0 0 en_fast2_n0
flabel comment s 9716 1877 9716 1877 0 FreeSans 300 0 0 0 en_fast_n1
flabel comment s 9697 2345 9697 2345 0 FreeSans 300 90 0 0 en_fast2_n1
flabel comment s 8428 957 8428 957 0 FreeSans 300 0 0 0 vcc_io
flabel comment s 8404 425 8404 425 0 FreeSans 300 0 0 0 vgnd_io
flabel comment s 7856 3276 7856 3276 0 FreeSans 300 0 0 0 pden_h_n
flabel comment s 8964 3921 8964 3921 0 FreeSans 300 90 0 0 pden_h_n
flabel comment s 8963 2297 8963 2297 0 FreeSans 300 90 0 0 pden_h_n
flabel metal1 s 151 861 191 1063 3 FreeSans 300 180 0 0 vcc_io
port 4 nsew
flabel metal1 s 151 2074 191 2204 3 FreeSans 300 180 0 0 vgnd_io
port 3 nsew
flabel metal1 s 11191 3012 11231 3214 7 FreeSans 300 180 0 0 vcc_io
port 4 nsew
flabel metal1 s 11367 2486 11407 2688 7 FreeSans 300 180 0 0 vgnd_io
port 3 nsew
flabel metal1 s 8617 1337 8617 1337 3 FreeSans 400 0 0 0 en_fast_h
flabel metal1 s 151 335 191 537 3 FreeSans 300 180 0 0 vgnd_io
port 3 nsew
flabel metal1 s 11367 3726 11407 3872 7 FreeSans 300 180 0 0 vcc_io
port 4 nsew
flabel metal1 s 11386 2587 11386 2587 7 FreeSans 300 180 0 0 vgnd_io
flabel metal1 s 11367 952 11407 1063 7 FreeSans 300 180 0 0 vcc_io
port 4 nsew
flabel metal1 s 11367 409 11407 537 7 FreeSans 300 180 0 0 vgnd_io
port 3 nsew
flabel metal1 s 11367 1458 11407 1588 7 FreeSans 300 180 0 0 vgnd_io
port 3 nsew
flabel metal1 s 13521 3457 13558 3489 3 FreeSans 300 0 0 0 pd_h<4>
port 2 nsew
flabel metal1 s 11367 2074 11407 2204 7 FreeSans 300 180 0 0 vgnd_io
port 3 nsew
flabel metal1 s 7106 255 7151 307 8 FreeSans 300 180 0 0 drvlo_h_n
port 5 nsew
flabel metal1 s 9272 1616 9318 1662 7 FreeSans 300 180 0 0 slow_h
port 6 nsew
flabel metal1 s 8947 787 8999 833 6 FreeSans 300 180 0 0 pden_h_n
port 7 nsew
flabel metal1 s 151 2486 191 2688 3 FreeSans 300 180 0 0 vgnd_io
port 3 nsew
flabel metal1 s 151 1458 191 1588 3 FreeSans 300 180 0 0 vgnd_io
port 3 nsew
flabel metal1 s 9229 1870 9229 1870 3 FreeSans 400 0 0 0 pbias_out
flabel locali s 14147 3945 14185 3976 3 FreeSans 300 0 0 0 i2c_mode_h_n
port 8 nsew
flabel metal2 s 10022 2312 10022 2312 3 FreeSans 400 0 0 0 en_fast2_n<0>
flabel metal2 s 9761 2295 9761 2295 3 FreeSans 400 0 0 0 en_fast2_n<1>
flabel metal2 s 9346 1249 9393 1301 3 FreeSans 300 180 0 0 pd_h<2>
port 9 nsew
flabel metal2 s 9815 2932 9873 2984 7 FreeSans 300 180 0 0 pd_h<3>
port 10 nsew
<< properties >>
string GDS_END 87975798
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 87934804
string path 221.775 111.675 224.975 111.675 
<< end >>
