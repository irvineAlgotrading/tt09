magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< pdiff >>
rect 8492 2224 8506 2258
rect 8506 2195 9104 2224
rect 8812 2041 9104 2195
rect 9085 1895 9104 2041
rect 8812 1874 9104 1895
rect 10092 2042 10805 2224
rect 10092 2020 10391 2042
rect 10447 2020 10805 2042
rect 10092 1874 10374 2020
rect 10473 1840 10805 2020
rect 10609 1797 10805 1840
rect 10609 1752 10779 1797
rect 11718 966 11752 992
<< metal1 >>
rect 0 39220 342 39272
rect 11610 39220 12410 39272
rect 0 38981 342 39027
rect 11504 38981 12410 39027
rect 1762 35344 1790 35408
tri 5522 21681 5594 21753 sw
rect 5522 21675 5594 21681
rect 5522 21623 5542 21675
rect 5522 21611 5594 21623
rect 5522 21559 5542 21611
rect 5522 21547 5594 21559
rect 5522 21495 5542 21547
rect 5522 21489 5594 21495
tri 5522 21417 5594 21489 nw
rect 16 4783 77 4835
rect 12184 4783 12394 4835
<< via1 >>
rect 5542 21623 5594 21675
rect 5542 21559 5594 21611
rect 5542 21495 5594 21547
<< metal2 >>
rect 345 39112 478 39372
rect 1793 39112 2022 39372
rect 4996 39300 5048 39352
tri 7356 39112 7500 39256 se
rect 8477 39112 8867 39372
tri 7176 38932 7356 39112 se
rect 7356 38932 7500 39112
tri 7419 26517 7444 26542 se
rect 7444 26517 7500 38932
rect 12038 26940 12349 39372
rect 7419 26449 7500 26517
tri 7419 26429 7439 26449 ne
rect 7439 26448 7500 26449
rect 7439 26429 7481 26448
tri 7481 26429 7500 26448 nw
rect 5542 21675 5594 21681
rect 5542 21611 5594 21623
rect 5542 21547 5594 21559
rect 5542 21489 5594 21495
tri 7478 11203 7492 11217 se
rect 7492 11203 7520 11659
tri 7446 11171 7478 11203 se
rect 7478 11171 7488 11203
tri 7488 11171 7520 11203 nw
tri 7404 11129 7446 11171 se
tri 7446 11129 7488 11171 nw
tri 7362 11087 7404 11129 se
tri 7404 11087 7446 11129 nw
tri 7306 11031 7362 11087 se
tri 7362 11045 7404 11087 nw
rect 7306 4757 7362 11031
tri 7362 4757 7578 4973 sw
tri 7306 4703 7360 4757 nw
rect 3680 0 3732 660
rect 3836 0 3888 660
rect 4111 0 4163 660
rect 6141 0 6193 660
rect 7650 0 7702 660
rect 7883 0 7935 660
rect 12080 0 12132 660
<< metal3 >>
rect 0 9677 12420 10873
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_0
timestamp 1704896540
transform 0 -1 5594 1 0 21489
box 0 0 1 1
use sky130_fd_io__opamp_1  sky130_fd_io__opamp_1_0
timestamp 1704896540
transform 1 0 4429 0 1 28170
box -130 -1600 7181 11182
use sky130_fd_io__opamp_stage_1  sky130_fd_io__opamp_stage_1_0
timestamp 1704896540
transform 1 0 345 0 1 28200
box -286 209 8707 11170
use sky130_fd_io__refgen_com_m2m3_strap  sky130_fd_io__refgen_com_m2m3_strap_0
timestamp 1704896540
transform 1 0 8124 0 1 5761
box 0 0 364 858
use sky130_fd_io__refgen_com_m2m3_strap  sky130_fd_io__refgen_com_m2m3_strap_1
timestamp 1704896540
transform 1 0 11642 0 1 11193
box 0 0 364 858
use sky130_fd_io__refgen_com_m2m3_strap  sky130_fd_io__refgen_com_m2m3_strap_2
timestamp 1704896540
transform 1 0 7338 0 1 5761
box 0 0 364 858
use sky130_fd_io__refgen_com_m2m3_strap  sky130_fd_io__refgen_com_m2m3_strap_3
timestamp 1704896540
transform 1 0 10044 0 1 8477
box 0 0 364 858
use sky130_fd_io__refgen_com_m2m3_strap  sky130_fd_io__refgen_com_m2m3_strap_4
timestamp 1704896540
transform 1 0 7152 0 1 11193
box 0 0 364 858
use sky130_fd_io__refgen_com_m2m3_strap  sky130_fd_io__refgen_com_m2m3_strap_5
timestamp 1704896540
transform 1 0 11012 0 1 1608
box 0 0 364 858
use sky130_fd_io__refgen_com_m2m3_strap  sky130_fd_io__refgen_com_m2m3_strap_6
timestamp 1704896540
transform 1 0 6225 0 1 9835
box 0 0 364 858
use sky130_fd_io__refgen_com_m2m3_strap  sky130_fd_io__refgen_com_m2m3_strap_7
timestamp 1704896540
transform 1 0 4604 0 1 4324
box 0 0 364 858
use sky130_fd_io__refgen_com_m2m3_strap  sky130_fd_io__refgen_com_m2m3_strap_8
timestamp 1704896540
transform 1 0 2097 0 1 4324
box 0 0 364 858
use sky130_fd_io__refgen_com_m2m3_strap  sky130_fd_io__refgen_com_m2m3_strap_9
timestamp 1704896540
transform 1 0 6777 0 1 4324
box 0 0 364 858
use sky130_fd_io__refgen_com_m2m3_strap  sky130_fd_io__refgen_com_m2m3_strap_10
timestamp 1704896540
transform 1 0 4072 0 1 5761
box 0 0 364 858
use sky130_fd_io__refgen_com_m2m3_strap  sky130_fd_io__refgen_com_m2m3_strap_11
timestamp 1704896540
transform 1 0 435 0 1 5761
box 0 0 364 858
use sky130_fd_io__refgen_com_m2m3_strap  sky130_fd_io__refgen_com_m2m3_strap_12
timestamp 1704896540
transform 1 0 942 0 1 5761
box 0 0 364 858
use sky130_fd_io__refgen_com_m2m3_strap  sky130_fd_io__refgen_com_m2m3_strap_13
timestamp 1704896540
transform 1 0 36 0 1 4324
box 0 0 364 858
use sky130_fd_io__refgen_com_m2m3_strap  sky130_fd_io__refgen_com_m2m3_strap_14
timestamp 1704896540
transform 1 0 8799 0 1 2966
box 0 0 364 858
use sky130_fd_io__refgen_com_m2m3_strap  sky130_fd_io__refgen_com_m2m3_strap_15
timestamp 1704896540
transform 1 0 9696 0 1 2966
box 0 0 364 858
use sky130_fd_io__refgen_com_m2m3_strap  sky130_fd_io__refgen_com_m2m3_strap_16
timestamp 1704896540
transform 1 0 5626 0 1 2966
box 0 0 364 858
use sky130_fd_io__refgen_com_m2m3_strap  sky130_fd_io__refgen_com_m2m3_strap_17
timestamp 1704896540
transform 1 0 3312 0 1 2966
box 0 0 364 858
use sky130_fd_io__refgen_com_m2m3_strap  sky130_fd_io__refgen_com_m2m3_strap_18
timestamp 1704896540
transform 1 0 2710 0 1 2966
box 0 0 364 858
use sky130_fd_io__refgen_com_m2m3_strap  sky130_fd_io__refgen_com_m2m3_strap_19
timestamp 1704896540
transform 1 0 942 0 1 2966
box 0 0 364 858
use sky130_fd_io__refgen_com_m2m3_strap  sky130_fd_io__refgen_com_m2m3_strap_20
timestamp 1704896540
transform 1 0 435 0 1 2966
box 0 0 364 858
use sky130_fd_io__refgen_com_m2m3_strap  sky130_fd_io__refgen_com_m2m3_strap_21
timestamp 1704896540
transform 1 0 38 0 1 11193
box 0 0 364 858
use sky130_fd_io__refgen_com_m2m3_strap  sky130_fd_io__refgen_com_m2m3_strap_22
timestamp 1704896540
transform 1 0 3433 0 1 5761
box 0 0 364 858
use sky130_fd_io__refgen_com_m2m3_strap  sky130_fd_io__refgen_com_m2m3_strap_23
timestamp 1704896540
transform 1 0 1453 0 1 11193
box 0 0 364 858
use sky130_fd_io__refgen_in_cswblk  sky130_fd_io__refgen_in_cswblk_0
timestamp 1704896540
transform 1 0 5682 0 1 4703
box 0 -14 4074 1730
use sky130_fd_io__refgen_in_logic  sky130_fd_io__refgen_in_logic_0
timestamp 1704896540
transform 1 0 7306 0 1 6392
box -160 0 5076 2350
use sky130_fd_io__refgen_in_xlators  sky130_fd_io__refgen_in_xlators_0
timestamp 1704896540
transform 1 0 3621 0 1 754
box -285 -134 8728 5669
use sky130_fd_io__refgen_out_resblk  sky130_fd_io__refgen_out_resblk_0
timestamp 1704896540
transform 1 0 8568 0 1 8742
box -1422 -41 4089 18198
use sky130_fd_io__refgen_out_sub  sky130_fd_io__refgen_out_sub_0
timestamp 1704896540
transform 1 0 2203 0 1 11318
box -242 110 14565 34922
use sky130_fd_io__res_ntwk_vinref_1  sky130_fd_io__res_ntwk_vinref_1_0
timestamp 1704896540
transform 1 0 0 0 1 642
box 0 -1056 7492 27937
use sky130_fd_io__sio_bus_slice  sky130_fd_io__sio_bus_slice_0
timestamp 1704896540
transform 1 0 11410 0 1 0
box 0 250 1000 13599
use sky130_fd_io__sio_bus_slice  sky130_fd_io__sio_bus_slice_1
timestamp 1704896540
transform 1 0 10410 0 1 0
box 0 250 1000 13599
use sky130_fd_io__sio_bus_slice  sky130_fd_io__sio_bus_slice_2
timestamp 1704896540
transform 1 0 9410 0 1 0
box 0 250 1000 13599
use sky130_fd_io__sio_bus_slice  sky130_fd_io__sio_bus_slice_3
timestamp 1704896540
transform 1 0 8410 0 1 0
box 0 250 1000 13599
use sky130_fd_io__sio_bus_slice  sky130_fd_io__sio_bus_slice_4
timestamp 1704896540
transform 1 0 7410 0 1 0
box 0 250 1000 13599
use sky130_fd_io__sio_bus_slice  sky130_fd_io__sio_bus_slice_5
timestamp 1704896540
transform 1 0 6410 0 1 0
box 0 250 1000 13599
use sky130_fd_io__sio_bus_slice  sky130_fd_io__sio_bus_slice_6
timestamp 1704896540
transform 1 0 5410 0 1 0
box 0 250 1000 13599
use sky130_fd_io__sio_bus_slice  sky130_fd_io__sio_bus_slice_7
timestamp 1704896540
transform 1 0 4410 0 1 0
box 0 250 1000 13599
use sky130_fd_io__sio_bus_slice  sky130_fd_io__sio_bus_slice_8
timestamp 1704896540
transform 1 0 3410 0 1 0
box 0 250 1000 13599
use sky130_fd_io__sio_bus_slice  sky130_fd_io__sio_bus_slice_9
timestamp 1704896540
transform 1 0 2410 0 1 0
box 0 250 1000 13599
use sky130_fd_io__sio_bus_slice  sky130_fd_io__sio_bus_slice_10
timestamp 1704896540
transform 1 0 1410 0 1 0
box 0 250 1000 13599
use sky130_fd_io__sio_bus_slice  sky130_fd_io__sio_bus_slice_11
timestamp 1704896540
transform 1 0 410 0 1 0
box 0 250 1000 13599
use sky130_fd_io__sio_bus_slice  sky130_fd_io__sio_bus_slice_12
timestamp 1704896540
transform 1 0 0 0 1 0
box 0 250 1000 13599
use sky130_fd_io__top_refgen_overlay  sky130_fd_io__top_refgen_overlay_0
timestamp 1704896540
transform 1 0 -32569 0 1 0
box 32759 -333 44800 38878
<< labels >>
flabel comment s 2411 38835 2411 38835 0 FreeSans 1000 0 0 0 condiode
flabel metal1 s 16 4783 77 4835 3 FreeSans 200 0 0 0 vinref
port 4 nsew
flabel metal1 s 12337 38981 12410 39027 3 FreeSans 200 180 0 0 refleak_bias
port 2 nsew
flabel metal1 s 12337 39220 12410 39272 3 FreeSans 200 180 0 0 voutref
port 3 nsew
flabel metal1 s 0 39220 73 39272 3 FreeSans 200 0 0 0 voutref
port 3 nsew
flabel metal1 s 0 38981 73 39027 3 FreeSans 200 0 0 0 refleak_bias
port 2 nsew
flabel metal1 s 12333 4783 12394 4835 3 FreeSans 200 180 0 0 vinref
port 4 nsew
flabel metal2 s 7883 0 7935 20 3 FreeSans 200 90 0 0 vref_sel
port 5 nsew
flabel metal2 s 12080 0 12132 20 3 FreeSans 200 90 0 0 vreg_en
port 6 nsew
flabel metal2 s 3680 0 3732 20 3 FreeSans 200 90 0 0 vtrip_sel
port 7 nsew
flabel metal2 s 4111 0 4163 20 3 FreeSans 200 90 0 0 hld_h_n
port 8 nsew
flabel metal2 s 3836 0 3888 20 3 FreeSans 200 90 0 0 od_h
port 9 nsew
flabel metal2 s 7650 0 7702 20 3 FreeSans 200 90 0 0 ibuf_sel
port 10 nsew
flabel metal2 s 6141 0 6193 20 3 FreeSans 200 90 0 0 vohref
port 11 nsew
flabel metal2 s 4996 39300 5048 39352 3 FreeSans 200 270 0 0 vohref
port 11 nsew
flabel metal2 s 12038 39330 12349 39372 7 FreeSans 600 90 0 0 vcc_a
port 12 nsew
flabel metal2 s 8477 39330 8867 39372 7 FreeSans 600 90 0 0 vcc_a
port 12 nsew
flabel metal2 s 1793 39330 2022 39372 7 FreeSans 600 90 0 0 vcc_a
port 12 nsew
flabel metal2 s 345 39330 478 39372 7 FreeSans 600 90 0 0 vcc_a
port 12 nsew
<< properties >>
string GDS_END 80496494
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 80489604
<< end >>
