magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< dnwell >>
rect 1102 8123 10046 11806
rect 1102 80 13186 8123
<< nwell >>
rect 1130 13148 11178 14301
rect 1131 13144 11178 13148
rect 1131 12286 11177 13144
rect 1022 11526 10126 11886
rect 1022 7126 1382 11526
rect 3554 7126 3914 11526
rect 1022 6766 3914 7126
rect 1022 2366 1382 6766
rect 3554 3850 3914 6766
rect 5394 3850 5754 11526
rect 7234 7126 7594 11526
rect 9766 8203 10126 11526
rect 9766 7843 13266 8203
rect 9766 7126 10126 7843
rect 7234 6766 10126 7126
rect 7234 3850 7594 6766
rect 3554 3490 7594 3850
rect 3554 2366 3914 3490
rect 1022 2006 3914 2366
rect 1022 360 1382 2006
rect 7234 2366 7594 3490
rect 9766 2366 10126 6766
rect 7234 2006 10126 2366
rect 9766 360 10126 2006
rect 12906 360 13266 7843
rect 1022 0 13266 360
<< pwell >>
rect 1178 11975 11144 12197
rect 1442 11361 3494 11447
rect 1442 7205 3494 7291
rect 1442 6601 3494 6687
rect 3974 11302 5334 11388
rect 3974 3996 4060 11302
rect 5248 3996 5334 11302
rect 3974 3910 5334 3996
rect 5814 11302 7174 11388
rect 5814 3996 5900 11302
rect 7088 3996 7174 11302
rect 5814 3910 7174 3996
rect 7654 11361 9706 11447
rect 7654 7205 9706 7291
rect 7654 6601 9706 6687
rect 1442 2445 3494 2531
rect 3974 1946 4060 3404
rect 1442 1860 4060 1946
rect 3586 506 4060 1860
rect 1504 420 4060 506
rect 5250 3274 5336 3404
rect 5812 3274 5898 3404
rect 5250 3188 5898 3274
rect 5250 2570 5336 3188
rect 5812 2570 5898 3188
rect 5250 422 5898 2570
rect 7088 1946 7174 3404
rect 7654 2445 9706 2531
rect 7088 1860 9706 1946
rect 7088 506 7562 1860
rect 7088 420 9644 506
rect 10186 7645 12825 7731
rect 10186 506 10272 7645
rect 10186 420 12825 506
<< mvpdiff >>
rect 5165 12839 5226 13839
rect 5868 12839 5929 13839
<< mvpsubdiff >>
rect 1204 12137 1228 12171
rect 1262 12137 1297 12171
rect 1331 12137 1366 12171
rect 1400 12137 1435 12171
rect 1469 12137 1504 12171
rect 1538 12137 1573 12171
rect 1607 12137 1642 12171
rect 1676 12137 1711 12171
rect 1745 12137 1780 12171
rect 1814 12137 1849 12171
rect 1883 12137 1918 12171
rect 1952 12137 1987 12171
rect 2021 12137 2056 12171
rect 2090 12137 2125 12171
rect 2159 12137 2194 12171
rect 2228 12137 2263 12171
rect 2297 12137 2332 12171
rect 2366 12137 2401 12171
rect 2435 12137 2470 12171
rect 2504 12137 2539 12171
rect 2573 12137 2608 12171
rect 2642 12137 2677 12171
rect 2711 12137 2746 12171
rect 2780 12137 2815 12171
rect 2849 12137 2884 12171
rect 2918 12137 2953 12171
rect 2987 12137 3022 12171
rect 3056 12137 3091 12171
rect 3125 12137 3160 12171
rect 3194 12137 3229 12171
rect 3263 12137 3298 12171
rect 3332 12137 3367 12171
rect 3401 12137 3436 12171
rect 3470 12137 3505 12171
rect 3539 12137 3574 12171
rect 3608 12137 3643 12171
rect 3677 12137 3712 12171
rect 3746 12137 3781 12171
rect 3815 12137 3850 12171
rect 3884 12137 3919 12171
rect 3953 12137 3988 12171
rect 1204 12103 3988 12137
rect 1204 12069 1228 12103
rect 1262 12069 1297 12103
rect 1331 12069 1366 12103
rect 1400 12069 1435 12103
rect 1469 12069 1504 12103
rect 1538 12069 1573 12103
rect 1607 12069 1642 12103
rect 1676 12069 1711 12103
rect 1745 12069 1780 12103
rect 1814 12069 1849 12103
rect 1883 12069 1918 12103
rect 1952 12069 1987 12103
rect 2021 12069 2056 12103
rect 2090 12069 2125 12103
rect 2159 12069 2194 12103
rect 2228 12069 2263 12103
rect 2297 12069 2332 12103
rect 2366 12069 2401 12103
rect 2435 12069 2470 12103
rect 2504 12069 2539 12103
rect 2573 12069 2608 12103
rect 2642 12069 2677 12103
rect 2711 12069 2746 12103
rect 2780 12069 2815 12103
rect 2849 12069 2884 12103
rect 2918 12069 2953 12103
rect 2987 12069 3022 12103
rect 3056 12069 3091 12103
rect 3125 12069 3160 12103
rect 3194 12069 3229 12103
rect 3263 12069 3298 12103
rect 3332 12069 3367 12103
rect 3401 12069 3436 12103
rect 3470 12069 3505 12103
rect 3539 12069 3574 12103
rect 3608 12069 3643 12103
rect 3677 12069 3712 12103
rect 3746 12069 3781 12103
rect 3815 12069 3850 12103
rect 3884 12069 3919 12103
rect 3953 12069 3988 12103
rect 1204 12035 3988 12069
rect 1204 12001 1228 12035
rect 1262 12001 1297 12035
rect 1331 12001 1366 12035
rect 1400 12001 1435 12035
rect 1469 12001 1504 12035
rect 1538 12001 1573 12035
rect 1607 12001 1642 12035
rect 1676 12001 1711 12035
rect 1745 12001 1780 12035
rect 1814 12001 1849 12035
rect 1883 12001 1918 12035
rect 1952 12001 1987 12035
rect 2021 12001 2056 12035
rect 2090 12001 2125 12035
rect 2159 12001 2194 12035
rect 2228 12001 2263 12035
rect 2297 12001 2332 12035
rect 2366 12001 2401 12035
rect 2435 12001 2470 12035
rect 2504 12001 2539 12035
rect 2573 12001 2608 12035
rect 2642 12001 2677 12035
rect 2711 12001 2746 12035
rect 2780 12001 2815 12035
rect 2849 12001 2884 12035
rect 2918 12001 2953 12035
rect 2987 12001 3022 12035
rect 3056 12001 3091 12035
rect 3125 12001 3160 12035
rect 3194 12001 3229 12035
rect 3263 12001 3298 12035
rect 3332 12001 3367 12035
rect 3401 12001 3436 12035
rect 3470 12001 3505 12035
rect 3539 12001 3574 12035
rect 3608 12001 3643 12035
rect 3677 12001 3712 12035
rect 3746 12001 3781 12035
rect 3815 12001 3850 12035
rect 3884 12001 3919 12035
rect 3953 12001 3988 12035
rect 11094 12001 11118 12171
rect 1468 11387 1492 11421
rect 1526 11387 1561 11421
rect 1595 11387 1630 11421
rect 1664 11387 1699 11421
rect 1733 11387 1768 11421
rect 1802 11387 1837 11421
rect 1871 11387 1906 11421
rect 1940 11387 1975 11421
rect 2009 11387 2044 11421
rect 2078 11387 2113 11421
rect 2147 11387 2182 11421
rect 2216 11387 2251 11421
rect 2285 11387 2320 11421
rect 2354 11387 2389 11421
rect 2423 11387 2458 11421
rect 2492 11387 2526 11421
rect 2560 11387 2594 11421
rect 2628 11387 2662 11421
rect 2696 11387 2730 11421
rect 2764 11387 2798 11421
rect 2832 11387 2866 11421
rect 2900 11387 2934 11421
rect 2968 11387 3002 11421
rect 3036 11387 3070 11421
rect 3104 11387 3138 11421
rect 3172 11387 3206 11421
rect 3240 11387 3274 11421
rect 3308 11387 3342 11421
rect 3376 11387 3410 11421
rect 3444 11387 3468 11421
rect 1468 7231 1492 7265
rect 1526 7231 1561 7265
rect 1595 7231 1630 7265
rect 1664 7231 1699 7265
rect 1733 7231 1768 7265
rect 1802 7231 1837 7265
rect 1871 7231 1906 7265
rect 1940 7231 1975 7265
rect 2009 7231 2044 7265
rect 2078 7231 2113 7265
rect 2147 7231 2182 7265
rect 2216 7231 2251 7265
rect 2285 7231 2320 7265
rect 2354 7231 2389 7265
rect 2423 7231 2458 7265
rect 2492 7231 2526 7265
rect 2560 7231 2594 7265
rect 2628 7231 2662 7265
rect 2696 7231 2730 7265
rect 2764 7231 2798 7265
rect 2832 7231 2866 7265
rect 2900 7231 2934 7265
rect 2968 7231 3002 7265
rect 3036 7231 3070 7265
rect 3104 7231 3138 7265
rect 3172 7231 3206 7265
rect 3240 7231 3274 7265
rect 3308 7231 3342 7265
rect 3376 7231 3410 7265
rect 3444 7231 3468 7265
rect 1468 6627 1492 6661
rect 1526 6627 1561 6661
rect 1595 6627 1630 6661
rect 1664 6627 1699 6661
rect 1733 6627 1768 6661
rect 1802 6627 1837 6661
rect 1871 6627 1906 6661
rect 1940 6627 1975 6661
rect 2009 6627 2044 6661
rect 2078 6627 2113 6661
rect 2147 6627 2182 6661
rect 2216 6627 2251 6661
rect 2285 6627 2320 6661
rect 2354 6627 2389 6661
rect 2423 6627 2458 6661
rect 2492 6627 2526 6661
rect 2560 6627 2594 6661
rect 2628 6627 2662 6661
rect 2696 6627 2730 6661
rect 2764 6627 2798 6661
rect 2832 6627 2866 6661
rect 2900 6627 2934 6661
rect 2968 6627 3002 6661
rect 3036 6627 3070 6661
rect 3104 6627 3138 6661
rect 3172 6627 3206 6661
rect 3240 6627 3274 6661
rect 3308 6627 3342 6661
rect 3376 6627 3410 6661
rect 3444 6627 3468 6661
rect 4000 11239 4034 11362
rect 4068 11328 4102 11362
rect 4136 11328 4170 11362
rect 4204 11328 4238 11362
rect 4272 11328 4306 11362
rect 4340 11328 4374 11362
rect 4408 11328 4442 11362
rect 4476 11328 4510 11362
rect 4544 11328 4578 11362
rect 4612 11328 4646 11362
rect 4680 11328 4714 11362
rect 4748 11328 4782 11362
rect 4816 11328 4850 11362
rect 4884 11328 4918 11362
rect 4952 11328 4986 11362
rect 5020 11328 5054 11362
rect 5088 11328 5122 11362
rect 5156 11328 5190 11362
rect 5224 11328 5308 11362
rect 4000 11170 4034 11205
rect 5274 11239 5308 11328
rect 4000 11101 4034 11136
rect 5274 11170 5308 11205
rect 5274 11101 5308 11136
rect 4000 11032 4034 11067
rect 4000 10963 4034 10998
rect 4000 10894 4034 10929
rect 4000 10825 4034 10860
rect 4000 10756 4034 10791
rect 4000 10687 4034 10722
rect 4000 10618 4034 10653
rect 4000 10549 4034 10584
rect 4000 10480 4034 10515
rect 4000 10411 4034 10446
rect 4000 10342 4034 10377
rect 4000 10273 4034 10308
rect 5274 11032 5308 11067
rect 5274 10963 5308 10998
rect 5274 10894 5308 10929
rect 5274 10825 5308 10860
rect 5274 10756 5308 10791
rect 5274 10687 5308 10722
rect 5274 10618 5308 10653
rect 5274 10549 5308 10584
rect 5274 10480 5308 10515
rect 5274 10411 5308 10446
rect 5274 10342 5308 10377
rect 5274 10273 5308 10308
rect 4000 10204 4034 10239
rect 5274 10204 5308 10239
rect 4000 10135 4034 10170
rect 4000 10066 4034 10101
rect 4000 9997 4034 10032
rect 4000 9928 4034 9963
rect 4000 9859 4034 9894
rect 4000 9790 4034 9825
rect 4000 9721 4034 9756
rect 4000 9652 4034 9687
rect 4000 9583 4034 9618
rect 4000 9514 4034 9549
rect 4000 9445 4034 9480
rect 4000 9376 4034 9411
rect 5274 10135 5308 10170
rect 5274 10066 5308 10101
rect 5274 9997 5308 10032
rect 5274 9928 5308 9963
rect 5274 9859 5308 9894
rect 5274 9790 5308 9825
rect 5274 9721 5308 9756
rect 5274 9652 5308 9687
rect 5274 9583 5308 9618
rect 5274 9514 5308 9549
rect 5274 9445 5308 9480
rect 4000 9307 4034 9342
rect 5274 9376 5308 9411
rect 4000 9238 4034 9273
rect 4000 9169 4034 9204
rect 4000 9100 4034 9135
rect 4000 9031 4034 9066
rect 4000 8962 4034 8997
rect 4000 8893 4034 8928
rect 4000 8824 4034 8859
rect 4000 8755 4034 8790
rect 4000 8686 4034 8721
rect 4000 8617 4034 8652
rect 4000 8548 4034 8583
rect 5274 9307 5308 9342
rect 5274 9238 5308 9273
rect 5274 9169 5308 9204
rect 5274 9100 5308 9135
rect 5274 9031 5308 9066
rect 5274 8962 5308 8997
rect 5274 8893 5308 8928
rect 5274 8824 5308 8859
rect 5274 8755 5308 8790
rect 5274 8686 5308 8721
rect 5274 8617 5308 8652
rect 5274 8548 5308 8583
rect 4000 8479 4034 8514
rect 5274 8479 5308 8514
rect 4000 8410 4034 8445
rect 4000 8341 4034 8376
rect 4000 8272 4034 8307
rect 4000 8203 4034 8238
rect 4000 8134 4034 8169
rect 4000 8065 4034 8100
rect 4000 7996 4034 8031
rect 4000 7927 4034 7962
rect 4000 7858 4034 7893
rect 4000 7789 4034 7824
rect 4000 7720 4034 7755
rect 4000 7651 4034 7686
rect 5274 8410 5308 8445
rect 5274 8341 5308 8376
rect 5274 8272 5308 8307
rect 5274 8203 5308 8238
rect 5274 8134 5308 8169
rect 5274 8065 5308 8100
rect 5274 7996 5308 8031
rect 5274 7927 5308 7962
rect 5274 7858 5308 7893
rect 5274 7789 5308 7824
rect 5274 7720 5308 7755
rect 5274 7651 5308 7686
rect 4000 7583 4034 7617
rect 4000 7515 4034 7549
rect 4000 7447 4034 7481
rect 4000 7379 4034 7413
rect 4000 7311 4034 7345
rect 4000 7243 4034 7277
rect 4000 7175 4034 7209
rect 4000 7107 4034 7141
rect 4000 7039 4034 7073
rect 4000 6971 4034 7005
rect 4000 6903 4034 6937
rect 4000 6835 4034 6869
rect 5274 7583 5308 7617
rect 5274 7515 5308 7549
rect 5274 7447 5308 7481
rect 5274 7379 5308 7413
rect 5274 7311 5308 7345
rect 5274 7243 5308 7277
rect 5274 7175 5308 7209
rect 5274 7107 5308 7141
rect 5274 7039 5308 7073
rect 5274 6971 5308 7005
rect 5274 6903 5308 6937
rect 5274 6835 5308 6869
rect 4000 6767 4034 6801
rect 5274 6767 5308 6801
rect 4000 6699 4034 6733
rect 4000 6631 4034 6665
rect 4000 6563 4034 6597
rect 4000 6495 4034 6529
rect 4000 6427 4034 6461
rect 4000 6359 4034 6393
rect 4000 6291 4034 6325
rect 4000 6223 4034 6257
rect 4000 6155 4034 6189
rect 4000 6087 4034 6121
rect 4000 6019 4034 6053
rect 4000 5951 4034 5985
rect 5274 6699 5308 6733
rect 5274 6631 5308 6665
rect 5274 6563 5308 6597
rect 5274 6495 5308 6529
rect 5274 6427 5308 6461
rect 5274 6359 5308 6393
rect 5274 6291 5308 6325
rect 5274 6223 5308 6257
rect 5274 6155 5308 6189
rect 5274 6087 5308 6121
rect 5274 6019 5308 6053
rect 4000 5883 4034 5917
rect 5274 5951 5308 5985
rect 4000 5815 4034 5849
rect 4000 5747 4034 5781
rect 4000 5679 4034 5713
rect 4000 5611 4034 5645
rect 4000 5543 4034 5577
rect 4000 5475 4034 5509
rect 4000 5407 4034 5441
rect 4000 5339 4034 5373
rect 4000 5271 4034 5305
rect 4000 5203 4034 5237
rect 4000 5135 4034 5169
rect 5274 5883 5308 5917
rect 5274 5815 5308 5849
rect 5274 5747 5308 5781
rect 5274 5679 5308 5713
rect 5274 5611 5308 5645
rect 5274 5543 5308 5577
rect 5274 5475 5308 5509
rect 5274 5407 5308 5441
rect 5274 5339 5308 5373
rect 5274 5271 5308 5305
rect 5274 5203 5308 5237
rect 5274 5135 5308 5169
rect 4000 5067 4034 5101
rect 5274 5067 5308 5101
rect 4000 4999 4034 5033
rect 4000 4931 4034 4965
rect 4000 4863 4034 4897
rect 4000 4795 4034 4829
rect 4000 4727 4034 4761
rect 4000 4659 4034 4693
rect 4000 4591 4034 4625
rect 4000 4523 4034 4557
rect 4000 4455 4034 4489
rect 4000 4387 4034 4421
rect 4000 4319 4034 4353
rect 4000 4251 4034 4285
rect 5274 4999 5308 5033
rect 5274 4931 5308 4965
rect 5274 4863 5308 4897
rect 5274 4795 5308 4829
rect 5274 4727 5308 4761
rect 5274 4659 5308 4693
rect 5274 4591 5308 4625
rect 5274 4523 5308 4557
rect 5274 4455 5308 4489
rect 5274 4387 5308 4421
rect 5274 4319 5308 4353
rect 4000 4183 4034 4217
rect 5274 4251 5308 4285
rect 4000 4115 4034 4149
rect 5274 4183 5308 4217
rect 5274 4115 5308 4149
rect 4000 3936 4034 4081
rect 5274 4004 5308 4081
rect 4068 3936 4102 3970
rect 4136 3936 4170 3970
rect 4204 3936 4238 3970
rect 4272 3936 4306 3970
rect 4340 3936 4374 3970
rect 4408 3936 4442 3970
rect 4476 3936 4510 3970
rect 4544 3936 4578 3970
rect 4612 3936 4646 3970
rect 4680 3936 4714 3970
rect 4748 3936 4782 3970
rect 4816 3936 4850 3970
rect 4884 3936 4918 3970
rect 4952 3936 4986 3970
rect 5020 3936 5054 3970
rect 5088 3936 5122 3970
rect 5156 3936 5190 3970
rect 5224 3936 5308 3970
rect 7680 11387 7704 11421
rect 7738 11387 7772 11421
rect 7806 11387 7840 11421
rect 7874 11387 7908 11421
rect 7942 11387 7976 11421
rect 8010 11387 8044 11421
rect 8078 11387 8112 11421
rect 8146 11387 8180 11421
rect 8214 11387 8248 11421
rect 8282 11387 8316 11421
rect 8350 11387 8384 11421
rect 8418 11387 8452 11421
rect 8486 11387 8520 11421
rect 8554 11387 8588 11421
rect 8622 11387 8656 11421
rect 8690 11387 8725 11421
rect 8759 11387 8794 11421
rect 8828 11387 8863 11421
rect 8897 11387 8932 11421
rect 8966 11387 9001 11421
rect 9035 11387 9070 11421
rect 9104 11387 9139 11421
rect 9173 11387 9208 11421
rect 9242 11387 9277 11421
rect 9311 11387 9346 11421
rect 9380 11387 9415 11421
rect 9449 11387 9484 11421
rect 9518 11387 9553 11421
rect 9587 11387 9622 11421
rect 9656 11387 9680 11421
rect 5840 11239 5874 11362
rect 5908 11328 5942 11362
rect 5976 11328 6010 11362
rect 6044 11328 6078 11362
rect 6112 11328 6146 11362
rect 6180 11328 6214 11362
rect 6248 11328 6282 11362
rect 6316 11328 6350 11362
rect 6384 11328 6418 11362
rect 6452 11328 6486 11362
rect 6520 11328 6554 11362
rect 6588 11328 6622 11362
rect 6656 11328 6690 11362
rect 6724 11328 6758 11362
rect 6792 11328 6826 11362
rect 6860 11328 6894 11362
rect 6928 11328 6962 11362
rect 6996 11328 7030 11362
rect 7064 11328 7148 11362
rect 5840 11170 5874 11205
rect 7114 11239 7148 11328
rect 5840 11101 5874 11136
rect 7114 11170 7148 11205
rect 7114 11101 7148 11136
rect 5840 11032 5874 11067
rect 5840 10963 5874 10998
rect 5840 10894 5874 10929
rect 5840 10825 5874 10860
rect 5840 10756 5874 10791
rect 5840 10687 5874 10722
rect 5840 10618 5874 10653
rect 5840 10549 5874 10584
rect 5840 10480 5874 10515
rect 5840 10411 5874 10446
rect 5840 10342 5874 10377
rect 5840 10273 5874 10308
rect 7114 11032 7148 11067
rect 7114 10963 7148 10998
rect 7114 10894 7148 10929
rect 7114 10825 7148 10860
rect 7114 10756 7148 10791
rect 7114 10687 7148 10722
rect 7114 10618 7148 10653
rect 7114 10549 7148 10584
rect 7114 10480 7148 10515
rect 7114 10411 7148 10446
rect 7114 10342 7148 10377
rect 7114 10273 7148 10308
rect 5840 10204 5874 10239
rect 7114 10204 7148 10239
rect 5840 10135 5874 10170
rect 5840 10066 5874 10101
rect 5840 9997 5874 10032
rect 5840 9928 5874 9963
rect 5840 9859 5874 9894
rect 5840 9790 5874 9825
rect 5840 9721 5874 9756
rect 5840 9652 5874 9687
rect 5840 9583 5874 9618
rect 5840 9514 5874 9549
rect 5840 9445 5874 9480
rect 5840 9376 5874 9411
rect 7114 10135 7148 10170
rect 7114 10066 7148 10101
rect 7114 9997 7148 10032
rect 7114 9928 7148 9963
rect 7114 9859 7148 9894
rect 7114 9790 7148 9825
rect 7114 9721 7148 9756
rect 7114 9652 7148 9687
rect 7114 9583 7148 9618
rect 7114 9514 7148 9549
rect 7114 9445 7148 9480
rect 5840 9307 5874 9342
rect 7114 9376 7148 9411
rect 5840 9238 5874 9273
rect 5840 9169 5874 9204
rect 5840 9100 5874 9135
rect 5840 9031 5874 9066
rect 5840 8962 5874 8997
rect 5840 8893 5874 8928
rect 5840 8824 5874 8859
rect 5840 8755 5874 8790
rect 5840 8686 5874 8721
rect 5840 8617 5874 8652
rect 5840 8548 5874 8583
rect 7114 9307 7148 9342
rect 7114 9238 7148 9273
rect 7114 9169 7148 9204
rect 7114 9100 7148 9135
rect 7114 9031 7148 9066
rect 7114 8962 7148 8997
rect 7114 8893 7148 8928
rect 7114 8824 7148 8859
rect 7114 8755 7148 8790
rect 7114 8686 7148 8721
rect 7114 8617 7148 8652
rect 7114 8548 7148 8583
rect 5840 8479 5874 8514
rect 7114 8479 7148 8514
rect 5840 8410 5874 8445
rect 5840 8341 5874 8376
rect 5840 8272 5874 8307
rect 5840 8203 5874 8238
rect 5840 8134 5874 8169
rect 5840 8065 5874 8100
rect 5840 7996 5874 8031
rect 5840 7927 5874 7962
rect 5840 7858 5874 7893
rect 5840 7789 5874 7824
rect 5840 7720 5874 7755
rect 5840 7651 5874 7686
rect 7114 8410 7148 8445
rect 7114 8341 7148 8376
rect 7114 8272 7148 8307
rect 7114 8203 7148 8238
rect 7114 8134 7148 8169
rect 7114 8065 7148 8100
rect 7114 7996 7148 8031
rect 7114 7927 7148 7962
rect 7114 7858 7148 7893
rect 7114 7789 7148 7824
rect 7114 7720 7148 7755
rect 7114 7651 7148 7686
rect 5840 7583 5874 7617
rect 5840 7515 5874 7549
rect 5840 7447 5874 7481
rect 5840 7379 5874 7413
rect 5840 7311 5874 7345
rect 5840 7243 5874 7277
rect 5840 7175 5874 7209
rect 5840 7107 5874 7141
rect 5840 7039 5874 7073
rect 5840 6971 5874 7005
rect 5840 6903 5874 6937
rect 5840 6835 5874 6869
rect 7114 7583 7148 7617
rect 7114 7515 7148 7549
rect 7114 7447 7148 7481
rect 7114 7379 7148 7413
rect 7114 7311 7148 7345
rect 7114 7243 7148 7277
rect 7114 7175 7148 7209
rect 7114 7107 7148 7141
rect 7114 7039 7148 7073
rect 7114 6971 7148 7005
rect 7114 6903 7148 6937
rect 7114 6835 7148 6869
rect 5840 6767 5874 6801
rect 7114 6767 7148 6801
rect 5840 6699 5874 6733
rect 5840 6631 5874 6665
rect 5840 6563 5874 6597
rect 5840 6495 5874 6529
rect 5840 6427 5874 6461
rect 5840 6359 5874 6393
rect 5840 6291 5874 6325
rect 5840 6223 5874 6257
rect 5840 6155 5874 6189
rect 5840 6087 5874 6121
rect 5840 6019 5874 6053
rect 5840 5951 5874 5985
rect 7114 6699 7148 6733
rect 7114 6631 7148 6665
rect 7114 6563 7148 6597
rect 7114 6495 7148 6529
rect 7114 6427 7148 6461
rect 7114 6359 7148 6393
rect 7114 6291 7148 6325
rect 7114 6223 7148 6257
rect 7114 6155 7148 6189
rect 7114 6087 7148 6121
rect 7114 6019 7148 6053
rect 5840 5883 5874 5917
rect 7114 5951 7148 5985
rect 5840 5815 5874 5849
rect 5840 5747 5874 5781
rect 5840 5679 5874 5713
rect 5840 5611 5874 5645
rect 5840 5543 5874 5577
rect 5840 5475 5874 5509
rect 5840 5407 5874 5441
rect 5840 5339 5874 5373
rect 5840 5271 5874 5305
rect 5840 5203 5874 5237
rect 5840 5135 5874 5169
rect 7114 5883 7148 5917
rect 7114 5815 7148 5849
rect 7114 5747 7148 5781
rect 7114 5679 7148 5713
rect 7114 5611 7148 5645
rect 7114 5543 7148 5577
rect 7114 5475 7148 5509
rect 7114 5407 7148 5441
rect 7114 5339 7148 5373
rect 7114 5271 7148 5305
rect 7114 5203 7148 5237
rect 7114 5135 7148 5169
rect 5840 5067 5874 5101
rect 7114 5067 7148 5101
rect 5840 4999 5874 5033
rect 5840 4931 5874 4965
rect 5840 4863 5874 4897
rect 5840 4795 5874 4829
rect 5840 4727 5874 4761
rect 5840 4659 5874 4693
rect 5840 4591 5874 4625
rect 5840 4523 5874 4557
rect 5840 4455 5874 4489
rect 5840 4387 5874 4421
rect 5840 4319 5874 4353
rect 5840 4251 5874 4285
rect 7114 4999 7148 5033
rect 7114 4931 7148 4965
rect 7114 4863 7148 4897
rect 7114 4795 7148 4829
rect 7114 4727 7148 4761
rect 7114 4659 7148 4693
rect 7114 4591 7148 4625
rect 7114 4523 7148 4557
rect 7114 4455 7148 4489
rect 7114 4387 7148 4421
rect 7114 4319 7148 4353
rect 5840 4183 5874 4217
rect 7114 4251 7148 4285
rect 5840 4115 5874 4149
rect 7114 4183 7148 4217
rect 7114 4115 7148 4149
rect 5840 3936 5874 4081
rect 7114 4004 7148 4081
rect 5908 3936 5942 3970
rect 5976 3936 6010 3970
rect 6044 3936 6078 3970
rect 6112 3936 6146 3970
rect 6180 3936 6214 3970
rect 6248 3936 6282 3970
rect 6316 3936 6350 3970
rect 6384 3936 6418 3970
rect 6452 3936 6486 3970
rect 6520 3936 6554 3970
rect 6588 3936 6622 3970
rect 6656 3936 6690 3970
rect 6724 3936 6758 3970
rect 6792 3936 6826 3970
rect 6860 3936 6894 3970
rect 6928 3936 6962 3970
rect 6996 3936 7030 3970
rect 7064 3936 7148 3970
rect 7680 7231 7704 7265
rect 7738 7231 7772 7265
rect 7806 7231 7840 7265
rect 7874 7231 7908 7265
rect 7942 7231 7976 7265
rect 8010 7231 8044 7265
rect 8078 7231 8112 7265
rect 8146 7231 8180 7265
rect 8214 7231 8248 7265
rect 8282 7231 8316 7265
rect 8350 7231 8384 7265
rect 8418 7231 8452 7265
rect 8486 7231 8520 7265
rect 8554 7231 8588 7265
rect 8622 7231 8656 7265
rect 8690 7231 8725 7265
rect 8759 7231 8794 7265
rect 8828 7231 8863 7265
rect 8897 7231 8932 7265
rect 8966 7231 9001 7265
rect 9035 7231 9070 7265
rect 9104 7231 9139 7265
rect 9173 7231 9208 7265
rect 9242 7231 9277 7265
rect 9311 7231 9346 7265
rect 9380 7231 9415 7265
rect 9449 7231 9484 7265
rect 9518 7231 9553 7265
rect 9587 7231 9622 7265
rect 9656 7231 9680 7265
rect 7680 6627 7704 6661
rect 7738 6627 7772 6661
rect 7806 6627 7840 6661
rect 7874 6627 7908 6661
rect 7942 6627 7976 6661
rect 8010 6627 8044 6661
rect 8078 6627 8112 6661
rect 8146 6627 8180 6661
rect 8214 6627 8248 6661
rect 8282 6627 8316 6661
rect 8350 6627 8384 6661
rect 8418 6627 8452 6661
rect 8486 6627 8520 6661
rect 8554 6627 8588 6661
rect 8622 6627 8656 6661
rect 8690 6627 8725 6661
rect 8759 6627 8794 6661
rect 8828 6627 8863 6661
rect 8897 6627 8932 6661
rect 8966 6627 9001 6661
rect 9035 6627 9070 6661
rect 9104 6627 9139 6661
rect 9173 6627 9208 6661
rect 9242 6627 9277 6661
rect 9311 6627 9346 6661
rect 9380 6627 9415 6661
rect 9449 6627 9484 6661
rect 9518 6627 9553 6661
rect 9587 6627 9622 6661
rect 9656 6627 9680 6661
rect 1468 2471 1492 2505
rect 1526 2471 1561 2505
rect 1595 2471 1630 2505
rect 1664 2471 1699 2505
rect 1733 2471 1768 2505
rect 1802 2471 1837 2505
rect 1871 2471 1906 2505
rect 1940 2471 1975 2505
rect 2009 2471 2044 2505
rect 2078 2471 2113 2505
rect 2147 2471 2182 2505
rect 2216 2471 2251 2505
rect 2285 2471 2320 2505
rect 2354 2471 2389 2505
rect 2423 2471 2458 2505
rect 2492 2471 2526 2505
rect 2560 2471 2594 2505
rect 2628 2471 2662 2505
rect 2696 2471 2730 2505
rect 2764 2471 2798 2505
rect 2832 2471 2866 2505
rect 2900 2471 2934 2505
rect 2968 2471 3002 2505
rect 3036 2471 3070 2505
rect 3104 2471 3138 2505
rect 3172 2471 3206 2505
rect 3240 2471 3274 2505
rect 3308 2471 3342 2505
rect 3376 2471 3410 2505
rect 3444 2471 3468 2505
rect 4000 3354 4034 3378
rect 5276 3354 5310 3378
rect 4000 3285 4034 3320
rect 4000 3216 4034 3251
rect 4000 3147 4034 3182
rect 5276 3285 5310 3320
rect 5276 3248 5310 3251
rect 5838 3354 5872 3378
rect 7114 3354 7148 3378
rect 5838 3285 5872 3320
rect 5838 3248 5872 3251
rect 5276 3216 5344 3248
rect 5310 3214 5344 3216
rect 5378 3214 5415 3248
rect 5449 3214 5486 3248
rect 5520 3214 5557 3248
rect 5591 3214 5628 3248
rect 5662 3214 5699 3248
rect 5733 3214 5770 3248
rect 5804 3216 5872 3248
rect 5804 3214 5838 3216
rect 5276 3147 5310 3182
rect 4000 3078 4034 3113
rect 5276 3078 5310 3113
rect 5838 3147 5872 3182
rect 7114 3285 7148 3320
rect 7114 3216 7148 3251
rect 7114 3147 7148 3182
rect 4000 3009 4034 3044
rect 4000 2940 4034 2975
rect 4000 2871 4034 2906
rect 5276 3009 5310 3044
rect 5276 2940 5310 2975
rect 5276 2871 5310 2906
rect 4000 2802 4034 2837
rect 4000 2733 4034 2768
rect 4000 2664 4034 2699
rect 4000 2595 4034 2630
rect 5276 2802 5310 2837
rect 5276 2733 5310 2768
rect 5276 2664 5310 2699
rect 5838 3078 5872 3113
rect 7114 3078 7148 3113
rect 5838 3009 5872 3044
rect 5838 2940 5872 2975
rect 5838 2871 5872 2906
rect 7114 3009 7148 3044
rect 7114 2940 7148 2975
rect 7114 2871 7148 2906
rect 5838 2802 5872 2837
rect 5838 2733 5872 2768
rect 4000 2526 4034 2561
rect 5276 2595 5310 2630
rect 4000 2457 4034 2492
rect 4000 2388 4034 2423
rect 5276 2544 5310 2561
rect 5838 2664 5872 2699
rect 5838 2595 5872 2630
rect 7114 2802 7148 2837
rect 7114 2733 7148 2768
rect 7114 2664 7148 2699
rect 5838 2544 5872 2561
rect 7114 2595 7148 2630
rect 5276 2526 5872 2544
rect 5310 2520 5838 2526
rect 5310 2492 5359 2520
rect 5276 2486 5359 2492
rect 5393 2486 5427 2520
rect 5461 2486 5495 2520
rect 5529 2486 5563 2520
rect 5597 2486 5631 2520
rect 5665 2486 5699 2520
rect 5733 2486 5767 2520
rect 5801 2492 5838 2520
rect 5801 2486 5872 2492
rect 5276 2457 5872 2486
rect 5310 2451 5838 2457
rect 5310 2423 5359 2451
rect 5276 2417 5359 2423
rect 5393 2417 5427 2451
rect 5461 2417 5495 2451
rect 5529 2417 5563 2451
rect 5597 2417 5631 2451
rect 5665 2417 5699 2451
rect 5733 2417 5767 2451
rect 5801 2423 5838 2451
rect 5801 2417 5872 2423
rect 5276 2388 5872 2417
rect 4000 2319 4034 2354
rect 5310 2382 5838 2388
rect 5310 2354 5359 2382
rect 5276 2348 5359 2354
rect 5393 2348 5427 2382
rect 5461 2348 5495 2382
rect 5529 2348 5563 2382
rect 5597 2348 5631 2382
rect 5665 2348 5699 2382
rect 5733 2348 5767 2382
rect 5801 2354 5838 2382
rect 7114 2526 7148 2561
rect 7114 2457 7148 2492
rect 7114 2388 7148 2423
rect 5801 2348 5872 2354
rect 5276 2319 5872 2348
rect 4000 2250 4034 2285
rect 4000 2181 4034 2216
rect 4000 2112 4034 2147
rect 5310 2313 5838 2319
rect 5310 2285 5359 2313
rect 5276 2279 5359 2285
rect 5393 2279 5427 2313
rect 5461 2279 5495 2313
rect 5529 2279 5563 2313
rect 5597 2279 5631 2313
rect 5665 2279 5699 2313
rect 5733 2279 5767 2313
rect 5801 2285 5838 2313
rect 7114 2319 7148 2354
rect 5801 2279 5872 2285
rect 5276 2250 5872 2279
rect 5310 2244 5838 2250
rect 5310 2216 5359 2244
rect 5276 2210 5359 2216
rect 5393 2210 5427 2244
rect 5461 2210 5495 2244
rect 5529 2210 5563 2244
rect 5597 2210 5631 2244
rect 5665 2210 5699 2244
rect 5733 2210 5767 2244
rect 5801 2216 5838 2244
rect 5801 2210 5872 2216
rect 5276 2181 5872 2210
rect 5310 2175 5838 2181
rect 5310 2147 5359 2175
rect 5276 2141 5359 2147
rect 5393 2141 5427 2175
rect 5461 2141 5495 2175
rect 5529 2141 5563 2175
rect 5597 2141 5631 2175
rect 5665 2141 5699 2175
rect 5733 2141 5767 2175
rect 5801 2147 5838 2175
rect 5801 2141 5872 2147
rect 5276 2112 5872 2141
rect 4000 2043 4034 2078
rect 5310 2106 5838 2112
rect 5310 2078 5359 2106
rect 5276 2072 5359 2078
rect 5393 2072 5427 2106
rect 5461 2072 5495 2106
rect 5529 2072 5563 2106
rect 5597 2072 5631 2106
rect 5665 2072 5699 2106
rect 5733 2072 5767 2106
rect 5801 2078 5838 2106
rect 7114 2250 7148 2285
rect 7114 2181 7148 2216
rect 7680 2471 7704 2505
rect 7738 2471 7772 2505
rect 7806 2471 7840 2505
rect 7874 2471 7908 2505
rect 7942 2471 7976 2505
rect 8010 2471 8044 2505
rect 8078 2471 8112 2505
rect 8146 2471 8180 2505
rect 8214 2471 8248 2505
rect 8282 2471 8316 2505
rect 8350 2471 8384 2505
rect 8418 2471 8452 2505
rect 8486 2471 8520 2505
rect 8554 2471 8588 2505
rect 8622 2471 8656 2505
rect 8690 2471 8725 2505
rect 8759 2471 8794 2505
rect 8828 2471 8863 2505
rect 8897 2471 8932 2505
rect 8966 2471 9001 2505
rect 9035 2471 9070 2505
rect 9104 2471 9139 2505
rect 9173 2471 9208 2505
rect 9242 2471 9277 2505
rect 9311 2471 9346 2505
rect 9380 2471 9415 2505
rect 9449 2471 9484 2505
rect 9518 2471 9553 2505
rect 9587 2471 9622 2505
rect 9656 2471 9680 2505
rect 7114 2112 7148 2147
rect 5801 2072 5872 2078
rect 4000 1974 4034 2009
rect 4000 1920 4034 1940
rect 1468 1886 1492 1920
rect 1526 1886 1562 1920
rect 1596 1886 1632 1920
rect 1666 1886 1702 1920
rect 1736 1886 1772 1920
rect 1806 1886 1842 1920
rect 1876 1886 1912 1920
rect 1946 1886 1982 1920
rect 2016 1886 2052 1920
rect 2086 1886 2122 1920
rect 2156 1886 2192 1920
rect 2226 1886 2262 1920
rect 2296 1886 2332 1920
rect 2366 1886 2402 1920
rect 2436 1886 2472 1920
rect 2506 1886 2542 1920
rect 2576 1886 2611 1920
rect 2645 1886 2680 1920
rect 2714 1886 2749 1920
rect 2783 1886 2818 1920
rect 2852 1886 2887 1920
rect 2921 1886 2956 1920
rect 2990 1886 3025 1920
rect 3059 1886 3094 1920
rect 3128 1886 3163 1920
rect 3197 1886 3232 1920
rect 3266 1886 3301 1920
rect 3335 1886 3370 1920
rect 3404 1886 3439 1920
rect 3473 1886 3508 1920
rect 3542 1904 4034 1920
rect 3542 1896 4000 1904
rect 3542 1886 3709 1896
rect 3646 1862 3709 1886
rect 3743 1862 3777 1896
rect 3811 1862 3845 1896
rect 3879 1862 3913 1896
rect 3947 1870 4000 1896
rect 3947 1862 4034 1870
rect 3646 1852 4034 1862
rect 3612 1834 4034 1852
rect 5276 2043 5872 2072
rect 5310 2037 5838 2043
rect 5310 2009 5359 2037
rect 5276 2003 5359 2009
rect 5393 2003 5427 2037
rect 5461 2003 5495 2037
rect 5529 2003 5563 2037
rect 5597 2003 5631 2037
rect 5665 2003 5699 2037
rect 5733 2003 5767 2037
rect 5801 2009 5838 2037
rect 5801 2003 5872 2009
rect 5276 1974 5872 2003
rect 5310 1968 5838 1974
rect 5310 1940 5359 1968
rect 5276 1934 5359 1940
rect 5393 1934 5427 1968
rect 5461 1934 5495 1968
rect 5529 1934 5563 1968
rect 5597 1934 5631 1968
rect 5665 1934 5699 1968
rect 5733 1934 5767 1968
rect 5801 1940 5838 1968
rect 5801 1934 5872 1940
rect 5276 1905 5872 1934
rect 5310 1899 5838 1905
rect 5310 1871 5359 1899
rect 5276 1865 5359 1871
rect 5393 1865 5427 1899
rect 5461 1865 5495 1899
rect 5529 1865 5563 1899
rect 5597 1865 5631 1899
rect 5665 1865 5699 1899
rect 5733 1865 5767 1899
rect 5801 1871 5838 1899
rect 5801 1865 5872 1871
rect 3612 1827 4000 1834
rect 3612 1816 3709 1827
rect 3646 1793 3709 1816
rect 3743 1793 3777 1827
rect 3811 1793 3845 1827
rect 3879 1793 3913 1827
rect 3947 1800 4000 1827
rect 3947 1793 4034 1800
rect 3646 1782 4034 1793
rect 5276 1836 5872 1865
rect 7114 2043 7148 2078
rect 7114 1974 7148 2009
rect 7114 1920 7148 1940
rect 7114 1904 7606 1920
rect 7148 1896 7606 1904
rect 7148 1870 7207 1896
rect 7114 1862 7207 1870
rect 7241 1862 7275 1896
rect 7309 1862 7343 1896
rect 7377 1862 7411 1896
rect 7445 1886 7606 1896
rect 7640 1886 7675 1920
rect 7709 1886 7744 1920
rect 7778 1886 7813 1920
rect 7847 1886 7882 1920
rect 7916 1886 7951 1920
rect 7985 1886 8020 1920
rect 8054 1886 8089 1920
rect 8123 1886 8158 1920
rect 8192 1886 8227 1920
rect 8261 1886 8296 1920
rect 8330 1886 8365 1920
rect 8399 1886 8434 1920
rect 8468 1886 8503 1920
rect 8537 1886 8572 1920
rect 8606 1886 8642 1920
rect 8676 1886 8712 1920
rect 8746 1886 8782 1920
rect 8816 1886 8852 1920
rect 8886 1886 8922 1920
rect 8956 1886 8992 1920
rect 9026 1886 9062 1920
rect 9096 1886 9132 1920
rect 9166 1886 9202 1920
rect 9236 1886 9272 1920
rect 9306 1886 9342 1920
rect 9376 1886 9412 1920
rect 9446 1886 9482 1920
rect 9516 1886 9552 1920
rect 9586 1886 9622 1920
rect 9656 1886 9680 1920
rect 7445 1862 7502 1886
rect 7114 1852 7502 1862
rect 5310 1830 5838 1836
rect 5310 1802 5359 1830
rect 5276 1796 5359 1802
rect 5393 1796 5427 1830
rect 5461 1796 5495 1830
rect 5529 1796 5563 1830
rect 5597 1796 5631 1830
rect 5665 1796 5699 1830
rect 5733 1796 5767 1830
rect 5801 1802 5838 1830
rect 5801 1796 5872 1802
rect 3612 1764 4034 1782
rect 3612 1758 4000 1764
rect 3612 1746 3709 1758
rect 3646 1724 3709 1746
rect 3743 1724 3777 1758
rect 3811 1724 3845 1758
rect 3879 1724 3913 1758
rect 3947 1730 4000 1758
rect 3947 1724 4034 1730
rect 3646 1712 4034 1724
rect 3612 1694 4034 1712
rect 3612 1689 4000 1694
rect 3612 1676 3709 1689
rect 3646 1655 3709 1676
rect 3743 1655 3777 1689
rect 3811 1655 3845 1689
rect 3879 1655 3913 1689
rect 3947 1660 4000 1689
rect 3947 1655 4034 1660
rect 3646 1642 4034 1655
rect 3612 1624 4034 1642
rect 3612 1620 4000 1624
rect 3612 1606 3709 1620
rect 3646 1586 3709 1606
rect 3743 1586 3777 1620
rect 3811 1586 3845 1620
rect 3879 1586 3913 1620
rect 3947 1590 4000 1620
rect 3947 1586 4034 1590
rect 5276 1766 5872 1796
rect 7114 1834 7536 1852
rect 7148 1827 7536 1834
rect 7148 1800 7207 1827
rect 7114 1793 7207 1800
rect 7241 1793 7275 1827
rect 7309 1793 7343 1827
rect 7377 1793 7411 1827
rect 7445 1816 7536 1827
rect 7445 1793 7502 1816
rect 5310 1761 5838 1766
rect 5310 1732 5359 1761
rect 5276 1727 5359 1732
rect 5393 1727 5427 1761
rect 5461 1727 5495 1761
rect 5529 1727 5563 1761
rect 5597 1727 5631 1761
rect 5665 1727 5699 1761
rect 5733 1727 5767 1761
rect 5801 1732 5838 1761
rect 5801 1727 5872 1732
rect 5276 1696 5872 1727
rect 5310 1692 5838 1696
rect 5310 1662 5359 1692
rect 5276 1658 5359 1662
rect 5393 1658 5427 1692
rect 5461 1658 5495 1692
rect 5529 1658 5563 1692
rect 5597 1658 5631 1692
rect 5665 1658 5699 1692
rect 5733 1658 5767 1692
rect 5801 1662 5838 1692
rect 5801 1658 5872 1662
rect 5276 1626 5872 1658
rect 5310 1623 5838 1626
rect 5310 1592 5359 1623
rect 5276 1589 5359 1592
rect 5393 1589 5427 1623
rect 5461 1589 5495 1623
rect 5529 1589 5563 1623
rect 5597 1589 5631 1623
rect 5665 1589 5699 1623
rect 5733 1589 5767 1623
rect 5801 1592 5838 1623
rect 5801 1589 5872 1592
rect 7114 1782 7502 1793
rect 7114 1764 7536 1782
rect 7148 1758 7536 1764
rect 7148 1730 7207 1758
rect 7114 1724 7207 1730
rect 7241 1724 7275 1758
rect 7309 1724 7343 1758
rect 7377 1724 7411 1758
rect 7445 1746 7536 1758
rect 7445 1724 7502 1746
rect 7114 1712 7502 1724
rect 7114 1694 7536 1712
rect 7148 1689 7536 1694
rect 7148 1660 7207 1689
rect 7114 1655 7207 1660
rect 7241 1655 7275 1689
rect 7309 1655 7343 1689
rect 7377 1655 7411 1689
rect 7445 1676 7536 1689
rect 7445 1655 7502 1676
rect 7114 1642 7502 1655
rect 7114 1624 7536 1642
rect 7148 1620 7536 1624
rect 7148 1590 7207 1620
rect 3646 1572 4034 1586
rect 3612 1554 4034 1572
rect 3612 1551 4000 1554
rect 3612 1536 3709 1551
rect 3646 1517 3709 1536
rect 3743 1517 3777 1551
rect 3811 1517 3845 1551
rect 3879 1517 3913 1551
rect 3947 1520 4000 1551
rect 5276 1556 5872 1589
rect 3947 1517 4034 1520
rect 3646 1502 4034 1517
rect 3612 1484 4034 1502
rect 3612 1482 4000 1484
rect 3612 1466 3709 1482
rect 3646 1448 3709 1466
rect 3743 1448 3777 1482
rect 3811 1448 3845 1482
rect 3879 1448 3913 1482
rect 3947 1450 4000 1482
rect 3947 1448 4034 1450
rect 3646 1432 4034 1448
rect 3612 1414 4034 1432
rect 3612 1413 4000 1414
rect 3612 1396 3709 1413
rect 3646 1379 3709 1396
rect 3743 1379 3777 1413
rect 3811 1379 3845 1413
rect 3879 1379 3913 1413
rect 3947 1380 4000 1413
rect 3947 1379 4034 1380
rect 3646 1362 4034 1379
rect 3612 1344 4034 1362
rect 3612 1326 3709 1344
rect 3646 1310 3709 1326
rect 3743 1310 3777 1344
rect 3811 1310 3845 1344
rect 3879 1310 3913 1344
rect 3947 1310 4000 1344
rect 5310 1554 5838 1556
rect 5310 1522 5359 1554
rect 5276 1520 5359 1522
rect 5393 1520 5427 1554
rect 5461 1520 5495 1554
rect 5529 1520 5563 1554
rect 5597 1520 5631 1554
rect 5665 1520 5699 1554
rect 5733 1520 5767 1554
rect 5801 1522 5838 1554
rect 7114 1586 7207 1590
rect 7241 1586 7275 1620
rect 7309 1586 7343 1620
rect 7377 1586 7411 1620
rect 7445 1606 7536 1620
rect 7445 1586 7502 1606
rect 7114 1572 7502 1586
rect 7114 1554 7536 1572
rect 5801 1520 5872 1522
rect 5276 1486 5872 1520
rect 5310 1485 5838 1486
rect 5310 1452 5359 1485
rect 5276 1451 5359 1452
rect 5393 1451 5427 1485
rect 5461 1451 5495 1485
rect 5529 1451 5563 1485
rect 5597 1451 5631 1485
rect 5665 1451 5699 1485
rect 5733 1451 5767 1485
rect 5801 1452 5838 1485
rect 5801 1451 5872 1452
rect 5276 1416 5872 1451
rect 5310 1382 5359 1416
rect 5393 1382 5427 1416
rect 5461 1382 5495 1416
rect 5529 1382 5563 1416
rect 5597 1382 5631 1416
rect 5665 1382 5699 1416
rect 5733 1382 5767 1416
rect 5801 1382 5838 1416
rect 5276 1346 5872 1382
rect 3646 1292 4034 1310
rect 3612 1274 4034 1292
rect 5310 1312 5359 1346
rect 5393 1312 5427 1346
rect 5461 1312 5495 1346
rect 5529 1312 5563 1346
rect 5597 1312 5631 1346
rect 5665 1312 5699 1346
rect 5733 1312 5767 1346
rect 5801 1312 5838 1346
rect 7148 1551 7536 1554
rect 7148 1520 7207 1551
rect 7114 1517 7207 1520
rect 7241 1517 7275 1551
rect 7309 1517 7343 1551
rect 7377 1517 7411 1551
rect 7445 1536 7536 1551
rect 7445 1517 7502 1536
rect 7114 1502 7502 1517
rect 7114 1484 7536 1502
rect 7148 1482 7536 1484
rect 7148 1450 7207 1482
rect 7114 1448 7207 1450
rect 7241 1448 7275 1482
rect 7309 1448 7343 1482
rect 7377 1448 7411 1482
rect 7445 1466 7536 1482
rect 7445 1448 7502 1466
rect 7114 1432 7502 1448
rect 7114 1414 7536 1432
rect 7148 1413 7536 1414
rect 7148 1380 7207 1413
rect 7114 1379 7207 1380
rect 7241 1379 7275 1413
rect 7309 1379 7343 1413
rect 7377 1379 7411 1413
rect 7445 1396 7536 1413
rect 7445 1379 7502 1396
rect 7114 1362 7502 1379
rect 7114 1344 7536 1362
rect 3612 1257 3709 1274
rect 3646 1240 3709 1257
rect 3743 1240 3777 1274
rect 3811 1240 3845 1274
rect 3879 1240 3913 1274
rect 3947 1240 4000 1274
rect 3646 1223 4034 1240
rect 3612 1204 4034 1223
rect 3612 1188 3709 1204
rect 3646 1170 3709 1188
rect 3743 1170 3777 1204
rect 3811 1170 3845 1204
rect 3879 1170 3913 1204
rect 3947 1170 4000 1204
rect 3646 1154 4034 1170
rect 3612 1134 4034 1154
rect 3612 1119 3709 1134
rect 3646 1100 3709 1119
rect 3743 1100 3777 1134
rect 3811 1100 3845 1134
rect 3879 1100 3913 1134
rect 3947 1100 4000 1134
rect 3646 1085 4034 1100
rect 3612 1064 4034 1085
rect 5276 1276 5872 1312
rect 7148 1310 7207 1344
rect 7241 1310 7275 1344
rect 7309 1310 7343 1344
rect 7377 1310 7411 1344
rect 7445 1326 7536 1344
rect 7445 1310 7502 1326
rect 7114 1292 7502 1310
rect 5310 1242 5359 1276
rect 5393 1242 5427 1276
rect 5461 1242 5495 1276
rect 5529 1242 5563 1276
rect 5597 1242 5631 1276
rect 5665 1242 5699 1276
rect 5733 1242 5767 1276
rect 5801 1242 5838 1276
rect 5276 1206 5872 1242
rect 5310 1172 5359 1206
rect 5393 1172 5427 1206
rect 5461 1172 5495 1206
rect 5529 1172 5563 1206
rect 5597 1172 5631 1206
rect 5665 1172 5699 1206
rect 5733 1172 5767 1206
rect 5801 1172 5838 1206
rect 5276 1136 5872 1172
rect 5310 1102 5359 1136
rect 5393 1102 5427 1136
rect 5461 1102 5495 1136
rect 5529 1102 5563 1136
rect 5597 1102 5631 1136
rect 5665 1102 5699 1136
rect 5733 1102 5767 1136
rect 5801 1102 5838 1136
rect 3612 1050 3709 1064
rect 3646 1030 3709 1050
rect 3743 1030 3777 1064
rect 3811 1030 3845 1064
rect 3879 1030 3913 1064
rect 3947 1030 4000 1064
rect 3646 1016 4034 1030
rect 5276 1066 5872 1102
rect 7114 1274 7536 1292
rect 7148 1240 7207 1274
rect 7241 1240 7275 1274
rect 7309 1240 7343 1274
rect 7377 1240 7411 1274
rect 7445 1257 7536 1274
rect 7445 1240 7502 1257
rect 7114 1223 7502 1240
rect 7114 1204 7536 1223
rect 7148 1170 7207 1204
rect 7241 1170 7275 1204
rect 7309 1170 7343 1204
rect 7377 1170 7411 1204
rect 7445 1188 7536 1204
rect 7445 1170 7502 1188
rect 7114 1154 7502 1170
rect 7114 1134 7536 1154
rect 7148 1100 7207 1134
rect 7241 1100 7275 1134
rect 7309 1100 7343 1134
rect 7377 1100 7411 1134
rect 7445 1119 7536 1134
rect 7445 1100 7502 1119
rect 7114 1085 7502 1100
rect 5310 1032 5359 1066
rect 5393 1032 5427 1066
rect 5461 1032 5495 1066
rect 5529 1032 5563 1066
rect 5597 1032 5631 1066
rect 5665 1032 5699 1066
rect 5733 1032 5767 1066
rect 5801 1032 5838 1066
rect 3612 994 4034 1016
rect 3612 981 3709 994
rect 3646 960 3709 981
rect 3743 960 3777 994
rect 3811 960 3845 994
rect 3879 960 3913 994
rect 3947 960 4000 994
rect 3646 947 4034 960
rect 3612 924 4034 947
rect 3612 912 3709 924
rect 3646 890 3709 912
rect 3743 890 3777 924
rect 3811 890 3845 924
rect 3879 890 3913 924
rect 3947 890 4000 924
rect 3646 878 4034 890
rect 5276 996 5872 1032
rect 7114 1064 7536 1085
rect 7148 1030 7207 1064
rect 7241 1030 7275 1064
rect 7309 1030 7343 1064
rect 7377 1030 7411 1064
rect 7445 1050 7536 1064
rect 7445 1030 7502 1050
rect 5310 962 5359 996
rect 5393 962 5427 996
rect 5461 962 5495 996
rect 5529 962 5563 996
rect 5597 962 5631 996
rect 5665 962 5699 996
rect 5733 962 5767 996
rect 5801 962 5838 996
rect 5276 926 5872 962
rect 5310 892 5359 926
rect 5393 892 5427 926
rect 5461 892 5495 926
rect 5529 892 5563 926
rect 5597 892 5631 926
rect 5665 892 5699 926
rect 5733 892 5767 926
rect 5801 892 5838 926
rect 3612 854 4034 878
rect 3612 843 3709 854
rect 3646 820 3709 843
rect 3743 820 3777 854
rect 3811 820 3845 854
rect 3879 820 3913 854
rect 3947 820 4000 854
rect 3646 809 4034 820
rect 3612 784 4034 809
rect 3612 774 3709 784
rect 3646 750 3709 774
rect 3743 750 3777 784
rect 3811 750 3845 784
rect 3879 750 3913 784
rect 3947 750 4000 784
rect 5276 856 5872 892
rect 7114 1016 7502 1030
rect 7114 994 7536 1016
rect 7148 960 7207 994
rect 7241 960 7275 994
rect 7309 960 7343 994
rect 7377 960 7411 994
rect 7445 981 7536 994
rect 7445 960 7502 981
rect 7114 947 7502 960
rect 7114 924 7536 947
rect 7148 890 7207 924
rect 7241 890 7275 924
rect 7309 890 7343 924
rect 7377 890 7411 924
rect 7445 912 7536 924
rect 7445 890 7502 912
rect 5310 822 5359 856
rect 5393 822 5427 856
rect 5461 822 5495 856
rect 5529 822 5563 856
rect 5597 822 5631 856
rect 5665 822 5699 856
rect 5733 822 5767 856
rect 5801 822 5838 856
rect 5276 786 5872 822
rect 3646 740 4034 750
rect 3612 714 4034 740
rect 3612 705 3709 714
rect 3646 680 3709 705
rect 3743 680 3777 714
rect 3811 680 3845 714
rect 3879 680 3913 714
rect 3947 680 4000 714
rect 3646 671 4034 680
rect 3612 644 4034 671
rect 3612 636 3709 644
rect 3646 610 3709 636
rect 3743 610 3777 644
rect 3811 610 3845 644
rect 3879 610 3913 644
rect 3947 610 4000 644
rect 3646 602 4034 610
rect 3612 574 4034 602
rect 3612 540 3709 574
rect 3743 540 3777 574
rect 3811 540 3845 574
rect 3879 540 3913 574
rect 3947 540 4000 574
rect 3612 504 4034 540
rect 1530 446 1554 480
rect 1588 446 1623 480
rect 1657 446 1692 480
rect 1726 446 1761 480
rect 1795 446 1830 480
rect 1864 446 1899 480
rect 1933 446 1968 480
rect 2002 446 2038 480
rect 2072 446 2108 480
rect 2142 446 2178 480
rect 2212 446 2248 480
rect 2282 446 2318 480
rect 2352 446 2388 480
rect 2422 446 2458 480
rect 2492 446 2528 480
rect 2562 446 2598 480
rect 2632 446 2668 480
rect 2702 446 2738 480
rect 2772 446 2808 480
rect 2842 446 2878 480
rect 2912 446 2948 480
rect 2982 446 3018 480
rect 3052 446 3088 480
rect 3122 446 3158 480
rect 3192 446 3228 480
rect 3262 446 3298 480
rect 3332 446 3368 480
rect 3402 446 3438 480
rect 3472 446 3508 480
rect 3542 446 3578 480
rect 3612 470 3709 504
rect 3743 470 3777 504
rect 3811 470 3845 504
rect 3879 470 3913 504
rect 3947 470 4000 504
rect 5310 752 5359 786
rect 5393 752 5427 786
rect 5461 752 5495 786
rect 5529 752 5563 786
rect 5597 752 5631 786
rect 5665 752 5699 786
rect 5733 752 5767 786
rect 5801 752 5838 786
rect 7114 878 7502 890
rect 7114 854 7536 878
rect 7148 820 7207 854
rect 7241 820 7275 854
rect 7309 820 7343 854
rect 7377 820 7411 854
rect 7445 843 7536 854
rect 7445 820 7502 843
rect 7114 809 7502 820
rect 7114 784 7536 809
rect 5276 716 5872 752
rect 5310 682 5359 716
rect 5393 682 5427 716
rect 5461 682 5495 716
rect 5529 682 5563 716
rect 5597 682 5631 716
rect 5665 682 5699 716
rect 5733 682 5767 716
rect 5801 682 5838 716
rect 5276 646 5872 682
rect 5310 612 5359 646
rect 5393 612 5427 646
rect 5461 612 5495 646
rect 5529 612 5563 646
rect 5597 612 5631 646
rect 5665 612 5699 646
rect 5733 612 5767 646
rect 5801 612 5838 646
rect 5276 576 5872 612
rect 5310 542 5359 576
rect 5393 542 5427 576
rect 5461 542 5495 576
rect 5529 542 5563 576
rect 5597 542 5631 576
rect 5665 542 5699 576
rect 5733 542 5767 576
rect 5801 542 5838 576
rect 5276 506 5872 542
rect 3612 446 4034 470
rect 5310 472 5359 506
rect 5393 472 5427 506
rect 5461 472 5495 506
rect 5529 472 5563 506
rect 5597 472 5631 506
rect 5665 472 5699 506
rect 5733 472 5767 506
rect 5801 472 5838 506
rect 7148 750 7207 784
rect 7241 750 7275 784
rect 7309 750 7343 784
rect 7377 750 7411 784
rect 7445 774 7536 784
rect 7445 750 7502 774
rect 7114 740 7502 750
rect 7114 714 7536 740
rect 7148 680 7207 714
rect 7241 680 7275 714
rect 7309 680 7343 714
rect 7377 680 7411 714
rect 7445 705 7536 714
rect 7445 680 7502 705
rect 7114 671 7502 680
rect 7114 644 7536 671
rect 7148 610 7207 644
rect 7241 610 7275 644
rect 7309 610 7343 644
rect 7377 610 7411 644
rect 7445 636 7536 644
rect 7445 610 7502 636
rect 7114 602 7502 610
rect 7114 574 7536 602
rect 7148 540 7207 574
rect 7241 540 7275 574
rect 7309 540 7343 574
rect 7377 540 7411 574
rect 7445 540 7536 574
rect 7114 504 7536 540
rect 5276 448 5872 472
rect 7148 470 7207 504
rect 7241 470 7275 504
rect 7309 470 7343 504
rect 7377 470 7411 504
rect 7445 470 7536 504
rect 7114 446 7536 470
rect 7570 446 7606 480
rect 7640 446 7676 480
rect 7710 446 7746 480
rect 7780 446 7816 480
rect 7850 446 7886 480
rect 7920 446 7956 480
rect 7990 446 8026 480
rect 8060 446 8096 480
rect 8130 446 8166 480
rect 8200 446 8236 480
rect 8270 446 8306 480
rect 8340 446 8376 480
rect 8410 446 8446 480
rect 8480 446 8516 480
rect 8550 446 8586 480
rect 8620 446 8656 480
rect 8690 446 8726 480
rect 8760 446 8796 480
rect 8830 446 8866 480
rect 8900 446 8936 480
rect 8970 446 9006 480
rect 9040 446 9076 480
rect 9110 446 9146 480
rect 9180 446 9215 480
rect 9249 446 9284 480
rect 9318 446 9353 480
rect 9387 446 9422 480
rect 9456 446 9491 480
rect 9525 446 9560 480
rect 9594 446 9618 480
rect 10212 7671 10283 7705
rect 10317 7671 10351 7705
rect 10385 7671 10419 7705
rect 10453 7671 10487 7705
rect 10521 7671 10555 7705
rect 10589 7671 10623 7705
rect 10657 7671 10691 7705
rect 10725 7671 10759 7705
rect 10793 7671 10827 7705
rect 10861 7671 10895 7705
rect 10929 7671 10963 7705
rect 10997 7671 11031 7705
rect 11065 7671 11099 7705
rect 11133 7671 11167 7705
rect 11201 7671 11235 7705
rect 11269 7671 11303 7705
rect 11337 7671 11371 7705
rect 11405 7671 11439 7705
rect 11473 7671 11507 7705
rect 11541 7671 11575 7705
rect 11609 7671 11643 7705
rect 11677 7671 11711 7705
rect 11745 7671 11779 7705
rect 11813 7671 11847 7705
rect 11881 7671 11915 7705
rect 11949 7671 11983 7705
rect 12017 7671 12051 7705
rect 12085 7671 12119 7705
rect 12153 7671 12187 7705
rect 12221 7671 12255 7705
rect 12289 7671 12323 7705
rect 12357 7671 12391 7705
rect 12425 7671 12459 7705
rect 12493 7671 12527 7705
rect 12561 7671 12595 7705
rect 12629 7671 12663 7705
rect 12697 7671 12731 7705
rect 12765 7671 12799 7705
rect 10212 7603 10246 7637
rect 10212 7535 10246 7569
rect 10212 7467 10246 7501
rect 10212 7399 10246 7433
rect 10212 7331 10246 7365
rect 10212 7263 10246 7297
rect 10212 7195 10246 7229
rect 10212 7127 10246 7161
rect 10212 7059 10246 7093
rect 10212 6991 10246 7025
rect 10212 6923 10246 6957
rect 10212 6855 10246 6889
rect 10212 6787 10246 6821
rect 10212 6719 10246 6753
rect 10212 6651 10246 6685
rect 10212 6583 10246 6617
rect 10212 6515 10246 6549
rect 10212 6447 10246 6481
rect 10212 6379 10246 6413
rect 10212 6311 10246 6345
rect 10212 6243 10246 6277
rect 10212 6175 10246 6209
rect 10212 6107 10246 6141
rect 10212 6039 10246 6073
rect 10212 5971 10246 6005
rect 10212 5903 10246 5937
rect 10212 5835 10246 5869
rect 10212 5767 10246 5801
rect 10212 5699 10246 5733
rect 10212 5631 10246 5665
rect 10212 5563 10246 5597
rect 10212 5495 10246 5529
rect 10212 5427 10246 5461
rect 10212 5359 10246 5393
rect 10212 5291 10246 5325
rect 10212 5223 10246 5257
rect 10212 5155 10246 5189
rect 10212 5087 10246 5121
rect 10212 5019 10246 5053
rect 10212 4951 10246 4985
rect 10212 4883 10246 4917
rect 10212 4815 10246 4849
rect 10212 4747 10246 4781
rect 10212 4679 10246 4713
rect 10212 4611 10246 4645
rect 10212 4543 10246 4577
rect 10212 4475 10246 4509
rect 10212 4407 10246 4441
rect 10212 4339 10246 4373
rect 10212 4271 10246 4305
rect 10212 4203 10246 4237
rect 10212 4135 10246 4169
rect 10212 4067 10246 4101
rect 10212 3999 10246 4033
rect 10212 3931 10246 3965
rect 10212 3863 10246 3897
rect 10212 3795 10246 3829
rect 10212 3727 10246 3761
rect 10212 3659 10246 3693
rect 10212 3591 10246 3625
rect 10212 3523 10246 3557
rect 10212 3455 10246 3489
rect 10212 3387 10246 3421
rect 10212 3319 10246 3353
rect 10212 3251 10246 3285
rect 10212 3183 10246 3217
rect 10212 3115 10246 3149
rect 10212 3047 10246 3081
rect 10212 2979 10246 3013
rect 10212 2911 10246 2945
rect 10212 2843 10246 2877
rect 10212 2775 10246 2809
rect 10212 2707 10246 2741
rect 10212 2639 10246 2673
rect 10212 2571 10246 2605
rect 10212 2503 10246 2537
rect 10212 2435 10246 2469
rect 10212 2367 10246 2401
rect 10212 2299 10246 2333
rect 10212 2231 10246 2265
rect 10212 2163 10246 2197
rect 10212 2095 10246 2129
rect 10212 2027 10246 2061
rect 10212 1959 10246 1993
rect 10212 1891 10246 1925
rect 10212 1823 10246 1857
rect 10212 1755 10246 1789
rect 10212 1687 10246 1721
rect 10212 1619 10246 1653
rect 10212 1551 10246 1585
rect 10212 1483 10246 1517
rect 10212 1415 10246 1449
rect 10212 1347 10246 1381
rect 10212 1279 10246 1313
rect 10212 1211 10246 1245
rect 10212 1143 10246 1177
rect 10212 1075 10246 1109
rect 10212 1007 10246 1041
rect 10212 939 10246 973
rect 10212 871 10246 905
rect 10212 803 10246 837
rect 10212 735 10246 769
rect 10212 667 10246 701
rect 10212 599 10246 633
rect 10212 446 10246 565
rect 10280 446 10314 480
rect 10348 446 10382 480
rect 10416 446 10450 480
rect 10484 446 10518 480
rect 10552 446 10586 480
rect 10620 446 10690 480
rect 10724 446 10758 480
rect 10792 446 10826 480
rect 10860 446 10894 480
rect 10928 446 10962 480
rect 10996 446 11030 480
rect 11064 446 11098 480
rect 11132 446 11166 480
rect 11200 446 11234 480
rect 11268 446 11302 480
rect 11336 446 11370 480
rect 11404 446 11438 480
rect 11472 446 11506 480
rect 11540 446 11574 480
rect 11608 446 11642 480
rect 11676 446 11710 480
rect 11744 446 11778 480
rect 11812 446 11846 480
rect 11880 446 11914 480
rect 11948 446 11982 480
rect 12016 446 12050 480
rect 12084 446 12118 480
rect 12152 446 12186 480
rect 12220 446 12254 480
rect 12288 446 12322 480
rect 12356 446 12390 480
rect 12424 446 12458 480
rect 12492 446 12526 480
rect 12560 446 12594 480
rect 12628 446 12662 480
rect 12696 446 12730 480
rect 12764 446 12799 480
<< mvnsubdiff >>
rect 1197 14200 1231 14234
rect 1265 14200 1299 14234
rect 1333 14200 1367 14234
rect 1401 14200 1435 14234
rect 1469 14200 1503 14234
rect 1537 14200 1571 14234
rect 1605 14200 1639 14234
rect 1673 14200 1707 14234
rect 1741 14200 1775 14234
rect 1809 14200 1843 14234
rect 1877 14200 1911 14234
rect 1945 14200 1979 14234
rect 2013 14200 2047 14234
rect 2081 14200 2115 14234
rect 2149 14200 2183 14234
rect 2217 14200 2251 14234
rect 2285 14200 2319 14234
rect 2353 14200 2387 14234
rect 2421 14200 2455 14234
rect 2489 14200 2523 14234
rect 2557 14200 2591 14234
rect 2625 14200 2659 14234
rect 2693 14200 2727 14234
rect 2761 14200 2795 14234
rect 2829 14200 2863 14234
rect 2897 14200 2931 14234
rect 2965 14200 2999 14234
rect 3033 14200 3067 14234
rect 3101 14200 3135 14234
rect 3169 14200 3203 14234
rect 3237 14200 3271 14234
rect 3305 14200 3339 14234
rect 3373 14200 3407 14234
rect 3441 14200 3475 14234
rect 3509 14200 3543 14234
rect 3577 14200 3611 14234
rect 3645 14200 3679 14234
rect 3713 14200 3747 14234
rect 3781 14200 3815 14234
rect 3849 14200 3883 14234
rect 3917 14200 3951 14234
rect 3985 14200 4019 14234
rect 4053 14200 4087 14234
rect 4121 14200 4155 14234
rect 4189 14200 4223 14234
rect 4257 14200 4291 14234
rect 4325 14200 4359 14234
rect 4393 14200 4427 14234
rect 4461 14200 4495 14234
rect 4529 14200 4563 14234
rect 4597 14200 4631 14234
rect 4665 14200 4699 14234
rect 4733 14200 4767 14234
rect 4801 14200 4835 14234
rect 4869 14200 4903 14234
rect 4937 14200 4971 14234
rect 5005 14200 5039 14234
rect 5073 14200 5107 14234
rect 5141 14200 5175 14234
rect 5209 14200 5243 14234
rect 5277 14200 5311 14234
rect 5345 14200 5379 14234
rect 5413 14200 5447 14234
rect 5481 14200 5515 14234
rect 5549 14200 5583 14234
rect 5617 14200 5651 14234
rect 5685 14200 5719 14234
rect 5753 14200 5787 14234
rect 5821 14200 5855 14234
rect 5889 14200 5923 14234
rect 5957 14200 5991 14234
rect 6025 14200 6059 14234
rect 6093 14200 6127 14234
rect 6161 14200 6195 14234
rect 6229 14200 6263 14234
rect 6297 14200 6331 14234
rect 6365 14200 6399 14234
rect 6433 14200 6467 14234
rect 6501 14200 6535 14234
rect 6569 14200 6603 14234
rect 6637 14200 6671 14234
rect 6705 14200 6739 14234
rect 6773 14200 6807 14234
rect 6841 14200 6875 14234
rect 6909 14200 6943 14234
rect 6977 14200 7011 14234
rect 7045 14200 7079 14234
rect 7113 14200 7147 14234
rect 7181 14200 7215 14234
rect 7249 14200 7283 14234
rect 7317 14200 7351 14234
rect 7385 14200 7419 14234
rect 7453 14200 7487 14234
rect 7521 14200 7555 14234
rect 7589 14200 7623 14234
rect 7657 14200 7691 14234
rect 7725 14200 7759 14234
rect 7793 14200 7827 14234
rect 7861 14200 7895 14234
rect 7929 14200 7963 14234
rect 7997 14200 8031 14234
rect 8065 14200 8099 14234
rect 8133 14200 8167 14234
rect 8201 14200 8235 14234
rect 8269 14200 8303 14234
rect 8337 14200 8371 14234
rect 8405 14200 8439 14234
rect 8473 14200 8507 14234
rect 8541 14200 8575 14234
rect 8609 14200 8643 14234
rect 8677 14200 8711 14234
rect 8745 14200 8779 14234
rect 8813 14200 8847 14234
rect 8881 14200 8915 14234
rect 8949 14200 8983 14234
rect 9017 14200 9051 14234
rect 9085 14200 9119 14234
rect 9153 14200 9187 14234
rect 9221 14200 9255 14234
rect 9289 14200 9323 14234
rect 9357 14200 9391 14234
rect 9425 14200 9459 14234
rect 9493 14200 9527 14234
rect 9561 14200 9595 14234
rect 9629 14200 9663 14234
rect 9697 14200 9731 14234
rect 9765 14200 9799 14234
rect 9833 14200 9867 14234
rect 9901 14200 9935 14234
rect 9969 14200 10003 14234
rect 10037 14200 10071 14234
rect 10105 14200 10139 14234
rect 10173 14200 10207 14234
rect 10241 14200 10275 14234
rect 10309 14200 10343 14234
rect 10377 14200 10411 14234
rect 10445 14200 10479 14234
rect 10513 14200 10547 14234
rect 10581 14200 10615 14234
rect 10649 14200 10683 14234
rect 10717 14200 10751 14234
rect 10785 14200 10819 14234
rect 10853 14200 10887 14234
rect 10921 14200 10955 14234
rect 10989 14200 11111 14234
rect 1197 14166 1560 14200
rect 1197 14132 1371 14166
rect 1405 14132 1443 14166
rect 1477 14132 1515 14166
rect 1549 14132 1560 14166
rect 1197 14100 1560 14132
rect 1231 14094 1560 14100
rect 1231 14066 1371 14094
rect 1197 14060 1371 14066
rect 1405 14060 1443 14094
rect 1477 14060 1515 14094
rect 1549 14060 1560 14094
rect 5165 14155 5929 14200
rect 5165 14121 5189 14155
rect 5223 14121 5265 14155
rect 5299 14121 5341 14155
rect 5375 14121 5417 14155
rect 5451 14121 5493 14155
rect 5527 14121 5569 14155
rect 5603 14121 5645 14155
rect 5679 14121 5721 14155
rect 5755 14121 5796 14155
rect 5830 14121 5871 14155
rect 5905 14121 5929 14155
rect 1197 14032 1560 14060
rect 1231 14021 1560 14032
rect 1231 13998 1371 14021
rect 1197 13987 1371 13998
rect 1405 13987 1443 14021
rect 1477 13987 1515 14021
rect 1549 13987 1560 14021
rect 1197 13964 1560 13987
rect 1231 13948 1560 13964
rect 1231 13930 1371 13948
rect 1197 13914 1371 13930
rect 1405 13914 1443 13948
rect 1477 13914 1515 13948
rect 1549 13914 1560 13948
rect 1197 13896 1560 13914
rect 1231 13875 1560 13896
rect 1231 13862 1371 13875
rect 1197 13841 1371 13862
rect 1405 13841 1443 13875
rect 1477 13841 1515 13875
rect 1549 13841 1560 13875
rect 1197 13828 1560 13841
rect 1231 13802 1560 13828
rect 1231 13794 1371 13802
rect 1197 13768 1371 13794
rect 1405 13768 1443 13802
rect 1477 13768 1515 13802
rect 1549 13768 1560 13802
rect 1197 13760 1560 13768
rect 1231 13729 1560 13760
rect 1231 13726 1371 13729
rect 1197 13695 1371 13726
rect 1405 13695 1443 13729
rect 1477 13695 1515 13729
rect 1549 13695 1560 13729
rect 1197 13692 1560 13695
rect 1231 13658 1560 13692
rect 1197 13656 1560 13658
rect 1197 13624 1371 13656
rect 1231 13622 1371 13624
rect 1405 13622 1443 13656
rect 1477 13622 1515 13656
rect 1549 13622 1560 13656
rect 1231 13590 1560 13622
rect 1197 13583 1560 13590
rect 1197 13556 1371 13583
rect 1231 13549 1371 13556
rect 1405 13549 1443 13583
rect 1477 13549 1515 13583
rect 1549 13549 1560 13583
rect 1231 13522 1560 13549
rect 1197 13510 1560 13522
rect 1197 13488 1371 13510
rect 1231 13476 1371 13488
rect 1405 13476 1443 13510
rect 1477 13476 1515 13510
rect 1549 13476 1560 13510
rect 1231 13454 1560 13476
rect 1197 13437 1560 13454
rect 1197 13420 1371 13437
rect 1231 13403 1371 13420
rect 1405 13403 1443 13437
rect 1477 13403 1515 13437
rect 1549 13403 1560 13437
rect 1231 13386 1560 13403
rect 1197 13364 1560 13386
rect 1197 13352 1371 13364
rect 1231 13330 1371 13352
rect 1405 13330 1443 13364
rect 1477 13330 1515 13364
rect 1549 13330 1560 13364
rect 1231 13318 1560 13330
rect 1197 13291 1560 13318
rect 1197 13284 1371 13291
rect 1231 13257 1371 13284
rect 1405 13257 1443 13291
rect 1477 13257 1515 13291
rect 1549 13257 1560 13291
rect 1231 13250 1560 13257
rect 1197 13218 1560 13250
rect 1197 13216 1371 13218
rect 1231 13184 1371 13216
rect 1405 13184 1443 13218
rect 1477 13184 1515 13218
rect 1549 13184 1560 13218
rect 1231 13182 1560 13184
rect 1197 13160 1560 13182
rect 1197 13124 1231 13160
rect 1197 13054 1231 13090
rect 1197 12984 1231 13020
rect 1197 12914 1231 12950
rect 1197 12844 1231 12880
rect 1197 12774 1231 12810
rect 1197 12704 1231 12740
rect 1197 12633 1231 12670
rect 1197 12562 1231 12599
rect 1197 12491 1231 12528
rect 5165 14083 5929 14121
rect 9365 14153 9903 14200
rect 9365 14119 9399 14153
rect 9433 14119 9472 14153
rect 9506 14119 9545 14153
rect 9579 14119 9618 14153
rect 9652 14119 9691 14153
rect 9725 14119 9763 14153
rect 9797 14119 9835 14153
rect 9869 14119 9903 14153
rect 5165 14049 5189 14083
rect 5223 14049 5265 14083
rect 5299 14049 5341 14083
rect 5375 14049 5417 14083
rect 5451 14049 5493 14083
rect 5527 14049 5569 14083
rect 5603 14049 5645 14083
rect 5679 14049 5721 14083
rect 5755 14049 5796 14083
rect 5830 14049 5871 14083
rect 5905 14049 5929 14083
rect 5165 14011 5929 14049
rect 5165 13977 5189 14011
rect 5223 13977 5265 14011
rect 5299 13977 5341 14011
rect 5375 13977 5417 14011
rect 5451 13977 5493 14011
rect 5527 13977 5569 14011
rect 5603 13977 5645 14011
rect 5679 13977 5721 14011
rect 5755 13977 5796 14011
rect 5830 13977 5871 14011
rect 5905 13977 5929 14011
rect 5165 13966 5929 13977
rect 5165 12668 5384 12708
rect 5165 12634 5219 12668
rect 5253 12634 5287 12668
rect 5321 12634 5384 12668
rect 1197 12420 1231 12457
rect 5165 12569 5384 12634
rect 5165 12535 5219 12569
rect 5253 12535 5287 12569
rect 5321 12535 5384 12569
rect 5165 12469 5384 12535
rect 5710 12668 5929 12708
rect 5710 12634 5764 12668
rect 5798 12634 5832 12668
rect 5866 12634 5929 12668
rect 5710 12569 5929 12634
rect 5710 12535 5764 12569
rect 5798 12535 5832 12569
rect 5866 12535 5929 12569
rect 5165 12435 5219 12469
rect 5253 12435 5287 12469
rect 5321 12435 5384 12469
rect 5165 12386 5384 12435
rect 5710 12469 5929 12535
rect 5710 12435 5764 12469
rect 5798 12435 5832 12469
rect 5866 12435 5929 12469
rect 9365 14085 9903 14119
rect 9365 14051 9399 14085
rect 9433 14051 9472 14085
rect 9506 14051 9545 14085
rect 9579 14051 9618 14085
rect 9652 14051 9691 14085
rect 9725 14051 9763 14085
rect 9797 14051 9835 14085
rect 9869 14051 9903 14085
rect 9365 14012 9903 14051
rect 9365 13978 9495 14012
rect 9529 13978 9563 14012
rect 9597 13978 9631 14012
rect 9665 13978 9699 14012
rect 9733 13978 9767 14012
rect 9801 13978 9835 14012
rect 9365 13910 9399 13944
rect 9365 13842 9399 13876
rect 9869 13907 9903 14012
rect 9365 13774 9399 13808
rect 9365 13706 9399 13740
rect 9365 13638 9399 13672
rect 9365 13570 9399 13604
rect 9365 13502 9399 13536
rect 9365 13434 9399 13468
rect 9365 13366 9399 13400
rect 9365 13298 9399 13332
rect 9365 13230 9399 13264
rect 9365 13162 9399 13196
rect 9365 13094 9399 13128
rect 9365 13026 9399 13060
rect 9365 12958 9399 12992
rect 9365 12751 9399 12924
rect 9869 13839 9903 13873
rect 9869 13771 9903 13805
rect 9869 13703 9903 13737
rect 9869 13635 9903 13669
rect 9869 13567 9903 13601
rect 9869 13499 9903 13533
rect 9869 13431 9903 13465
rect 9869 13363 9903 13397
rect 9869 13295 9903 13329
rect 9869 13227 9903 13261
rect 9869 13159 9903 13193
rect 9869 13091 9903 13125
rect 9869 13023 9903 13057
rect 9869 12955 9903 12989
rect 9869 12887 9903 12921
rect 9869 12819 9903 12853
rect 9433 12751 9467 12785
rect 9501 12751 9535 12785
rect 9569 12751 9603 12785
rect 9637 12751 9671 12785
rect 9705 12751 9739 12785
rect 9773 12751 9903 12785
rect 9365 12690 9903 12751
rect 9365 12656 9419 12690
rect 9453 12656 9487 12690
rect 9521 12656 9747 12690
rect 9781 12656 9815 12690
rect 9849 12656 9903 12690
rect 9365 12617 9903 12656
rect 9365 12583 9419 12617
rect 9453 12583 9487 12617
rect 9521 12583 9747 12617
rect 9781 12583 9815 12617
rect 9849 12583 9903 12617
rect 9365 12543 9903 12583
rect 9365 12509 9419 12543
rect 9453 12509 9487 12543
rect 9521 12509 9747 12543
rect 9781 12509 9815 12543
rect 9849 12509 9903 12543
rect 9365 12469 9903 12509
rect 5710 12386 5929 12435
rect 9365 12435 9419 12469
rect 9453 12435 9487 12469
rect 9521 12435 9747 12469
rect 9781 12435 9815 12469
rect 9849 12435 9903 12469
rect 9365 12386 9903 12435
rect 11077 14132 11111 14166
rect 11077 14064 11111 14098
rect 11077 13996 11111 14030
rect 11077 13928 11111 13962
rect 11077 13860 11111 13894
rect 11077 13792 11111 13826
rect 11077 13724 11111 13758
rect 11077 13656 11111 13690
rect 11077 13588 11111 13622
rect 11077 13520 11111 13554
rect 11077 13452 11111 13486
rect 11077 13384 11111 13418
rect 11077 13316 11111 13350
rect 11077 13248 11111 13282
rect 11077 13120 11111 13214
rect 11077 13050 11111 13086
rect 11077 12980 11111 13016
rect 11077 12910 11111 12946
rect 11077 12840 11111 12876
rect 11077 12770 11111 12806
rect 11077 12700 11111 12736
rect 11077 12630 11111 12666
rect 11077 12560 11111 12596
rect 11077 12490 11111 12526
rect 11077 12420 11111 12456
rect 1197 12352 1299 12386
rect 1333 12352 1367 12386
rect 1401 12352 1435 12386
rect 1469 12352 1503 12386
rect 1537 12352 1571 12386
rect 1605 12352 1639 12386
rect 1673 12352 1707 12386
rect 1741 12352 1775 12386
rect 1809 12352 1843 12386
rect 1877 12352 1911 12386
rect 1945 12352 1979 12386
rect 2013 12352 2047 12386
rect 2081 12352 2115 12386
rect 2149 12352 2183 12386
rect 2217 12352 2251 12386
rect 2285 12352 2319 12386
rect 2353 12352 2387 12386
rect 2421 12352 2455 12386
rect 2489 12352 2523 12386
rect 2557 12352 2591 12386
rect 2625 12352 2659 12386
rect 2693 12352 2727 12386
rect 2761 12352 2795 12386
rect 2829 12352 2863 12386
rect 2897 12352 2931 12386
rect 2965 12352 2999 12386
rect 3033 12352 3067 12386
rect 3101 12352 3135 12386
rect 3169 12352 3203 12386
rect 3237 12352 3271 12386
rect 3305 12352 3339 12386
rect 3373 12352 3407 12386
rect 3441 12352 3475 12386
rect 3509 12352 3543 12386
rect 3577 12352 3611 12386
rect 3645 12352 3679 12386
rect 3713 12352 3747 12386
rect 3781 12352 3815 12386
rect 3849 12352 3883 12386
rect 3917 12352 3951 12386
rect 3985 12352 4019 12386
rect 4053 12352 4087 12386
rect 4121 12352 4155 12386
rect 4189 12352 4223 12386
rect 4257 12352 4291 12386
rect 4325 12352 4359 12386
rect 4393 12352 4427 12386
rect 4461 12352 4495 12386
rect 4529 12352 4563 12386
rect 4597 12352 4631 12386
rect 4665 12352 4699 12386
rect 4733 12352 4767 12386
rect 4801 12352 4835 12386
rect 4869 12352 4903 12386
rect 4937 12352 4971 12386
rect 5005 12352 5039 12386
rect 5073 12352 5107 12386
rect 5141 12352 5175 12386
rect 5209 12352 5243 12386
rect 5277 12352 5311 12386
rect 5345 12352 5379 12386
rect 5413 12352 5447 12386
rect 5481 12352 5515 12386
rect 5549 12352 5583 12386
rect 5617 12352 5651 12386
rect 5685 12352 5719 12386
rect 5753 12352 5787 12386
rect 5821 12352 5855 12386
rect 5889 12352 5923 12386
rect 5957 12352 5991 12386
rect 6025 12352 6059 12386
rect 6093 12352 6127 12386
rect 6161 12352 6195 12386
rect 6229 12352 6263 12386
rect 6297 12352 6331 12386
rect 6365 12352 6399 12386
rect 6433 12352 6467 12386
rect 6501 12352 6535 12386
rect 6569 12352 6603 12386
rect 6637 12352 6671 12386
rect 6705 12352 6739 12386
rect 6773 12352 6807 12386
rect 6841 12352 6875 12386
rect 6909 12352 6943 12386
rect 6977 12352 7011 12386
rect 7045 12352 7079 12386
rect 7113 12352 7147 12386
rect 7181 12352 7215 12386
rect 7249 12352 7283 12386
rect 7317 12352 7351 12386
rect 7385 12352 7419 12386
rect 7453 12352 7487 12386
rect 7521 12352 7555 12386
rect 7589 12352 7623 12386
rect 7657 12352 7691 12386
rect 7725 12352 7759 12386
rect 7793 12352 7827 12386
rect 7861 12352 7895 12386
rect 7929 12352 7963 12386
rect 7997 12352 8031 12386
rect 8065 12352 8099 12386
rect 8133 12352 8167 12386
rect 8201 12352 8235 12386
rect 8269 12352 8303 12386
rect 8337 12352 8371 12386
rect 8405 12352 8439 12386
rect 8473 12352 8507 12386
rect 8541 12352 8575 12386
rect 8609 12352 8643 12386
rect 8677 12352 8711 12386
rect 8745 12352 8779 12386
rect 8813 12352 8847 12386
rect 8881 12352 8915 12386
rect 8949 12352 8983 12386
rect 9017 12352 9052 12386
rect 9086 12352 9121 12386
rect 9155 12352 9190 12386
rect 9224 12352 9259 12386
rect 9293 12352 9328 12386
rect 9362 12352 9397 12386
rect 9431 12352 9466 12386
rect 9500 12352 9535 12386
rect 9569 12352 9604 12386
rect 9638 12352 9673 12386
rect 9707 12352 9742 12386
rect 9776 12352 9811 12386
rect 9845 12352 9880 12386
rect 9914 12352 9949 12386
rect 9983 12352 10018 12386
rect 10052 12352 10087 12386
rect 10121 12352 10156 12386
rect 10190 12352 10225 12386
rect 10259 12352 10294 12386
rect 10328 12352 10363 12386
rect 10397 12352 10432 12386
rect 10466 12352 10501 12386
rect 10535 12352 10583 12386
rect 10617 12352 10659 12386
rect 10693 12352 10735 12386
rect 10769 12352 10811 12386
rect 10845 12352 10886 12386
rect 10920 12352 10961 12386
rect 10995 12352 11111 12386
rect 1117 11699 1219 11723
rect 1151 11665 1219 11699
rect 1321 11689 1355 11723
rect 1389 11689 1423 11723
rect 1457 11689 1491 11723
rect 1525 11689 1559 11723
rect 1593 11689 1627 11723
rect 1661 11689 1695 11723
rect 1729 11689 1763 11723
rect 1797 11689 1831 11723
rect 1865 11689 1899 11723
rect 1933 11689 1967 11723
rect 2001 11689 2035 11723
rect 2069 11689 2103 11723
rect 2137 11689 2171 11723
rect 2205 11689 2239 11723
rect 2273 11689 2307 11723
rect 2341 11689 2375 11723
rect 2409 11689 2443 11723
rect 2477 11689 2511 11723
rect 2545 11689 2579 11723
rect 2613 11689 2647 11723
rect 2681 11689 2715 11723
rect 2749 11689 2841 11723
rect 2875 11689 2909 11723
rect 2943 11689 2977 11723
rect 3011 11689 3045 11723
rect 3079 11689 3113 11723
rect 3147 11689 3181 11723
rect 3215 11689 3249 11723
rect 3283 11689 3317 11723
rect 3351 11689 3385 11723
rect 3419 11689 3453 11723
rect 3487 11689 3521 11723
rect 3555 11689 3589 11723
rect 3623 11689 3657 11723
rect 3691 11689 3725 11723
rect 3759 11689 3793 11723
rect 3827 11689 3861 11723
rect 3895 11689 3929 11723
rect 3963 11689 3997 11723
rect 4031 11689 4065 11723
rect 4099 11689 4133 11723
rect 4167 11689 4201 11723
rect 4235 11689 4269 11723
rect 4303 11689 4337 11723
rect 4371 11689 4405 11723
rect 4439 11689 4473 11723
rect 4507 11689 4541 11723
rect 4575 11689 4609 11723
rect 4643 11689 4677 11723
rect 4711 11689 4745 11723
rect 4779 11689 4813 11723
rect 4847 11689 4881 11723
rect 4915 11689 4949 11723
rect 4983 11689 5017 11723
rect 5051 11689 5085 11723
rect 5119 11689 5153 11723
rect 5187 11689 5221 11723
rect 5255 11689 5289 11723
rect 5323 11689 5357 11723
rect 5391 11689 5425 11723
rect 5459 11689 5688 11723
rect 5722 11689 5756 11723
rect 5790 11689 5824 11723
rect 5858 11689 5892 11723
rect 5926 11689 5960 11723
rect 5994 11689 6028 11723
rect 6062 11689 6096 11723
rect 6130 11689 6164 11723
rect 6198 11689 6232 11723
rect 6266 11689 6300 11723
rect 6334 11689 6368 11723
rect 6402 11689 6436 11723
rect 6470 11689 6504 11723
rect 6538 11689 6572 11723
rect 6606 11689 6640 11723
rect 6674 11689 6708 11723
rect 6742 11689 6776 11723
rect 6810 11689 6844 11723
rect 6878 11689 6912 11723
rect 6946 11689 6980 11723
rect 7014 11689 7048 11723
rect 7082 11689 7116 11723
rect 7150 11689 7184 11723
rect 7218 11689 7252 11723
rect 7286 11689 7320 11723
rect 7354 11689 7388 11723
rect 7422 11689 7456 11723
rect 7490 11689 7524 11723
rect 7558 11689 7592 11723
rect 7626 11689 7660 11723
rect 7694 11689 7728 11723
rect 7762 11689 7796 11723
rect 7830 11689 7923 11723
rect 7957 11689 7991 11723
rect 8025 11689 8059 11723
rect 8093 11689 8127 11723
rect 8161 11689 8195 11723
rect 8229 11689 8263 11723
rect 8297 11689 8331 11723
rect 8365 11689 8399 11723
rect 8433 11689 8467 11723
rect 8501 11689 8535 11723
rect 8569 11689 8603 11723
rect 8637 11689 8671 11723
rect 8705 11689 8739 11723
rect 8773 11689 8807 11723
rect 8841 11689 8875 11723
rect 8909 11689 8943 11723
rect 8977 11689 9011 11723
rect 9045 11689 9079 11723
rect 9113 11689 9147 11723
rect 9181 11689 9215 11723
rect 9249 11689 9283 11723
rect 9317 11689 9351 11723
rect 9385 11689 9419 11723
rect 9453 11689 9487 11723
rect 9521 11689 9555 11723
rect 9589 11689 9623 11723
rect 9657 11689 9691 11723
rect 9725 11689 9759 11723
rect 9793 11689 9827 11723
rect 9861 11689 9895 11723
rect 1117 11655 1219 11665
rect 3717 11655 3751 11689
rect 3717 11587 3751 11621
rect 3717 11519 3751 11553
rect 3717 11451 3751 11485
rect 1219 11246 1287 11281
rect 1219 11212 1253 11246
rect 3717 11383 3751 11417
rect 5557 11621 5591 11655
rect 5557 11553 5591 11587
rect 5557 11485 5591 11519
rect 5557 11417 5591 11451
rect 3717 11315 3751 11349
rect 3717 11247 3751 11281
rect 1219 11177 1287 11212
rect 1219 11143 1253 11177
rect 1219 11108 1287 11143
rect 1219 11074 1253 11108
rect 1219 11039 1287 11074
rect 1219 11005 1253 11039
rect 1219 10970 1287 11005
rect 1219 10936 1253 10970
rect 1219 10901 1287 10936
rect 1219 10867 1253 10901
rect 1219 10832 1287 10867
rect 1219 10798 1253 10832
rect 1219 10763 1287 10798
rect 1219 10729 1253 10763
rect 1219 10694 1287 10729
rect 1219 10660 1253 10694
rect 1219 10625 1287 10660
rect 1219 10591 1253 10625
rect 1219 10556 1287 10591
rect 1219 10522 1253 10556
rect 1219 10487 1287 10522
rect 1219 10453 1253 10487
rect 1219 10418 1287 10453
rect 3717 11179 3751 11213
rect 3717 11111 3751 11145
rect 3717 11043 3751 11077
rect 3717 10975 3751 11009
rect 3717 10907 3751 10941
rect 3717 10839 3751 10873
rect 3717 10771 3751 10805
rect 3717 10703 3751 10737
rect 3717 10635 3751 10669
rect 3717 10567 3751 10601
rect 3717 10499 3751 10533
rect 1219 10384 1253 10418
rect 1219 10349 1287 10384
rect 1219 10315 1253 10349
rect 1219 10280 1287 10315
rect 1219 10246 1253 10280
rect 1219 10211 1287 10246
rect 1219 10177 1253 10211
rect 1219 10142 1287 10177
rect 3717 10431 3751 10465
rect 3717 10363 3751 10397
rect 3717 10295 3751 10329
rect 3717 10227 3751 10261
rect 3717 10159 3751 10193
rect 1219 10108 1253 10142
rect 1219 10073 1287 10108
rect 1219 10039 1253 10073
rect 1219 10004 1287 10039
rect 1219 9970 1253 10004
rect 1219 9935 1287 9970
rect 1219 9901 1253 9935
rect 1219 9866 1287 9901
rect 1219 9832 1253 9866
rect 1219 9797 1287 9832
rect 1219 9763 1253 9797
rect 1219 9728 1287 9763
rect 1219 9694 1253 9728
rect 1219 9659 1287 9694
rect 1219 9625 1253 9659
rect 1219 9590 1287 9625
rect 1219 9556 1253 9590
rect 1219 9521 1287 9556
rect 1219 9487 1253 9521
rect 1219 9452 1287 9487
rect 1219 9418 1253 9452
rect 1219 9383 1287 9418
rect 1219 9349 1253 9383
rect 3717 10091 3751 10125
rect 3717 10023 3751 10057
rect 3717 9955 3751 9989
rect 3717 9887 3751 9921
rect 3717 9819 3751 9853
rect 3717 9751 3751 9785
rect 3717 9683 3751 9717
rect 3717 9615 3751 9649
rect 3717 9547 3751 9581
rect 3717 9479 3751 9513
rect 3717 9411 3751 9445
rect 1219 9314 1287 9349
rect 1219 9280 1253 9314
rect 3717 9343 3751 9377
rect 1219 9245 1287 9280
rect 1219 9211 1253 9245
rect 1219 9176 1287 9211
rect 1219 9142 1253 9176
rect 1219 9107 1287 9142
rect 1219 9073 1253 9107
rect 1219 9038 1287 9073
rect 1219 9004 1253 9038
rect 1219 8969 1287 9004
rect 1219 8935 1253 8969
rect 1219 8900 1287 8935
rect 1219 8866 1253 8900
rect 1219 8831 1287 8866
rect 1219 8797 1253 8831
rect 1219 8762 1287 8797
rect 1219 8728 1253 8762
rect 1219 8693 1287 8728
rect 1219 8659 1253 8693
rect 1219 8624 1287 8659
rect 1219 8590 1253 8624
rect 1219 8555 1287 8590
rect 1219 8521 1253 8555
rect 1219 8486 1287 8521
rect 3717 9275 3751 9309
rect 3717 9207 3751 9241
rect 3717 9139 3751 9173
rect 3717 9071 3751 9105
rect 3717 9003 3751 9037
rect 3717 8935 3751 8969
rect 3717 8867 3751 8901
rect 3717 8799 3751 8833
rect 3717 8731 3751 8765
rect 3717 8663 3751 8697
rect 3717 8595 3751 8629
rect 3717 8527 3751 8561
rect 1219 8452 1253 8486
rect 1219 8417 1287 8452
rect 1219 8383 1253 8417
rect 1219 8348 1287 8383
rect 1219 8314 1253 8348
rect 1219 8279 1287 8314
rect 1219 8245 1253 8279
rect 1219 8210 1287 8245
rect 3717 8459 3751 8493
rect 3717 8391 3751 8425
rect 3717 8323 3751 8357
rect 3717 8255 3751 8289
rect 1219 8176 1253 8210
rect 1219 8141 1287 8176
rect 1219 8107 1253 8141
rect 1219 8072 1287 8107
rect 1219 8038 1253 8072
rect 1219 8003 1287 8038
rect 1219 7969 1253 8003
rect 1219 7934 1287 7969
rect 1219 7900 1253 7934
rect 1219 7865 1287 7900
rect 1219 7831 1253 7865
rect 1219 7796 1287 7831
rect 1219 7762 1253 7796
rect 1219 7727 1287 7762
rect 1219 7693 1253 7727
rect 1219 7658 1287 7693
rect 1219 7624 1253 7658
rect 1219 7589 1287 7624
rect 1219 7555 1253 7589
rect 1219 7520 1287 7555
rect 1219 7486 1253 7520
rect 1219 7451 1287 7486
rect 1219 7417 1253 7451
rect 1219 7382 1287 7417
rect 3717 8187 3751 8221
rect 3717 8119 3751 8153
rect 3717 8051 3751 8085
rect 3717 7983 3751 8017
rect 3717 7915 3751 7949
rect 3717 7847 3751 7881
rect 3717 7779 3751 7813
rect 3717 7711 3751 7745
rect 3717 7643 3751 7677
rect 3717 7575 3751 7609
rect 3717 7507 3751 7541
rect 3717 7439 3751 7473
rect 1219 7348 1253 7382
rect 1219 7313 1287 7348
rect 1219 7279 1253 7313
rect 1219 7244 1287 7279
rect 3717 7371 3751 7405
rect 3717 7303 3751 7337
rect 1219 7210 1253 7244
rect 3717 7235 3751 7269
rect 1219 7175 1287 7210
rect 1219 7141 1253 7175
rect 1219 7106 1287 7141
rect 1219 7072 1253 7106
rect 1219 7037 1287 7072
rect 1219 7003 1253 7037
rect 1219 6963 1287 7003
rect 3717 7167 3751 7201
rect 3717 7099 3751 7133
rect 3717 7031 3751 7065
rect 3717 6963 3751 6997
rect 1287 6929 1321 6963
rect 1355 6929 1389 6963
rect 1423 6929 1457 6963
rect 1491 6929 1525 6963
rect 1559 6929 1593 6963
rect 1627 6929 1661 6963
rect 1695 6929 1729 6963
rect 1763 6929 1797 6963
rect 1831 6929 1865 6963
rect 1899 6929 1933 6963
rect 1967 6929 2001 6963
rect 2035 6929 2069 6963
rect 2103 6929 2137 6963
rect 2171 6929 2205 6963
rect 2239 6929 2273 6963
rect 2307 6929 2341 6963
rect 2375 6929 2409 6963
rect 2443 6929 2477 6963
rect 2511 6929 2545 6963
rect 2579 6929 2613 6963
rect 2647 6929 2681 6963
rect 2715 6929 2749 6963
rect 2783 6929 2817 6963
rect 2851 6929 2885 6963
rect 2919 6929 2953 6963
rect 2987 6929 3021 6963
rect 3055 6929 3089 6963
rect 3123 6929 3157 6963
rect 3191 6929 3225 6963
rect 3259 6929 3293 6963
rect 3327 6929 3361 6963
rect 3395 6929 3429 6963
rect 3463 6929 3497 6963
rect 3531 6929 3565 6963
rect 3599 6929 3633 6963
rect 3667 6929 3717 6963
rect 3717 6895 3751 6929
rect 3717 6827 3751 6861
rect 3717 6759 3751 6793
rect 3717 6691 3751 6725
rect 3717 6623 3751 6657
rect 3717 6555 3751 6589
rect 3717 6487 3751 6521
rect 3717 6419 3751 6453
rect 3717 6351 3751 6385
rect 3717 6283 3751 6317
rect 3717 6215 3751 6249
rect 3717 6147 3751 6181
rect 3717 6079 3751 6113
rect 3717 6011 3751 6045
rect 3717 5943 3751 5977
rect 3717 5875 3751 5909
rect 3717 5807 3751 5841
rect 3717 5739 3751 5773
rect 3717 5671 3751 5705
rect 3717 5603 3751 5637
rect 3717 5535 3751 5569
rect 3717 5467 3751 5501
rect 3717 5399 3751 5433
rect 3717 5331 3751 5365
rect 3717 5263 3751 5297
rect 3717 5195 3751 5229
rect 3717 5127 3751 5161
rect 3717 5059 3751 5093
rect 3717 4991 3751 5025
rect 3717 4923 3751 4957
rect 3717 4855 3751 4889
rect 3717 4787 3751 4821
rect 3717 4719 3751 4753
rect 3717 4651 3751 4685
rect 3717 4583 3751 4617
rect 1117 3878 1185 3913
rect 1151 3844 1185 3878
rect 1117 3809 1185 3844
rect 1151 3775 1185 3809
rect 1117 3740 1185 3775
rect 1151 3706 1185 3740
rect 1117 3671 1185 3706
rect 1151 3637 1185 3671
rect 1117 3602 1185 3637
rect 1151 3568 1185 3602
rect 1117 3533 1185 3568
rect 1151 3499 1185 3533
rect 1117 3464 1185 3499
rect 1151 3430 1185 3464
rect 1117 3395 1185 3430
rect 1151 3361 1185 3395
rect 1117 3326 1185 3361
rect 1151 3292 1185 3326
rect 1117 3257 1185 3292
rect 1151 3223 1185 3257
rect 1117 3188 1185 3223
rect 1151 3154 1185 3188
rect 1117 3119 1185 3154
rect 1151 3085 1185 3119
rect 1117 3050 1185 3085
rect 1151 3016 1185 3050
rect 1117 2981 1185 3016
rect 1151 2947 1185 2981
rect 1117 2912 1185 2947
rect 1151 2878 1185 2912
rect 1117 2843 1185 2878
rect 1151 2809 1185 2843
rect 1117 2774 1185 2809
rect 1151 2740 1185 2774
rect 1117 2705 1185 2740
rect 1151 2671 1185 2705
rect 1117 2636 1185 2671
rect 1151 2602 1185 2636
rect 1117 2577 1185 2602
rect 3717 4515 3751 4549
rect 3717 4447 3751 4481
rect 3717 4379 3751 4413
rect 3717 4311 3751 4345
rect 3717 4243 3751 4277
rect 3717 4175 3751 4209
rect 3717 4107 3751 4141
rect 3717 4039 3751 4073
rect 3717 3971 3751 4005
rect 3717 3903 3751 3937
rect 5557 11349 5591 11383
rect 7397 11655 7431 11689
rect 7397 11587 7431 11621
rect 7397 11519 7431 11553
rect 7397 11451 7431 11485
rect 9929 11655 9963 11723
rect 9929 11587 9963 11621
rect 9929 11519 9963 11553
rect 9929 11451 9963 11485
rect 7397 11383 7431 11417
rect 5557 11281 5591 11315
rect 5557 11213 5591 11247
rect 5557 11145 5591 11179
rect 5557 11077 5591 11111
rect 5557 11009 5591 11043
rect 5557 10941 5591 10975
rect 5557 10873 5591 10907
rect 5557 10805 5591 10839
rect 5557 10737 5591 10771
rect 5557 10669 5591 10703
rect 5557 10601 5591 10635
rect 5557 10533 5591 10567
rect 5557 10465 5591 10499
rect 5557 10397 5591 10431
rect 5557 10329 5591 10363
rect 5557 10261 5591 10295
rect 5557 10193 5591 10227
rect 5557 10125 5591 10159
rect 5557 10057 5591 10091
rect 5557 9989 5591 10023
rect 5557 9921 5591 9955
rect 5557 9853 5591 9887
rect 5557 9785 5591 9819
rect 5557 9717 5591 9751
rect 5557 9649 5591 9683
rect 5557 9581 5591 9615
rect 5557 9513 5591 9547
rect 5557 9445 5591 9479
rect 5557 9377 5591 9411
rect 5557 9309 5591 9343
rect 5557 9241 5591 9275
rect 5557 9173 5591 9207
rect 5557 9105 5591 9139
rect 5557 9037 5591 9071
rect 5557 8969 5591 9003
rect 5557 8901 5591 8935
rect 5557 8833 5591 8867
rect 5557 8765 5591 8799
rect 5557 8697 5591 8731
rect 5557 8629 5591 8663
rect 5557 8561 5591 8595
rect 5557 8493 5591 8527
rect 5557 8425 5591 8459
rect 5557 8357 5591 8391
rect 5557 8289 5591 8323
rect 5557 8221 5591 8255
rect 5557 8153 5591 8187
rect 5557 8085 5591 8119
rect 5557 8017 5591 8051
rect 5557 7949 5591 7983
rect 5557 7881 5591 7915
rect 5557 7813 5591 7847
rect 5557 7745 5591 7779
rect 5557 7677 5591 7711
rect 5557 7609 5591 7643
rect 5557 7541 5591 7575
rect 5557 7473 5591 7507
rect 5557 7405 5591 7439
rect 5557 7337 5591 7371
rect 5557 7269 5591 7303
rect 5557 7201 5591 7235
rect 5557 7133 5591 7167
rect 5557 7065 5591 7099
rect 5557 6997 5591 7031
rect 5557 6929 5591 6963
rect 5557 6861 5591 6895
rect 5557 6793 5591 6827
rect 5557 6725 5591 6759
rect 5557 6657 5591 6691
rect 5557 6589 5591 6623
rect 5557 6521 5591 6555
rect 5557 6453 5591 6487
rect 5557 6385 5591 6419
rect 5557 6317 5591 6351
rect 5557 6249 5591 6283
rect 5557 6181 5591 6215
rect 5557 6113 5591 6147
rect 5557 6045 5591 6079
rect 5557 5977 5591 6011
rect 5557 5909 5591 5943
rect 5557 5841 5591 5875
rect 5557 5773 5591 5807
rect 5557 5705 5591 5739
rect 5557 5637 5591 5671
rect 5557 5569 5591 5603
rect 5557 5501 5591 5535
rect 5557 5433 5591 5467
rect 5557 5365 5591 5399
rect 5557 5297 5591 5331
rect 5557 5229 5591 5263
rect 5557 5161 5591 5195
rect 5557 5093 5591 5127
rect 5557 5025 5591 5059
rect 5557 4957 5591 4991
rect 5557 4889 5591 4923
rect 5557 4821 5591 4855
rect 5557 4753 5591 4787
rect 5557 4685 5591 4719
rect 5557 4617 5591 4651
rect 5557 4549 5591 4583
rect 5557 4481 5591 4515
rect 5557 4413 5591 4447
rect 5557 4345 5591 4379
rect 5557 4277 5591 4311
rect 5557 4209 5591 4243
rect 5557 4141 5591 4175
rect 5557 4073 5591 4107
rect 5557 4005 5591 4039
rect 5557 3937 5591 3971
rect 3717 3835 3751 3869
rect 3717 3767 3751 3801
rect 3717 3699 3751 3733
rect 7397 11315 7431 11349
rect 7397 11247 7431 11281
rect 9929 11383 9963 11417
rect 9929 11315 9963 11349
rect 9929 11247 9963 11281
rect 7397 11179 7431 11213
rect 7397 11111 7431 11145
rect 7397 11043 7431 11077
rect 7397 10975 7431 11009
rect 7397 10907 7431 10941
rect 7397 10839 7431 10873
rect 7397 10771 7431 10805
rect 7397 10703 7431 10737
rect 7397 10635 7431 10669
rect 7397 10567 7431 10601
rect 7397 10499 7431 10533
rect 7397 10431 7431 10465
rect 9929 11179 9963 11213
rect 9929 11111 9963 11145
rect 9929 11043 9963 11077
rect 9929 10975 9963 11009
rect 9929 10907 9963 10941
rect 9929 10839 9963 10873
rect 9929 10771 9963 10805
rect 9929 10703 9963 10737
rect 9929 10635 9963 10669
rect 9929 10567 9963 10601
rect 9929 10499 9963 10533
rect 7397 10363 7431 10397
rect 7397 10295 7431 10329
rect 7397 10227 7431 10261
rect 7397 10159 7431 10193
rect 9929 10431 9963 10465
rect 9929 10363 9963 10397
rect 9929 10295 9963 10329
rect 9929 10227 9963 10261
rect 9929 10159 9963 10193
rect 7397 10091 7431 10125
rect 7397 10023 7431 10057
rect 7397 9955 7431 9989
rect 7397 9887 7431 9921
rect 7397 9819 7431 9853
rect 7397 9751 7431 9785
rect 7397 9683 7431 9717
rect 7397 9615 7431 9649
rect 7397 9547 7431 9581
rect 7397 9479 7431 9513
rect 7397 9411 7431 9445
rect 7397 9343 7431 9377
rect 9929 10091 9963 10125
rect 9929 10023 9963 10057
rect 9929 9955 9963 9989
rect 9929 9887 9963 9921
rect 9929 9819 9963 9853
rect 9929 9751 9963 9785
rect 9929 9683 9963 9717
rect 9929 9615 9963 9649
rect 9929 9547 9963 9581
rect 9929 9479 9963 9513
rect 9929 9411 9963 9445
rect 7397 9275 7431 9309
rect 9929 9343 9963 9377
rect 7397 9207 7431 9241
rect 7397 9139 7431 9173
rect 7397 9071 7431 9105
rect 7397 9003 7431 9037
rect 7397 8935 7431 8969
rect 7397 8867 7431 8901
rect 7397 8799 7431 8833
rect 7397 8731 7431 8765
rect 7397 8663 7431 8697
rect 7397 8595 7431 8629
rect 7397 8527 7431 8561
rect 9929 9275 9963 9309
rect 9929 9207 9963 9241
rect 9929 9139 9963 9173
rect 9929 9071 9963 9105
rect 9929 9003 9963 9037
rect 9929 8935 9963 8969
rect 9929 8867 9963 8901
rect 9929 8799 9963 8833
rect 9929 8731 9963 8765
rect 9929 8663 9963 8697
rect 9929 8595 9963 8629
rect 9929 8527 9963 8561
rect 7397 8459 7431 8493
rect 7397 8391 7431 8425
rect 7397 8323 7431 8357
rect 7397 8255 7431 8289
rect 7397 8187 7431 8221
rect 9929 8459 9963 8493
rect 9929 8391 9963 8425
rect 9929 8323 9963 8357
rect 9929 8255 9963 8289
rect 7397 8119 7431 8153
rect 7397 8051 7431 8085
rect 7397 7983 7431 8017
rect 7397 7915 7431 7949
rect 7397 7847 7431 7881
rect 7397 7779 7431 7813
rect 7397 7711 7431 7745
rect 7397 7643 7431 7677
rect 7397 7575 7431 7609
rect 7397 7507 7431 7541
rect 7397 7439 7431 7473
rect 9929 8187 9963 8221
rect 9929 8119 9963 8153
rect 9929 8051 9963 8085
rect 9963 8017 9997 8040
rect 9929 8006 9997 8017
rect 10031 8006 10065 8040
rect 10099 8006 10133 8040
rect 10167 8006 10201 8040
rect 10235 8006 10269 8040
rect 10303 8006 10337 8040
rect 10371 8006 10405 8040
rect 10439 8006 10473 8040
rect 10507 8006 10541 8040
rect 10575 8006 10609 8040
rect 10643 8006 10677 8040
rect 10711 8006 10745 8040
rect 10779 8006 10813 8040
rect 10847 8006 10881 8040
rect 10915 8006 10949 8040
rect 10983 8006 11017 8040
rect 11051 8006 11085 8040
rect 11119 8006 11153 8040
rect 11187 8006 11221 8040
rect 11255 8006 11289 8040
rect 11323 8006 11357 8040
rect 11391 8006 11425 8040
rect 11459 8006 11493 8040
rect 11527 8006 11561 8040
rect 11595 8006 11629 8040
rect 11663 8006 11697 8040
rect 11731 8006 11765 8040
rect 11799 8006 11833 8040
rect 11867 8006 11901 8040
rect 11935 8006 11969 8040
rect 12003 8006 12037 8040
rect 12071 8006 12105 8040
rect 12139 8006 12173 8040
rect 12207 8006 12241 8040
rect 12275 8006 12309 8040
rect 12343 8006 12377 8040
rect 12411 8006 12445 8040
rect 12479 8006 12513 8040
rect 12547 8006 12581 8040
rect 12615 8006 12649 8040
rect 12683 8006 12717 8040
rect 12751 8006 12785 8040
rect 12819 8006 12853 8040
rect 12887 8006 12921 8040
rect 12955 8006 12989 8040
rect 13023 8006 13103 8040
rect 9929 7983 9963 8006
rect 9929 7915 9963 7949
rect 9929 7847 9963 7881
rect 9929 7779 9963 7813
rect 9929 7711 9963 7745
rect 13069 7938 13103 7972
rect 13069 7870 13103 7904
rect 13069 7802 13103 7836
rect 13069 7734 13103 7768
rect 9929 7643 9963 7677
rect 9929 7575 9963 7609
rect 9929 7507 9963 7541
rect 9929 7439 9963 7473
rect 7397 7371 7431 7405
rect 7397 7303 7431 7337
rect 7397 7235 7431 7269
rect 9929 7371 9963 7405
rect 9929 7303 9963 7337
rect 9929 7235 9963 7269
rect 7397 7167 7431 7201
rect 7397 7099 7431 7133
rect 7397 7031 7431 7065
rect 7397 6963 7431 6997
rect 9929 7167 9963 7201
rect 9929 7099 9963 7133
rect 9929 7031 9963 7065
rect 9929 6963 9963 6997
rect 7431 6929 7481 6963
rect 7515 6929 7549 6963
rect 7583 6929 7617 6963
rect 7651 6929 7685 6963
rect 7719 6929 7753 6963
rect 7787 6929 7821 6963
rect 7855 6929 7889 6963
rect 7923 6929 7957 6963
rect 7991 6929 8025 6963
rect 8059 6929 8093 6963
rect 8127 6929 8161 6963
rect 8195 6929 8229 6963
rect 8263 6929 8297 6963
rect 8331 6929 8365 6963
rect 8399 6929 8433 6963
rect 8467 6929 8501 6963
rect 8535 6929 8569 6963
rect 8603 6929 8637 6963
rect 8671 6929 8705 6963
rect 8739 6929 8773 6963
rect 8807 6929 8841 6963
rect 8875 6929 8909 6963
rect 8943 6929 8977 6963
rect 9011 6929 9045 6963
rect 9079 6929 9113 6963
rect 9147 6929 9181 6963
rect 9215 6929 9249 6963
rect 9283 6929 9317 6963
rect 9351 6929 9385 6963
rect 9419 6929 9453 6963
rect 9487 6929 9521 6963
rect 9555 6929 9589 6963
rect 9623 6929 9657 6963
rect 9691 6929 9725 6963
rect 9759 6929 9793 6963
rect 9827 6929 9861 6963
rect 9895 6929 9929 6963
rect 7397 6895 7431 6929
rect 7397 6827 7431 6861
rect 7397 6759 7431 6793
rect 7397 6691 7431 6725
rect 9929 6895 9963 6929
rect 9929 6827 9963 6861
rect 9929 6759 9963 6793
rect 9929 6691 9963 6725
rect 7397 6623 7431 6657
rect 7397 6555 7431 6589
rect 7397 6487 7431 6521
rect 9929 6623 9963 6657
rect 9929 6555 9963 6589
rect 9929 6487 9963 6521
rect 7397 6419 7431 6453
rect 7397 6351 7431 6385
rect 7397 6283 7431 6317
rect 7397 6215 7431 6249
rect 7397 6147 7431 6181
rect 7397 6079 7431 6113
rect 7397 6011 7431 6045
rect 7397 5943 7431 5977
rect 7397 5875 7431 5909
rect 7397 5807 7431 5841
rect 7397 5739 7431 5773
rect 7397 5671 7431 5705
rect 9929 6419 9963 6453
rect 9929 6351 9963 6385
rect 9929 6283 9963 6317
rect 9929 6215 9963 6249
rect 9929 6147 9963 6181
rect 9929 6079 9963 6113
rect 9929 6011 9963 6045
rect 9929 5943 9963 5977
rect 9929 5875 9963 5909
rect 9929 5807 9963 5841
rect 9929 5739 9963 5773
rect 9929 5671 9963 5705
rect 7397 5603 7431 5637
rect 7397 5535 7431 5569
rect 7397 5467 7431 5501
rect 7397 5399 7431 5433
rect 9929 5603 9963 5637
rect 9929 5535 9963 5569
rect 9929 5467 9963 5501
rect 9929 5399 9963 5433
rect 7397 5331 7431 5365
rect 7397 5263 7431 5297
rect 7397 5195 7431 5229
rect 7397 5127 7431 5161
rect 7397 5059 7431 5093
rect 7397 4991 7431 5025
rect 7397 4923 7431 4957
rect 7397 4855 7431 4889
rect 7397 4787 7431 4821
rect 7397 4719 7431 4753
rect 7397 4651 7431 4685
rect 7397 4583 7431 4617
rect 9929 5331 9963 5365
rect 9929 5263 9963 5297
rect 9929 5195 9963 5229
rect 9929 5127 9963 5161
rect 9929 5059 9963 5093
rect 9929 4991 9963 5025
rect 9929 4923 9963 4957
rect 9929 4855 9963 4889
rect 9929 4787 9963 4821
rect 9929 4719 9963 4753
rect 9929 4651 9963 4685
rect 7397 4515 7431 4549
rect 9929 4583 9963 4617
rect 7397 4447 7431 4481
rect 7397 4379 7431 4413
rect 7397 4311 7431 4345
rect 7397 4243 7431 4277
rect 7397 4175 7431 4209
rect 7397 4107 7431 4141
rect 7397 4039 7431 4073
rect 7397 3971 7431 4005
rect 5557 3869 5591 3903
rect 5557 3801 5591 3835
rect 5557 3687 5591 3767
rect 7397 3903 7431 3937
rect 7397 3835 7431 3869
rect 7397 3767 7431 3801
rect 9929 4515 9963 4549
rect 9929 4447 9963 4481
rect 9929 4379 9963 4413
rect 9929 4311 9963 4345
rect 9929 4243 9963 4277
rect 9929 4175 9963 4209
rect 9929 4107 9963 4141
rect 9929 4039 9963 4073
rect 9929 3971 9963 4005
rect 9929 3903 9963 3937
rect 9929 3835 9963 3869
rect 9929 3767 9963 3801
rect 7397 3699 7431 3733
rect 3751 3665 3785 3687
rect 3717 3653 3785 3665
rect 3819 3653 3853 3687
rect 3887 3653 3921 3687
rect 3955 3653 3989 3687
rect 4023 3653 4057 3687
rect 4091 3653 4125 3687
rect 4159 3653 4193 3687
rect 4227 3653 4261 3687
rect 4295 3653 4329 3687
rect 4363 3653 4397 3687
rect 4431 3653 4465 3687
rect 4499 3653 4533 3687
rect 4567 3653 4601 3687
rect 4635 3653 4669 3687
rect 4703 3653 4737 3687
rect 4771 3653 4805 3687
rect 4839 3653 4873 3687
rect 4907 3653 4941 3687
rect 4975 3653 5009 3687
rect 5043 3653 5077 3687
rect 5111 3653 5145 3687
rect 5179 3653 5213 3687
rect 5247 3653 5281 3687
rect 5315 3653 5349 3687
rect 5383 3653 5417 3687
rect 5451 3653 5485 3687
rect 5519 3653 5625 3687
rect 5659 3653 5693 3687
rect 5727 3653 5761 3687
rect 5795 3653 5829 3687
rect 5863 3653 5897 3687
rect 5931 3653 5965 3687
rect 5999 3653 6033 3687
rect 6067 3653 6101 3687
rect 6135 3653 6169 3687
rect 6203 3653 6237 3687
rect 6271 3653 6305 3687
rect 6339 3653 6373 3687
rect 6407 3653 6441 3687
rect 6475 3653 6509 3687
rect 6543 3653 6577 3687
rect 6611 3653 6645 3687
rect 6679 3653 6713 3687
rect 6747 3653 6781 3687
rect 6815 3653 6849 3687
rect 6883 3653 6917 3687
rect 6951 3653 6985 3687
rect 7019 3653 7053 3687
rect 7087 3653 7121 3687
rect 7155 3653 7189 3687
rect 7223 3653 7257 3687
rect 7291 3653 7325 3687
rect 7359 3665 7397 3687
rect 7359 3653 7431 3665
rect 3717 3631 3751 3653
rect 3717 3563 3751 3597
rect 3717 3495 3751 3529
rect 3717 3427 3751 3461
rect 3717 3359 3751 3393
rect 7397 3631 7431 3653
rect 7397 3563 7431 3597
rect 7397 3495 7431 3529
rect 7397 3427 7431 3461
rect 9929 3699 9963 3733
rect 9929 3631 9963 3665
rect 9929 3563 9963 3597
rect 9929 3495 9963 3529
rect 3717 3291 3751 3325
rect 3717 3223 3751 3257
rect 3717 3155 3751 3189
rect 3717 3087 3751 3121
rect 3717 3019 3751 3053
rect 3717 2951 3751 2985
rect 3717 2883 3751 2917
rect 3717 2815 3751 2849
rect 3717 2747 3751 2781
rect 3717 2679 3751 2713
rect 1117 2567 1287 2577
rect 1151 2543 1287 2567
rect 1151 2533 1185 2543
rect 1117 2509 1185 2533
rect 1219 2542 1287 2543
rect 1219 2509 1253 2542
rect 1117 2508 1253 2509
rect 1117 2498 1287 2508
rect 3717 2611 3751 2645
rect 3717 2543 3751 2577
rect 1151 2475 1287 2498
rect 1151 2464 1185 2475
rect 1117 2441 1185 2464
rect 1219 2473 1287 2475
rect 1219 2441 1253 2473
rect 1117 2439 1253 2441
rect 3717 2475 3751 2509
rect 1117 2429 1287 2439
rect 1151 2407 1287 2429
rect 1151 2395 1185 2407
rect 1117 2373 1185 2395
rect 1219 2404 1287 2407
rect 1219 2373 1253 2404
rect 1117 2370 1253 2373
rect 1117 2360 1287 2370
rect 1151 2339 1287 2360
rect 1151 2326 1185 2339
rect 1117 2305 1185 2326
rect 1219 2335 1287 2339
rect 1219 2305 1253 2335
rect 1117 2301 1253 2305
rect 1117 2291 1287 2301
rect 1151 2271 1287 2291
rect 1151 2257 1185 2271
rect 1117 2237 1185 2257
rect 1219 2266 1287 2271
rect 1219 2237 1253 2266
rect 1117 2232 1253 2237
rect 1117 2222 1287 2232
rect 1151 2203 1287 2222
rect 3717 2407 3751 2441
rect 3717 2339 3751 2373
rect 3717 2271 3751 2305
rect 1151 2188 1185 2203
rect 1117 2169 1185 2188
rect 1219 2197 1371 2203
rect 1219 2169 1253 2197
rect 1117 2163 1253 2169
rect 1287 2169 1371 2197
rect 1405 2169 1439 2203
rect 1473 2169 1507 2203
rect 1541 2169 1575 2203
rect 1609 2169 1643 2203
rect 1677 2169 1711 2203
rect 1745 2169 1779 2203
rect 1813 2169 1847 2203
rect 1881 2169 1915 2203
rect 1949 2169 1983 2203
rect 2017 2169 2051 2203
rect 2085 2169 2119 2203
rect 2153 2169 2187 2203
rect 2221 2169 2255 2203
rect 2289 2169 2323 2203
rect 2357 2169 2391 2203
rect 2425 2169 2459 2203
rect 2493 2169 2527 2203
rect 2561 2169 2595 2203
rect 2629 2169 2663 2203
rect 2697 2169 2731 2203
rect 2765 2169 2799 2203
rect 2833 2169 2867 2203
rect 2901 2169 2935 2203
rect 2969 2169 3003 2203
rect 3037 2169 3071 2203
rect 3105 2169 3139 2203
rect 3173 2169 3207 2203
rect 3241 2169 3275 2203
rect 3309 2169 3343 2203
rect 3377 2169 3411 2203
rect 3445 2169 3479 2203
rect 3513 2169 3547 2203
rect 3581 2169 3615 2203
rect 3649 2169 3683 2203
rect 3717 2169 3751 2237
rect 1117 2153 1287 2163
rect 1151 2135 1287 2153
rect 1151 2119 1185 2135
rect 1117 2101 1185 2119
rect 1219 2128 1287 2135
rect 1219 2101 1253 2128
rect 1117 2094 1253 2101
rect 1117 2084 1287 2094
rect 1151 2067 1287 2084
rect 1151 2050 1185 2067
rect 1117 2033 1185 2050
rect 1219 2059 1287 2067
rect 1219 2033 1253 2059
rect 1117 2025 1253 2033
rect 1117 2015 1287 2025
rect 1151 1999 1287 2015
rect 1151 1981 1185 1999
rect 1117 1965 1185 1981
rect 1219 1990 1287 1999
rect 1219 1965 1253 1990
rect 1117 1956 1253 1965
rect 1117 1946 1287 1956
rect 1151 1931 1287 1946
rect 1151 1912 1185 1931
rect 1117 1897 1185 1912
rect 1219 1921 1287 1931
rect 1219 1897 1253 1921
rect 1117 1887 1253 1897
rect 7397 3359 7431 3393
rect 7397 3291 7431 3325
rect 7397 3223 7431 3257
rect 7397 3155 7431 3189
rect 7397 3087 7431 3121
rect 7397 3019 7431 3053
rect 7397 2951 7431 2985
rect 7397 2883 7431 2917
rect 7397 2815 7431 2849
rect 7397 2747 7431 2781
rect 7397 2679 7431 2713
rect 9929 3427 9963 3461
rect 9929 3359 9963 3393
rect 9929 3291 9963 3325
rect 9929 3223 9963 3257
rect 9929 3155 9963 3189
rect 9929 3087 9963 3121
rect 9929 3019 9963 3053
rect 9929 2951 9963 2985
rect 9929 2883 9963 2917
rect 9929 2815 9963 2849
rect 9929 2747 9963 2781
rect 9929 2679 9963 2713
rect 7397 2611 7431 2645
rect 7397 2543 7431 2577
rect 7397 2475 7431 2509
rect 9929 2611 9963 2645
rect 9929 2543 9963 2577
rect 9929 2475 9963 2509
rect 7397 2407 7431 2441
rect 7397 2339 7431 2373
rect 7397 2271 7431 2305
rect 7397 2169 7431 2237
rect 9929 2407 9963 2441
rect 9929 2339 9963 2373
rect 9929 2271 9963 2305
rect 9929 2203 9963 2237
rect 7465 2169 7499 2203
rect 7533 2169 7567 2203
rect 7601 2169 7635 2203
rect 7669 2169 7703 2203
rect 7737 2169 7771 2203
rect 7805 2169 7839 2203
rect 7873 2169 7907 2203
rect 7941 2169 7975 2203
rect 8009 2169 8043 2203
rect 8077 2169 8111 2203
rect 8145 2169 8179 2203
rect 8213 2169 8247 2203
rect 8281 2169 8315 2203
rect 8349 2169 8383 2203
rect 8417 2169 8451 2203
rect 8485 2169 8519 2203
rect 8553 2169 8587 2203
rect 8621 2169 8655 2203
rect 8689 2169 8723 2203
rect 8757 2169 8791 2203
rect 8825 2169 8859 2203
rect 8893 2169 8927 2203
rect 8961 2169 8995 2203
rect 9029 2169 9063 2203
rect 9097 2169 9131 2203
rect 9165 2169 9199 2203
rect 9233 2169 9267 2203
rect 9301 2169 9335 2203
rect 9369 2169 9403 2203
rect 9437 2169 9471 2203
rect 9505 2169 9539 2203
rect 9573 2169 9607 2203
rect 9641 2169 9675 2203
rect 9709 2169 9743 2203
rect 9777 2169 9811 2203
rect 9845 2169 9929 2203
rect 1117 1877 1287 1887
rect 1151 1863 1287 1877
rect 1151 1843 1185 1863
rect 1117 1829 1185 1843
rect 1219 1852 1287 1863
rect 1219 1829 1253 1852
rect 1117 1818 1253 1829
rect 1117 1808 1287 1818
rect 1151 1795 1287 1808
rect 1151 1774 1185 1795
rect 1117 1761 1185 1774
rect 1219 1783 1287 1795
rect 1219 1761 1253 1783
rect 1117 1749 1253 1761
rect 9929 2135 9963 2169
rect 9929 2067 9963 2101
rect 9929 1999 9963 2033
rect 9929 1931 9963 1965
rect 1117 1739 1287 1749
rect 1151 1727 1287 1739
rect 1151 1705 1185 1727
rect 1117 1693 1185 1705
rect 1219 1714 1287 1727
rect 1219 1693 1253 1714
rect 1117 1680 1253 1693
rect 1117 1670 1287 1680
rect 1151 1659 1287 1670
rect 1151 1636 1185 1659
rect 1117 1625 1185 1636
rect 1219 1645 1287 1659
rect 1219 1625 1253 1645
rect 1117 1611 1253 1625
rect 1117 1601 1287 1611
rect 1151 1591 1287 1601
rect 1151 1567 1185 1591
rect 1117 1557 1185 1567
rect 1219 1576 1287 1591
rect 1219 1557 1253 1576
rect 1117 1542 1253 1557
rect 1117 1532 1287 1542
rect 1151 1523 1287 1532
rect 1151 1498 1185 1523
rect 1117 1489 1185 1498
rect 1219 1507 1287 1523
rect 1219 1489 1253 1507
rect 1117 1473 1253 1489
rect 1117 1463 1287 1473
rect 1151 1455 1287 1463
rect 1151 1429 1185 1455
rect 1117 1421 1185 1429
rect 1219 1438 1287 1455
rect 1219 1421 1253 1438
rect 1117 1404 1253 1421
rect 1117 1394 1287 1404
rect 1151 1387 1287 1394
rect 1151 1360 1185 1387
rect 1117 1353 1185 1360
rect 1219 1369 1287 1387
rect 1219 1353 1253 1369
rect 1117 1335 1253 1353
rect 1117 1325 1287 1335
rect 1151 1319 1287 1325
rect 1151 1291 1185 1319
rect 1117 1285 1185 1291
rect 1219 1300 1287 1319
rect 1219 1285 1253 1300
rect 1117 1266 1253 1285
rect 1117 1256 1287 1266
rect 1151 1251 1287 1256
rect 1151 1222 1185 1251
rect 1117 1217 1185 1222
rect 1219 1231 1287 1251
rect 1219 1217 1253 1231
rect 1117 1197 1253 1217
rect 1117 1187 1287 1197
rect 1151 1183 1287 1187
rect 1151 1153 1185 1183
rect 1117 1149 1185 1153
rect 1219 1162 1287 1183
rect 1219 1149 1253 1162
rect 1117 1128 1253 1149
rect 1117 1118 1287 1128
rect 1151 1115 1287 1118
rect 1151 1084 1185 1115
rect 1117 1081 1185 1084
rect 1219 1093 1287 1115
rect 1219 1081 1253 1093
rect 1117 1059 1253 1081
rect 1117 1049 1287 1059
rect 1151 1047 1287 1049
rect 1151 1015 1185 1047
rect 1117 1013 1185 1015
rect 1219 1024 1287 1047
rect 1219 1013 1253 1024
rect 1117 990 1253 1013
rect 1117 980 1287 990
rect 1151 979 1287 980
rect 1151 946 1185 979
rect 1117 945 1185 946
rect 1219 955 1287 979
rect 9929 1863 9963 1897
rect 9929 1795 9963 1829
rect 1219 945 1253 955
rect 1117 921 1253 945
rect 1117 911 1287 921
rect 1151 877 1185 911
rect 1219 886 1287 911
rect 1219 877 1253 886
rect 1117 852 1253 877
rect 1117 843 1287 852
rect 1117 842 1185 843
rect 1151 809 1185 842
rect 1219 817 1287 843
rect 1219 809 1253 817
rect 1151 808 1253 809
rect 1117 783 1253 808
rect 1117 775 1287 783
rect 1117 773 1185 775
rect 1151 741 1185 773
rect 1219 748 1287 775
rect 1219 741 1253 748
rect 1151 739 1253 741
rect 1117 714 1253 739
rect 1117 707 1287 714
rect 1117 704 1185 707
rect 1151 673 1185 704
rect 1219 679 1287 707
rect 1219 673 1253 679
rect 1151 670 1253 673
rect 1117 645 1253 670
rect 1117 639 1287 645
rect 1117 635 1185 639
rect 1151 605 1185 635
rect 1219 610 1287 639
rect 1219 605 1253 610
rect 1151 601 1253 605
rect 1117 576 1253 601
rect 9929 1727 9963 1761
rect 9929 1659 9963 1693
rect 9929 1591 9963 1625
rect 9929 1523 9963 1557
rect 9929 1455 9963 1489
rect 9929 1387 9963 1421
rect 9929 1319 9963 1353
rect 9929 1251 9963 1285
rect 9929 1183 9963 1217
rect 9929 1115 9963 1149
rect 9929 1047 9963 1081
rect 9929 979 9963 1013
rect 1117 571 1287 576
rect 1117 566 1185 571
rect 1151 537 1185 566
rect 1219 541 1287 571
rect 1219 537 1253 541
rect 1151 532 1253 537
rect 1117 507 1253 532
rect 1117 503 1287 507
rect 1117 497 1185 503
rect 1151 469 1185 497
rect 1219 472 1287 503
rect 1219 469 1253 472
rect 1151 463 1253 469
rect 1117 438 1253 463
rect 9929 911 9963 945
rect 9929 843 9963 877
rect 9929 775 9963 809
rect 9929 707 9963 741
rect 9929 639 9963 673
rect 9929 571 9963 605
rect 9929 503 9963 537
rect 1117 435 1287 438
rect 1117 428 1185 435
rect 1151 401 1185 428
rect 1219 403 1287 435
rect 1219 401 1253 403
rect 1151 394 1253 401
rect 1117 369 1253 394
rect 1117 367 1287 369
rect 1117 359 1185 367
rect 1151 333 1185 359
rect 1219 334 1287 367
rect 1219 333 1253 334
rect 1151 325 1253 333
rect 1117 300 1253 325
rect 1117 299 1287 300
rect 1117 290 1185 299
rect 1151 265 1185 290
rect 1219 265 1287 299
rect 1151 256 1253 265
rect 1117 231 1253 256
rect 1117 221 1185 231
rect 1151 197 1185 221
rect 1219 197 1287 231
rect 9929 435 9963 469
rect 13069 7666 13103 7700
rect 13069 7598 13103 7632
rect 13069 7530 13103 7564
rect 13069 7462 13103 7496
rect 13069 7394 13103 7428
rect 13069 7326 13103 7360
rect 13069 7258 13103 7292
rect 13069 7190 13103 7224
rect 13069 7122 13103 7156
rect 13069 7054 13103 7088
rect 13069 6986 13103 7020
rect 13069 6918 13103 6952
rect 13069 6850 13103 6884
rect 13069 6782 13103 6816
rect 13069 6714 13103 6748
rect 13069 6646 13103 6680
rect 13069 6578 13103 6612
rect 13069 6510 13103 6544
rect 13069 6442 13103 6476
rect 13069 6374 13103 6408
rect 13069 6306 13103 6340
rect 13069 6238 13103 6272
rect 13069 6170 13103 6204
rect 13069 6102 13103 6136
rect 13069 6034 13103 6068
rect 13069 5966 13103 6000
rect 13069 5898 13103 5932
rect 13069 5830 13103 5864
rect 13069 5762 13103 5796
rect 13069 5694 13103 5728
rect 13069 5626 13103 5660
rect 13069 5558 13103 5592
rect 13069 5490 13103 5524
rect 13069 5422 13103 5456
rect 13069 5354 13103 5388
rect 13069 5286 13103 5320
rect 13069 5218 13103 5252
rect 13069 5150 13103 5184
rect 13069 5082 13103 5116
rect 13069 5014 13103 5048
rect 13069 4946 13103 4980
rect 13069 4878 13103 4912
rect 13069 4810 13103 4844
rect 13069 4742 13103 4776
rect 13069 4674 13103 4708
rect 13069 4606 13103 4640
rect 13069 4538 13103 4572
rect 13069 4470 13103 4504
rect 13069 4402 13103 4436
rect 13069 4334 13103 4368
rect 13069 4266 13103 4300
rect 13069 4198 13103 4232
rect 13069 4130 13103 4164
rect 13069 4062 13103 4096
rect 13069 3994 13103 4028
rect 13069 3926 13103 3960
rect 13069 3858 13103 3892
rect 13069 3790 13103 3824
rect 13069 3722 13103 3756
rect 13069 3654 13103 3688
rect 13069 3586 13103 3620
rect 13069 3518 13103 3552
rect 13069 3450 13103 3484
rect 13069 3382 13103 3416
rect 13069 3314 13103 3348
rect 13069 3246 13103 3280
rect 13069 3178 13103 3212
rect 13069 3110 13103 3144
rect 13069 3042 13103 3076
rect 13069 2974 13103 3008
rect 13069 2906 13103 2940
rect 13069 2838 13103 2872
rect 13069 2770 13103 2804
rect 13069 2702 13103 2736
rect 13069 2634 13103 2668
rect 13069 2566 13103 2600
rect 13069 2498 13103 2532
rect 13069 2430 13103 2464
rect 13069 2362 13103 2396
rect 13069 2294 13103 2328
rect 13069 2226 13103 2260
rect 13069 2158 13103 2192
rect 13069 2090 13103 2124
rect 13069 2022 13103 2056
rect 13069 1954 13103 1988
rect 13069 1886 13103 1920
rect 13069 1818 13103 1852
rect 13069 1750 13103 1784
rect 13069 1682 13103 1716
rect 13069 1614 13103 1648
rect 13069 1546 13103 1580
rect 13069 1478 13103 1512
rect 13069 1410 13103 1444
rect 13069 1342 13103 1376
rect 13069 1274 13103 1308
rect 13069 1206 13103 1240
rect 13069 1138 13103 1172
rect 13069 1070 13103 1104
rect 13069 1002 13103 1036
rect 13069 934 13103 968
rect 13069 866 13103 900
rect 13069 798 13103 832
rect 13069 730 13103 764
rect 13069 662 13103 696
rect 13069 594 13103 628
rect 13069 526 13103 560
rect 13069 458 13103 492
rect 9929 367 9963 401
rect 9929 299 9963 333
rect 9929 231 9963 265
rect 13069 390 13103 424
rect 13069 322 13103 356
rect 1151 187 1282 197
rect 1117 163 1282 187
rect 1316 163 1350 197
rect 1384 163 1418 197
rect 1452 163 1486 197
rect 1520 163 1554 197
rect 1588 163 1622 197
rect 1656 163 1690 197
rect 1724 163 1758 197
rect 1792 163 1826 197
rect 1860 163 1894 197
rect 1928 163 1962 197
rect 1996 163 2030 197
rect 2064 163 2098 197
rect 2132 163 2166 197
rect 2200 163 2234 197
rect 2268 163 2302 197
rect 2336 163 2370 197
rect 2404 163 2438 197
rect 2472 163 2506 197
rect 2540 163 2574 197
rect 2608 163 2642 197
rect 2676 163 2710 197
rect 2744 163 2778 197
rect 2812 163 2846 197
rect 2880 163 2914 197
rect 2948 163 2982 197
rect 3016 163 3050 197
rect 3084 163 3118 197
rect 3152 163 3186 197
rect 3220 163 3254 197
rect 3288 163 3322 197
rect 3356 163 3390 197
rect 3424 163 3458 197
rect 3492 163 3526 197
rect 3560 163 3594 197
rect 3628 163 3662 197
rect 3696 163 3730 197
rect 3764 163 3798 197
rect 3832 163 3866 197
rect 3900 163 3934 197
rect 3968 163 4002 197
rect 4036 163 4070 197
rect 4104 163 4138 197
rect 4172 163 4206 197
rect 4240 163 4274 197
rect 4308 163 4342 197
rect 4376 163 4410 197
rect 4444 163 4478 197
rect 4512 163 4546 197
rect 4580 163 4614 197
rect 4648 163 4682 197
rect 4716 163 4750 197
rect 4784 163 4818 197
rect 4852 163 4886 197
rect 4920 163 4954 197
rect 4988 163 5022 197
rect 5056 163 5090 197
rect 5124 163 5158 197
rect 5192 163 5226 197
rect 5260 163 5294 197
rect 5328 163 5362 197
rect 5396 163 5430 197
rect 5464 163 5498 197
rect 5532 163 5566 197
rect 5600 163 5668 197
rect 5702 163 5736 197
rect 5770 163 5804 197
rect 5838 163 5872 197
rect 5906 163 5940 197
rect 5974 163 6008 197
rect 6042 163 6076 197
rect 6110 163 6144 197
rect 6178 163 6212 197
rect 6246 163 6280 197
rect 6314 163 6348 197
rect 6382 163 6416 197
rect 6450 163 6484 197
rect 6518 163 6552 197
rect 6586 163 6620 197
rect 6654 163 6688 197
rect 6722 163 6756 197
rect 6790 163 6824 197
rect 6858 163 6892 197
rect 6926 163 6960 197
rect 6994 163 7028 197
rect 7062 163 7096 197
rect 7130 163 7164 197
rect 7198 163 7232 197
rect 7266 163 7300 197
rect 7334 163 7368 197
rect 7402 163 7436 197
rect 7470 163 7504 197
rect 7538 163 7572 197
rect 7606 163 7640 197
rect 7674 163 7708 197
rect 7742 163 7776 197
rect 7810 163 7844 197
rect 7878 163 7912 197
rect 7946 163 7980 197
rect 8014 163 8048 197
rect 8082 163 8116 197
rect 8150 163 8184 197
rect 8218 163 8252 197
rect 8286 163 8320 197
rect 8354 163 8388 197
rect 8422 163 8456 197
rect 8490 163 8524 197
rect 8558 163 8592 197
rect 8626 163 8660 197
rect 8694 163 8728 197
rect 8762 163 8796 197
rect 8830 163 8864 197
rect 8898 163 8932 197
rect 8966 163 9000 197
rect 9034 163 9068 197
rect 9102 163 9136 197
rect 9170 163 9204 197
rect 9238 163 9272 197
rect 9306 163 9340 197
rect 9374 163 9408 197
rect 9442 163 9476 197
rect 9510 163 9544 197
rect 9578 163 9612 197
rect 9646 163 9680 197
rect 9714 163 9748 197
rect 9782 163 9816 197
rect 9850 163 10043 197
rect 10077 163 10111 197
rect 10145 163 10179 197
rect 10213 163 10247 197
rect 10281 163 10315 197
rect 10349 163 10383 197
rect 10417 163 10451 197
rect 10485 163 10519 197
rect 10553 163 10587 197
rect 10621 163 10655 197
rect 10689 163 10723 197
rect 10757 163 10791 197
rect 10825 163 10859 197
rect 10893 163 10927 197
rect 10961 163 10995 197
rect 11029 163 11063 197
rect 11097 163 11131 197
rect 11165 163 11199 197
rect 11233 163 11267 197
rect 11301 163 11335 197
rect 11369 163 11403 197
rect 11437 163 11471 197
rect 11505 163 11539 197
rect 11573 163 11607 197
rect 11641 163 11675 197
rect 11709 163 11743 197
rect 11777 163 11811 197
rect 11845 163 11879 197
rect 11913 163 11947 197
rect 11981 163 12015 197
rect 12049 163 12083 197
rect 12117 163 12151 197
rect 12185 163 12219 197
rect 12253 163 12287 197
rect 12321 163 12355 197
rect 12389 163 12423 197
rect 12457 163 12491 197
rect 12525 163 12559 197
rect 12593 163 12627 197
rect 12661 163 12695 197
rect 12729 163 12763 197
rect 12797 163 12831 197
rect 12865 163 12899 197
rect 12933 163 12967 197
rect 13001 163 13035 197
rect 13069 163 13103 288
<< psubdiffcont >>
rect 1492 11387 1526 11421
rect 1561 11387 1595 11421
rect 1630 11387 1664 11421
rect 1699 11387 1733 11421
rect 1768 11387 1802 11421
rect 1837 11387 1871 11421
rect 1906 11387 1940 11421
rect 1975 11387 2009 11421
rect 2044 11387 2078 11421
rect 2113 11387 2147 11421
rect 2182 11387 2216 11421
rect 2251 11387 2285 11421
rect 2320 11387 2354 11421
rect 2389 11387 2423 11421
rect 2458 11387 2492 11421
rect 2526 11387 2560 11421
rect 2594 11387 2628 11421
rect 2662 11387 2696 11421
rect 2730 11387 2764 11421
rect 2798 11387 2832 11421
rect 2866 11387 2900 11421
rect 2934 11387 2968 11421
rect 3002 11387 3036 11421
rect 3070 11387 3104 11421
rect 3138 11387 3172 11421
rect 3206 11387 3240 11421
rect 3274 11387 3308 11421
rect 3342 11387 3376 11421
rect 3410 11387 3444 11421
rect 1492 7231 1526 7265
rect 1561 7231 1595 7265
rect 1630 7231 1664 7265
rect 1699 7231 1733 7265
rect 1768 7231 1802 7265
rect 1837 7231 1871 7265
rect 1906 7231 1940 7265
rect 1975 7231 2009 7265
rect 2044 7231 2078 7265
rect 2113 7231 2147 7265
rect 2182 7231 2216 7265
rect 2251 7231 2285 7265
rect 2320 7231 2354 7265
rect 2389 7231 2423 7265
rect 2458 7231 2492 7265
rect 2526 7231 2560 7265
rect 2594 7231 2628 7265
rect 2662 7231 2696 7265
rect 2730 7231 2764 7265
rect 2798 7231 2832 7265
rect 2866 7231 2900 7265
rect 2934 7231 2968 7265
rect 3002 7231 3036 7265
rect 3070 7231 3104 7265
rect 3138 7231 3172 7265
rect 3206 7231 3240 7265
rect 3274 7231 3308 7265
rect 3342 7231 3376 7265
rect 3410 7231 3444 7265
rect 1492 6627 1526 6661
rect 1561 6627 1595 6661
rect 1630 6627 1664 6661
rect 1699 6627 1733 6661
rect 1768 6627 1802 6661
rect 1837 6627 1871 6661
rect 1906 6627 1940 6661
rect 1975 6627 2009 6661
rect 2044 6627 2078 6661
rect 2113 6627 2147 6661
rect 2182 6627 2216 6661
rect 2251 6627 2285 6661
rect 2320 6627 2354 6661
rect 2389 6627 2423 6661
rect 2458 6627 2492 6661
rect 2526 6627 2560 6661
rect 2594 6627 2628 6661
rect 2662 6627 2696 6661
rect 2730 6627 2764 6661
rect 2798 6627 2832 6661
rect 2866 6627 2900 6661
rect 2934 6627 2968 6661
rect 3002 6627 3036 6661
rect 3070 6627 3104 6661
rect 3138 6627 3172 6661
rect 3206 6627 3240 6661
rect 3274 6627 3308 6661
rect 3342 6627 3376 6661
rect 3410 6627 3444 6661
rect 7704 11387 7738 11421
rect 7772 11387 7806 11421
rect 7840 11387 7874 11421
rect 7908 11387 7942 11421
rect 7976 11387 8010 11421
rect 8044 11387 8078 11421
rect 8112 11387 8146 11421
rect 8180 11387 8214 11421
rect 8248 11387 8282 11421
rect 8316 11387 8350 11421
rect 8384 11387 8418 11421
rect 8452 11387 8486 11421
rect 8520 11387 8554 11421
rect 8588 11387 8622 11421
rect 8656 11387 8690 11421
rect 8725 11387 8759 11421
rect 8794 11387 8828 11421
rect 8863 11387 8897 11421
rect 8932 11387 8966 11421
rect 9001 11387 9035 11421
rect 9070 11387 9104 11421
rect 9139 11387 9173 11421
rect 9208 11387 9242 11421
rect 9277 11387 9311 11421
rect 9346 11387 9380 11421
rect 9415 11387 9449 11421
rect 9484 11387 9518 11421
rect 9553 11387 9587 11421
rect 9622 11387 9656 11421
rect 7704 7231 7738 7265
rect 7772 7231 7806 7265
rect 7840 7231 7874 7265
rect 7908 7231 7942 7265
rect 7976 7231 8010 7265
rect 8044 7231 8078 7265
rect 8112 7231 8146 7265
rect 8180 7231 8214 7265
rect 8248 7231 8282 7265
rect 8316 7231 8350 7265
rect 8384 7231 8418 7265
rect 8452 7231 8486 7265
rect 8520 7231 8554 7265
rect 8588 7231 8622 7265
rect 8656 7231 8690 7265
rect 8725 7231 8759 7265
rect 8794 7231 8828 7265
rect 8863 7231 8897 7265
rect 8932 7231 8966 7265
rect 9001 7231 9035 7265
rect 9070 7231 9104 7265
rect 9139 7231 9173 7265
rect 9208 7231 9242 7265
rect 9277 7231 9311 7265
rect 9346 7231 9380 7265
rect 9415 7231 9449 7265
rect 9484 7231 9518 7265
rect 9553 7231 9587 7265
rect 9622 7231 9656 7265
rect 7704 6627 7738 6661
rect 7772 6627 7806 6661
rect 7840 6627 7874 6661
rect 7908 6627 7942 6661
rect 7976 6627 8010 6661
rect 8044 6627 8078 6661
rect 8112 6627 8146 6661
rect 8180 6627 8214 6661
rect 8248 6627 8282 6661
rect 8316 6627 8350 6661
rect 8384 6627 8418 6661
rect 8452 6627 8486 6661
rect 8520 6627 8554 6661
rect 8588 6627 8622 6661
rect 8656 6627 8690 6661
rect 8725 6627 8759 6661
rect 8794 6627 8828 6661
rect 8863 6627 8897 6661
rect 8932 6627 8966 6661
rect 9001 6627 9035 6661
rect 9070 6627 9104 6661
rect 9139 6627 9173 6661
rect 9208 6627 9242 6661
rect 9277 6627 9311 6661
rect 9346 6627 9380 6661
rect 9415 6627 9449 6661
rect 9484 6627 9518 6661
rect 9553 6627 9587 6661
rect 9622 6627 9656 6661
rect 1492 2471 1526 2505
rect 1561 2471 1595 2505
rect 1630 2471 1664 2505
rect 1699 2471 1733 2505
rect 1768 2471 1802 2505
rect 1837 2471 1871 2505
rect 1906 2471 1940 2505
rect 1975 2471 2009 2505
rect 2044 2471 2078 2505
rect 2113 2471 2147 2505
rect 2182 2471 2216 2505
rect 2251 2471 2285 2505
rect 2320 2471 2354 2505
rect 2389 2471 2423 2505
rect 2458 2471 2492 2505
rect 2526 2471 2560 2505
rect 2594 2471 2628 2505
rect 2662 2471 2696 2505
rect 2730 2471 2764 2505
rect 2798 2471 2832 2505
rect 2866 2471 2900 2505
rect 2934 2471 2968 2505
rect 3002 2471 3036 2505
rect 3070 2471 3104 2505
rect 3138 2471 3172 2505
rect 3206 2471 3240 2505
rect 3274 2471 3308 2505
rect 3342 2471 3376 2505
rect 3410 2471 3444 2505
rect 7704 2471 7738 2505
rect 7772 2471 7806 2505
rect 7840 2471 7874 2505
rect 7908 2471 7942 2505
rect 7976 2471 8010 2505
rect 8044 2471 8078 2505
rect 8112 2471 8146 2505
rect 8180 2471 8214 2505
rect 8248 2471 8282 2505
rect 8316 2471 8350 2505
rect 8384 2471 8418 2505
rect 8452 2471 8486 2505
rect 8520 2471 8554 2505
rect 8588 2471 8622 2505
rect 8656 2471 8690 2505
rect 8725 2471 8759 2505
rect 8794 2471 8828 2505
rect 8863 2471 8897 2505
rect 8932 2471 8966 2505
rect 9001 2471 9035 2505
rect 9070 2471 9104 2505
rect 9139 2471 9173 2505
rect 9208 2471 9242 2505
rect 9277 2471 9311 2505
rect 9346 2471 9380 2505
rect 9415 2471 9449 2505
rect 9484 2471 9518 2505
rect 9553 2471 9587 2505
rect 9622 2471 9656 2505
<< mvpsubdiffcont >>
rect 1228 12137 1262 12171
rect 1297 12137 1331 12171
rect 1366 12137 1400 12171
rect 1435 12137 1469 12171
rect 1504 12137 1538 12171
rect 1573 12137 1607 12171
rect 1642 12137 1676 12171
rect 1711 12137 1745 12171
rect 1780 12137 1814 12171
rect 1849 12137 1883 12171
rect 1918 12137 1952 12171
rect 1987 12137 2021 12171
rect 2056 12137 2090 12171
rect 2125 12137 2159 12171
rect 2194 12137 2228 12171
rect 2263 12137 2297 12171
rect 2332 12137 2366 12171
rect 2401 12137 2435 12171
rect 2470 12137 2504 12171
rect 2539 12137 2573 12171
rect 2608 12137 2642 12171
rect 2677 12137 2711 12171
rect 2746 12137 2780 12171
rect 2815 12137 2849 12171
rect 2884 12137 2918 12171
rect 2953 12137 2987 12171
rect 3022 12137 3056 12171
rect 3091 12137 3125 12171
rect 3160 12137 3194 12171
rect 3229 12137 3263 12171
rect 3298 12137 3332 12171
rect 3367 12137 3401 12171
rect 3436 12137 3470 12171
rect 3505 12137 3539 12171
rect 3574 12137 3608 12171
rect 3643 12137 3677 12171
rect 3712 12137 3746 12171
rect 3781 12137 3815 12171
rect 3850 12137 3884 12171
rect 3919 12137 3953 12171
rect 1228 12069 1262 12103
rect 1297 12069 1331 12103
rect 1366 12069 1400 12103
rect 1435 12069 1469 12103
rect 1504 12069 1538 12103
rect 1573 12069 1607 12103
rect 1642 12069 1676 12103
rect 1711 12069 1745 12103
rect 1780 12069 1814 12103
rect 1849 12069 1883 12103
rect 1918 12069 1952 12103
rect 1987 12069 2021 12103
rect 2056 12069 2090 12103
rect 2125 12069 2159 12103
rect 2194 12069 2228 12103
rect 2263 12069 2297 12103
rect 2332 12069 2366 12103
rect 2401 12069 2435 12103
rect 2470 12069 2504 12103
rect 2539 12069 2573 12103
rect 2608 12069 2642 12103
rect 2677 12069 2711 12103
rect 2746 12069 2780 12103
rect 2815 12069 2849 12103
rect 2884 12069 2918 12103
rect 2953 12069 2987 12103
rect 3022 12069 3056 12103
rect 3091 12069 3125 12103
rect 3160 12069 3194 12103
rect 3229 12069 3263 12103
rect 3298 12069 3332 12103
rect 3367 12069 3401 12103
rect 3436 12069 3470 12103
rect 3505 12069 3539 12103
rect 3574 12069 3608 12103
rect 3643 12069 3677 12103
rect 3712 12069 3746 12103
rect 3781 12069 3815 12103
rect 3850 12069 3884 12103
rect 3919 12069 3953 12103
rect 1228 12001 1262 12035
rect 1297 12001 1331 12035
rect 1366 12001 1400 12035
rect 1435 12001 1469 12035
rect 1504 12001 1538 12035
rect 1573 12001 1607 12035
rect 1642 12001 1676 12035
rect 1711 12001 1745 12035
rect 1780 12001 1814 12035
rect 1849 12001 1883 12035
rect 1918 12001 1952 12035
rect 1987 12001 2021 12035
rect 2056 12001 2090 12035
rect 2125 12001 2159 12035
rect 2194 12001 2228 12035
rect 2263 12001 2297 12035
rect 2332 12001 2366 12035
rect 2401 12001 2435 12035
rect 2470 12001 2504 12035
rect 2539 12001 2573 12035
rect 2608 12001 2642 12035
rect 2677 12001 2711 12035
rect 2746 12001 2780 12035
rect 2815 12001 2849 12035
rect 2884 12001 2918 12035
rect 2953 12001 2987 12035
rect 3022 12001 3056 12035
rect 3091 12001 3125 12035
rect 3160 12001 3194 12035
rect 3229 12001 3263 12035
rect 3298 12001 3332 12035
rect 3367 12001 3401 12035
rect 3436 12001 3470 12035
rect 3505 12001 3539 12035
rect 3574 12001 3608 12035
rect 3643 12001 3677 12035
rect 3712 12001 3746 12035
rect 3781 12001 3815 12035
rect 3850 12001 3884 12035
rect 3919 12001 3953 12035
rect 3988 12001 11094 12171
rect 4034 11328 4068 11362
rect 4102 11328 4136 11362
rect 4170 11328 4204 11362
rect 4238 11328 4272 11362
rect 4306 11328 4340 11362
rect 4374 11328 4408 11362
rect 4442 11328 4476 11362
rect 4510 11328 4544 11362
rect 4578 11328 4612 11362
rect 4646 11328 4680 11362
rect 4714 11328 4748 11362
rect 4782 11328 4816 11362
rect 4850 11328 4884 11362
rect 4918 11328 4952 11362
rect 4986 11328 5020 11362
rect 5054 11328 5088 11362
rect 5122 11328 5156 11362
rect 5190 11328 5224 11362
rect 4000 11205 4034 11239
rect 5274 11205 5308 11239
rect 4000 11136 4034 11170
rect 5274 11136 5308 11170
rect 4000 11067 4034 11101
rect 5274 11067 5308 11101
rect 4000 10998 4034 11032
rect 4000 10929 4034 10963
rect 4000 10860 4034 10894
rect 4000 10791 4034 10825
rect 4000 10722 4034 10756
rect 4000 10653 4034 10687
rect 4000 10584 4034 10618
rect 4000 10515 4034 10549
rect 4000 10446 4034 10480
rect 4000 10377 4034 10411
rect 4000 10308 4034 10342
rect 4000 10239 4034 10273
rect 5274 10998 5308 11032
rect 5274 10929 5308 10963
rect 5274 10860 5308 10894
rect 5274 10791 5308 10825
rect 5274 10722 5308 10756
rect 5274 10653 5308 10687
rect 5274 10584 5308 10618
rect 5274 10515 5308 10549
rect 5274 10446 5308 10480
rect 5274 10377 5308 10411
rect 5274 10308 5308 10342
rect 4000 10170 4034 10204
rect 5274 10239 5308 10273
rect 4000 10101 4034 10135
rect 4000 10032 4034 10066
rect 4000 9963 4034 9997
rect 4000 9894 4034 9928
rect 4000 9825 4034 9859
rect 4000 9756 4034 9790
rect 4000 9687 4034 9721
rect 4000 9618 4034 9652
rect 4000 9549 4034 9583
rect 4000 9480 4034 9514
rect 4000 9411 4034 9445
rect 5274 10170 5308 10204
rect 5274 10101 5308 10135
rect 5274 10032 5308 10066
rect 5274 9963 5308 9997
rect 5274 9894 5308 9928
rect 5274 9825 5308 9859
rect 5274 9756 5308 9790
rect 5274 9687 5308 9721
rect 5274 9618 5308 9652
rect 5274 9549 5308 9583
rect 5274 9480 5308 9514
rect 5274 9411 5308 9445
rect 4000 9342 4034 9376
rect 5274 9342 5308 9376
rect 4000 9273 4034 9307
rect 4000 9204 4034 9238
rect 4000 9135 4034 9169
rect 4000 9066 4034 9100
rect 4000 8997 4034 9031
rect 4000 8928 4034 8962
rect 4000 8859 4034 8893
rect 4000 8790 4034 8824
rect 4000 8721 4034 8755
rect 4000 8652 4034 8686
rect 4000 8583 4034 8617
rect 4000 8514 4034 8548
rect 5274 9273 5308 9307
rect 5274 9204 5308 9238
rect 5274 9135 5308 9169
rect 5274 9066 5308 9100
rect 5274 8997 5308 9031
rect 5274 8928 5308 8962
rect 5274 8859 5308 8893
rect 5274 8790 5308 8824
rect 5274 8721 5308 8755
rect 5274 8652 5308 8686
rect 5274 8583 5308 8617
rect 4000 8445 4034 8479
rect 5274 8514 5308 8548
rect 4000 8376 4034 8410
rect 4000 8307 4034 8341
rect 4000 8238 4034 8272
rect 4000 8169 4034 8203
rect 4000 8100 4034 8134
rect 4000 8031 4034 8065
rect 4000 7962 4034 7996
rect 4000 7893 4034 7927
rect 4000 7824 4034 7858
rect 4000 7755 4034 7789
rect 4000 7686 4034 7720
rect 5274 8445 5308 8479
rect 5274 8376 5308 8410
rect 5274 8307 5308 8341
rect 5274 8238 5308 8272
rect 5274 8169 5308 8203
rect 5274 8100 5308 8134
rect 5274 8031 5308 8065
rect 5274 7962 5308 7996
rect 5274 7893 5308 7927
rect 5274 7824 5308 7858
rect 5274 7755 5308 7789
rect 5274 7686 5308 7720
rect 4000 7617 4034 7651
rect 4000 7549 4034 7583
rect 4000 7481 4034 7515
rect 4000 7413 4034 7447
rect 4000 7345 4034 7379
rect 4000 7277 4034 7311
rect 4000 7209 4034 7243
rect 4000 7141 4034 7175
rect 4000 7073 4034 7107
rect 4000 7005 4034 7039
rect 4000 6937 4034 6971
rect 4000 6869 4034 6903
rect 4000 6801 4034 6835
rect 5274 7617 5308 7651
rect 5274 7549 5308 7583
rect 5274 7481 5308 7515
rect 5274 7413 5308 7447
rect 5274 7345 5308 7379
rect 5274 7277 5308 7311
rect 5274 7209 5308 7243
rect 5274 7141 5308 7175
rect 5274 7073 5308 7107
rect 5274 7005 5308 7039
rect 5274 6937 5308 6971
rect 5274 6869 5308 6903
rect 4000 6733 4034 6767
rect 5274 6801 5308 6835
rect 4000 6665 4034 6699
rect 4000 6597 4034 6631
rect 4000 6529 4034 6563
rect 4000 6461 4034 6495
rect 4000 6393 4034 6427
rect 4000 6325 4034 6359
rect 4000 6257 4034 6291
rect 4000 6189 4034 6223
rect 4000 6121 4034 6155
rect 4000 6053 4034 6087
rect 4000 5985 4034 6019
rect 5274 6733 5308 6767
rect 5274 6665 5308 6699
rect 5274 6597 5308 6631
rect 5274 6529 5308 6563
rect 5274 6461 5308 6495
rect 5274 6393 5308 6427
rect 5274 6325 5308 6359
rect 5274 6257 5308 6291
rect 5274 6189 5308 6223
rect 5274 6121 5308 6155
rect 5274 6053 5308 6087
rect 5274 5985 5308 6019
rect 4000 5917 4034 5951
rect 5274 5917 5308 5951
rect 4000 5849 4034 5883
rect 4000 5781 4034 5815
rect 4000 5713 4034 5747
rect 4000 5645 4034 5679
rect 4000 5577 4034 5611
rect 4000 5509 4034 5543
rect 4000 5441 4034 5475
rect 4000 5373 4034 5407
rect 4000 5305 4034 5339
rect 4000 5237 4034 5271
rect 4000 5169 4034 5203
rect 4000 5101 4034 5135
rect 5274 5849 5308 5883
rect 5274 5781 5308 5815
rect 5274 5713 5308 5747
rect 5274 5645 5308 5679
rect 5274 5577 5308 5611
rect 5274 5509 5308 5543
rect 5274 5441 5308 5475
rect 5274 5373 5308 5407
rect 5274 5305 5308 5339
rect 5274 5237 5308 5271
rect 5274 5169 5308 5203
rect 4000 5033 4034 5067
rect 5274 5101 5308 5135
rect 4000 4965 4034 4999
rect 4000 4897 4034 4931
rect 4000 4829 4034 4863
rect 4000 4761 4034 4795
rect 4000 4693 4034 4727
rect 4000 4625 4034 4659
rect 4000 4557 4034 4591
rect 4000 4489 4034 4523
rect 4000 4421 4034 4455
rect 4000 4353 4034 4387
rect 4000 4285 4034 4319
rect 5274 5033 5308 5067
rect 5274 4965 5308 4999
rect 5274 4897 5308 4931
rect 5274 4829 5308 4863
rect 5274 4761 5308 4795
rect 5274 4693 5308 4727
rect 5274 4625 5308 4659
rect 5274 4557 5308 4591
rect 5274 4489 5308 4523
rect 5274 4421 5308 4455
rect 5274 4353 5308 4387
rect 5274 4285 5308 4319
rect 4000 4217 4034 4251
rect 5274 4217 5308 4251
rect 4000 4149 4034 4183
rect 4000 4081 4034 4115
rect 5274 4149 5308 4183
rect 5274 4081 5308 4115
rect 5274 3970 5308 4004
rect 4034 3936 4068 3970
rect 4102 3936 4136 3970
rect 4170 3936 4204 3970
rect 4238 3936 4272 3970
rect 4306 3936 4340 3970
rect 4374 3936 4408 3970
rect 4442 3936 4476 3970
rect 4510 3936 4544 3970
rect 4578 3936 4612 3970
rect 4646 3936 4680 3970
rect 4714 3936 4748 3970
rect 4782 3936 4816 3970
rect 4850 3936 4884 3970
rect 4918 3936 4952 3970
rect 4986 3936 5020 3970
rect 5054 3936 5088 3970
rect 5122 3936 5156 3970
rect 5190 3936 5224 3970
rect 5874 11328 5908 11362
rect 5942 11328 5976 11362
rect 6010 11328 6044 11362
rect 6078 11328 6112 11362
rect 6146 11328 6180 11362
rect 6214 11328 6248 11362
rect 6282 11328 6316 11362
rect 6350 11328 6384 11362
rect 6418 11328 6452 11362
rect 6486 11328 6520 11362
rect 6554 11328 6588 11362
rect 6622 11328 6656 11362
rect 6690 11328 6724 11362
rect 6758 11328 6792 11362
rect 6826 11328 6860 11362
rect 6894 11328 6928 11362
rect 6962 11328 6996 11362
rect 7030 11328 7064 11362
rect 5840 11205 5874 11239
rect 7114 11205 7148 11239
rect 5840 11136 5874 11170
rect 7114 11136 7148 11170
rect 5840 11067 5874 11101
rect 7114 11067 7148 11101
rect 5840 10998 5874 11032
rect 5840 10929 5874 10963
rect 5840 10860 5874 10894
rect 5840 10791 5874 10825
rect 5840 10722 5874 10756
rect 5840 10653 5874 10687
rect 5840 10584 5874 10618
rect 5840 10515 5874 10549
rect 5840 10446 5874 10480
rect 5840 10377 5874 10411
rect 5840 10308 5874 10342
rect 5840 10239 5874 10273
rect 7114 10998 7148 11032
rect 7114 10929 7148 10963
rect 7114 10860 7148 10894
rect 7114 10791 7148 10825
rect 7114 10722 7148 10756
rect 7114 10653 7148 10687
rect 7114 10584 7148 10618
rect 7114 10515 7148 10549
rect 7114 10446 7148 10480
rect 7114 10377 7148 10411
rect 7114 10308 7148 10342
rect 5840 10170 5874 10204
rect 7114 10239 7148 10273
rect 5840 10101 5874 10135
rect 5840 10032 5874 10066
rect 5840 9963 5874 9997
rect 5840 9894 5874 9928
rect 5840 9825 5874 9859
rect 5840 9756 5874 9790
rect 5840 9687 5874 9721
rect 5840 9618 5874 9652
rect 5840 9549 5874 9583
rect 5840 9480 5874 9514
rect 5840 9411 5874 9445
rect 7114 10170 7148 10204
rect 7114 10101 7148 10135
rect 7114 10032 7148 10066
rect 7114 9963 7148 9997
rect 7114 9894 7148 9928
rect 7114 9825 7148 9859
rect 7114 9756 7148 9790
rect 7114 9687 7148 9721
rect 7114 9618 7148 9652
rect 7114 9549 7148 9583
rect 7114 9480 7148 9514
rect 7114 9411 7148 9445
rect 5840 9342 5874 9376
rect 7114 9342 7148 9376
rect 5840 9273 5874 9307
rect 5840 9204 5874 9238
rect 5840 9135 5874 9169
rect 5840 9066 5874 9100
rect 5840 8997 5874 9031
rect 5840 8928 5874 8962
rect 5840 8859 5874 8893
rect 5840 8790 5874 8824
rect 5840 8721 5874 8755
rect 5840 8652 5874 8686
rect 5840 8583 5874 8617
rect 5840 8514 5874 8548
rect 7114 9273 7148 9307
rect 7114 9204 7148 9238
rect 7114 9135 7148 9169
rect 7114 9066 7148 9100
rect 7114 8997 7148 9031
rect 7114 8928 7148 8962
rect 7114 8859 7148 8893
rect 7114 8790 7148 8824
rect 7114 8721 7148 8755
rect 7114 8652 7148 8686
rect 7114 8583 7148 8617
rect 5840 8445 5874 8479
rect 7114 8514 7148 8548
rect 5840 8376 5874 8410
rect 5840 8307 5874 8341
rect 5840 8238 5874 8272
rect 5840 8169 5874 8203
rect 5840 8100 5874 8134
rect 5840 8031 5874 8065
rect 5840 7962 5874 7996
rect 5840 7893 5874 7927
rect 5840 7824 5874 7858
rect 5840 7755 5874 7789
rect 5840 7686 5874 7720
rect 7114 8445 7148 8479
rect 7114 8376 7148 8410
rect 7114 8307 7148 8341
rect 7114 8238 7148 8272
rect 7114 8169 7148 8203
rect 7114 8100 7148 8134
rect 7114 8031 7148 8065
rect 7114 7962 7148 7996
rect 7114 7893 7148 7927
rect 7114 7824 7148 7858
rect 7114 7755 7148 7789
rect 7114 7686 7148 7720
rect 5840 7617 5874 7651
rect 5840 7549 5874 7583
rect 5840 7481 5874 7515
rect 5840 7413 5874 7447
rect 5840 7345 5874 7379
rect 5840 7277 5874 7311
rect 5840 7209 5874 7243
rect 5840 7141 5874 7175
rect 5840 7073 5874 7107
rect 5840 7005 5874 7039
rect 5840 6937 5874 6971
rect 5840 6869 5874 6903
rect 5840 6801 5874 6835
rect 7114 7617 7148 7651
rect 7114 7549 7148 7583
rect 7114 7481 7148 7515
rect 7114 7413 7148 7447
rect 7114 7345 7148 7379
rect 7114 7277 7148 7311
rect 7114 7209 7148 7243
rect 7114 7141 7148 7175
rect 7114 7073 7148 7107
rect 7114 7005 7148 7039
rect 7114 6937 7148 6971
rect 7114 6869 7148 6903
rect 5840 6733 5874 6767
rect 7114 6801 7148 6835
rect 5840 6665 5874 6699
rect 5840 6597 5874 6631
rect 5840 6529 5874 6563
rect 5840 6461 5874 6495
rect 5840 6393 5874 6427
rect 5840 6325 5874 6359
rect 5840 6257 5874 6291
rect 5840 6189 5874 6223
rect 5840 6121 5874 6155
rect 5840 6053 5874 6087
rect 5840 5985 5874 6019
rect 7114 6733 7148 6767
rect 7114 6665 7148 6699
rect 7114 6597 7148 6631
rect 7114 6529 7148 6563
rect 7114 6461 7148 6495
rect 7114 6393 7148 6427
rect 7114 6325 7148 6359
rect 7114 6257 7148 6291
rect 7114 6189 7148 6223
rect 7114 6121 7148 6155
rect 7114 6053 7148 6087
rect 7114 5985 7148 6019
rect 5840 5917 5874 5951
rect 7114 5917 7148 5951
rect 5840 5849 5874 5883
rect 5840 5781 5874 5815
rect 5840 5713 5874 5747
rect 5840 5645 5874 5679
rect 5840 5577 5874 5611
rect 5840 5509 5874 5543
rect 5840 5441 5874 5475
rect 5840 5373 5874 5407
rect 5840 5305 5874 5339
rect 5840 5237 5874 5271
rect 5840 5169 5874 5203
rect 5840 5101 5874 5135
rect 7114 5849 7148 5883
rect 7114 5781 7148 5815
rect 7114 5713 7148 5747
rect 7114 5645 7148 5679
rect 7114 5577 7148 5611
rect 7114 5509 7148 5543
rect 7114 5441 7148 5475
rect 7114 5373 7148 5407
rect 7114 5305 7148 5339
rect 7114 5237 7148 5271
rect 7114 5169 7148 5203
rect 5840 5033 5874 5067
rect 7114 5101 7148 5135
rect 5840 4965 5874 4999
rect 5840 4897 5874 4931
rect 5840 4829 5874 4863
rect 5840 4761 5874 4795
rect 5840 4693 5874 4727
rect 5840 4625 5874 4659
rect 5840 4557 5874 4591
rect 5840 4489 5874 4523
rect 5840 4421 5874 4455
rect 5840 4353 5874 4387
rect 5840 4285 5874 4319
rect 7114 5033 7148 5067
rect 7114 4965 7148 4999
rect 7114 4897 7148 4931
rect 7114 4829 7148 4863
rect 7114 4761 7148 4795
rect 7114 4693 7148 4727
rect 7114 4625 7148 4659
rect 7114 4557 7148 4591
rect 7114 4489 7148 4523
rect 7114 4421 7148 4455
rect 7114 4353 7148 4387
rect 7114 4285 7148 4319
rect 5840 4217 5874 4251
rect 7114 4217 7148 4251
rect 5840 4149 5874 4183
rect 5840 4081 5874 4115
rect 7114 4149 7148 4183
rect 7114 4081 7148 4115
rect 7114 3970 7148 4004
rect 5874 3936 5908 3970
rect 5942 3936 5976 3970
rect 6010 3936 6044 3970
rect 6078 3936 6112 3970
rect 6146 3936 6180 3970
rect 6214 3936 6248 3970
rect 6282 3936 6316 3970
rect 6350 3936 6384 3970
rect 6418 3936 6452 3970
rect 6486 3936 6520 3970
rect 6554 3936 6588 3970
rect 6622 3936 6656 3970
rect 6690 3936 6724 3970
rect 6758 3936 6792 3970
rect 6826 3936 6860 3970
rect 6894 3936 6928 3970
rect 6962 3936 6996 3970
rect 7030 3936 7064 3970
rect 4000 3320 4034 3354
rect 4000 3251 4034 3285
rect 4000 3182 4034 3216
rect 4000 3113 4034 3147
rect 5276 3320 5310 3354
rect 5276 3251 5310 3285
rect 5838 3320 5872 3354
rect 5838 3251 5872 3285
rect 5276 3182 5310 3216
rect 5344 3214 5378 3248
rect 5415 3214 5449 3248
rect 5486 3214 5520 3248
rect 5557 3214 5591 3248
rect 5628 3214 5662 3248
rect 5699 3214 5733 3248
rect 5770 3214 5804 3248
rect 4000 3044 4034 3078
rect 5276 3113 5310 3147
rect 5838 3182 5872 3216
rect 5838 3113 5872 3147
rect 7114 3320 7148 3354
rect 7114 3251 7148 3285
rect 7114 3182 7148 3216
rect 4000 2975 4034 3009
rect 4000 2906 4034 2940
rect 4000 2837 4034 2871
rect 5276 3044 5310 3078
rect 5276 2975 5310 3009
rect 5276 2906 5310 2940
rect 5276 2837 5310 2871
rect 4000 2768 4034 2802
rect 4000 2699 4034 2733
rect 4000 2630 4034 2664
rect 5276 2768 5310 2802
rect 5276 2699 5310 2733
rect 5838 3044 5872 3078
rect 7114 3113 7148 3147
rect 5838 2975 5872 3009
rect 5838 2906 5872 2940
rect 5838 2837 5872 2871
rect 7114 3044 7148 3078
rect 7114 2975 7148 3009
rect 7114 2906 7148 2940
rect 7114 2837 7148 2871
rect 5838 2768 5872 2802
rect 5838 2699 5872 2733
rect 5276 2630 5310 2664
rect 4000 2561 4034 2595
rect 5276 2561 5310 2595
rect 4000 2492 4034 2526
rect 4000 2423 4034 2457
rect 4000 2354 4034 2388
rect 5838 2630 5872 2664
rect 7114 2768 7148 2802
rect 7114 2699 7148 2733
rect 7114 2630 7148 2664
rect 5838 2561 5872 2595
rect 7114 2561 7148 2595
rect 5276 2492 5310 2526
rect 5359 2486 5393 2520
rect 5427 2486 5461 2520
rect 5495 2486 5529 2520
rect 5563 2486 5597 2520
rect 5631 2486 5665 2520
rect 5699 2486 5733 2520
rect 5767 2486 5801 2520
rect 5838 2492 5872 2526
rect 5276 2423 5310 2457
rect 5359 2417 5393 2451
rect 5427 2417 5461 2451
rect 5495 2417 5529 2451
rect 5563 2417 5597 2451
rect 5631 2417 5665 2451
rect 5699 2417 5733 2451
rect 5767 2417 5801 2451
rect 5838 2423 5872 2457
rect 4000 2285 4034 2319
rect 5276 2354 5310 2388
rect 5359 2348 5393 2382
rect 5427 2348 5461 2382
rect 5495 2348 5529 2382
rect 5563 2348 5597 2382
rect 5631 2348 5665 2382
rect 5699 2348 5733 2382
rect 5767 2348 5801 2382
rect 5838 2354 5872 2388
rect 7114 2492 7148 2526
rect 7114 2423 7148 2457
rect 4000 2216 4034 2250
rect 4000 2147 4034 2181
rect 4000 2078 4034 2112
rect 5276 2285 5310 2319
rect 5359 2279 5393 2313
rect 5427 2279 5461 2313
rect 5495 2279 5529 2313
rect 5563 2279 5597 2313
rect 5631 2279 5665 2313
rect 5699 2279 5733 2313
rect 5767 2279 5801 2313
rect 5838 2285 5872 2319
rect 7114 2354 7148 2388
rect 5276 2216 5310 2250
rect 5359 2210 5393 2244
rect 5427 2210 5461 2244
rect 5495 2210 5529 2244
rect 5563 2210 5597 2244
rect 5631 2210 5665 2244
rect 5699 2210 5733 2244
rect 5767 2210 5801 2244
rect 5838 2216 5872 2250
rect 5276 2147 5310 2181
rect 5359 2141 5393 2175
rect 5427 2141 5461 2175
rect 5495 2141 5529 2175
rect 5563 2141 5597 2175
rect 5631 2141 5665 2175
rect 5699 2141 5733 2175
rect 5767 2141 5801 2175
rect 5838 2147 5872 2181
rect 5276 2078 5310 2112
rect 5359 2072 5393 2106
rect 5427 2072 5461 2106
rect 5495 2072 5529 2106
rect 5563 2072 5597 2106
rect 5631 2072 5665 2106
rect 5699 2072 5733 2106
rect 5767 2072 5801 2106
rect 5838 2078 5872 2112
rect 7114 2285 7148 2319
rect 7114 2216 7148 2250
rect 7114 2147 7148 2181
rect 4000 2009 4034 2043
rect 4000 1940 4034 1974
rect 1492 1886 1526 1920
rect 1562 1886 1596 1920
rect 1632 1886 1666 1920
rect 1702 1886 1736 1920
rect 1772 1886 1806 1920
rect 1842 1886 1876 1920
rect 1912 1886 1946 1920
rect 1982 1886 2016 1920
rect 2052 1886 2086 1920
rect 2122 1886 2156 1920
rect 2192 1886 2226 1920
rect 2262 1886 2296 1920
rect 2332 1886 2366 1920
rect 2402 1886 2436 1920
rect 2472 1886 2506 1920
rect 2542 1886 2576 1920
rect 2611 1886 2645 1920
rect 2680 1886 2714 1920
rect 2749 1886 2783 1920
rect 2818 1886 2852 1920
rect 2887 1886 2921 1920
rect 2956 1886 2990 1920
rect 3025 1886 3059 1920
rect 3094 1886 3128 1920
rect 3163 1886 3197 1920
rect 3232 1886 3266 1920
rect 3301 1886 3335 1920
rect 3370 1886 3404 1920
rect 3439 1886 3473 1920
rect 3508 1886 3542 1920
rect 3612 1852 3646 1886
rect 3709 1862 3743 1896
rect 3777 1862 3811 1896
rect 3845 1862 3879 1896
rect 3913 1862 3947 1896
rect 4000 1870 4034 1904
rect 7114 2078 7148 2112
rect 5276 2009 5310 2043
rect 5359 2003 5393 2037
rect 5427 2003 5461 2037
rect 5495 2003 5529 2037
rect 5563 2003 5597 2037
rect 5631 2003 5665 2037
rect 5699 2003 5733 2037
rect 5767 2003 5801 2037
rect 5838 2009 5872 2043
rect 5276 1940 5310 1974
rect 5359 1934 5393 1968
rect 5427 1934 5461 1968
rect 5495 1934 5529 1968
rect 5563 1934 5597 1968
rect 5631 1934 5665 1968
rect 5699 1934 5733 1968
rect 5767 1934 5801 1968
rect 5838 1940 5872 1974
rect 5276 1871 5310 1905
rect 5359 1865 5393 1899
rect 5427 1865 5461 1899
rect 5495 1865 5529 1899
rect 5563 1865 5597 1899
rect 5631 1865 5665 1899
rect 5699 1865 5733 1899
rect 5767 1865 5801 1899
rect 5838 1871 5872 1905
rect 3612 1782 3646 1816
rect 3709 1793 3743 1827
rect 3777 1793 3811 1827
rect 3845 1793 3879 1827
rect 3913 1793 3947 1827
rect 4000 1800 4034 1834
rect 7114 2009 7148 2043
rect 7114 1940 7148 1974
rect 7114 1870 7148 1904
rect 7207 1862 7241 1896
rect 7275 1862 7309 1896
rect 7343 1862 7377 1896
rect 7411 1862 7445 1896
rect 7606 1886 7640 1920
rect 7675 1886 7709 1920
rect 7744 1886 7778 1920
rect 7813 1886 7847 1920
rect 7882 1886 7916 1920
rect 7951 1886 7985 1920
rect 8020 1886 8054 1920
rect 8089 1886 8123 1920
rect 8158 1886 8192 1920
rect 8227 1886 8261 1920
rect 8296 1886 8330 1920
rect 8365 1886 8399 1920
rect 8434 1886 8468 1920
rect 8503 1886 8537 1920
rect 8572 1886 8606 1920
rect 8642 1886 8676 1920
rect 8712 1886 8746 1920
rect 8782 1886 8816 1920
rect 8852 1886 8886 1920
rect 8922 1886 8956 1920
rect 8992 1886 9026 1920
rect 9062 1886 9096 1920
rect 9132 1886 9166 1920
rect 9202 1886 9236 1920
rect 9272 1886 9306 1920
rect 9342 1886 9376 1920
rect 9412 1886 9446 1920
rect 9482 1886 9516 1920
rect 9552 1886 9586 1920
rect 9622 1886 9656 1920
rect 7502 1852 7536 1886
rect 5276 1802 5310 1836
rect 5359 1796 5393 1830
rect 5427 1796 5461 1830
rect 5495 1796 5529 1830
rect 5563 1796 5597 1830
rect 5631 1796 5665 1830
rect 5699 1796 5733 1830
rect 5767 1796 5801 1830
rect 5838 1802 5872 1836
rect 3612 1712 3646 1746
rect 3709 1724 3743 1758
rect 3777 1724 3811 1758
rect 3845 1724 3879 1758
rect 3913 1724 3947 1758
rect 4000 1730 4034 1764
rect 3612 1642 3646 1676
rect 3709 1655 3743 1689
rect 3777 1655 3811 1689
rect 3845 1655 3879 1689
rect 3913 1655 3947 1689
rect 4000 1660 4034 1694
rect 3612 1572 3646 1606
rect 3709 1586 3743 1620
rect 3777 1586 3811 1620
rect 3845 1586 3879 1620
rect 3913 1586 3947 1620
rect 4000 1590 4034 1624
rect 7114 1800 7148 1834
rect 7207 1793 7241 1827
rect 7275 1793 7309 1827
rect 7343 1793 7377 1827
rect 7411 1793 7445 1827
rect 5276 1732 5310 1766
rect 5359 1727 5393 1761
rect 5427 1727 5461 1761
rect 5495 1727 5529 1761
rect 5563 1727 5597 1761
rect 5631 1727 5665 1761
rect 5699 1727 5733 1761
rect 5767 1727 5801 1761
rect 5838 1732 5872 1766
rect 5276 1662 5310 1696
rect 5359 1658 5393 1692
rect 5427 1658 5461 1692
rect 5495 1658 5529 1692
rect 5563 1658 5597 1692
rect 5631 1658 5665 1692
rect 5699 1658 5733 1692
rect 5767 1658 5801 1692
rect 5838 1662 5872 1696
rect 5276 1592 5310 1626
rect 5359 1589 5393 1623
rect 5427 1589 5461 1623
rect 5495 1589 5529 1623
rect 5563 1589 5597 1623
rect 5631 1589 5665 1623
rect 5699 1589 5733 1623
rect 5767 1589 5801 1623
rect 5838 1592 5872 1626
rect 7502 1782 7536 1816
rect 7114 1730 7148 1764
rect 7207 1724 7241 1758
rect 7275 1724 7309 1758
rect 7343 1724 7377 1758
rect 7411 1724 7445 1758
rect 7502 1712 7536 1746
rect 7114 1660 7148 1694
rect 7207 1655 7241 1689
rect 7275 1655 7309 1689
rect 7343 1655 7377 1689
rect 7411 1655 7445 1689
rect 7502 1642 7536 1676
rect 7114 1590 7148 1624
rect 3612 1502 3646 1536
rect 3709 1517 3743 1551
rect 3777 1517 3811 1551
rect 3845 1517 3879 1551
rect 3913 1517 3947 1551
rect 4000 1520 4034 1554
rect 3612 1432 3646 1466
rect 3709 1448 3743 1482
rect 3777 1448 3811 1482
rect 3845 1448 3879 1482
rect 3913 1448 3947 1482
rect 4000 1450 4034 1484
rect 3612 1362 3646 1396
rect 3709 1379 3743 1413
rect 3777 1379 3811 1413
rect 3845 1379 3879 1413
rect 3913 1379 3947 1413
rect 4000 1380 4034 1414
rect 3612 1292 3646 1326
rect 3709 1310 3743 1344
rect 3777 1310 3811 1344
rect 3845 1310 3879 1344
rect 3913 1310 3947 1344
rect 4000 1310 4034 1344
rect 5276 1522 5310 1556
rect 5359 1520 5393 1554
rect 5427 1520 5461 1554
rect 5495 1520 5529 1554
rect 5563 1520 5597 1554
rect 5631 1520 5665 1554
rect 5699 1520 5733 1554
rect 5767 1520 5801 1554
rect 5838 1522 5872 1556
rect 7207 1586 7241 1620
rect 7275 1586 7309 1620
rect 7343 1586 7377 1620
rect 7411 1586 7445 1620
rect 7502 1572 7536 1606
rect 5276 1452 5310 1486
rect 5359 1451 5393 1485
rect 5427 1451 5461 1485
rect 5495 1451 5529 1485
rect 5563 1451 5597 1485
rect 5631 1451 5665 1485
rect 5699 1451 5733 1485
rect 5767 1451 5801 1485
rect 5838 1452 5872 1486
rect 5276 1382 5310 1416
rect 5359 1382 5393 1416
rect 5427 1382 5461 1416
rect 5495 1382 5529 1416
rect 5563 1382 5597 1416
rect 5631 1382 5665 1416
rect 5699 1382 5733 1416
rect 5767 1382 5801 1416
rect 5838 1382 5872 1416
rect 5276 1312 5310 1346
rect 5359 1312 5393 1346
rect 5427 1312 5461 1346
rect 5495 1312 5529 1346
rect 5563 1312 5597 1346
rect 5631 1312 5665 1346
rect 5699 1312 5733 1346
rect 5767 1312 5801 1346
rect 5838 1312 5872 1346
rect 7114 1520 7148 1554
rect 7207 1517 7241 1551
rect 7275 1517 7309 1551
rect 7343 1517 7377 1551
rect 7411 1517 7445 1551
rect 7502 1502 7536 1536
rect 7114 1450 7148 1484
rect 7207 1448 7241 1482
rect 7275 1448 7309 1482
rect 7343 1448 7377 1482
rect 7411 1448 7445 1482
rect 7502 1432 7536 1466
rect 7114 1380 7148 1414
rect 7207 1379 7241 1413
rect 7275 1379 7309 1413
rect 7343 1379 7377 1413
rect 7411 1379 7445 1413
rect 7502 1362 7536 1396
rect 3612 1223 3646 1257
rect 3709 1240 3743 1274
rect 3777 1240 3811 1274
rect 3845 1240 3879 1274
rect 3913 1240 3947 1274
rect 4000 1240 4034 1274
rect 3612 1154 3646 1188
rect 3709 1170 3743 1204
rect 3777 1170 3811 1204
rect 3845 1170 3879 1204
rect 3913 1170 3947 1204
rect 4000 1170 4034 1204
rect 3612 1085 3646 1119
rect 3709 1100 3743 1134
rect 3777 1100 3811 1134
rect 3845 1100 3879 1134
rect 3913 1100 3947 1134
rect 4000 1100 4034 1134
rect 7114 1310 7148 1344
rect 7207 1310 7241 1344
rect 7275 1310 7309 1344
rect 7343 1310 7377 1344
rect 7411 1310 7445 1344
rect 7502 1292 7536 1326
rect 5276 1242 5310 1276
rect 5359 1242 5393 1276
rect 5427 1242 5461 1276
rect 5495 1242 5529 1276
rect 5563 1242 5597 1276
rect 5631 1242 5665 1276
rect 5699 1242 5733 1276
rect 5767 1242 5801 1276
rect 5838 1242 5872 1276
rect 5276 1172 5310 1206
rect 5359 1172 5393 1206
rect 5427 1172 5461 1206
rect 5495 1172 5529 1206
rect 5563 1172 5597 1206
rect 5631 1172 5665 1206
rect 5699 1172 5733 1206
rect 5767 1172 5801 1206
rect 5838 1172 5872 1206
rect 5276 1102 5310 1136
rect 5359 1102 5393 1136
rect 5427 1102 5461 1136
rect 5495 1102 5529 1136
rect 5563 1102 5597 1136
rect 5631 1102 5665 1136
rect 5699 1102 5733 1136
rect 5767 1102 5801 1136
rect 5838 1102 5872 1136
rect 3612 1016 3646 1050
rect 3709 1030 3743 1064
rect 3777 1030 3811 1064
rect 3845 1030 3879 1064
rect 3913 1030 3947 1064
rect 4000 1030 4034 1064
rect 7114 1240 7148 1274
rect 7207 1240 7241 1274
rect 7275 1240 7309 1274
rect 7343 1240 7377 1274
rect 7411 1240 7445 1274
rect 7502 1223 7536 1257
rect 7114 1170 7148 1204
rect 7207 1170 7241 1204
rect 7275 1170 7309 1204
rect 7343 1170 7377 1204
rect 7411 1170 7445 1204
rect 7502 1154 7536 1188
rect 7114 1100 7148 1134
rect 7207 1100 7241 1134
rect 7275 1100 7309 1134
rect 7343 1100 7377 1134
rect 7411 1100 7445 1134
rect 7502 1085 7536 1119
rect 5276 1032 5310 1066
rect 5359 1032 5393 1066
rect 5427 1032 5461 1066
rect 5495 1032 5529 1066
rect 5563 1032 5597 1066
rect 5631 1032 5665 1066
rect 5699 1032 5733 1066
rect 5767 1032 5801 1066
rect 5838 1032 5872 1066
rect 3612 947 3646 981
rect 3709 960 3743 994
rect 3777 960 3811 994
rect 3845 960 3879 994
rect 3913 960 3947 994
rect 4000 960 4034 994
rect 3612 878 3646 912
rect 3709 890 3743 924
rect 3777 890 3811 924
rect 3845 890 3879 924
rect 3913 890 3947 924
rect 4000 890 4034 924
rect 7114 1030 7148 1064
rect 7207 1030 7241 1064
rect 7275 1030 7309 1064
rect 7343 1030 7377 1064
rect 7411 1030 7445 1064
rect 5276 962 5310 996
rect 5359 962 5393 996
rect 5427 962 5461 996
rect 5495 962 5529 996
rect 5563 962 5597 996
rect 5631 962 5665 996
rect 5699 962 5733 996
rect 5767 962 5801 996
rect 5838 962 5872 996
rect 5276 892 5310 926
rect 5359 892 5393 926
rect 5427 892 5461 926
rect 5495 892 5529 926
rect 5563 892 5597 926
rect 5631 892 5665 926
rect 5699 892 5733 926
rect 5767 892 5801 926
rect 5838 892 5872 926
rect 3612 809 3646 843
rect 3709 820 3743 854
rect 3777 820 3811 854
rect 3845 820 3879 854
rect 3913 820 3947 854
rect 4000 820 4034 854
rect 3612 740 3646 774
rect 3709 750 3743 784
rect 3777 750 3811 784
rect 3845 750 3879 784
rect 3913 750 3947 784
rect 4000 750 4034 784
rect 7502 1016 7536 1050
rect 7114 960 7148 994
rect 7207 960 7241 994
rect 7275 960 7309 994
rect 7343 960 7377 994
rect 7411 960 7445 994
rect 7502 947 7536 981
rect 7114 890 7148 924
rect 7207 890 7241 924
rect 7275 890 7309 924
rect 7343 890 7377 924
rect 7411 890 7445 924
rect 5276 822 5310 856
rect 5359 822 5393 856
rect 5427 822 5461 856
rect 5495 822 5529 856
rect 5563 822 5597 856
rect 5631 822 5665 856
rect 5699 822 5733 856
rect 5767 822 5801 856
rect 5838 822 5872 856
rect 3612 671 3646 705
rect 3709 680 3743 714
rect 3777 680 3811 714
rect 3845 680 3879 714
rect 3913 680 3947 714
rect 4000 680 4034 714
rect 3612 602 3646 636
rect 3709 610 3743 644
rect 3777 610 3811 644
rect 3845 610 3879 644
rect 3913 610 3947 644
rect 4000 610 4034 644
rect 3709 540 3743 574
rect 3777 540 3811 574
rect 3845 540 3879 574
rect 3913 540 3947 574
rect 4000 540 4034 574
rect 1554 446 1588 480
rect 1623 446 1657 480
rect 1692 446 1726 480
rect 1761 446 1795 480
rect 1830 446 1864 480
rect 1899 446 1933 480
rect 1968 446 2002 480
rect 2038 446 2072 480
rect 2108 446 2142 480
rect 2178 446 2212 480
rect 2248 446 2282 480
rect 2318 446 2352 480
rect 2388 446 2422 480
rect 2458 446 2492 480
rect 2528 446 2562 480
rect 2598 446 2632 480
rect 2668 446 2702 480
rect 2738 446 2772 480
rect 2808 446 2842 480
rect 2878 446 2912 480
rect 2948 446 2982 480
rect 3018 446 3052 480
rect 3088 446 3122 480
rect 3158 446 3192 480
rect 3228 446 3262 480
rect 3298 446 3332 480
rect 3368 446 3402 480
rect 3438 446 3472 480
rect 3508 446 3542 480
rect 3578 446 3612 480
rect 3709 470 3743 504
rect 3777 470 3811 504
rect 3845 470 3879 504
rect 3913 470 3947 504
rect 4000 470 4034 504
rect 5276 752 5310 786
rect 5359 752 5393 786
rect 5427 752 5461 786
rect 5495 752 5529 786
rect 5563 752 5597 786
rect 5631 752 5665 786
rect 5699 752 5733 786
rect 5767 752 5801 786
rect 5838 752 5872 786
rect 7502 878 7536 912
rect 7114 820 7148 854
rect 7207 820 7241 854
rect 7275 820 7309 854
rect 7343 820 7377 854
rect 7411 820 7445 854
rect 7502 809 7536 843
rect 5276 682 5310 716
rect 5359 682 5393 716
rect 5427 682 5461 716
rect 5495 682 5529 716
rect 5563 682 5597 716
rect 5631 682 5665 716
rect 5699 682 5733 716
rect 5767 682 5801 716
rect 5838 682 5872 716
rect 5276 612 5310 646
rect 5359 612 5393 646
rect 5427 612 5461 646
rect 5495 612 5529 646
rect 5563 612 5597 646
rect 5631 612 5665 646
rect 5699 612 5733 646
rect 5767 612 5801 646
rect 5838 612 5872 646
rect 5276 542 5310 576
rect 5359 542 5393 576
rect 5427 542 5461 576
rect 5495 542 5529 576
rect 5563 542 5597 576
rect 5631 542 5665 576
rect 5699 542 5733 576
rect 5767 542 5801 576
rect 5838 542 5872 576
rect 5276 472 5310 506
rect 5359 472 5393 506
rect 5427 472 5461 506
rect 5495 472 5529 506
rect 5563 472 5597 506
rect 5631 472 5665 506
rect 5699 472 5733 506
rect 5767 472 5801 506
rect 5838 472 5872 506
rect 7114 750 7148 784
rect 7207 750 7241 784
rect 7275 750 7309 784
rect 7343 750 7377 784
rect 7411 750 7445 784
rect 7502 740 7536 774
rect 7114 680 7148 714
rect 7207 680 7241 714
rect 7275 680 7309 714
rect 7343 680 7377 714
rect 7411 680 7445 714
rect 7502 671 7536 705
rect 7114 610 7148 644
rect 7207 610 7241 644
rect 7275 610 7309 644
rect 7343 610 7377 644
rect 7411 610 7445 644
rect 7502 602 7536 636
rect 7114 540 7148 574
rect 7207 540 7241 574
rect 7275 540 7309 574
rect 7343 540 7377 574
rect 7411 540 7445 574
rect 7114 470 7148 504
rect 7207 470 7241 504
rect 7275 470 7309 504
rect 7343 470 7377 504
rect 7411 470 7445 504
rect 7536 446 7570 480
rect 7606 446 7640 480
rect 7676 446 7710 480
rect 7746 446 7780 480
rect 7816 446 7850 480
rect 7886 446 7920 480
rect 7956 446 7990 480
rect 8026 446 8060 480
rect 8096 446 8130 480
rect 8166 446 8200 480
rect 8236 446 8270 480
rect 8306 446 8340 480
rect 8376 446 8410 480
rect 8446 446 8480 480
rect 8516 446 8550 480
rect 8586 446 8620 480
rect 8656 446 8690 480
rect 8726 446 8760 480
rect 8796 446 8830 480
rect 8866 446 8900 480
rect 8936 446 8970 480
rect 9006 446 9040 480
rect 9076 446 9110 480
rect 9146 446 9180 480
rect 9215 446 9249 480
rect 9284 446 9318 480
rect 9353 446 9387 480
rect 9422 446 9456 480
rect 9491 446 9525 480
rect 9560 446 9594 480
rect 10283 7671 10317 7705
rect 10351 7671 10385 7705
rect 10419 7671 10453 7705
rect 10487 7671 10521 7705
rect 10555 7671 10589 7705
rect 10623 7671 10657 7705
rect 10691 7671 10725 7705
rect 10759 7671 10793 7705
rect 10827 7671 10861 7705
rect 10895 7671 10929 7705
rect 10963 7671 10997 7705
rect 11031 7671 11065 7705
rect 11099 7671 11133 7705
rect 11167 7671 11201 7705
rect 11235 7671 11269 7705
rect 11303 7671 11337 7705
rect 11371 7671 11405 7705
rect 11439 7671 11473 7705
rect 11507 7671 11541 7705
rect 11575 7671 11609 7705
rect 11643 7671 11677 7705
rect 11711 7671 11745 7705
rect 11779 7671 11813 7705
rect 11847 7671 11881 7705
rect 11915 7671 11949 7705
rect 11983 7671 12017 7705
rect 12051 7671 12085 7705
rect 12119 7671 12153 7705
rect 12187 7671 12221 7705
rect 12255 7671 12289 7705
rect 12323 7671 12357 7705
rect 12391 7671 12425 7705
rect 12459 7671 12493 7705
rect 12527 7671 12561 7705
rect 12595 7671 12629 7705
rect 12663 7671 12697 7705
rect 12731 7671 12765 7705
rect 10212 7637 10246 7671
rect 10212 7569 10246 7603
rect 10212 7501 10246 7535
rect 10212 7433 10246 7467
rect 10212 7365 10246 7399
rect 10212 7297 10246 7331
rect 10212 7229 10246 7263
rect 10212 7161 10246 7195
rect 10212 7093 10246 7127
rect 10212 7025 10246 7059
rect 10212 6957 10246 6991
rect 10212 6889 10246 6923
rect 10212 6821 10246 6855
rect 10212 6753 10246 6787
rect 10212 6685 10246 6719
rect 10212 6617 10246 6651
rect 10212 6549 10246 6583
rect 10212 6481 10246 6515
rect 10212 6413 10246 6447
rect 10212 6345 10246 6379
rect 10212 6277 10246 6311
rect 10212 6209 10246 6243
rect 10212 6141 10246 6175
rect 10212 6073 10246 6107
rect 10212 6005 10246 6039
rect 10212 5937 10246 5971
rect 10212 5869 10246 5903
rect 10212 5801 10246 5835
rect 10212 5733 10246 5767
rect 10212 5665 10246 5699
rect 10212 5597 10246 5631
rect 10212 5529 10246 5563
rect 10212 5461 10246 5495
rect 10212 5393 10246 5427
rect 10212 5325 10246 5359
rect 10212 5257 10246 5291
rect 10212 5189 10246 5223
rect 10212 5121 10246 5155
rect 10212 5053 10246 5087
rect 10212 4985 10246 5019
rect 10212 4917 10246 4951
rect 10212 4849 10246 4883
rect 10212 4781 10246 4815
rect 10212 4713 10246 4747
rect 10212 4645 10246 4679
rect 10212 4577 10246 4611
rect 10212 4509 10246 4543
rect 10212 4441 10246 4475
rect 10212 4373 10246 4407
rect 10212 4305 10246 4339
rect 10212 4237 10246 4271
rect 10212 4169 10246 4203
rect 10212 4101 10246 4135
rect 10212 4033 10246 4067
rect 10212 3965 10246 3999
rect 10212 3897 10246 3931
rect 10212 3829 10246 3863
rect 10212 3761 10246 3795
rect 10212 3693 10246 3727
rect 10212 3625 10246 3659
rect 10212 3557 10246 3591
rect 10212 3489 10246 3523
rect 10212 3421 10246 3455
rect 10212 3353 10246 3387
rect 10212 3285 10246 3319
rect 10212 3217 10246 3251
rect 10212 3149 10246 3183
rect 10212 3081 10246 3115
rect 10212 3013 10246 3047
rect 10212 2945 10246 2979
rect 10212 2877 10246 2911
rect 10212 2809 10246 2843
rect 10212 2741 10246 2775
rect 10212 2673 10246 2707
rect 10212 2605 10246 2639
rect 10212 2537 10246 2571
rect 10212 2469 10246 2503
rect 10212 2401 10246 2435
rect 10212 2333 10246 2367
rect 10212 2265 10246 2299
rect 10212 2197 10246 2231
rect 10212 2129 10246 2163
rect 10212 2061 10246 2095
rect 10212 1993 10246 2027
rect 10212 1925 10246 1959
rect 10212 1857 10246 1891
rect 10212 1789 10246 1823
rect 10212 1721 10246 1755
rect 10212 1653 10246 1687
rect 10212 1585 10246 1619
rect 10212 1517 10246 1551
rect 10212 1449 10246 1483
rect 10212 1381 10246 1415
rect 10212 1313 10246 1347
rect 10212 1245 10246 1279
rect 10212 1177 10246 1211
rect 10212 1109 10246 1143
rect 10212 1041 10246 1075
rect 10212 973 10246 1007
rect 10212 905 10246 939
rect 10212 837 10246 871
rect 10212 769 10246 803
rect 10212 701 10246 735
rect 10212 633 10246 667
rect 10212 565 10246 599
rect 10246 446 10280 480
rect 10314 446 10348 480
rect 10382 446 10416 480
rect 10450 446 10484 480
rect 10518 446 10552 480
rect 10586 446 10620 480
rect 10690 446 10724 480
rect 10758 446 10792 480
rect 10826 446 10860 480
rect 10894 446 10928 480
rect 10962 446 10996 480
rect 11030 446 11064 480
rect 11098 446 11132 480
rect 11166 446 11200 480
rect 11234 446 11268 480
rect 11302 446 11336 480
rect 11370 446 11404 480
rect 11438 446 11472 480
rect 11506 446 11540 480
rect 11574 446 11608 480
rect 11642 446 11676 480
rect 11710 446 11744 480
rect 11778 446 11812 480
rect 11846 446 11880 480
rect 11914 446 11948 480
rect 11982 446 12016 480
rect 12050 446 12084 480
rect 12118 446 12152 480
rect 12186 446 12220 480
rect 12254 446 12288 480
rect 12322 446 12356 480
rect 12390 446 12424 480
rect 12458 446 12492 480
rect 12526 446 12560 480
rect 12594 446 12628 480
rect 12662 446 12696 480
rect 12730 446 12764 480
<< mvnsubdiffcont >>
rect 1231 14200 1265 14234
rect 1299 14200 1333 14234
rect 1367 14200 1401 14234
rect 1435 14200 1469 14234
rect 1503 14200 1537 14234
rect 1571 14200 1605 14234
rect 1639 14200 1673 14234
rect 1707 14200 1741 14234
rect 1775 14200 1809 14234
rect 1843 14200 1877 14234
rect 1911 14200 1945 14234
rect 1979 14200 2013 14234
rect 2047 14200 2081 14234
rect 2115 14200 2149 14234
rect 2183 14200 2217 14234
rect 2251 14200 2285 14234
rect 2319 14200 2353 14234
rect 2387 14200 2421 14234
rect 2455 14200 2489 14234
rect 2523 14200 2557 14234
rect 2591 14200 2625 14234
rect 2659 14200 2693 14234
rect 2727 14200 2761 14234
rect 2795 14200 2829 14234
rect 2863 14200 2897 14234
rect 2931 14200 2965 14234
rect 2999 14200 3033 14234
rect 3067 14200 3101 14234
rect 3135 14200 3169 14234
rect 3203 14200 3237 14234
rect 3271 14200 3305 14234
rect 3339 14200 3373 14234
rect 3407 14200 3441 14234
rect 3475 14200 3509 14234
rect 3543 14200 3577 14234
rect 3611 14200 3645 14234
rect 3679 14200 3713 14234
rect 3747 14200 3781 14234
rect 3815 14200 3849 14234
rect 3883 14200 3917 14234
rect 3951 14200 3985 14234
rect 4019 14200 4053 14234
rect 4087 14200 4121 14234
rect 4155 14200 4189 14234
rect 4223 14200 4257 14234
rect 4291 14200 4325 14234
rect 4359 14200 4393 14234
rect 4427 14200 4461 14234
rect 4495 14200 4529 14234
rect 4563 14200 4597 14234
rect 4631 14200 4665 14234
rect 4699 14200 4733 14234
rect 4767 14200 4801 14234
rect 4835 14200 4869 14234
rect 4903 14200 4937 14234
rect 4971 14200 5005 14234
rect 5039 14200 5073 14234
rect 5107 14200 5141 14234
rect 5175 14200 5209 14234
rect 5243 14200 5277 14234
rect 5311 14200 5345 14234
rect 5379 14200 5413 14234
rect 5447 14200 5481 14234
rect 5515 14200 5549 14234
rect 5583 14200 5617 14234
rect 5651 14200 5685 14234
rect 5719 14200 5753 14234
rect 5787 14200 5821 14234
rect 5855 14200 5889 14234
rect 5923 14200 5957 14234
rect 5991 14200 6025 14234
rect 6059 14200 6093 14234
rect 6127 14200 6161 14234
rect 6195 14200 6229 14234
rect 6263 14200 6297 14234
rect 6331 14200 6365 14234
rect 6399 14200 6433 14234
rect 6467 14200 6501 14234
rect 6535 14200 6569 14234
rect 6603 14200 6637 14234
rect 6671 14200 6705 14234
rect 6739 14200 6773 14234
rect 6807 14200 6841 14234
rect 6875 14200 6909 14234
rect 6943 14200 6977 14234
rect 7011 14200 7045 14234
rect 7079 14200 7113 14234
rect 7147 14200 7181 14234
rect 7215 14200 7249 14234
rect 7283 14200 7317 14234
rect 7351 14200 7385 14234
rect 7419 14200 7453 14234
rect 7487 14200 7521 14234
rect 7555 14200 7589 14234
rect 7623 14200 7657 14234
rect 7691 14200 7725 14234
rect 7759 14200 7793 14234
rect 7827 14200 7861 14234
rect 7895 14200 7929 14234
rect 7963 14200 7997 14234
rect 8031 14200 8065 14234
rect 8099 14200 8133 14234
rect 8167 14200 8201 14234
rect 8235 14200 8269 14234
rect 8303 14200 8337 14234
rect 8371 14200 8405 14234
rect 8439 14200 8473 14234
rect 8507 14200 8541 14234
rect 8575 14200 8609 14234
rect 8643 14200 8677 14234
rect 8711 14200 8745 14234
rect 8779 14200 8813 14234
rect 8847 14200 8881 14234
rect 8915 14200 8949 14234
rect 8983 14200 9017 14234
rect 9051 14200 9085 14234
rect 9119 14200 9153 14234
rect 9187 14200 9221 14234
rect 9255 14200 9289 14234
rect 9323 14200 9357 14234
rect 9391 14200 9425 14234
rect 9459 14200 9493 14234
rect 9527 14200 9561 14234
rect 9595 14200 9629 14234
rect 9663 14200 9697 14234
rect 9731 14200 9765 14234
rect 9799 14200 9833 14234
rect 9867 14200 9901 14234
rect 9935 14200 9969 14234
rect 10003 14200 10037 14234
rect 10071 14200 10105 14234
rect 10139 14200 10173 14234
rect 10207 14200 10241 14234
rect 10275 14200 10309 14234
rect 10343 14200 10377 14234
rect 10411 14200 10445 14234
rect 10479 14200 10513 14234
rect 10547 14200 10581 14234
rect 10615 14200 10649 14234
rect 10683 14200 10717 14234
rect 10751 14200 10785 14234
rect 10819 14200 10853 14234
rect 10887 14200 10921 14234
rect 10955 14200 10989 14234
rect 1371 14132 1405 14166
rect 1443 14132 1477 14166
rect 1515 14132 1549 14166
rect 1197 14066 1231 14100
rect 1371 14060 1405 14094
rect 1443 14060 1477 14094
rect 1515 14060 1549 14094
rect 5189 14121 5223 14155
rect 5265 14121 5299 14155
rect 5341 14121 5375 14155
rect 5417 14121 5451 14155
rect 5493 14121 5527 14155
rect 5569 14121 5603 14155
rect 5645 14121 5679 14155
rect 5721 14121 5755 14155
rect 5796 14121 5830 14155
rect 5871 14121 5905 14155
rect 1197 13998 1231 14032
rect 1371 13987 1405 14021
rect 1443 13987 1477 14021
rect 1515 13987 1549 14021
rect 1197 13930 1231 13964
rect 1371 13914 1405 13948
rect 1443 13914 1477 13948
rect 1515 13914 1549 13948
rect 1197 13862 1231 13896
rect 1371 13841 1405 13875
rect 1443 13841 1477 13875
rect 1515 13841 1549 13875
rect 1197 13794 1231 13828
rect 1371 13768 1405 13802
rect 1443 13768 1477 13802
rect 1515 13768 1549 13802
rect 1197 13726 1231 13760
rect 1371 13695 1405 13729
rect 1443 13695 1477 13729
rect 1515 13695 1549 13729
rect 1197 13658 1231 13692
rect 1197 13590 1231 13624
rect 1371 13622 1405 13656
rect 1443 13622 1477 13656
rect 1515 13622 1549 13656
rect 1197 13522 1231 13556
rect 1371 13549 1405 13583
rect 1443 13549 1477 13583
rect 1515 13549 1549 13583
rect 1197 13454 1231 13488
rect 1371 13476 1405 13510
rect 1443 13476 1477 13510
rect 1515 13476 1549 13510
rect 1197 13386 1231 13420
rect 1371 13403 1405 13437
rect 1443 13403 1477 13437
rect 1515 13403 1549 13437
rect 1197 13318 1231 13352
rect 1371 13330 1405 13364
rect 1443 13330 1477 13364
rect 1515 13330 1549 13364
rect 1197 13250 1231 13284
rect 1371 13257 1405 13291
rect 1443 13257 1477 13291
rect 1515 13257 1549 13291
rect 1197 13182 1231 13216
rect 1371 13184 1405 13218
rect 1443 13184 1477 13218
rect 1515 13184 1549 13218
rect 1197 13090 1231 13124
rect 1197 13020 1231 13054
rect 1197 12950 1231 12984
rect 1197 12880 1231 12914
rect 1197 12810 1231 12844
rect 1197 12740 1231 12774
rect 1197 12670 1231 12704
rect 1197 12599 1231 12633
rect 1197 12528 1231 12562
rect 9399 14119 9433 14153
rect 9472 14119 9506 14153
rect 9545 14119 9579 14153
rect 9618 14119 9652 14153
rect 9691 14119 9725 14153
rect 9763 14119 9797 14153
rect 9835 14119 9869 14153
rect 5189 14049 5223 14083
rect 5265 14049 5299 14083
rect 5341 14049 5375 14083
rect 5417 14049 5451 14083
rect 5493 14049 5527 14083
rect 5569 14049 5603 14083
rect 5645 14049 5679 14083
rect 5721 14049 5755 14083
rect 5796 14049 5830 14083
rect 5871 14049 5905 14083
rect 5189 13977 5223 14011
rect 5265 13977 5299 14011
rect 5341 13977 5375 14011
rect 5417 13977 5451 14011
rect 5493 13977 5527 14011
rect 5569 13977 5603 14011
rect 5645 13977 5679 14011
rect 5721 13977 5755 14011
rect 5796 13977 5830 14011
rect 5871 13977 5905 14011
rect 5219 12634 5253 12668
rect 5287 12634 5321 12668
rect 1197 12457 1231 12491
rect 1197 12386 1231 12420
rect 5219 12535 5253 12569
rect 5287 12535 5321 12569
rect 5764 12634 5798 12668
rect 5832 12634 5866 12668
rect 5764 12535 5798 12569
rect 5832 12535 5866 12569
rect 5219 12435 5253 12469
rect 5287 12435 5321 12469
rect 5764 12435 5798 12469
rect 5832 12435 5866 12469
rect 9399 14051 9433 14085
rect 9472 14051 9506 14085
rect 9545 14051 9579 14085
rect 9618 14051 9652 14085
rect 9691 14051 9725 14085
rect 9763 14051 9797 14085
rect 9835 14051 9869 14085
rect 9495 13978 9529 14012
rect 9563 13978 9597 14012
rect 9631 13978 9665 14012
rect 9699 13978 9733 14012
rect 9767 13978 9801 14012
rect 9835 13978 9869 14012
rect 9365 13944 9399 13978
rect 9365 13876 9399 13910
rect 9869 13873 9903 13907
rect 9365 13808 9399 13842
rect 9365 13740 9399 13774
rect 9365 13672 9399 13706
rect 9365 13604 9399 13638
rect 9365 13536 9399 13570
rect 9365 13468 9399 13502
rect 9365 13400 9399 13434
rect 9365 13332 9399 13366
rect 9365 13264 9399 13298
rect 9365 13196 9399 13230
rect 9365 13128 9399 13162
rect 9365 13060 9399 13094
rect 9365 12992 9399 13026
rect 9365 12924 9399 12958
rect 9869 13805 9903 13839
rect 9869 13737 9903 13771
rect 9869 13669 9903 13703
rect 9869 13601 9903 13635
rect 9869 13533 9903 13567
rect 9869 13465 9903 13499
rect 9869 13397 9903 13431
rect 9869 13329 9903 13363
rect 9869 13261 9903 13295
rect 9869 13193 9903 13227
rect 9869 13125 9903 13159
rect 9869 13057 9903 13091
rect 9869 12989 9903 13023
rect 9869 12921 9903 12955
rect 9869 12853 9903 12887
rect 9869 12785 9903 12819
rect 9399 12751 9433 12785
rect 9467 12751 9501 12785
rect 9535 12751 9569 12785
rect 9603 12751 9637 12785
rect 9671 12751 9705 12785
rect 9739 12751 9773 12785
rect 9419 12656 9453 12690
rect 9487 12656 9521 12690
rect 9747 12656 9781 12690
rect 9815 12656 9849 12690
rect 9419 12583 9453 12617
rect 9487 12583 9521 12617
rect 9747 12583 9781 12617
rect 9815 12583 9849 12617
rect 9419 12509 9453 12543
rect 9487 12509 9521 12543
rect 9747 12509 9781 12543
rect 9815 12509 9849 12543
rect 9419 12435 9453 12469
rect 9487 12435 9521 12469
rect 9747 12435 9781 12469
rect 9815 12435 9849 12469
rect 11077 14166 11111 14200
rect 11077 14098 11111 14132
rect 11077 14030 11111 14064
rect 11077 13962 11111 13996
rect 11077 13894 11111 13928
rect 11077 13826 11111 13860
rect 11077 13758 11111 13792
rect 11077 13690 11111 13724
rect 11077 13622 11111 13656
rect 11077 13554 11111 13588
rect 11077 13486 11111 13520
rect 11077 13418 11111 13452
rect 11077 13350 11111 13384
rect 11077 13282 11111 13316
rect 11077 13214 11111 13248
rect 11077 13086 11111 13120
rect 11077 13016 11111 13050
rect 11077 12946 11111 12980
rect 11077 12876 11111 12910
rect 11077 12806 11111 12840
rect 11077 12736 11111 12770
rect 11077 12666 11111 12700
rect 11077 12596 11111 12630
rect 11077 12526 11111 12560
rect 11077 12456 11111 12490
rect 11077 12386 11111 12420
rect 1299 12352 1333 12386
rect 1367 12352 1401 12386
rect 1435 12352 1469 12386
rect 1503 12352 1537 12386
rect 1571 12352 1605 12386
rect 1639 12352 1673 12386
rect 1707 12352 1741 12386
rect 1775 12352 1809 12386
rect 1843 12352 1877 12386
rect 1911 12352 1945 12386
rect 1979 12352 2013 12386
rect 2047 12352 2081 12386
rect 2115 12352 2149 12386
rect 2183 12352 2217 12386
rect 2251 12352 2285 12386
rect 2319 12352 2353 12386
rect 2387 12352 2421 12386
rect 2455 12352 2489 12386
rect 2523 12352 2557 12386
rect 2591 12352 2625 12386
rect 2659 12352 2693 12386
rect 2727 12352 2761 12386
rect 2795 12352 2829 12386
rect 2863 12352 2897 12386
rect 2931 12352 2965 12386
rect 2999 12352 3033 12386
rect 3067 12352 3101 12386
rect 3135 12352 3169 12386
rect 3203 12352 3237 12386
rect 3271 12352 3305 12386
rect 3339 12352 3373 12386
rect 3407 12352 3441 12386
rect 3475 12352 3509 12386
rect 3543 12352 3577 12386
rect 3611 12352 3645 12386
rect 3679 12352 3713 12386
rect 3747 12352 3781 12386
rect 3815 12352 3849 12386
rect 3883 12352 3917 12386
rect 3951 12352 3985 12386
rect 4019 12352 4053 12386
rect 4087 12352 4121 12386
rect 4155 12352 4189 12386
rect 4223 12352 4257 12386
rect 4291 12352 4325 12386
rect 4359 12352 4393 12386
rect 4427 12352 4461 12386
rect 4495 12352 4529 12386
rect 4563 12352 4597 12386
rect 4631 12352 4665 12386
rect 4699 12352 4733 12386
rect 4767 12352 4801 12386
rect 4835 12352 4869 12386
rect 4903 12352 4937 12386
rect 4971 12352 5005 12386
rect 5039 12352 5073 12386
rect 5107 12352 5141 12386
rect 5175 12352 5209 12386
rect 5243 12352 5277 12386
rect 5311 12352 5345 12386
rect 5379 12352 5413 12386
rect 5447 12352 5481 12386
rect 5515 12352 5549 12386
rect 5583 12352 5617 12386
rect 5651 12352 5685 12386
rect 5719 12352 5753 12386
rect 5787 12352 5821 12386
rect 5855 12352 5889 12386
rect 5923 12352 5957 12386
rect 5991 12352 6025 12386
rect 6059 12352 6093 12386
rect 6127 12352 6161 12386
rect 6195 12352 6229 12386
rect 6263 12352 6297 12386
rect 6331 12352 6365 12386
rect 6399 12352 6433 12386
rect 6467 12352 6501 12386
rect 6535 12352 6569 12386
rect 6603 12352 6637 12386
rect 6671 12352 6705 12386
rect 6739 12352 6773 12386
rect 6807 12352 6841 12386
rect 6875 12352 6909 12386
rect 6943 12352 6977 12386
rect 7011 12352 7045 12386
rect 7079 12352 7113 12386
rect 7147 12352 7181 12386
rect 7215 12352 7249 12386
rect 7283 12352 7317 12386
rect 7351 12352 7385 12386
rect 7419 12352 7453 12386
rect 7487 12352 7521 12386
rect 7555 12352 7589 12386
rect 7623 12352 7657 12386
rect 7691 12352 7725 12386
rect 7759 12352 7793 12386
rect 7827 12352 7861 12386
rect 7895 12352 7929 12386
rect 7963 12352 7997 12386
rect 8031 12352 8065 12386
rect 8099 12352 8133 12386
rect 8167 12352 8201 12386
rect 8235 12352 8269 12386
rect 8303 12352 8337 12386
rect 8371 12352 8405 12386
rect 8439 12352 8473 12386
rect 8507 12352 8541 12386
rect 8575 12352 8609 12386
rect 8643 12352 8677 12386
rect 8711 12352 8745 12386
rect 8779 12352 8813 12386
rect 8847 12352 8881 12386
rect 8915 12352 8949 12386
rect 8983 12352 9017 12386
rect 9052 12352 9086 12386
rect 9121 12352 9155 12386
rect 9190 12352 9224 12386
rect 9259 12352 9293 12386
rect 9328 12352 9362 12386
rect 9397 12352 9431 12386
rect 9466 12352 9500 12386
rect 9535 12352 9569 12386
rect 9604 12352 9638 12386
rect 9673 12352 9707 12386
rect 9742 12352 9776 12386
rect 9811 12352 9845 12386
rect 9880 12352 9914 12386
rect 9949 12352 9983 12386
rect 10018 12352 10052 12386
rect 10087 12352 10121 12386
rect 10156 12352 10190 12386
rect 10225 12352 10259 12386
rect 10294 12352 10328 12386
rect 10363 12352 10397 12386
rect 10432 12352 10466 12386
rect 10501 12352 10535 12386
rect 10583 12352 10617 12386
rect 10659 12352 10693 12386
rect 10735 12352 10769 12386
rect 10811 12352 10845 12386
rect 10886 12352 10920 12386
rect 10961 12352 10995 12386
rect 1117 11665 1151 11699
rect 1219 11689 1321 11723
rect 1355 11689 1389 11723
rect 1423 11689 1457 11723
rect 1491 11689 1525 11723
rect 1559 11689 1593 11723
rect 1627 11689 1661 11723
rect 1695 11689 1729 11723
rect 1763 11689 1797 11723
rect 1831 11689 1865 11723
rect 1899 11689 1933 11723
rect 1967 11689 2001 11723
rect 2035 11689 2069 11723
rect 2103 11689 2137 11723
rect 2171 11689 2205 11723
rect 2239 11689 2273 11723
rect 2307 11689 2341 11723
rect 2375 11689 2409 11723
rect 2443 11689 2477 11723
rect 2511 11689 2545 11723
rect 2579 11689 2613 11723
rect 2647 11689 2681 11723
rect 2715 11689 2749 11723
rect 2841 11689 2875 11723
rect 2909 11689 2943 11723
rect 2977 11689 3011 11723
rect 3045 11689 3079 11723
rect 3113 11689 3147 11723
rect 3181 11689 3215 11723
rect 3249 11689 3283 11723
rect 3317 11689 3351 11723
rect 3385 11689 3419 11723
rect 3453 11689 3487 11723
rect 3521 11689 3555 11723
rect 3589 11689 3623 11723
rect 3657 11689 3691 11723
rect 3725 11689 3759 11723
rect 3793 11689 3827 11723
rect 3861 11689 3895 11723
rect 3929 11689 3963 11723
rect 3997 11689 4031 11723
rect 4065 11689 4099 11723
rect 4133 11689 4167 11723
rect 4201 11689 4235 11723
rect 4269 11689 4303 11723
rect 4337 11689 4371 11723
rect 4405 11689 4439 11723
rect 4473 11689 4507 11723
rect 4541 11689 4575 11723
rect 4609 11689 4643 11723
rect 4677 11689 4711 11723
rect 4745 11689 4779 11723
rect 4813 11689 4847 11723
rect 4881 11689 4915 11723
rect 4949 11689 4983 11723
rect 5017 11689 5051 11723
rect 5085 11689 5119 11723
rect 5153 11689 5187 11723
rect 5221 11689 5255 11723
rect 5289 11689 5323 11723
rect 5357 11689 5391 11723
rect 5425 11689 5459 11723
rect 5688 11689 5722 11723
rect 5756 11689 5790 11723
rect 5824 11689 5858 11723
rect 5892 11689 5926 11723
rect 5960 11689 5994 11723
rect 6028 11689 6062 11723
rect 6096 11689 6130 11723
rect 6164 11689 6198 11723
rect 6232 11689 6266 11723
rect 6300 11689 6334 11723
rect 6368 11689 6402 11723
rect 6436 11689 6470 11723
rect 6504 11689 6538 11723
rect 6572 11689 6606 11723
rect 6640 11689 6674 11723
rect 6708 11689 6742 11723
rect 6776 11689 6810 11723
rect 6844 11689 6878 11723
rect 6912 11689 6946 11723
rect 6980 11689 7014 11723
rect 7048 11689 7082 11723
rect 7116 11689 7150 11723
rect 7184 11689 7218 11723
rect 7252 11689 7286 11723
rect 7320 11689 7354 11723
rect 7388 11689 7422 11723
rect 7456 11689 7490 11723
rect 7524 11689 7558 11723
rect 7592 11689 7626 11723
rect 7660 11689 7694 11723
rect 7728 11689 7762 11723
rect 7796 11689 7830 11723
rect 7923 11689 7957 11723
rect 7991 11689 8025 11723
rect 8059 11689 8093 11723
rect 8127 11689 8161 11723
rect 8195 11689 8229 11723
rect 8263 11689 8297 11723
rect 8331 11689 8365 11723
rect 8399 11689 8433 11723
rect 8467 11689 8501 11723
rect 8535 11689 8569 11723
rect 8603 11689 8637 11723
rect 8671 11689 8705 11723
rect 8739 11689 8773 11723
rect 8807 11689 8841 11723
rect 8875 11689 8909 11723
rect 8943 11689 8977 11723
rect 9011 11689 9045 11723
rect 9079 11689 9113 11723
rect 9147 11689 9181 11723
rect 9215 11689 9249 11723
rect 9283 11689 9317 11723
rect 9351 11689 9385 11723
rect 9419 11689 9453 11723
rect 9487 11689 9521 11723
rect 9555 11689 9589 11723
rect 9623 11689 9657 11723
rect 9691 11689 9725 11723
rect 9759 11689 9793 11723
rect 9827 11689 9861 11723
rect 9895 11689 9929 11723
rect 1219 11655 1287 11689
rect 1117 11281 1287 11655
rect 3717 11621 3751 11655
rect 3717 11553 3751 11587
rect 3717 11485 3751 11519
rect 3717 11417 3751 11451
rect 1117 6963 1219 11281
rect 1253 11212 1287 11246
rect 3717 11349 3751 11383
rect 5557 11655 5591 11689
rect 5557 11587 5591 11621
rect 5557 11519 5591 11553
rect 5557 11451 5591 11485
rect 5557 11383 5591 11417
rect 3717 11281 3751 11315
rect 1253 11143 1287 11177
rect 1253 11074 1287 11108
rect 1253 11005 1287 11039
rect 1253 10936 1287 10970
rect 1253 10867 1287 10901
rect 1253 10798 1287 10832
rect 1253 10729 1287 10763
rect 1253 10660 1287 10694
rect 1253 10591 1287 10625
rect 1253 10522 1287 10556
rect 1253 10453 1287 10487
rect 3717 11213 3751 11247
rect 3717 11145 3751 11179
rect 3717 11077 3751 11111
rect 3717 11009 3751 11043
rect 3717 10941 3751 10975
rect 3717 10873 3751 10907
rect 3717 10805 3751 10839
rect 3717 10737 3751 10771
rect 3717 10669 3751 10703
rect 3717 10601 3751 10635
rect 3717 10533 3751 10567
rect 3717 10465 3751 10499
rect 1253 10384 1287 10418
rect 1253 10315 1287 10349
rect 1253 10246 1287 10280
rect 1253 10177 1287 10211
rect 3717 10397 3751 10431
rect 3717 10329 3751 10363
rect 3717 10261 3751 10295
rect 3717 10193 3751 10227
rect 1253 10108 1287 10142
rect 1253 10039 1287 10073
rect 1253 9970 1287 10004
rect 1253 9901 1287 9935
rect 1253 9832 1287 9866
rect 1253 9763 1287 9797
rect 1253 9694 1287 9728
rect 1253 9625 1287 9659
rect 1253 9556 1287 9590
rect 1253 9487 1287 9521
rect 1253 9418 1287 9452
rect 1253 9349 1287 9383
rect 3717 10125 3751 10159
rect 3717 10057 3751 10091
rect 3717 9989 3751 10023
rect 3717 9921 3751 9955
rect 3717 9853 3751 9887
rect 3717 9785 3751 9819
rect 3717 9717 3751 9751
rect 3717 9649 3751 9683
rect 3717 9581 3751 9615
rect 3717 9513 3751 9547
rect 3717 9445 3751 9479
rect 3717 9377 3751 9411
rect 1253 9280 1287 9314
rect 3717 9309 3751 9343
rect 1253 9211 1287 9245
rect 1253 9142 1287 9176
rect 1253 9073 1287 9107
rect 1253 9004 1287 9038
rect 1253 8935 1287 8969
rect 1253 8866 1287 8900
rect 1253 8797 1287 8831
rect 1253 8728 1287 8762
rect 1253 8659 1287 8693
rect 1253 8590 1287 8624
rect 1253 8521 1287 8555
rect 3717 9241 3751 9275
rect 3717 9173 3751 9207
rect 3717 9105 3751 9139
rect 3717 9037 3751 9071
rect 3717 8969 3751 9003
rect 3717 8901 3751 8935
rect 3717 8833 3751 8867
rect 3717 8765 3751 8799
rect 3717 8697 3751 8731
rect 3717 8629 3751 8663
rect 3717 8561 3751 8595
rect 1253 8452 1287 8486
rect 1253 8383 1287 8417
rect 1253 8314 1287 8348
rect 1253 8245 1287 8279
rect 3717 8493 3751 8527
rect 3717 8425 3751 8459
rect 3717 8357 3751 8391
rect 3717 8289 3751 8323
rect 1253 8176 1287 8210
rect 1253 8107 1287 8141
rect 1253 8038 1287 8072
rect 1253 7969 1287 8003
rect 1253 7900 1287 7934
rect 1253 7831 1287 7865
rect 1253 7762 1287 7796
rect 1253 7693 1287 7727
rect 1253 7624 1287 7658
rect 1253 7555 1287 7589
rect 1253 7486 1287 7520
rect 1253 7417 1287 7451
rect 3717 8221 3751 8255
rect 3717 8153 3751 8187
rect 3717 8085 3751 8119
rect 3717 8017 3751 8051
rect 3717 7949 3751 7983
rect 3717 7881 3751 7915
rect 3717 7813 3751 7847
rect 3717 7745 3751 7779
rect 3717 7677 3751 7711
rect 3717 7609 3751 7643
rect 3717 7541 3751 7575
rect 3717 7473 3751 7507
rect 1253 7348 1287 7382
rect 1253 7279 1287 7313
rect 3717 7405 3751 7439
rect 3717 7337 3751 7371
rect 3717 7269 3751 7303
rect 1253 7210 1287 7244
rect 1253 7141 1287 7175
rect 1253 7072 1287 7106
rect 1253 7003 1287 7037
rect 3717 7201 3751 7235
rect 3717 7133 3751 7167
rect 3717 7065 3751 7099
rect 3717 6997 3751 7031
rect 1117 3913 1287 6963
rect 1321 6929 1355 6963
rect 1389 6929 1423 6963
rect 1457 6929 1491 6963
rect 1525 6929 1559 6963
rect 1593 6929 1627 6963
rect 1661 6929 1695 6963
rect 1729 6929 1763 6963
rect 1797 6929 1831 6963
rect 1865 6929 1899 6963
rect 1933 6929 1967 6963
rect 2001 6929 2035 6963
rect 2069 6929 2103 6963
rect 2137 6929 2171 6963
rect 2205 6929 2239 6963
rect 2273 6929 2307 6963
rect 2341 6929 2375 6963
rect 2409 6929 2443 6963
rect 2477 6929 2511 6963
rect 2545 6929 2579 6963
rect 2613 6929 2647 6963
rect 2681 6929 2715 6963
rect 2749 6929 2783 6963
rect 2817 6929 2851 6963
rect 2885 6929 2919 6963
rect 2953 6929 2987 6963
rect 3021 6929 3055 6963
rect 3089 6929 3123 6963
rect 3157 6929 3191 6963
rect 3225 6929 3259 6963
rect 3293 6929 3327 6963
rect 3361 6929 3395 6963
rect 3429 6929 3463 6963
rect 3497 6929 3531 6963
rect 3565 6929 3599 6963
rect 3633 6929 3667 6963
rect 3717 6929 3751 6963
rect 3717 6861 3751 6895
rect 3717 6793 3751 6827
rect 3717 6725 3751 6759
rect 3717 6657 3751 6691
rect 3717 6589 3751 6623
rect 3717 6521 3751 6555
rect 3717 6453 3751 6487
rect 3717 6385 3751 6419
rect 3717 6317 3751 6351
rect 3717 6249 3751 6283
rect 3717 6181 3751 6215
rect 3717 6113 3751 6147
rect 3717 6045 3751 6079
rect 3717 5977 3751 6011
rect 3717 5909 3751 5943
rect 3717 5841 3751 5875
rect 3717 5773 3751 5807
rect 3717 5705 3751 5739
rect 3717 5637 3751 5671
rect 3717 5569 3751 5603
rect 3717 5501 3751 5535
rect 3717 5433 3751 5467
rect 3717 5365 3751 5399
rect 3717 5297 3751 5331
rect 3717 5229 3751 5263
rect 3717 5161 3751 5195
rect 3717 5093 3751 5127
rect 3717 5025 3751 5059
rect 3717 4957 3751 4991
rect 3717 4889 3751 4923
rect 3717 4821 3751 4855
rect 3717 4753 3751 4787
rect 3717 4685 3751 4719
rect 3717 4617 3751 4651
rect 3717 4549 3751 4583
rect 1117 3844 1151 3878
rect 1117 3775 1151 3809
rect 1117 3706 1151 3740
rect 1117 3637 1151 3671
rect 1117 3568 1151 3602
rect 1117 3499 1151 3533
rect 1117 3430 1151 3464
rect 1117 3361 1151 3395
rect 1117 3292 1151 3326
rect 1117 3223 1151 3257
rect 1117 3154 1151 3188
rect 1117 3085 1151 3119
rect 1117 3016 1151 3050
rect 1117 2947 1151 2981
rect 1117 2878 1151 2912
rect 1117 2809 1151 2843
rect 1117 2740 1151 2774
rect 1117 2671 1151 2705
rect 1117 2602 1151 2636
rect 1185 2577 1287 3913
rect 3717 4481 3751 4515
rect 3717 4413 3751 4447
rect 3717 4345 3751 4379
rect 3717 4277 3751 4311
rect 3717 4209 3751 4243
rect 3717 4141 3751 4175
rect 3717 4073 3751 4107
rect 3717 4005 3751 4039
rect 3717 3937 3751 3971
rect 7397 11621 7431 11655
rect 7397 11553 7431 11587
rect 7397 11485 7431 11519
rect 7397 11417 7431 11451
rect 9929 11621 9963 11655
rect 9929 11553 9963 11587
rect 9929 11485 9963 11519
rect 9929 11417 9963 11451
rect 5557 11315 5591 11349
rect 5557 11247 5591 11281
rect 5557 11179 5591 11213
rect 5557 11111 5591 11145
rect 5557 11043 5591 11077
rect 5557 10975 5591 11009
rect 5557 10907 5591 10941
rect 5557 10839 5591 10873
rect 5557 10771 5591 10805
rect 5557 10703 5591 10737
rect 5557 10635 5591 10669
rect 5557 10567 5591 10601
rect 5557 10499 5591 10533
rect 5557 10431 5591 10465
rect 5557 10363 5591 10397
rect 5557 10295 5591 10329
rect 5557 10227 5591 10261
rect 5557 10159 5591 10193
rect 5557 10091 5591 10125
rect 5557 10023 5591 10057
rect 5557 9955 5591 9989
rect 5557 9887 5591 9921
rect 5557 9819 5591 9853
rect 5557 9751 5591 9785
rect 5557 9683 5591 9717
rect 5557 9615 5591 9649
rect 5557 9547 5591 9581
rect 5557 9479 5591 9513
rect 5557 9411 5591 9445
rect 5557 9343 5591 9377
rect 5557 9275 5591 9309
rect 5557 9207 5591 9241
rect 5557 9139 5591 9173
rect 5557 9071 5591 9105
rect 5557 9003 5591 9037
rect 5557 8935 5591 8969
rect 5557 8867 5591 8901
rect 5557 8799 5591 8833
rect 5557 8731 5591 8765
rect 5557 8663 5591 8697
rect 5557 8595 5591 8629
rect 5557 8527 5591 8561
rect 5557 8459 5591 8493
rect 5557 8391 5591 8425
rect 5557 8323 5591 8357
rect 5557 8255 5591 8289
rect 5557 8187 5591 8221
rect 5557 8119 5591 8153
rect 5557 8051 5591 8085
rect 5557 7983 5591 8017
rect 5557 7915 5591 7949
rect 5557 7847 5591 7881
rect 5557 7779 5591 7813
rect 5557 7711 5591 7745
rect 5557 7643 5591 7677
rect 5557 7575 5591 7609
rect 5557 7507 5591 7541
rect 5557 7439 5591 7473
rect 5557 7371 5591 7405
rect 5557 7303 5591 7337
rect 5557 7235 5591 7269
rect 5557 7167 5591 7201
rect 5557 7099 5591 7133
rect 5557 7031 5591 7065
rect 5557 6963 5591 6997
rect 5557 6895 5591 6929
rect 5557 6827 5591 6861
rect 5557 6759 5591 6793
rect 5557 6691 5591 6725
rect 5557 6623 5591 6657
rect 5557 6555 5591 6589
rect 5557 6487 5591 6521
rect 5557 6419 5591 6453
rect 5557 6351 5591 6385
rect 5557 6283 5591 6317
rect 5557 6215 5591 6249
rect 5557 6147 5591 6181
rect 5557 6079 5591 6113
rect 5557 6011 5591 6045
rect 5557 5943 5591 5977
rect 5557 5875 5591 5909
rect 5557 5807 5591 5841
rect 5557 5739 5591 5773
rect 5557 5671 5591 5705
rect 5557 5603 5591 5637
rect 5557 5535 5591 5569
rect 5557 5467 5591 5501
rect 5557 5399 5591 5433
rect 5557 5331 5591 5365
rect 5557 5263 5591 5297
rect 5557 5195 5591 5229
rect 5557 5127 5591 5161
rect 5557 5059 5591 5093
rect 5557 4991 5591 5025
rect 5557 4923 5591 4957
rect 5557 4855 5591 4889
rect 5557 4787 5591 4821
rect 5557 4719 5591 4753
rect 5557 4651 5591 4685
rect 5557 4583 5591 4617
rect 5557 4515 5591 4549
rect 5557 4447 5591 4481
rect 5557 4379 5591 4413
rect 5557 4311 5591 4345
rect 5557 4243 5591 4277
rect 5557 4175 5591 4209
rect 5557 4107 5591 4141
rect 5557 4039 5591 4073
rect 5557 3971 5591 4005
rect 3717 3869 3751 3903
rect 3717 3801 3751 3835
rect 3717 3733 3751 3767
rect 3717 3665 3751 3699
rect 5557 3903 5591 3937
rect 7397 11349 7431 11383
rect 7397 11281 7431 11315
rect 7397 11213 7431 11247
rect 9929 11349 9963 11383
rect 9929 11281 9963 11315
rect 7397 11145 7431 11179
rect 7397 11077 7431 11111
rect 7397 11009 7431 11043
rect 7397 10941 7431 10975
rect 7397 10873 7431 10907
rect 7397 10805 7431 10839
rect 7397 10737 7431 10771
rect 7397 10669 7431 10703
rect 7397 10601 7431 10635
rect 7397 10533 7431 10567
rect 7397 10465 7431 10499
rect 9929 11213 9963 11247
rect 9929 11145 9963 11179
rect 9929 11077 9963 11111
rect 9929 11009 9963 11043
rect 9929 10941 9963 10975
rect 9929 10873 9963 10907
rect 9929 10805 9963 10839
rect 9929 10737 9963 10771
rect 9929 10669 9963 10703
rect 9929 10601 9963 10635
rect 9929 10533 9963 10567
rect 9929 10465 9963 10499
rect 7397 10397 7431 10431
rect 7397 10329 7431 10363
rect 7397 10261 7431 10295
rect 7397 10193 7431 10227
rect 7397 10125 7431 10159
rect 9929 10397 9963 10431
rect 9929 10329 9963 10363
rect 9929 10261 9963 10295
rect 9929 10193 9963 10227
rect 7397 10057 7431 10091
rect 7397 9989 7431 10023
rect 7397 9921 7431 9955
rect 7397 9853 7431 9887
rect 7397 9785 7431 9819
rect 7397 9717 7431 9751
rect 7397 9649 7431 9683
rect 7397 9581 7431 9615
rect 7397 9513 7431 9547
rect 7397 9445 7431 9479
rect 7397 9377 7431 9411
rect 9929 10125 9963 10159
rect 9929 10057 9963 10091
rect 9929 9989 9963 10023
rect 9929 9921 9963 9955
rect 9929 9853 9963 9887
rect 9929 9785 9963 9819
rect 9929 9717 9963 9751
rect 9929 9649 9963 9683
rect 9929 9581 9963 9615
rect 9929 9513 9963 9547
rect 9929 9445 9963 9479
rect 9929 9377 9963 9411
rect 7397 9309 7431 9343
rect 9929 9309 9963 9343
rect 7397 9241 7431 9275
rect 7397 9173 7431 9207
rect 7397 9105 7431 9139
rect 7397 9037 7431 9071
rect 7397 8969 7431 9003
rect 7397 8901 7431 8935
rect 7397 8833 7431 8867
rect 7397 8765 7431 8799
rect 7397 8697 7431 8731
rect 7397 8629 7431 8663
rect 7397 8561 7431 8595
rect 7397 8493 7431 8527
rect 9929 9241 9963 9275
rect 9929 9173 9963 9207
rect 9929 9105 9963 9139
rect 9929 9037 9963 9071
rect 9929 8969 9963 9003
rect 9929 8901 9963 8935
rect 9929 8833 9963 8867
rect 9929 8765 9963 8799
rect 9929 8697 9963 8731
rect 9929 8629 9963 8663
rect 9929 8561 9963 8595
rect 7397 8425 7431 8459
rect 7397 8357 7431 8391
rect 7397 8289 7431 8323
rect 7397 8221 7431 8255
rect 9929 8493 9963 8527
rect 9929 8425 9963 8459
rect 9929 8357 9963 8391
rect 9929 8289 9963 8323
rect 9929 8221 9963 8255
rect 7397 8153 7431 8187
rect 7397 8085 7431 8119
rect 7397 8017 7431 8051
rect 7397 7949 7431 7983
rect 7397 7881 7431 7915
rect 7397 7813 7431 7847
rect 7397 7745 7431 7779
rect 7397 7677 7431 7711
rect 7397 7609 7431 7643
rect 7397 7541 7431 7575
rect 7397 7473 7431 7507
rect 7397 7405 7431 7439
rect 9929 8153 9963 8187
rect 9929 8085 9963 8119
rect 9929 8017 9963 8051
rect 9997 8006 10031 8040
rect 10065 8006 10099 8040
rect 10133 8006 10167 8040
rect 10201 8006 10235 8040
rect 10269 8006 10303 8040
rect 10337 8006 10371 8040
rect 10405 8006 10439 8040
rect 10473 8006 10507 8040
rect 10541 8006 10575 8040
rect 10609 8006 10643 8040
rect 10677 8006 10711 8040
rect 10745 8006 10779 8040
rect 10813 8006 10847 8040
rect 10881 8006 10915 8040
rect 10949 8006 10983 8040
rect 11017 8006 11051 8040
rect 11085 8006 11119 8040
rect 11153 8006 11187 8040
rect 11221 8006 11255 8040
rect 11289 8006 11323 8040
rect 11357 8006 11391 8040
rect 11425 8006 11459 8040
rect 11493 8006 11527 8040
rect 11561 8006 11595 8040
rect 11629 8006 11663 8040
rect 11697 8006 11731 8040
rect 11765 8006 11799 8040
rect 11833 8006 11867 8040
rect 11901 8006 11935 8040
rect 11969 8006 12003 8040
rect 12037 8006 12071 8040
rect 12105 8006 12139 8040
rect 12173 8006 12207 8040
rect 12241 8006 12275 8040
rect 12309 8006 12343 8040
rect 12377 8006 12411 8040
rect 12445 8006 12479 8040
rect 12513 8006 12547 8040
rect 12581 8006 12615 8040
rect 12649 8006 12683 8040
rect 12717 8006 12751 8040
rect 12785 8006 12819 8040
rect 12853 8006 12887 8040
rect 12921 8006 12955 8040
rect 12989 8006 13023 8040
rect 9929 7949 9963 7983
rect 9929 7881 9963 7915
rect 9929 7813 9963 7847
rect 9929 7745 9963 7779
rect 9929 7677 9963 7711
rect 13069 7972 13103 8006
rect 13069 7904 13103 7938
rect 13069 7836 13103 7870
rect 13069 7768 13103 7802
rect 9929 7609 9963 7643
rect 9929 7541 9963 7575
rect 9929 7473 9963 7507
rect 7397 7337 7431 7371
rect 7397 7269 7431 7303
rect 9929 7405 9963 7439
rect 9929 7337 9963 7371
rect 9929 7269 9963 7303
rect 7397 7201 7431 7235
rect 7397 7133 7431 7167
rect 7397 7065 7431 7099
rect 7397 6997 7431 7031
rect 9929 7201 9963 7235
rect 9929 7133 9963 7167
rect 9929 7065 9963 7099
rect 9929 6997 9963 7031
rect 7397 6929 7431 6963
rect 7481 6929 7515 6963
rect 7549 6929 7583 6963
rect 7617 6929 7651 6963
rect 7685 6929 7719 6963
rect 7753 6929 7787 6963
rect 7821 6929 7855 6963
rect 7889 6929 7923 6963
rect 7957 6929 7991 6963
rect 8025 6929 8059 6963
rect 8093 6929 8127 6963
rect 8161 6929 8195 6963
rect 8229 6929 8263 6963
rect 8297 6929 8331 6963
rect 8365 6929 8399 6963
rect 8433 6929 8467 6963
rect 8501 6929 8535 6963
rect 8569 6929 8603 6963
rect 8637 6929 8671 6963
rect 8705 6929 8739 6963
rect 8773 6929 8807 6963
rect 8841 6929 8875 6963
rect 8909 6929 8943 6963
rect 8977 6929 9011 6963
rect 9045 6929 9079 6963
rect 9113 6929 9147 6963
rect 9181 6929 9215 6963
rect 9249 6929 9283 6963
rect 9317 6929 9351 6963
rect 9385 6929 9419 6963
rect 9453 6929 9487 6963
rect 9521 6929 9555 6963
rect 9589 6929 9623 6963
rect 9657 6929 9691 6963
rect 9725 6929 9759 6963
rect 9793 6929 9827 6963
rect 9861 6929 9895 6963
rect 9929 6929 9963 6963
rect 7397 6861 7431 6895
rect 7397 6793 7431 6827
rect 7397 6725 7431 6759
rect 7397 6657 7431 6691
rect 9929 6861 9963 6895
rect 9929 6793 9963 6827
rect 9929 6725 9963 6759
rect 9929 6657 9963 6691
rect 7397 6589 7431 6623
rect 7397 6521 7431 6555
rect 7397 6453 7431 6487
rect 9929 6589 9963 6623
rect 9929 6521 9963 6555
rect 7397 6385 7431 6419
rect 7397 6317 7431 6351
rect 7397 6249 7431 6283
rect 7397 6181 7431 6215
rect 7397 6113 7431 6147
rect 7397 6045 7431 6079
rect 7397 5977 7431 6011
rect 7397 5909 7431 5943
rect 7397 5841 7431 5875
rect 7397 5773 7431 5807
rect 7397 5705 7431 5739
rect 7397 5637 7431 5671
rect 9929 6453 9963 6487
rect 9929 6385 9963 6419
rect 9929 6317 9963 6351
rect 9929 6249 9963 6283
rect 9929 6181 9963 6215
rect 9929 6113 9963 6147
rect 9929 6045 9963 6079
rect 9929 5977 9963 6011
rect 9929 5909 9963 5943
rect 9929 5841 9963 5875
rect 9929 5773 9963 5807
rect 9929 5705 9963 5739
rect 7397 5569 7431 5603
rect 7397 5501 7431 5535
rect 7397 5433 7431 5467
rect 7397 5365 7431 5399
rect 9929 5637 9963 5671
rect 9929 5569 9963 5603
rect 9929 5501 9963 5535
rect 9929 5433 9963 5467
rect 7397 5297 7431 5331
rect 7397 5229 7431 5263
rect 7397 5161 7431 5195
rect 7397 5093 7431 5127
rect 7397 5025 7431 5059
rect 7397 4957 7431 4991
rect 7397 4889 7431 4923
rect 7397 4821 7431 4855
rect 7397 4753 7431 4787
rect 7397 4685 7431 4719
rect 7397 4617 7431 4651
rect 9929 5365 9963 5399
rect 9929 5297 9963 5331
rect 9929 5229 9963 5263
rect 9929 5161 9963 5195
rect 9929 5093 9963 5127
rect 9929 5025 9963 5059
rect 9929 4957 9963 4991
rect 9929 4889 9963 4923
rect 9929 4821 9963 4855
rect 9929 4753 9963 4787
rect 9929 4685 9963 4719
rect 9929 4617 9963 4651
rect 7397 4549 7431 4583
rect 9929 4549 9963 4583
rect 7397 4481 7431 4515
rect 7397 4413 7431 4447
rect 7397 4345 7431 4379
rect 7397 4277 7431 4311
rect 7397 4209 7431 4243
rect 7397 4141 7431 4175
rect 7397 4073 7431 4107
rect 7397 4005 7431 4039
rect 7397 3937 7431 3971
rect 5557 3835 5591 3869
rect 5557 3767 5591 3801
rect 7397 3869 7431 3903
rect 7397 3801 7431 3835
rect 7397 3733 7431 3767
rect 9929 4481 9963 4515
rect 9929 4413 9963 4447
rect 9929 4345 9963 4379
rect 9929 4277 9963 4311
rect 9929 4209 9963 4243
rect 9929 4141 9963 4175
rect 9929 4073 9963 4107
rect 9929 4005 9963 4039
rect 9929 3937 9963 3971
rect 9929 3869 9963 3903
rect 9929 3801 9963 3835
rect 3785 3653 3819 3687
rect 3853 3653 3887 3687
rect 3921 3653 3955 3687
rect 3989 3653 4023 3687
rect 4057 3653 4091 3687
rect 4125 3653 4159 3687
rect 4193 3653 4227 3687
rect 4261 3653 4295 3687
rect 4329 3653 4363 3687
rect 4397 3653 4431 3687
rect 4465 3653 4499 3687
rect 4533 3653 4567 3687
rect 4601 3653 4635 3687
rect 4669 3653 4703 3687
rect 4737 3653 4771 3687
rect 4805 3653 4839 3687
rect 4873 3653 4907 3687
rect 4941 3653 4975 3687
rect 5009 3653 5043 3687
rect 5077 3653 5111 3687
rect 5145 3653 5179 3687
rect 5213 3653 5247 3687
rect 5281 3653 5315 3687
rect 5349 3653 5383 3687
rect 5417 3653 5451 3687
rect 5485 3653 5519 3687
rect 5625 3653 5659 3687
rect 5693 3653 5727 3687
rect 5761 3653 5795 3687
rect 5829 3653 5863 3687
rect 5897 3653 5931 3687
rect 5965 3653 5999 3687
rect 6033 3653 6067 3687
rect 6101 3653 6135 3687
rect 6169 3653 6203 3687
rect 6237 3653 6271 3687
rect 6305 3653 6339 3687
rect 6373 3653 6407 3687
rect 6441 3653 6475 3687
rect 6509 3653 6543 3687
rect 6577 3653 6611 3687
rect 6645 3653 6679 3687
rect 6713 3653 6747 3687
rect 6781 3653 6815 3687
rect 6849 3653 6883 3687
rect 6917 3653 6951 3687
rect 6985 3653 7019 3687
rect 7053 3653 7087 3687
rect 7121 3653 7155 3687
rect 7189 3653 7223 3687
rect 7257 3653 7291 3687
rect 7325 3653 7359 3687
rect 7397 3665 7431 3699
rect 3717 3597 3751 3631
rect 3717 3529 3751 3563
rect 3717 3461 3751 3495
rect 3717 3393 3751 3427
rect 7397 3597 7431 3631
rect 7397 3529 7431 3563
rect 7397 3461 7431 3495
rect 9929 3733 9963 3767
rect 9929 3665 9963 3699
rect 9929 3597 9963 3631
rect 9929 3529 9963 3563
rect 9929 3461 9963 3495
rect 7397 3393 7431 3427
rect 3717 3325 3751 3359
rect 3717 3257 3751 3291
rect 3717 3189 3751 3223
rect 3717 3121 3751 3155
rect 3717 3053 3751 3087
rect 3717 2985 3751 3019
rect 3717 2917 3751 2951
rect 3717 2849 3751 2883
rect 3717 2781 3751 2815
rect 3717 2713 3751 2747
rect 1117 2533 1151 2567
rect 1185 2509 1219 2543
rect 1253 2508 1287 2542
rect 3717 2645 3751 2679
rect 3717 2577 3751 2611
rect 3717 2509 3751 2543
rect 1117 2464 1151 2498
rect 1185 2441 1219 2475
rect 1253 2439 1287 2473
rect 1117 2395 1151 2429
rect 1185 2373 1219 2407
rect 1253 2370 1287 2404
rect 1117 2326 1151 2360
rect 1185 2305 1219 2339
rect 1253 2301 1287 2335
rect 1117 2257 1151 2291
rect 1185 2237 1219 2271
rect 1253 2232 1287 2266
rect 1117 2188 1151 2222
rect 3717 2441 3751 2475
rect 3717 2373 3751 2407
rect 3717 2305 3751 2339
rect 3717 2237 3751 2271
rect 1185 2169 1219 2203
rect 1253 2163 1287 2197
rect 1371 2169 1405 2203
rect 1439 2169 1473 2203
rect 1507 2169 1541 2203
rect 1575 2169 1609 2203
rect 1643 2169 1677 2203
rect 1711 2169 1745 2203
rect 1779 2169 1813 2203
rect 1847 2169 1881 2203
rect 1915 2169 1949 2203
rect 1983 2169 2017 2203
rect 2051 2169 2085 2203
rect 2119 2169 2153 2203
rect 2187 2169 2221 2203
rect 2255 2169 2289 2203
rect 2323 2169 2357 2203
rect 2391 2169 2425 2203
rect 2459 2169 2493 2203
rect 2527 2169 2561 2203
rect 2595 2169 2629 2203
rect 2663 2169 2697 2203
rect 2731 2169 2765 2203
rect 2799 2169 2833 2203
rect 2867 2169 2901 2203
rect 2935 2169 2969 2203
rect 3003 2169 3037 2203
rect 3071 2169 3105 2203
rect 3139 2169 3173 2203
rect 3207 2169 3241 2203
rect 3275 2169 3309 2203
rect 3343 2169 3377 2203
rect 3411 2169 3445 2203
rect 3479 2169 3513 2203
rect 3547 2169 3581 2203
rect 3615 2169 3649 2203
rect 3683 2169 3717 2203
rect 1117 2119 1151 2153
rect 1185 2101 1219 2135
rect 1253 2094 1287 2128
rect 1117 2050 1151 2084
rect 1185 2033 1219 2067
rect 1253 2025 1287 2059
rect 1117 1981 1151 2015
rect 1185 1965 1219 1999
rect 1253 1956 1287 1990
rect 1117 1912 1151 1946
rect 1185 1897 1219 1931
rect 1253 1887 1287 1921
rect 7397 3325 7431 3359
rect 7397 3257 7431 3291
rect 7397 3189 7431 3223
rect 7397 3121 7431 3155
rect 7397 3053 7431 3087
rect 7397 2985 7431 3019
rect 7397 2917 7431 2951
rect 7397 2849 7431 2883
rect 7397 2781 7431 2815
rect 7397 2713 7431 2747
rect 7397 2645 7431 2679
rect 9929 3393 9963 3427
rect 9929 3325 9963 3359
rect 9929 3257 9963 3291
rect 9929 3189 9963 3223
rect 9929 3121 9963 3155
rect 9929 3053 9963 3087
rect 9929 2985 9963 3019
rect 9929 2917 9963 2951
rect 9929 2849 9963 2883
rect 9929 2781 9963 2815
rect 9929 2713 9963 2747
rect 7397 2577 7431 2611
rect 7397 2509 7431 2543
rect 9929 2645 9963 2679
rect 9929 2577 9963 2611
rect 9929 2509 9963 2543
rect 7397 2441 7431 2475
rect 7397 2373 7431 2407
rect 7397 2305 7431 2339
rect 7397 2237 7431 2271
rect 9929 2441 9963 2475
rect 9929 2373 9963 2407
rect 9929 2305 9963 2339
rect 9929 2237 9963 2271
rect 7431 2169 7465 2203
rect 7499 2169 7533 2203
rect 7567 2169 7601 2203
rect 7635 2169 7669 2203
rect 7703 2169 7737 2203
rect 7771 2169 7805 2203
rect 7839 2169 7873 2203
rect 7907 2169 7941 2203
rect 7975 2169 8009 2203
rect 8043 2169 8077 2203
rect 8111 2169 8145 2203
rect 8179 2169 8213 2203
rect 8247 2169 8281 2203
rect 8315 2169 8349 2203
rect 8383 2169 8417 2203
rect 8451 2169 8485 2203
rect 8519 2169 8553 2203
rect 8587 2169 8621 2203
rect 8655 2169 8689 2203
rect 8723 2169 8757 2203
rect 8791 2169 8825 2203
rect 8859 2169 8893 2203
rect 8927 2169 8961 2203
rect 8995 2169 9029 2203
rect 9063 2169 9097 2203
rect 9131 2169 9165 2203
rect 9199 2169 9233 2203
rect 9267 2169 9301 2203
rect 9335 2169 9369 2203
rect 9403 2169 9437 2203
rect 9471 2169 9505 2203
rect 9539 2169 9573 2203
rect 9607 2169 9641 2203
rect 9675 2169 9709 2203
rect 9743 2169 9777 2203
rect 9811 2169 9845 2203
rect 9929 2169 9963 2203
rect 1117 1843 1151 1877
rect 1185 1829 1219 1863
rect 1253 1818 1287 1852
rect 1117 1774 1151 1808
rect 1185 1761 1219 1795
rect 1253 1749 1287 1783
rect 9929 2101 9963 2135
rect 9929 2033 9963 2067
rect 9929 1965 9963 1999
rect 9929 1897 9963 1931
rect 1117 1705 1151 1739
rect 1185 1693 1219 1727
rect 1253 1680 1287 1714
rect 1117 1636 1151 1670
rect 1185 1625 1219 1659
rect 1253 1611 1287 1645
rect 1117 1567 1151 1601
rect 1185 1557 1219 1591
rect 1253 1542 1287 1576
rect 1117 1498 1151 1532
rect 1185 1489 1219 1523
rect 1253 1473 1287 1507
rect 1117 1429 1151 1463
rect 1185 1421 1219 1455
rect 1253 1404 1287 1438
rect 1117 1360 1151 1394
rect 1185 1353 1219 1387
rect 1253 1335 1287 1369
rect 1117 1291 1151 1325
rect 1185 1285 1219 1319
rect 1253 1266 1287 1300
rect 1117 1222 1151 1256
rect 1185 1217 1219 1251
rect 1253 1197 1287 1231
rect 1117 1153 1151 1187
rect 1185 1149 1219 1183
rect 1253 1128 1287 1162
rect 1117 1084 1151 1118
rect 1185 1081 1219 1115
rect 1253 1059 1287 1093
rect 1117 1015 1151 1049
rect 1185 1013 1219 1047
rect 1253 990 1287 1024
rect 1117 946 1151 980
rect 1185 945 1219 979
rect 9929 1829 9963 1863
rect 9929 1761 9963 1795
rect 1253 921 1287 955
rect 1117 877 1151 911
rect 1185 877 1219 911
rect 1253 852 1287 886
rect 1117 808 1151 842
rect 1185 809 1219 843
rect 1253 783 1287 817
rect 1117 739 1151 773
rect 1185 741 1219 775
rect 1253 714 1287 748
rect 1117 670 1151 704
rect 1185 673 1219 707
rect 1253 645 1287 679
rect 1117 601 1151 635
rect 1185 605 1219 639
rect 1253 576 1287 610
rect 9929 1693 9963 1727
rect 9929 1625 9963 1659
rect 9929 1557 9963 1591
rect 9929 1489 9963 1523
rect 9929 1421 9963 1455
rect 9929 1353 9963 1387
rect 9929 1285 9963 1319
rect 9929 1217 9963 1251
rect 9929 1149 9963 1183
rect 9929 1081 9963 1115
rect 9929 1013 9963 1047
rect 1117 532 1151 566
rect 1185 537 1219 571
rect 1253 507 1287 541
rect 1117 463 1151 497
rect 1185 469 1219 503
rect 1253 438 1287 472
rect 9929 945 9963 979
rect 9929 877 9963 911
rect 9929 809 9963 843
rect 9929 741 9963 775
rect 9929 673 9963 707
rect 9929 605 9963 639
rect 9929 537 9963 571
rect 9929 469 9963 503
rect 1117 394 1151 428
rect 1185 401 1219 435
rect 1253 369 1287 403
rect 1117 325 1151 359
rect 1185 333 1219 367
rect 1253 300 1287 334
rect 1117 256 1151 290
rect 1185 265 1219 299
rect 1253 231 1287 265
rect 1117 187 1151 221
rect 1185 197 1219 231
rect 13069 7700 13103 7734
rect 13069 7632 13103 7666
rect 13069 7564 13103 7598
rect 13069 7496 13103 7530
rect 13069 7428 13103 7462
rect 13069 7360 13103 7394
rect 13069 7292 13103 7326
rect 13069 7224 13103 7258
rect 13069 7156 13103 7190
rect 13069 7088 13103 7122
rect 13069 7020 13103 7054
rect 13069 6952 13103 6986
rect 13069 6884 13103 6918
rect 13069 6816 13103 6850
rect 13069 6748 13103 6782
rect 13069 6680 13103 6714
rect 13069 6612 13103 6646
rect 13069 6544 13103 6578
rect 13069 6476 13103 6510
rect 13069 6408 13103 6442
rect 13069 6340 13103 6374
rect 13069 6272 13103 6306
rect 13069 6204 13103 6238
rect 13069 6136 13103 6170
rect 13069 6068 13103 6102
rect 13069 6000 13103 6034
rect 13069 5932 13103 5966
rect 13069 5864 13103 5898
rect 13069 5796 13103 5830
rect 13069 5728 13103 5762
rect 13069 5660 13103 5694
rect 13069 5592 13103 5626
rect 13069 5524 13103 5558
rect 13069 5456 13103 5490
rect 13069 5388 13103 5422
rect 13069 5320 13103 5354
rect 13069 5252 13103 5286
rect 13069 5184 13103 5218
rect 13069 5116 13103 5150
rect 13069 5048 13103 5082
rect 13069 4980 13103 5014
rect 13069 4912 13103 4946
rect 13069 4844 13103 4878
rect 13069 4776 13103 4810
rect 13069 4708 13103 4742
rect 13069 4640 13103 4674
rect 13069 4572 13103 4606
rect 13069 4504 13103 4538
rect 13069 4436 13103 4470
rect 13069 4368 13103 4402
rect 13069 4300 13103 4334
rect 13069 4232 13103 4266
rect 13069 4164 13103 4198
rect 13069 4096 13103 4130
rect 13069 4028 13103 4062
rect 13069 3960 13103 3994
rect 13069 3892 13103 3926
rect 13069 3824 13103 3858
rect 13069 3756 13103 3790
rect 13069 3688 13103 3722
rect 13069 3620 13103 3654
rect 13069 3552 13103 3586
rect 13069 3484 13103 3518
rect 13069 3416 13103 3450
rect 13069 3348 13103 3382
rect 13069 3280 13103 3314
rect 13069 3212 13103 3246
rect 13069 3144 13103 3178
rect 13069 3076 13103 3110
rect 13069 3008 13103 3042
rect 13069 2940 13103 2974
rect 13069 2872 13103 2906
rect 13069 2804 13103 2838
rect 13069 2736 13103 2770
rect 13069 2668 13103 2702
rect 13069 2600 13103 2634
rect 13069 2532 13103 2566
rect 13069 2464 13103 2498
rect 13069 2396 13103 2430
rect 13069 2328 13103 2362
rect 13069 2260 13103 2294
rect 13069 2192 13103 2226
rect 13069 2124 13103 2158
rect 13069 2056 13103 2090
rect 13069 1988 13103 2022
rect 13069 1920 13103 1954
rect 13069 1852 13103 1886
rect 13069 1784 13103 1818
rect 13069 1716 13103 1750
rect 13069 1648 13103 1682
rect 13069 1580 13103 1614
rect 13069 1512 13103 1546
rect 13069 1444 13103 1478
rect 13069 1376 13103 1410
rect 13069 1308 13103 1342
rect 13069 1240 13103 1274
rect 13069 1172 13103 1206
rect 13069 1104 13103 1138
rect 13069 1036 13103 1070
rect 13069 968 13103 1002
rect 13069 900 13103 934
rect 13069 832 13103 866
rect 13069 764 13103 798
rect 13069 696 13103 730
rect 13069 628 13103 662
rect 13069 560 13103 594
rect 13069 492 13103 526
rect 9929 401 9963 435
rect 9929 333 9963 367
rect 9929 265 9963 299
rect 9929 197 9963 231
rect 13069 424 13103 458
rect 13069 356 13103 390
rect 13069 288 13103 322
rect 1282 163 1316 197
rect 1350 163 1384 197
rect 1418 163 1452 197
rect 1486 163 1520 197
rect 1554 163 1588 197
rect 1622 163 1656 197
rect 1690 163 1724 197
rect 1758 163 1792 197
rect 1826 163 1860 197
rect 1894 163 1928 197
rect 1962 163 1996 197
rect 2030 163 2064 197
rect 2098 163 2132 197
rect 2166 163 2200 197
rect 2234 163 2268 197
rect 2302 163 2336 197
rect 2370 163 2404 197
rect 2438 163 2472 197
rect 2506 163 2540 197
rect 2574 163 2608 197
rect 2642 163 2676 197
rect 2710 163 2744 197
rect 2778 163 2812 197
rect 2846 163 2880 197
rect 2914 163 2948 197
rect 2982 163 3016 197
rect 3050 163 3084 197
rect 3118 163 3152 197
rect 3186 163 3220 197
rect 3254 163 3288 197
rect 3322 163 3356 197
rect 3390 163 3424 197
rect 3458 163 3492 197
rect 3526 163 3560 197
rect 3594 163 3628 197
rect 3662 163 3696 197
rect 3730 163 3764 197
rect 3798 163 3832 197
rect 3866 163 3900 197
rect 3934 163 3968 197
rect 4002 163 4036 197
rect 4070 163 4104 197
rect 4138 163 4172 197
rect 4206 163 4240 197
rect 4274 163 4308 197
rect 4342 163 4376 197
rect 4410 163 4444 197
rect 4478 163 4512 197
rect 4546 163 4580 197
rect 4614 163 4648 197
rect 4682 163 4716 197
rect 4750 163 4784 197
rect 4818 163 4852 197
rect 4886 163 4920 197
rect 4954 163 4988 197
rect 5022 163 5056 197
rect 5090 163 5124 197
rect 5158 163 5192 197
rect 5226 163 5260 197
rect 5294 163 5328 197
rect 5362 163 5396 197
rect 5430 163 5464 197
rect 5498 163 5532 197
rect 5566 163 5600 197
rect 5668 163 5702 197
rect 5736 163 5770 197
rect 5804 163 5838 197
rect 5872 163 5906 197
rect 5940 163 5974 197
rect 6008 163 6042 197
rect 6076 163 6110 197
rect 6144 163 6178 197
rect 6212 163 6246 197
rect 6280 163 6314 197
rect 6348 163 6382 197
rect 6416 163 6450 197
rect 6484 163 6518 197
rect 6552 163 6586 197
rect 6620 163 6654 197
rect 6688 163 6722 197
rect 6756 163 6790 197
rect 6824 163 6858 197
rect 6892 163 6926 197
rect 6960 163 6994 197
rect 7028 163 7062 197
rect 7096 163 7130 197
rect 7164 163 7198 197
rect 7232 163 7266 197
rect 7300 163 7334 197
rect 7368 163 7402 197
rect 7436 163 7470 197
rect 7504 163 7538 197
rect 7572 163 7606 197
rect 7640 163 7674 197
rect 7708 163 7742 197
rect 7776 163 7810 197
rect 7844 163 7878 197
rect 7912 163 7946 197
rect 7980 163 8014 197
rect 8048 163 8082 197
rect 8116 163 8150 197
rect 8184 163 8218 197
rect 8252 163 8286 197
rect 8320 163 8354 197
rect 8388 163 8422 197
rect 8456 163 8490 197
rect 8524 163 8558 197
rect 8592 163 8626 197
rect 8660 163 8694 197
rect 8728 163 8762 197
rect 8796 163 8830 197
rect 8864 163 8898 197
rect 8932 163 8966 197
rect 9000 163 9034 197
rect 9068 163 9102 197
rect 9136 163 9170 197
rect 9204 163 9238 197
rect 9272 163 9306 197
rect 9340 163 9374 197
rect 9408 163 9442 197
rect 9476 163 9510 197
rect 9544 163 9578 197
rect 9612 163 9646 197
rect 9680 163 9714 197
rect 9748 163 9782 197
rect 9816 163 9850 197
rect 10043 163 10077 197
rect 10111 163 10145 197
rect 10179 163 10213 197
rect 10247 163 10281 197
rect 10315 163 10349 197
rect 10383 163 10417 197
rect 10451 163 10485 197
rect 10519 163 10553 197
rect 10587 163 10621 197
rect 10655 163 10689 197
rect 10723 163 10757 197
rect 10791 163 10825 197
rect 10859 163 10893 197
rect 10927 163 10961 197
rect 10995 163 11029 197
rect 11063 163 11097 197
rect 11131 163 11165 197
rect 11199 163 11233 197
rect 11267 163 11301 197
rect 11335 163 11369 197
rect 11403 163 11437 197
rect 11471 163 11505 197
rect 11539 163 11573 197
rect 11607 163 11641 197
rect 11675 163 11709 197
rect 11743 163 11777 197
rect 11811 163 11845 197
rect 11879 163 11913 197
rect 11947 163 11981 197
rect 12015 163 12049 197
rect 12083 163 12117 197
rect 12151 163 12185 197
rect 12219 163 12253 197
rect 12287 163 12321 197
rect 12355 163 12389 197
rect 12423 163 12457 197
rect 12491 163 12525 197
rect 12559 163 12593 197
rect 12627 163 12661 197
rect 12695 163 12729 197
rect 12763 163 12797 197
rect 12831 163 12865 197
rect 12899 163 12933 197
rect 12967 163 13001 197
rect 13035 163 13069 197
<< poly >>
rect 1741 14077 1813 14093
rect 1741 14043 1757 14077
rect 1791 14043 1813 14077
rect 1741 14007 1813 14043
rect 1741 13973 1757 14007
rect 1791 13973 1813 14007
rect 1741 13937 1813 13973
rect 1741 13903 1757 13937
rect 1791 13903 1813 13937
rect 1741 13867 1813 13903
rect 1741 13833 1757 13867
rect 1791 13833 1813 13867
rect 1741 13797 1813 13833
rect 1741 13763 1757 13797
rect 1791 13763 1813 13797
rect 1741 13727 1813 13763
rect 1741 13693 1757 13727
rect 1791 13693 1813 13727
rect 1741 13657 1813 13693
rect 1741 13623 1757 13657
rect 1791 13623 1813 13657
rect 1741 13587 1813 13623
rect 1741 13553 1757 13587
rect 1791 13553 1813 13587
rect 1741 13517 1813 13553
rect 1741 13483 1757 13517
rect 1791 13483 1813 13517
rect 1741 13447 1813 13483
rect 1741 13413 1757 13447
rect 1791 13413 1813 13447
rect 1741 13377 1813 13413
rect 1741 13343 1757 13377
rect 1791 13343 1813 13377
rect 1741 13307 1813 13343
rect 1741 13273 1757 13307
rect 1791 13273 1813 13307
rect 1741 13237 1813 13273
rect 1741 13203 1757 13237
rect 1791 13203 1813 13237
rect 1741 13167 1813 13203
rect 1741 13133 1757 13167
rect 1791 13133 1813 13167
rect 1741 13097 1813 13133
rect 1741 13063 1757 13097
rect 1791 13063 1813 13097
rect 1741 13027 1813 13063
rect 1741 12993 1757 13027
rect 1791 12993 1813 13027
rect 1741 12957 1813 12993
rect 1741 12923 1757 12957
rect 1791 12923 1813 12957
rect 1741 12888 1813 12923
rect 1741 12854 1757 12888
rect 1791 12854 1813 12888
rect 1741 12819 1813 12854
rect 1741 12785 1757 12819
rect 1791 12785 1813 12819
rect 1741 12750 1813 12785
rect 1741 12716 1757 12750
rect 1791 12716 1813 12750
rect 1741 12681 1813 12716
rect 1741 12647 1757 12681
rect 1791 12647 1813 12681
rect 1741 12612 1813 12647
rect 1741 12578 1757 12612
rect 1791 12578 1813 12612
rect 1741 12543 1813 12578
rect 1741 12509 1757 12543
rect 1791 12509 1813 12543
rect 1741 12493 1813 12509
rect 3265 14077 3337 14093
rect 3265 14043 3287 14077
rect 3321 14043 3337 14077
rect 3265 14007 3337 14043
rect 3265 13973 3287 14007
rect 3321 13973 3337 14007
rect 3265 13937 3337 13973
rect 4229 14047 4295 14063
rect 4229 14013 4245 14047
rect 4279 14013 4295 14047
rect 4229 13979 4295 14013
rect 3265 13903 3287 13937
rect 3321 13903 3337 13937
rect 3265 13867 3337 13903
rect 3265 13833 3287 13867
rect 3321 13833 3337 13867
rect 3391 13953 3457 13969
rect 3391 13919 3407 13953
rect 3441 13919 3457 13953
rect 3391 13885 3457 13919
rect 3391 13851 3407 13885
rect 3441 13851 3457 13885
rect 3391 13835 3457 13851
rect 4121 13953 4187 13969
rect 4121 13919 4137 13953
rect 4171 13919 4187 13953
rect 4229 13945 4245 13979
rect 4279 13945 4295 13979
rect 4229 13929 4295 13945
rect 4959 14047 5025 14063
rect 4959 14013 4975 14047
rect 5009 14013 5025 14047
rect 4959 13979 5025 14013
rect 4959 13945 4975 13979
rect 5009 13945 5025 13979
rect 7745 14077 7817 14093
rect 6069 14047 6135 14063
rect 6069 14013 6085 14047
rect 6119 14013 6135 14047
rect 7745 14043 7761 14077
rect 7795 14043 7817 14077
rect 6069 13979 6135 14013
rect 4959 13929 5025 13945
rect 6069 13945 6085 13979
rect 6119 13945 6135 13979
rect 4121 13885 4187 13919
rect 4121 13851 4137 13885
rect 4171 13851 4187 13885
rect 5268 13921 5836 13937
rect 6069 13929 6135 13945
rect 6819 13929 6862 14029
rect 7745 14007 7817 14043
rect 7745 13973 7761 14007
rect 7795 13973 7817 14007
rect 6907 13953 6973 13969
rect 5268 13887 5284 13921
rect 5318 13887 5356 13921
rect 5390 13887 5428 13921
rect 5462 13887 5500 13921
rect 5534 13887 5572 13921
rect 5606 13887 5644 13921
rect 5678 13887 5715 13921
rect 5749 13887 5786 13921
rect 5820 13887 5836 13921
rect 4121 13835 4187 13851
rect 4229 13850 4275 13873
rect 4979 13850 5025 13873
rect 5268 13871 5836 13887
rect 6907 13919 6923 13953
rect 6957 13919 6973 13953
rect 6907 13885 6973 13919
rect 3265 13797 3337 13833
rect 3265 13763 3287 13797
rect 3321 13763 3337 13797
rect 4229 13834 4295 13850
rect 4229 13800 4245 13834
rect 4279 13800 4295 13834
rect 3265 13727 3337 13763
rect 3265 13693 3287 13727
rect 3321 13693 3337 13727
rect 3265 13657 3337 13693
rect 3265 13623 3287 13657
rect 3321 13623 3337 13657
rect 3265 13587 3337 13623
rect 3265 13553 3287 13587
rect 3321 13553 3337 13587
rect 3391 13756 3437 13779
rect 4141 13756 4187 13779
rect 3391 13740 3457 13756
rect 3391 13706 3407 13740
rect 3441 13706 3457 13740
rect 3391 13652 3457 13706
rect 3391 13618 3407 13652
rect 3441 13618 3457 13652
rect 3391 13602 3457 13618
rect 4121 13740 4187 13756
rect 4121 13706 4137 13740
rect 4171 13706 4187 13740
rect 4121 13652 4187 13706
rect 4229 13746 4295 13800
rect 4229 13712 4245 13746
rect 4279 13712 4295 13746
rect 4229 13696 4295 13712
rect 4959 13834 5025 13850
rect 6069 13850 6115 13873
rect 6819 13850 6865 13873
rect 4959 13800 4975 13834
rect 5009 13800 5025 13834
rect 4959 13746 5025 13800
rect 4959 13712 4975 13746
rect 5009 13712 5025 13746
rect 4959 13696 5025 13712
rect 4229 13673 4275 13696
rect 4979 13673 5025 13696
rect 4121 13618 4137 13652
rect 4171 13618 4187 13652
rect 4121 13602 4187 13618
rect 3391 13579 3437 13602
rect 4141 13579 4187 13602
rect 4229 13594 4275 13617
rect 4979 13594 5025 13617
rect 3265 13517 3337 13553
rect 4229 13578 4295 13594
rect 4229 13544 4245 13578
rect 4279 13544 4295 13578
rect 3265 13483 3287 13517
rect 3321 13483 3337 13517
rect 3265 13447 3337 13483
rect 3265 13413 3287 13447
rect 3321 13413 3337 13447
rect 3265 13377 3337 13413
rect 3265 13343 3287 13377
rect 3321 13343 3337 13377
rect 3265 13307 3337 13343
rect 3391 13500 3437 13523
rect 4141 13500 4187 13523
rect 3391 13484 3457 13500
rect 3391 13450 3407 13484
rect 3441 13450 3457 13484
rect 3391 13396 3457 13450
rect 3391 13362 3407 13396
rect 3441 13362 3457 13396
rect 3391 13346 3457 13362
rect 4121 13484 4187 13500
rect 4121 13450 4137 13484
rect 4171 13450 4187 13484
rect 4121 13396 4187 13450
rect 4229 13490 4295 13544
rect 4229 13456 4245 13490
rect 4279 13456 4295 13490
rect 4229 13440 4295 13456
rect 4959 13578 5025 13594
rect 4959 13544 4975 13578
rect 5009 13544 5025 13578
rect 4959 13490 5025 13544
rect 4959 13456 4975 13490
rect 5009 13456 5025 13490
rect 4959 13440 5025 13456
rect 4229 13417 4275 13440
rect 4979 13417 5025 13440
rect 4121 13362 4137 13396
rect 4171 13362 4187 13396
rect 4121 13346 4187 13362
rect 3391 13323 3437 13346
rect 4141 13323 4187 13346
rect 4229 13338 4275 13361
rect 4979 13338 5025 13361
rect 3265 13273 3287 13307
rect 3321 13273 3337 13307
rect 3265 13237 3337 13273
rect 4229 13322 4295 13338
rect 4229 13288 4245 13322
rect 4279 13288 4295 13322
rect 3265 13203 3287 13237
rect 3321 13203 3337 13237
rect 3265 13167 3337 13203
rect 3265 13133 3287 13167
rect 3321 13133 3337 13167
rect 3265 13097 3337 13133
rect 3265 13063 3287 13097
rect 3321 13063 3337 13097
rect 3391 13244 3437 13267
rect 4141 13244 4187 13267
rect 3391 13228 3457 13244
rect 3391 13194 3407 13228
rect 3441 13194 3457 13228
rect 3391 13140 3457 13194
rect 3391 13106 3407 13140
rect 3441 13106 3457 13140
rect 3391 13090 3457 13106
rect 4121 13228 4187 13244
rect 4121 13194 4137 13228
rect 4171 13194 4187 13228
rect 4121 13140 4187 13194
rect 4229 13234 4295 13288
rect 4229 13200 4245 13234
rect 4279 13200 4295 13234
rect 4229 13184 4295 13200
rect 4959 13322 5025 13338
rect 4959 13288 4975 13322
rect 5009 13288 5025 13322
rect 4959 13234 5025 13288
rect 4959 13200 4975 13234
rect 5009 13200 5025 13234
rect 4959 13184 5025 13200
rect 4229 13161 4275 13184
rect 4979 13161 5025 13184
rect 4121 13106 4137 13140
rect 4171 13106 4187 13140
rect 4121 13090 4187 13106
rect 3391 13067 3437 13090
rect 4141 13067 4187 13090
rect 4229 13082 4275 13105
rect 3265 13027 3337 13063
rect 3265 12993 3287 13027
rect 3321 12993 3337 13027
rect 4229 13066 4295 13082
rect 4979 13081 5025 13105
rect 4229 13032 4245 13066
rect 4279 13032 4295 13066
rect 3265 12957 3337 12993
rect 3265 12923 3287 12957
rect 3321 12923 3337 12957
rect 3265 12888 3337 12923
rect 3265 12854 3287 12888
rect 3321 12854 3337 12888
rect 3265 12819 3337 12854
rect 3265 12785 3287 12819
rect 3321 12785 3337 12819
rect 3391 12988 3437 13011
rect 4141 12988 4187 13011
rect 3391 12972 3457 12988
rect 3391 12938 3407 12972
rect 3441 12938 3457 12972
rect 3391 12884 3457 12938
rect 3391 12850 3407 12884
rect 3441 12850 3457 12884
rect 3391 12834 3457 12850
rect 4121 12972 4187 12988
rect 4121 12938 4137 12972
rect 4171 12938 4187 12972
rect 4121 12884 4187 12938
rect 4229 12978 4295 13032
rect 4229 12944 4245 12978
rect 4279 12944 4295 12978
rect 4229 12928 4295 12944
rect 4959 13065 5025 13081
rect 4959 13031 4975 13065
rect 5009 13031 5025 13065
rect 4959 12977 5025 13031
rect 4959 12943 4975 12977
rect 5009 12943 5025 12977
rect 4229 12905 4275 12928
rect 4959 12927 5025 12943
rect 4979 12905 5025 12927
rect 4121 12850 4137 12884
rect 4171 12850 4187 12884
rect 4121 12834 4187 12850
rect 3391 12811 3437 12834
rect 4141 12811 4187 12834
rect 4229 12826 4275 12849
rect 4979 12826 5025 12849
rect 6069 13834 6135 13850
rect 6069 13800 6085 13834
rect 6119 13800 6135 13834
rect 6069 13746 6135 13800
rect 6069 13712 6085 13746
rect 6119 13712 6135 13746
rect 6069 13696 6135 13712
rect 6799 13834 6865 13850
rect 6907 13851 6923 13885
rect 6957 13851 6973 13885
rect 6907 13835 6973 13851
rect 7637 13953 7703 13969
rect 7637 13919 7653 13953
rect 7687 13919 7703 13953
rect 7637 13885 7703 13919
rect 7637 13851 7653 13885
rect 7687 13851 7703 13885
rect 7637 13835 7703 13851
rect 7745 13937 7817 13973
rect 7745 13903 7761 13937
rect 7795 13903 7817 13937
rect 7745 13867 7817 13903
rect 6799 13800 6815 13834
rect 6849 13800 6865 13834
rect 6799 13746 6865 13800
rect 7745 13833 7761 13867
rect 7795 13833 7817 13867
rect 7745 13797 7817 13833
rect 6799 13712 6815 13746
rect 6849 13712 6865 13746
rect 6799 13696 6865 13712
rect 6069 13673 6115 13696
rect 6819 13673 6865 13696
rect 6907 13756 6953 13779
rect 7657 13756 7703 13779
rect 6907 13740 6973 13756
rect 6907 13706 6923 13740
rect 6957 13706 6973 13740
rect 6907 13652 6973 13706
rect 6907 13618 6923 13652
rect 6957 13618 6973 13652
rect 6069 13594 6115 13617
rect 6819 13594 6865 13617
rect 6069 13578 6135 13594
rect 6069 13544 6085 13578
rect 6119 13544 6135 13578
rect 6069 13490 6135 13544
rect 6069 13456 6085 13490
rect 6119 13456 6135 13490
rect 6069 13440 6135 13456
rect 6799 13578 6865 13594
rect 6907 13602 6973 13618
rect 7637 13740 7703 13756
rect 7637 13706 7653 13740
rect 7687 13706 7703 13740
rect 7637 13652 7703 13706
rect 7637 13618 7653 13652
rect 7687 13618 7703 13652
rect 7637 13602 7703 13618
rect 6907 13579 6953 13602
rect 7657 13579 7703 13602
rect 7745 13763 7761 13797
rect 7795 13763 7817 13797
rect 7745 13727 7817 13763
rect 7745 13693 7761 13727
rect 7795 13693 7817 13727
rect 7745 13657 7817 13693
rect 7745 13623 7761 13657
rect 7795 13623 7817 13657
rect 7745 13587 7817 13623
rect 6799 13544 6815 13578
rect 6849 13544 6865 13578
rect 6799 13490 6865 13544
rect 7745 13553 7761 13587
rect 7795 13553 7817 13587
rect 6799 13456 6815 13490
rect 6849 13456 6865 13490
rect 6799 13440 6865 13456
rect 6069 13417 6115 13440
rect 6819 13417 6865 13440
rect 6907 13500 6953 13523
rect 7657 13500 7703 13523
rect 6907 13484 6973 13500
rect 6907 13450 6923 13484
rect 6957 13450 6973 13484
rect 6907 13396 6973 13450
rect 6907 13362 6923 13396
rect 6957 13362 6973 13396
rect 6069 13338 6115 13361
rect 6819 13338 6865 13361
rect 6069 13322 6135 13338
rect 6069 13288 6085 13322
rect 6119 13288 6135 13322
rect 6069 13234 6135 13288
rect 6069 13200 6085 13234
rect 6119 13200 6135 13234
rect 6069 13184 6135 13200
rect 6799 13322 6865 13338
rect 6907 13346 6973 13362
rect 7637 13484 7703 13500
rect 7637 13450 7653 13484
rect 7687 13450 7703 13484
rect 7637 13396 7703 13450
rect 7637 13362 7653 13396
rect 7687 13362 7703 13396
rect 7637 13346 7703 13362
rect 6907 13323 6953 13346
rect 7657 13323 7703 13346
rect 7745 13517 7817 13553
rect 7745 13483 7761 13517
rect 7795 13483 7817 13517
rect 7745 13447 7817 13483
rect 7745 13413 7761 13447
rect 7795 13413 7817 13447
rect 7745 13377 7817 13413
rect 7745 13343 7761 13377
rect 7795 13343 7817 13377
rect 6799 13288 6815 13322
rect 6849 13288 6865 13322
rect 6799 13234 6865 13288
rect 7745 13307 7817 13343
rect 7745 13273 7761 13307
rect 7795 13273 7817 13307
rect 6799 13200 6815 13234
rect 6849 13200 6865 13234
rect 6799 13184 6865 13200
rect 6069 13161 6115 13184
rect 6819 13161 6865 13184
rect 6907 13244 6953 13267
rect 7657 13244 7703 13267
rect 6907 13228 6973 13244
rect 6907 13194 6923 13228
rect 6957 13194 6973 13228
rect 6907 13140 6973 13194
rect 6907 13106 6923 13140
rect 6957 13106 6973 13140
rect 6069 13082 6115 13105
rect 6069 13066 6135 13082
rect 6819 13081 6865 13105
rect 6069 13032 6085 13066
rect 6119 13032 6135 13066
rect 6069 12978 6135 13032
rect 6069 12944 6085 12978
rect 6119 12944 6135 12978
rect 6069 12928 6135 12944
rect 6799 13065 6865 13081
rect 6907 13090 6973 13106
rect 7637 13228 7703 13244
rect 7637 13194 7653 13228
rect 7687 13194 7703 13228
rect 7637 13140 7703 13194
rect 7637 13106 7653 13140
rect 7687 13106 7703 13140
rect 7637 13090 7703 13106
rect 6907 13067 6953 13090
rect 7657 13067 7703 13090
rect 7745 13237 7817 13273
rect 7745 13203 7761 13237
rect 7795 13203 7817 13237
rect 7745 13167 7817 13203
rect 7745 13133 7761 13167
rect 7795 13133 7817 13167
rect 7745 13097 7817 13133
rect 6799 13031 6815 13065
rect 6849 13031 6865 13065
rect 6799 12977 6865 13031
rect 7745 13063 7761 13097
rect 7795 13063 7817 13097
rect 7745 13027 7817 13063
rect 6799 12943 6815 12977
rect 6849 12943 6865 12977
rect 6069 12905 6115 12928
rect 6799 12927 6865 12943
rect 6819 12905 6865 12927
rect 6907 12988 6953 13011
rect 7657 12988 7703 13011
rect 6907 12972 6973 12988
rect 6907 12938 6923 12972
rect 6957 12938 6973 12972
rect 6907 12884 6973 12938
rect 6907 12850 6923 12884
rect 6957 12850 6973 12884
rect 3265 12750 3337 12785
rect 4229 12810 4295 12826
rect 4229 12776 4245 12810
rect 4279 12776 4295 12810
rect 3265 12716 3287 12750
rect 3321 12716 3337 12750
rect 3265 12681 3337 12716
rect 3265 12647 3287 12681
rect 3321 12647 3337 12681
rect 3265 12612 3337 12647
rect 3391 12739 3457 12755
rect 3391 12705 3407 12739
rect 3441 12705 3457 12739
rect 3391 12671 3457 12705
rect 3391 12637 3407 12671
rect 3441 12637 3457 12671
rect 3391 12621 3457 12637
rect 4121 12739 4187 12755
rect 4121 12705 4137 12739
rect 4171 12705 4187 12739
rect 4121 12671 4187 12705
rect 4121 12637 4137 12671
rect 4171 12637 4187 12671
rect 4229 12722 4295 12776
rect 4229 12688 4245 12722
rect 4279 12688 4295 12722
rect 4229 12672 4295 12688
rect 4959 12810 5025 12826
rect 4959 12776 4975 12810
rect 5009 12776 5025 12810
rect 6069 12826 6115 12849
rect 6819 12826 6865 12849
rect 6069 12810 6135 12826
rect 4959 12722 5025 12776
rect 5257 12791 5837 12807
rect 5257 12757 5273 12791
rect 5307 12757 5347 12791
rect 5381 12757 5421 12791
rect 5455 12757 5495 12791
rect 5529 12757 5568 12791
rect 5602 12757 5641 12791
rect 5675 12757 5714 12791
rect 5748 12757 5787 12791
rect 5821 12757 5837 12791
rect 5257 12741 5837 12757
rect 6069 12776 6085 12810
rect 6119 12776 6135 12810
rect 4959 12688 4975 12722
rect 5009 12688 5025 12722
rect 6069 12722 6135 12776
rect 4959 12672 5025 12688
rect 4229 12649 4275 12672
rect 4979 12649 5025 12672
rect 4121 12621 4187 12637
rect 3265 12578 3287 12612
rect 3321 12578 3337 12612
rect 3265 12543 3337 12578
rect 3265 12509 3287 12543
rect 3321 12509 3337 12543
rect 3265 12493 3337 12509
rect 4229 12577 4295 12593
rect 4229 12543 4245 12577
rect 4279 12543 4295 12577
rect 4229 12509 4295 12543
rect 1402 12458 1602 12480
rect 4229 12475 4245 12509
rect 4279 12475 4295 12509
rect 4229 12459 4295 12475
rect 4959 12577 5025 12593
rect 4959 12543 4975 12577
rect 5009 12543 5025 12577
rect 4959 12509 5025 12543
rect 4959 12475 4975 12509
rect 5009 12475 5025 12509
rect 4959 12459 5025 12475
rect 6069 12688 6085 12722
rect 6119 12688 6135 12722
rect 6069 12672 6135 12688
rect 6799 12810 6865 12826
rect 6907 12834 6973 12850
rect 7637 12972 7703 12988
rect 7637 12938 7653 12972
rect 7687 12938 7703 12972
rect 7637 12884 7703 12938
rect 7637 12850 7653 12884
rect 7687 12850 7703 12884
rect 7637 12834 7703 12850
rect 6907 12811 6953 12834
rect 7657 12811 7703 12834
rect 7745 12993 7761 13027
rect 7795 12993 7817 13027
rect 7745 12957 7817 12993
rect 7745 12923 7761 12957
rect 7795 12923 7817 12957
rect 7745 12888 7817 12923
rect 7745 12854 7761 12888
rect 7795 12854 7817 12888
rect 7745 12819 7817 12854
rect 6799 12776 6815 12810
rect 6849 12776 6865 12810
rect 6799 12722 6865 12776
rect 7745 12785 7761 12819
rect 7795 12785 7817 12819
rect 6799 12688 6815 12722
rect 6849 12688 6865 12722
rect 6799 12672 6865 12688
rect 6069 12649 6115 12672
rect 6819 12649 6865 12672
rect 6907 12739 6973 12755
rect 6907 12705 6923 12739
rect 6957 12705 6973 12739
rect 6907 12671 6973 12705
rect 6907 12637 6923 12671
rect 6957 12637 6973 12671
rect 6907 12621 6973 12637
rect 7637 12739 7703 12755
rect 7637 12705 7653 12739
rect 7687 12705 7703 12739
rect 7637 12671 7703 12705
rect 7637 12637 7653 12671
rect 7687 12637 7703 12671
rect 7637 12621 7703 12637
rect 7745 12750 7817 12785
rect 7745 12716 7761 12750
rect 7795 12716 7817 12750
rect 7745 12681 7817 12716
rect 7745 12647 7761 12681
rect 7795 12647 7817 12681
rect 7745 12612 7817 12647
rect 5503 12474 5603 12480
rect 1402 12424 1422 12458
rect 1456 12424 1552 12458
rect 1586 12424 1602 12458
rect 1402 12408 1602 12424
rect 5486 12458 5620 12474
rect 5486 12424 5502 12458
rect 5536 12424 5570 12458
rect 5604 12424 5620 12458
rect 5486 12408 5620 12424
rect 6799 12577 6865 12593
rect 6799 12543 6815 12577
rect 6849 12543 6865 12577
rect 6799 12509 6865 12543
rect 6799 12475 6815 12509
rect 6849 12475 6865 12509
rect 7745 12578 7761 12612
rect 7795 12578 7817 12612
rect 7745 12543 7817 12578
rect 7745 12509 7761 12543
rect 7795 12509 7817 12543
rect 7745 12493 7817 12509
rect 9269 14077 9341 14093
rect 9269 14043 9291 14077
rect 9325 14043 9341 14077
rect 9269 14007 9341 14043
rect 9269 13973 9291 14007
rect 9325 13973 9341 14007
rect 9269 13937 9341 13973
rect 9269 13903 9291 13937
rect 9325 13903 9341 13937
rect 9269 13867 9341 13903
rect 9269 13833 9291 13867
rect 9325 13833 9341 13867
rect 9269 13797 9341 13833
rect 9269 13763 9291 13797
rect 9325 13763 9341 13797
rect 9269 13727 9341 13763
rect 9269 13693 9291 13727
rect 9325 13693 9341 13727
rect 9269 13657 9341 13693
rect 9269 13623 9291 13657
rect 9325 13623 9341 13657
rect 9269 13587 9341 13623
rect 9269 13553 9291 13587
rect 9325 13553 9341 13587
rect 9269 13517 9341 13553
rect 9269 13483 9291 13517
rect 9325 13483 9341 13517
rect 9269 13447 9341 13483
rect 9269 13413 9291 13447
rect 9325 13413 9341 13447
rect 9269 13377 9341 13413
rect 9269 13343 9291 13377
rect 9325 13343 9341 13377
rect 9269 13307 9341 13343
rect 9269 13273 9291 13307
rect 9325 13273 9341 13307
rect 9269 13237 9341 13273
rect 9269 13203 9291 13237
rect 9325 13203 9341 13237
rect 9269 13167 9341 13203
rect 9269 13133 9291 13167
rect 9325 13133 9341 13167
rect 9269 13097 9341 13133
rect 9269 13063 9291 13097
rect 9325 13063 9341 13097
rect 9269 13027 9341 13063
rect 9269 12993 9291 13027
rect 9325 12993 9341 13027
rect 9269 12957 9341 12993
rect 9269 12923 9291 12957
rect 9325 12923 9341 12957
rect 9269 12888 9341 12923
rect 9269 12854 9291 12888
rect 9325 12854 9341 12888
rect 9269 12819 9341 12854
rect 9269 12785 9291 12819
rect 9325 12785 9341 12819
rect 9269 12750 9341 12785
rect 9269 12716 9291 12750
rect 9325 12716 9341 12750
rect 9269 12681 9341 12716
rect 9269 12647 9291 12681
rect 9325 12647 9341 12681
rect 9269 12612 9341 12647
rect 9269 12578 9291 12612
rect 9325 12578 9341 12612
rect 9269 12543 9341 12578
rect 9269 12509 9291 12543
rect 9325 12509 9341 12543
rect 9269 12493 9341 12509
rect 9506 13921 9762 13937
rect 9506 13887 9522 13921
rect 9556 13887 9617 13921
rect 9651 13887 9712 13921
rect 9746 13887 9762 13921
rect 9506 13871 9762 13887
rect 9506 13865 9606 13871
rect 9662 13865 9762 13871
rect 6799 12459 6865 12475
rect 1380 11224 1446 11240
rect 1380 11190 1396 11224
rect 1430 11190 1446 11224
rect 1380 11151 1446 11190
rect 1380 11117 1396 11151
rect 1430 11117 1446 11151
rect 1380 11078 1446 11117
rect 1380 11044 1396 11078
rect 1430 11044 1446 11078
rect 1380 11005 1446 11044
rect 1380 10971 1396 11005
rect 1430 10971 1446 11005
rect 1380 10932 1446 10971
rect 1380 10898 1396 10932
rect 1430 10898 1446 10932
rect 1380 10859 1446 10898
rect 1380 10825 1396 10859
rect 1430 10825 1446 10859
rect 1380 10786 1446 10825
rect 1380 10752 1396 10786
rect 1430 10752 1446 10786
rect 1380 10712 1446 10752
rect 1380 10678 1396 10712
rect 1430 10678 1446 10712
rect 1380 10638 1446 10678
rect 1380 10604 1396 10638
rect 1430 10604 1446 10638
rect 1380 10564 1446 10604
rect 1380 10530 1396 10564
rect 1430 10530 1446 10564
rect 1380 10490 1446 10530
rect 1380 10456 1396 10490
rect 1430 10456 1446 10490
rect 1380 10440 1446 10456
rect 3490 11224 3556 11240
rect 3490 11190 3506 11224
rect 3540 11190 3556 11224
rect 3490 11151 3556 11190
rect 3490 11117 3506 11151
rect 3540 11117 3556 11151
rect 3490 11078 3556 11117
rect 3490 11044 3506 11078
rect 3540 11044 3556 11078
rect 3490 11005 3556 11044
rect 3490 10971 3506 11005
rect 3540 10971 3556 11005
rect 3490 10932 3556 10971
rect 3490 10898 3506 10932
rect 3540 10898 3556 10932
rect 3490 10859 3556 10898
rect 3490 10825 3506 10859
rect 3540 10825 3556 10859
rect 3490 10786 3556 10825
rect 3490 10752 3506 10786
rect 3540 10752 3556 10786
rect 3490 10712 3556 10752
rect 3490 10678 3506 10712
rect 3540 10678 3556 10712
rect 3490 10638 3556 10678
rect 3490 10604 3506 10638
rect 3540 10604 3556 10638
rect 3490 10564 3556 10604
rect 3490 10530 3506 10564
rect 3540 10530 3556 10564
rect 3490 10490 3556 10530
rect 3490 10456 3506 10490
rect 3540 10456 3556 10490
rect 3490 10440 3556 10456
rect 1380 10138 1446 10154
rect 1380 10104 1396 10138
rect 1430 10104 1446 10138
rect 1380 10065 1446 10104
rect 1380 10031 1396 10065
rect 1430 10031 1446 10065
rect 1380 9992 1446 10031
rect 1380 9958 1396 9992
rect 1430 9958 1446 9992
rect 1380 9919 1446 9958
rect 1380 9885 1396 9919
rect 1430 9885 1446 9919
rect 1380 9846 1446 9885
rect 1380 9812 1396 9846
rect 1430 9812 1446 9846
rect 1380 9773 1446 9812
rect 1380 9739 1396 9773
rect 1430 9739 1446 9773
rect 1380 9700 1446 9739
rect 1380 9666 1396 9700
rect 1430 9666 1446 9700
rect 1380 9626 1446 9666
rect 1380 9592 1396 9626
rect 1430 9592 1446 9626
rect 1380 9552 1446 9592
rect 1380 9518 1396 9552
rect 1430 9518 1446 9552
rect 1380 9478 1446 9518
rect 1380 9444 1396 9478
rect 1430 9444 1446 9478
rect 1380 9404 1446 9444
rect 1380 9370 1396 9404
rect 1430 9370 1446 9404
rect 1380 9354 1446 9370
rect 3490 10138 3556 10154
rect 3490 10104 3506 10138
rect 3540 10104 3556 10138
rect 3490 10065 3556 10104
rect 3490 10031 3506 10065
rect 3540 10031 3556 10065
rect 3490 9992 3556 10031
rect 3490 9958 3506 9992
rect 3540 9958 3556 9992
rect 3490 9919 3556 9958
rect 3490 9885 3506 9919
rect 3540 9885 3556 9919
rect 3490 9846 3556 9885
rect 3490 9812 3506 9846
rect 3540 9812 3556 9846
rect 3490 9773 3556 9812
rect 3490 9739 3506 9773
rect 3540 9739 3556 9773
rect 3490 9700 3556 9739
rect 3490 9666 3506 9700
rect 3540 9666 3556 9700
rect 3490 9626 3556 9666
rect 3490 9592 3506 9626
rect 3540 9592 3556 9626
rect 3490 9552 3556 9592
rect 3490 9518 3506 9552
rect 3540 9518 3556 9552
rect 3490 9478 3556 9518
rect 3490 9444 3506 9478
rect 3540 9444 3556 9478
rect 3490 9404 3556 9444
rect 3490 9370 3506 9404
rect 3540 9370 3556 9404
rect 3490 9354 3556 9370
rect 1380 9282 1446 9298
rect 1380 9248 1396 9282
rect 1430 9248 1446 9282
rect 1380 9209 1446 9248
rect 1380 9175 1396 9209
rect 1430 9175 1446 9209
rect 1380 9136 1446 9175
rect 1380 9102 1396 9136
rect 1430 9102 1446 9136
rect 1380 9063 1446 9102
rect 1380 9029 1396 9063
rect 1430 9029 1446 9063
rect 1380 8990 1446 9029
rect 1380 8956 1396 8990
rect 1430 8956 1446 8990
rect 1380 8917 1446 8956
rect 1380 8883 1396 8917
rect 1430 8883 1446 8917
rect 1380 8844 1446 8883
rect 1380 8810 1396 8844
rect 1430 8810 1446 8844
rect 1380 8770 1446 8810
rect 1380 8736 1396 8770
rect 1430 8736 1446 8770
rect 1380 8696 1446 8736
rect 1380 8662 1396 8696
rect 1430 8662 1446 8696
rect 1380 8622 1446 8662
rect 1380 8588 1396 8622
rect 1430 8588 1446 8622
rect 1380 8548 1446 8588
rect 1380 8514 1396 8548
rect 1430 8514 1446 8548
rect 1380 8498 1446 8514
rect 3490 9282 3556 9298
rect 3490 9248 3506 9282
rect 3540 9248 3556 9282
rect 3490 9209 3556 9248
rect 3490 9175 3506 9209
rect 3540 9175 3556 9209
rect 3490 9136 3556 9175
rect 3490 9102 3506 9136
rect 3540 9102 3556 9136
rect 3490 9063 3556 9102
rect 3490 9029 3506 9063
rect 3540 9029 3556 9063
rect 3490 8990 3556 9029
rect 3490 8956 3506 8990
rect 3540 8956 3556 8990
rect 3490 8917 3556 8956
rect 3490 8883 3506 8917
rect 3540 8883 3556 8917
rect 3490 8844 3556 8883
rect 3490 8810 3506 8844
rect 3540 8810 3556 8844
rect 3490 8770 3556 8810
rect 3490 8736 3506 8770
rect 3540 8736 3556 8770
rect 3490 8696 3556 8736
rect 3490 8662 3506 8696
rect 3540 8662 3556 8696
rect 3490 8622 3556 8662
rect 3490 8588 3506 8622
rect 3540 8588 3556 8622
rect 3490 8548 3556 8588
rect 3490 8514 3506 8548
rect 3540 8514 3556 8548
rect 3490 8498 3556 8514
rect 1380 8222 1446 8238
rect 1380 8188 1396 8222
rect 1430 8188 1446 8222
rect 1380 8153 1446 8188
rect 1380 8119 1396 8153
rect 1430 8119 1446 8153
rect 1380 8084 1446 8119
rect 1380 8050 1396 8084
rect 1430 8050 1446 8084
rect 1380 8015 1446 8050
rect 1380 7981 1396 8015
rect 1430 7981 1446 8015
rect 1380 7946 1446 7981
rect 1380 7912 1396 7946
rect 1430 7912 1446 7946
rect 1380 7877 1446 7912
rect 1380 7843 1396 7877
rect 1430 7843 1446 7877
rect 1380 7808 1446 7843
rect 1380 7774 1396 7808
rect 1430 7774 1446 7808
rect 1380 7739 1446 7774
rect 1380 7705 1396 7739
rect 1430 7705 1446 7739
rect 1380 7670 1446 7705
rect 1380 7636 1396 7670
rect 1430 7636 1446 7670
rect 1380 7601 1446 7636
rect 1380 7567 1396 7601
rect 1430 7567 1446 7601
rect 1380 7532 1446 7567
rect 1380 7498 1396 7532
rect 1430 7498 1446 7532
rect 1380 7462 1446 7498
rect 1380 7428 1396 7462
rect 1430 7428 1446 7462
rect 1380 7412 1446 7428
rect 3490 8222 3556 8238
rect 3490 8188 3506 8222
rect 3540 8188 3556 8222
rect 3490 8153 3556 8188
rect 3490 8119 3506 8153
rect 3540 8119 3556 8153
rect 3490 8084 3556 8119
rect 3490 8050 3506 8084
rect 3540 8050 3556 8084
rect 3490 8015 3556 8050
rect 3490 7981 3506 8015
rect 3540 7981 3556 8015
rect 3490 7946 3556 7981
rect 3490 7912 3506 7946
rect 3540 7912 3556 7946
rect 3490 7877 3556 7912
rect 3490 7843 3506 7877
rect 3540 7843 3556 7877
rect 3490 7808 3556 7843
rect 3490 7774 3506 7808
rect 3540 7774 3556 7808
rect 3490 7739 3556 7774
rect 3490 7705 3506 7739
rect 3540 7705 3556 7739
rect 3490 7670 3556 7705
rect 3490 7636 3506 7670
rect 3540 7636 3556 7670
rect 3490 7601 3556 7636
rect 3490 7567 3506 7601
rect 3540 7567 3556 7601
rect 3490 7532 3556 7567
rect 3490 7498 3506 7532
rect 3540 7498 3556 7532
rect 3490 7462 3556 7498
rect 3490 7428 3506 7462
rect 3540 7428 3556 7462
rect 3490 7412 3556 7428
rect 1380 6464 1446 6480
rect 1380 6430 1396 6464
rect 1430 6430 1446 6464
rect 1380 6391 1446 6430
rect 1380 6357 1396 6391
rect 1430 6357 1446 6391
rect 1380 6318 1446 6357
rect 1380 6284 1396 6318
rect 1430 6284 1446 6318
rect 1380 6245 1446 6284
rect 1380 6211 1396 6245
rect 1430 6211 1446 6245
rect 1380 6172 1446 6211
rect 1380 6138 1396 6172
rect 1430 6138 1446 6172
rect 1380 6099 1446 6138
rect 1380 6065 1396 6099
rect 1430 6065 1446 6099
rect 1380 6026 1446 6065
rect 1380 5992 1396 6026
rect 1430 5992 1446 6026
rect 1380 5952 1446 5992
rect 1380 5918 1396 5952
rect 1430 5918 1446 5952
rect 1380 5878 1446 5918
rect 1380 5844 1396 5878
rect 1430 5844 1446 5878
rect 1380 5804 1446 5844
rect 1380 5770 1396 5804
rect 1430 5770 1446 5804
rect 1380 5730 1446 5770
rect 1380 5696 1396 5730
rect 1430 5696 1446 5730
rect 1380 5680 1446 5696
rect 3490 6464 3556 6480
rect 3490 6430 3506 6464
rect 3540 6430 3556 6464
rect 3490 6391 3556 6430
rect 3490 6357 3506 6391
rect 3540 6357 3556 6391
rect 3490 6318 3556 6357
rect 3490 6284 3506 6318
rect 3540 6284 3556 6318
rect 3490 6245 3556 6284
rect 3490 6211 3506 6245
rect 3540 6211 3556 6245
rect 3490 6172 3556 6211
rect 3490 6138 3506 6172
rect 3540 6138 3556 6172
rect 3490 6099 3556 6138
rect 3490 6065 3506 6099
rect 3540 6065 3556 6099
rect 3490 6026 3556 6065
rect 3490 5992 3506 6026
rect 3540 5992 3556 6026
rect 3490 5952 3556 5992
rect 3490 5918 3506 5952
rect 3540 5918 3556 5952
rect 3490 5878 3556 5918
rect 3490 5844 3506 5878
rect 3540 5844 3556 5878
rect 3490 5804 3556 5844
rect 3490 5770 3506 5804
rect 3540 5770 3556 5804
rect 3490 5730 3556 5770
rect 3490 5696 3506 5730
rect 3540 5696 3556 5730
rect 3490 5680 3556 5696
rect 1380 5378 1446 5394
rect 1380 5344 1396 5378
rect 1430 5344 1446 5378
rect 1380 5305 1446 5344
rect 1380 5271 1396 5305
rect 1430 5271 1446 5305
rect 1380 5232 1446 5271
rect 1380 5198 1396 5232
rect 1430 5198 1446 5232
rect 1380 5159 1446 5198
rect 1380 5125 1396 5159
rect 1430 5125 1446 5159
rect 1380 5086 1446 5125
rect 1380 5052 1396 5086
rect 1430 5052 1446 5086
rect 1380 5013 1446 5052
rect 1380 4979 1396 5013
rect 1430 4979 1446 5013
rect 1380 4940 1446 4979
rect 1380 4906 1396 4940
rect 1430 4906 1446 4940
rect 1380 4866 1446 4906
rect 1380 4832 1396 4866
rect 1430 4832 1446 4866
rect 1380 4792 1446 4832
rect 1380 4758 1396 4792
rect 1430 4758 1446 4792
rect 1380 4718 1446 4758
rect 1380 4684 1396 4718
rect 1430 4684 1446 4718
rect 1380 4644 1446 4684
rect 1380 4610 1396 4644
rect 1430 4610 1446 4644
rect 1380 4594 1446 4610
rect 3490 5378 3556 5394
rect 3490 5344 3506 5378
rect 3540 5344 3556 5378
rect 3490 5305 3556 5344
rect 3490 5271 3506 5305
rect 3540 5271 3556 5305
rect 3490 5232 3556 5271
rect 3490 5198 3506 5232
rect 3540 5198 3556 5232
rect 3490 5159 3556 5198
rect 3490 5125 3506 5159
rect 3540 5125 3556 5159
rect 3490 5086 3556 5125
rect 3490 5052 3506 5086
rect 3540 5052 3556 5086
rect 3490 5013 3556 5052
rect 3490 4979 3506 5013
rect 3540 4979 3556 5013
rect 3490 4940 3556 4979
rect 3490 4906 3506 4940
rect 3540 4906 3556 4940
rect 3490 4866 3556 4906
rect 3490 4832 3506 4866
rect 3540 4832 3556 4866
rect 3490 4792 3556 4832
rect 3490 4758 3506 4792
rect 3540 4758 3556 4792
rect 3490 4718 3556 4758
rect 3490 4684 3506 4718
rect 3540 4684 3556 4718
rect 3490 4644 3556 4684
rect 3490 4610 3506 4644
rect 3540 4610 3556 4644
rect 3490 4594 3556 4610
rect 1380 4522 1446 4538
rect 1380 4488 1396 4522
rect 1430 4488 1446 4522
rect 1380 4449 1446 4488
rect 1380 4415 1396 4449
rect 1430 4415 1446 4449
rect 1380 4376 1446 4415
rect 1380 4342 1396 4376
rect 1430 4342 1446 4376
rect 1380 4303 1446 4342
rect 1380 4269 1396 4303
rect 1430 4269 1446 4303
rect 1380 4230 1446 4269
rect 1380 4196 1396 4230
rect 1430 4196 1446 4230
rect 1380 4157 1446 4196
rect 1380 4123 1396 4157
rect 1430 4123 1446 4157
rect 1380 4084 1446 4123
rect 1380 4050 1396 4084
rect 1430 4050 1446 4084
rect 1380 4010 1446 4050
rect 1380 3976 1396 4010
rect 1430 3976 1446 4010
rect 1380 3936 1446 3976
rect 1380 3902 1396 3936
rect 1430 3902 1446 3936
rect 1380 3862 1446 3902
rect 1380 3828 1396 3862
rect 1430 3828 1446 3862
rect 1380 3788 1446 3828
rect 1380 3754 1396 3788
rect 1430 3754 1446 3788
rect 1380 3738 1446 3754
rect 3490 4522 3556 4538
rect 3490 4488 3506 4522
rect 3540 4488 3556 4522
rect 3490 4449 3556 4488
rect 3490 4415 3506 4449
rect 3540 4415 3556 4449
rect 3490 4376 3556 4415
rect 3490 4342 3506 4376
rect 3540 4342 3556 4376
rect 3490 4303 3556 4342
rect 3490 4269 3506 4303
rect 3540 4269 3556 4303
rect 3490 4230 3556 4269
rect 3490 4196 3506 4230
rect 3540 4196 3556 4230
rect 3490 4157 3556 4196
rect 3490 4123 3506 4157
rect 3540 4123 3556 4157
rect 3490 4084 3556 4123
rect 3490 4050 3506 4084
rect 3540 4050 3556 4084
rect 3490 4010 3556 4050
rect 3490 3976 3506 4010
rect 3540 3976 3556 4010
rect 3490 3936 3556 3976
rect 3490 3902 3506 3936
rect 3540 3902 3556 3936
rect 3490 3862 3556 3902
rect 3490 3828 3506 3862
rect 3540 3828 3556 3862
rect 3490 3788 3556 3828
rect 3490 3754 3506 3788
rect 3540 3754 3556 3788
rect 3490 3738 3556 3754
rect 4066 11170 5242 11201
rect 4066 11136 4082 11170
rect 4116 11136 5192 11170
rect 5226 11136 5242 11170
rect 4066 11101 5242 11136
rect 4066 11029 4132 11045
rect 4066 10995 4082 11029
rect 4116 10995 4132 11029
rect 4066 10956 4132 10995
rect 4066 10922 4082 10956
rect 4116 10922 4132 10956
rect 4066 10883 4132 10922
rect 4066 10849 4082 10883
rect 4116 10849 4132 10883
rect 4066 10810 4132 10849
rect 4066 10776 4082 10810
rect 4116 10776 4132 10810
rect 4066 10737 4132 10776
rect 4066 10703 4082 10737
rect 4116 10703 4132 10737
rect 4066 10664 4132 10703
rect 4066 10630 4082 10664
rect 4116 10630 4132 10664
rect 4066 10591 4132 10630
rect 4066 10557 4082 10591
rect 4116 10557 4132 10591
rect 4066 10517 4132 10557
rect 4066 10483 4082 10517
rect 4116 10483 4132 10517
rect 4066 10443 4132 10483
rect 4066 10409 4082 10443
rect 4116 10409 4132 10443
rect 4066 10369 4132 10409
rect 4066 10335 4082 10369
rect 4116 10335 4132 10369
rect 4066 10295 4132 10335
rect 4066 10261 4082 10295
rect 4116 10261 4132 10295
rect 4066 10245 4132 10261
rect 5176 11029 5242 11045
rect 5176 10995 5192 11029
rect 5226 10995 5242 11029
rect 5176 10956 5242 10995
rect 5176 10922 5192 10956
rect 5226 10922 5242 10956
rect 5176 10883 5242 10922
rect 5176 10849 5192 10883
rect 5226 10849 5242 10883
rect 5176 10810 5242 10849
rect 5176 10776 5192 10810
rect 5226 10776 5242 10810
rect 5176 10737 5242 10776
rect 5176 10703 5192 10737
rect 5226 10703 5242 10737
rect 5176 10664 5242 10703
rect 5176 10630 5192 10664
rect 5226 10630 5242 10664
rect 5176 10591 5242 10630
rect 5176 10557 5192 10591
rect 5226 10557 5242 10591
rect 5176 10517 5242 10557
rect 5176 10483 5192 10517
rect 5226 10483 5242 10517
rect 5176 10443 5242 10483
rect 5176 10409 5192 10443
rect 5226 10409 5242 10443
rect 5176 10369 5242 10409
rect 5176 10335 5192 10369
rect 5226 10335 5242 10369
rect 5176 10295 5242 10335
rect 5176 10261 5192 10295
rect 5226 10261 5242 10295
rect 5176 10245 5242 10261
rect 4066 10173 4132 10189
rect 4066 10139 4082 10173
rect 4116 10139 4132 10173
rect 4066 10100 4132 10139
rect 4066 10066 4082 10100
rect 4116 10066 4132 10100
rect 4066 10027 4132 10066
rect 4066 9993 4082 10027
rect 4116 9993 4132 10027
rect 4066 9954 4132 9993
rect 4066 9920 4082 9954
rect 4116 9920 4132 9954
rect 4066 9881 4132 9920
rect 4066 9847 4082 9881
rect 4116 9847 4132 9881
rect 4066 9808 4132 9847
rect 4066 9774 4082 9808
rect 4116 9774 4132 9808
rect 4066 9735 4132 9774
rect 4066 9701 4082 9735
rect 4116 9701 4132 9735
rect 4066 9661 4132 9701
rect 4066 9627 4082 9661
rect 4116 9627 4132 9661
rect 4066 9587 4132 9627
rect 4066 9553 4082 9587
rect 4116 9553 4132 9587
rect 4066 9513 4132 9553
rect 4066 9479 4082 9513
rect 4116 9479 4132 9513
rect 4066 9439 4132 9479
rect 4066 9405 4082 9439
rect 4116 9405 4132 9439
rect 4066 9389 4132 9405
rect 5176 10173 5242 10189
rect 5176 10139 5192 10173
rect 5226 10139 5242 10173
rect 5176 10100 5242 10139
rect 5176 10066 5192 10100
rect 5226 10066 5242 10100
rect 5176 10027 5242 10066
rect 5176 9993 5192 10027
rect 5226 9993 5242 10027
rect 5176 9954 5242 9993
rect 5176 9920 5192 9954
rect 5226 9920 5242 9954
rect 5176 9881 5242 9920
rect 5176 9847 5192 9881
rect 5226 9847 5242 9881
rect 5176 9808 5242 9847
rect 5176 9774 5192 9808
rect 5226 9774 5242 9808
rect 5176 9735 5242 9774
rect 5176 9701 5192 9735
rect 5226 9701 5242 9735
rect 5176 9661 5242 9701
rect 5176 9627 5192 9661
rect 5226 9627 5242 9661
rect 5176 9587 5242 9627
rect 5176 9553 5192 9587
rect 5226 9553 5242 9587
rect 5176 9513 5242 9553
rect 5176 9479 5192 9513
rect 5226 9479 5242 9513
rect 5176 9439 5242 9479
rect 5176 9405 5192 9439
rect 5226 9405 5242 9439
rect 5176 9389 5242 9405
rect 4066 9317 4132 9333
rect 4066 9283 4082 9317
rect 4116 9283 4132 9317
rect 4066 9244 4132 9283
rect 4066 9210 4082 9244
rect 4116 9210 4132 9244
rect 4066 9171 4132 9210
rect 4066 9137 4082 9171
rect 4116 9137 4132 9171
rect 4066 9098 4132 9137
rect 4066 9064 4082 9098
rect 4116 9064 4132 9098
rect 4066 9025 4132 9064
rect 4066 8991 4082 9025
rect 4116 8991 4132 9025
rect 4066 8952 4132 8991
rect 4066 8918 4082 8952
rect 4116 8918 4132 8952
rect 4066 8879 4132 8918
rect 4066 8845 4082 8879
rect 4116 8845 4132 8879
rect 4066 8805 4132 8845
rect 4066 8771 4082 8805
rect 4116 8771 4132 8805
rect 4066 8731 4132 8771
rect 4066 8697 4082 8731
rect 4116 8697 4132 8731
rect 4066 8657 4132 8697
rect 4066 8623 4082 8657
rect 4116 8623 4132 8657
rect 4066 8583 4132 8623
rect 4066 8549 4082 8583
rect 4116 8549 4132 8583
rect 4066 8533 4132 8549
rect 5176 9317 5242 9333
rect 5176 9283 5192 9317
rect 5226 9283 5242 9317
rect 5176 9244 5242 9283
rect 5176 9210 5192 9244
rect 5226 9210 5242 9244
rect 5176 9171 5242 9210
rect 5176 9137 5192 9171
rect 5226 9137 5242 9171
rect 5176 9098 5242 9137
rect 5176 9064 5192 9098
rect 5226 9064 5242 9098
rect 5176 9025 5242 9064
rect 5176 8991 5192 9025
rect 5226 8991 5242 9025
rect 5176 8952 5242 8991
rect 5176 8918 5192 8952
rect 5226 8918 5242 8952
rect 5176 8879 5242 8918
rect 5176 8845 5192 8879
rect 5226 8845 5242 8879
rect 5176 8805 5242 8845
rect 5176 8771 5192 8805
rect 5226 8771 5242 8805
rect 5176 8731 5242 8771
rect 5176 8697 5192 8731
rect 5226 8697 5242 8731
rect 5176 8657 5242 8697
rect 5176 8623 5192 8657
rect 5226 8623 5242 8657
rect 5176 8583 5242 8623
rect 5176 8549 5192 8583
rect 5226 8549 5242 8583
rect 5176 8533 5242 8549
rect 4066 8461 4132 8477
rect 4066 8427 4082 8461
rect 4116 8427 4132 8461
rect 4066 8388 4132 8427
rect 4066 8354 4082 8388
rect 4116 8354 4132 8388
rect 4066 8315 4132 8354
rect 4066 8281 4082 8315
rect 4116 8281 4132 8315
rect 4066 8242 4132 8281
rect 4066 8208 4082 8242
rect 4116 8208 4132 8242
rect 4066 8169 4132 8208
rect 4066 8135 4082 8169
rect 4116 8135 4132 8169
rect 4066 8096 4132 8135
rect 4066 8062 4082 8096
rect 4116 8062 4132 8096
rect 4066 8023 4132 8062
rect 4066 7989 4082 8023
rect 4116 7989 4132 8023
rect 4066 7949 4132 7989
rect 4066 7915 4082 7949
rect 4116 7915 4132 7949
rect 4066 7875 4132 7915
rect 4066 7841 4082 7875
rect 4116 7841 4132 7875
rect 4066 7801 4132 7841
rect 4066 7767 4082 7801
rect 4116 7767 4132 7801
rect 4066 7727 4132 7767
rect 4066 7693 4082 7727
rect 4116 7693 4132 7727
rect 4066 7677 4132 7693
rect 5176 8461 5242 8477
rect 5176 8427 5192 8461
rect 5226 8427 5242 8461
rect 5176 8388 5242 8427
rect 5176 8354 5192 8388
rect 5226 8354 5242 8388
rect 5176 8315 5242 8354
rect 5176 8281 5192 8315
rect 5226 8281 5242 8315
rect 5176 8242 5242 8281
rect 5176 8208 5192 8242
rect 5226 8208 5242 8242
rect 5176 8169 5242 8208
rect 5176 8135 5192 8169
rect 5226 8135 5242 8169
rect 5176 8096 5242 8135
rect 5176 8062 5192 8096
rect 5226 8062 5242 8096
rect 5176 8023 5242 8062
rect 5176 7989 5192 8023
rect 5226 7989 5242 8023
rect 5176 7949 5242 7989
rect 5176 7915 5192 7949
rect 5226 7915 5242 7949
rect 5176 7875 5242 7915
rect 5176 7841 5192 7875
rect 5226 7841 5242 7875
rect 5176 7801 5242 7841
rect 5176 7767 5192 7801
rect 5226 7767 5242 7801
rect 5176 7727 5242 7767
rect 5176 7693 5192 7727
rect 5226 7693 5242 7727
rect 5176 7677 5242 7693
rect 4066 7605 4132 7621
rect 4066 7571 4082 7605
rect 4116 7571 4132 7605
rect 4066 7532 4132 7571
rect 4066 7498 4082 7532
rect 4116 7498 4132 7532
rect 4066 7459 4132 7498
rect 4066 7425 4082 7459
rect 4116 7425 4132 7459
rect 4066 7386 4132 7425
rect 4066 7352 4082 7386
rect 4116 7352 4132 7386
rect 4066 7313 4132 7352
rect 4066 7279 4082 7313
rect 4116 7279 4132 7313
rect 4066 7240 4132 7279
rect 4066 7206 4082 7240
rect 4116 7206 4132 7240
rect 4066 7167 4132 7206
rect 4066 7133 4082 7167
rect 4116 7133 4132 7167
rect 4066 7093 4132 7133
rect 4066 7059 4082 7093
rect 4116 7059 4132 7093
rect 4066 7019 4132 7059
rect 4066 6985 4082 7019
rect 4116 6985 4132 7019
rect 4066 6945 4132 6985
rect 4066 6911 4082 6945
rect 4116 6911 4132 6945
rect 4066 6871 4132 6911
rect 4066 6837 4082 6871
rect 4116 6837 4132 6871
rect 4066 6821 4132 6837
rect 5176 7605 5242 7621
rect 5176 7571 5192 7605
rect 5226 7571 5242 7605
rect 5176 7532 5242 7571
rect 5176 7498 5192 7532
rect 5226 7498 5242 7532
rect 5176 7459 5242 7498
rect 5176 7425 5192 7459
rect 5226 7425 5242 7459
rect 5176 7386 5242 7425
rect 5176 7352 5192 7386
rect 5226 7352 5242 7386
rect 5176 7313 5242 7352
rect 5176 7279 5192 7313
rect 5226 7279 5242 7313
rect 5176 7240 5242 7279
rect 5176 7206 5192 7240
rect 5226 7206 5242 7240
rect 5176 7167 5242 7206
rect 5176 7133 5192 7167
rect 5226 7133 5242 7167
rect 5176 7093 5242 7133
rect 5176 7059 5192 7093
rect 5226 7059 5242 7093
rect 5176 7019 5242 7059
rect 5176 6985 5192 7019
rect 5226 6985 5242 7019
rect 5176 6945 5242 6985
rect 5176 6911 5192 6945
rect 5226 6911 5242 6945
rect 5176 6871 5242 6911
rect 5176 6837 5192 6871
rect 5226 6837 5242 6871
rect 5176 6821 5242 6837
rect 4066 6749 4132 6765
rect 4066 6715 4082 6749
rect 4116 6715 4132 6749
rect 4066 6676 4132 6715
rect 4066 6642 4082 6676
rect 4116 6642 4132 6676
rect 4066 6603 4132 6642
rect 4066 6569 4082 6603
rect 4116 6569 4132 6603
rect 4066 6530 4132 6569
rect 4066 6496 4082 6530
rect 4116 6496 4132 6530
rect 4066 6457 4132 6496
rect 4066 6423 4082 6457
rect 4116 6423 4132 6457
rect 4066 6384 4132 6423
rect 4066 6350 4082 6384
rect 4116 6350 4132 6384
rect 4066 6311 4132 6350
rect 4066 6277 4082 6311
rect 4116 6277 4132 6311
rect 4066 6237 4132 6277
rect 4066 6203 4082 6237
rect 4116 6203 4132 6237
rect 4066 6163 4132 6203
rect 4066 6129 4082 6163
rect 4116 6129 4132 6163
rect 4066 6089 4132 6129
rect 4066 6055 4082 6089
rect 4116 6055 4132 6089
rect 4066 6015 4132 6055
rect 4066 5981 4082 6015
rect 4116 5981 4132 6015
rect 4066 5965 4132 5981
rect 5176 6749 5242 6765
rect 5176 6715 5192 6749
rect 5226 6715 5242 6749
rect 5176 6676 5242 6715
rect 5176 6642 5192 6676
rect 5226 6642 5242 6676
rect 5176 6603 5242 6642
rect 5176 6569 5192 6603
rect 5226 6569 5242 6603
rect 5176 6530 5242 6569
rect 5176 6496 5192 6530
rect 5226 6496 5242 6530
rect 5176 6457 5242 6496
rect 5176 6423 5192 6457
rect 5226 6423 5242 6457
rect 5176 6384 5242 6423
rect 5176 6350 5192 6384
rect 5226 6350 5242 6384
rect 5176 6311 5242 6350
rect 5176 6277 5192 6311
rect 5226 6277 5242 6311
rect 5176 6237 5242 6277
rect 5176 6203 5192 6237
rect 5226 6203 5242 6237
rect 5176 6163 5242 6203
rect 5176 6129 5192 6163
rect 5226 6129 5242 6163
rect 5176 6089 5242 6129
rect 5176 6055 5192 6089
rect 5226 6055 5242 6089
rect 5176 6015 5242 6055
rect 5176 5981 5192 6015
rect 5226 5981 5242 6015
rect 5176 5965 5242 5981
rect 4066 5893 4132 5909
rect 4066 5859 4082 5893
rect 4116 5859 4132 5893
rect 4066 5820 4132 5859
rect 4066 5786 4082 5820
rect 4116 5786 4132 5820
rect 4066 5747 4132 5786
rect 4066 5713 4082 5747
rect 4116 5713 4132 5747
rect 4066 5674 4132 5713
rect 4066 5640 4082 5674
rect 4116 5640 4132 5674
rect 4066 5601 4132 5640
rect 4066 5567 4082 5601
rect 4116 5567 4132 5601
rect 4066 5528 4132 5567
rect 4066 5494 4082 5528
rect 4116 5494 4132 5528
rect 4066 5455 4132 5494
rect 4066 5421 4082 5455
rect 4116 5421 4132 5455
rect 4066 5381 4132 5421
rect 4066 5347 4082 5381
rect 4116 5347 4132 5381
rect 4066 5307 4132 5347
rect 4066 5273 4082 5307
rect 4116 5273 4132 5307
rect 4066 5233 4132 5273
rect 4066 5199 4082 5233
rect 4116 5199 4132 5233
rect 4066 5159 4132 5199
rect 4066 5125 4082 5159
rect 4116 5125 4132 5159
rect 4066 5109 4132 5125
rect 5176 5893 5242 5909
rect 5176 5859 5192 5893
rect 5226 5859 5242 5893
rect 5176 5820 5242 5859
rect 5176 5786 5192 5820
rect 5226 5786 5242 5820
rect 5176 5747 5242 5786
rect 5176 5713 5192 5747
rect 5226 5713 5242 5747
rect 5176 5674 5242 5713
rect 5176 5640 5192 5674
rect 5226 5640 5242 5674
rect 5176 5601 5242 5640
rect 5176 5567 5192 5601
rect 5226 5567 5242 5601
rect 5176 5528 5242 5567
rect 5176 5494 5192 5528
rect 5226 5494 5242 5528
rect 5176 5455 5242 5494
rect 5176 5421 5192 5455
rect 5226 5421 5242 5455
rect 5176 5381 5242 5421
rect 5176 5347 5192 5381
rect 5226 5347 5242 5381
rect 5176 5307 5242 5347
rect 5176 5273 5192 5307
rect 5226 5273 5242 5307
rect 5176 5233 5242 5273
rect 5176 5199 5192 5233
rect 5226 5199 5242 5233
rect 5176 5159 5242 5199
rect 5176 5125 5192 5159
rect 5226 5125 5242 5159
rect 5176 5109 5242 5125
rect 4066 5037 4132 5053
rect 4066 5003 4082 5037
rect 4116 5003 4132 5037
rect 4066 4964 4132 5003
rect 4066 4930 4082 4964
rect 4116 4930 4132 4964
rect 4066 4891 4132 4930
rect 4066 4857 4082 4891
rect 4116 4857 4132 4891
rect 4066 4818 4132 4857
rect 4066 4784 4082 4818
rect 4116 4784 4132 4818
rect 4066 4745 4132 4784
rect 4066 4711 4082 4745
rect 4116 4711 4132 4745
rect 4066 4672 4132 4711
rect 4066 4638 4082 4672
rect 4116 4638 4132 4672
rect 4066 4599 4132 4638
rect 4066 4565 4082 4599
rect 4116 4565 4132 4599
rect 4066 4525 4132 4565
rect 4066 4491 4082 4525
rect 4116 4491 4132 4525
rect 4066 4451 4132 4491
rect 4066 4417 4082 4451
rect 4116 4417 4132 4451
rect 4066 4377 4132 4417
rect 4066 4343 4082 4377
rect 4116 4343 4132 4377
rect 4066 4303 4132 4343
rect 4066 4269 4082 4303
rect 4116 4269 4132 4303
rect 4066 4253 4132 4269
rect 5176 5037 5242 5053
rect 5176 5003 5192 5037
rect 5226 5003 5242 5037
rect 5176 4964 5242 5003
rect 5176 4930 5192 4964
rect 5226 4930 5242 4964
rect 5176 4891 5242 4930
rect 5176 4857 5192 4891
rect 5226 4857 5242 4891
rect 5176 4818 5242 4857
rect 5176 4784 5192 4818
rect 5226 4784 5242 4818
rect 5176 4745 5242 4784
rect 5176 4711 5192 4745
rect 5226 4711 5242 4745
rect 5176 4672 5242 4711
rect 5176 4638 5192 4672
rect 5226 4638 5242 4672
rect 5176 4599 5242 4638
rect 5176 4565 5192 4599
rect 5226 4565 5242 4599
rect 5176 4525 5242 4565
rect 5176 4491 5192 4525
rect 5226 4491 5242 4525
rect 5176 4451 5242 4491
rect 5176 4417 5192 4451
rect 5226 4417 5242 4451
rect 5176 4377 5242 4417
rect 5176 4343 5192 4377
rect 5226 4343 5242 4377
rect 5176 4303 5242 4343
rect 5176 4269 5192 4303
rect 5226 4269 5242 4303
rect 5176 4253 5242 4269
rect 4066 4166 5242 4197
rect 4066 4132 4082 4166
rect 4116 4132 5192 4166
rect 5226 4132 5242 4166
rect 4066 4097 5242 4132
rect 5906 11170 7082 11201
rect 5906 11136 5922 11170
rect 5956 11136 7032 11170
rect 7066 11136 7082 11170
rect 5906 11101 7082 11136
rect 5906 11029 5972 11045
rect 5906 10995 5922 11029
rect 5956 10995 5972 11029
rect 5906 10956 5972 10995
rect 5906 10922 5922 10956
rect 5956 10922 5972 10956
rect 5906 10883 5972 10922
rect 5906 10849 5922 10883
rect 5956 10849 5972 10883
rect 5906 10810 5972 10849
rect 5906 10776 5922 10810
rect 5956 10776 5972 10810
rect 5906 10737 5972 10776
rect 5906 10703 5922 10737
rect 5956 10703 5972 10737
rect 5906 10664 5972 10703
rect 5906 10630 5922 10664
rect 5956 10630 5972 10664
rect 5906 10591 5972 10630
rect 5906 10557 5922 10591
rect 5956 10557 5972 10591
rect 5906 10517 5972 10557
rect 5906 10483 5922 10517
rect 5956 10483 5972 10517
rect 5906 10443 5972 10483
rect 5906 10409 5922 10443
rect 5956 10409 5972 10443
rect 5906 10369 5972 10409
rect 5906 10335 5922 10369
rect 5956 10335 5972 10369
rect 5906 10295 5972 10335
rect 5906 10261 5922 10295
rect 5956 10261 5972 10295
rect 5906 10245 5972 10261
rect 7016 11029 7082 11045
rect 7016 10995 7032 11029
rect 7066 10995 7082 11029
rect 7016 10956 7082 10995
rect 7016 10922 7032 10956
rect 7066 10922 7082 10956
rect 7016 10883 7082 10922
rect 7016 10849 7032 10883
rect 7066 10849 7082 10883
rect 7016 10810 7082 10849
rect 7016 10776 7032 10810
rect 7066 10776 7082 10810
rect 7016 10737 7082 10776
rect 7016 10703 7032 10737
rect 7066 10703 7082 10737
rect 7016 10664 7082 10703
rect 7016 10630 7032 10664
rect 7066 10630 7082 10664
rect 7016 10591 7082 10630
rect 7016 10557 7032 10591
rect 7066 10557 7082 10591
rect 7016 10517 7082 10557
rect 7016 10483 7032 10517
rect 7066 10483 7082 10517
rect 7016 10443 7082 10483
rect 7016 10409 7032 10443
rect 7066 10409 7082 10443
rect 7016 10369 7082 10409
rect 7016 10335 7032 10369
rect 7066 10335 7082 10369
rect 7016 10295 7082 10335
rect 7016 10261 7032 10295
rect 7066 10261 7082 10295
rect 7016 10245 7082 10261
rect 5906 10173 5972 10189
rect 5906 10139 5922 10173
rect 5956 10139 5972 10173
rect 5906 10100 5972 10139
rect 5906 10066 5922 10100
rect 5956 10066 5972 10100
rect 5906 10027 5972 10066
rect 5906 9993 5922 10027
rect 5956 9993 5972 10027
rect 5906 9954 5972 9993
rect 5906 9920 5922 9954
rect 5956 9920 5972 9954
rect 5906 9881 5972 9920
rect 5906 9847 5922 9881
rect 5956 9847 5972 9881
rect 5906 9808 5972 9847
rect 5906 9774 5922 9808
rect 5956 9774 5972 9808
rect 5906 9735 5972 9774
rect 5906 9701 5922 9735
rect 5956 9701 5972 9735
rect 5906 9661 5972 9701
rect 5906 9627 5922 9661
rect 5956 9627 5972 9661
rect 5906 9587 5972 9627
rect 5906 9553 5922 9587
rect 5956 9553 5972 9587
rect 5906 9513 5972 9553
rect 5906 9479 5922 9513
rect 5956 9479 5972 9513
rect 5906 9439 5972 9479
rect 5906 9405 5922 9439
rect 5956 9405 5972 9439
rect 5906 9389 5972 9405
rect 7016 10173 7082 10189
rect 7016 10139 7032 10173
rect 7066 10139 7082 10173
rect 7016 10100 7082 10139
rect 7016 10066 7032 10100
rect 7066 10066 7082 10100
rect 7016 10027 7082 10066
rect 7016 9993 7032 10027
rect 7066 9993 7082 10027
rect 7016 9954 7082 9993
rect 7016 9920 7032 9954
rect 7066 9920 7082 9954
rect 7016 9881 7082 9920
rect 7016 9847 7032 9881
rect 7066 9847 7082 9881
rect 7016 9808 7082 9847
rect 7016 9774 7032 9808
rect 7066 9774 7082 9808
rect 7016 9735 7082 9774
rect 7016 9701 7032 9735
rect 7066 9701 7082 9735
rect 7016 9661 7082 9701
rect 7016 9627 7032 9661
rect 7066 9627 7082 9661
rect 7016 9587 7082 9627
rect 7016 9553 7032 9587
rect 7066 9553 7082 9587
rect 7016 9513 7082 9553
rect 7016 9479 7032 9513
rect 7066 9479 7082 9513
rect 7016 9439 7082 9479
rect 7016 9405 7032 9439
rect 7066 9405 7082 9439
rect 7016 9389 7082 9405
rect 5906 9317 5972 9333
rect 5906 9283 5922 9317
rect 5956 9283 5972 9317
rect 5906 9244 5972 9283
rect 5906 9210 5922 9244
rect 5956 9210 5972 9244
rect 5906 9171 5972 9210
rect 5906 9137 5922 9171
rect 5956 9137 5972 9171
rect 5906 9098 5972 9137
rect 5906 9064 5922 9098
rect 5956 9064 5972 9098
rect 5906 9025 5972 9064
rect 5906 8991 5922 9025
rect 5956 8991 5972 9025
rect 5906 8952 5972 8991
rect 5906 8918 5922 8952
rect 5956 8918 5972 8952
rect 5906 8879 5972 8918
rect 5906 8845 5922 8879
rect 5956 8845 5972 8879
rect 5906 8805 5972 8845
rect 5906 8771 5922 8805
rect 5956 8771 5972 8805
rect 5906 8731 5972 8771
rect 5906 8697 5922 8731
rect 5956 8697 5972 8731
rect 5906 8657 5972 8697
rect 5906 8623 5922 8657
rect 5956 8623 5972 8657
rect 5906 8583 5972 8623
rect 5906 8549 5922 8583
rect 5956 8549 5972 8583
rect 5906 8533 5972 8549
rect 7016 9317 7082 9333
rect 7016 9283 7032 9317
rect 7066 9283 7082 9317
rect 7016 9244 7082 9283
rect 7016 9210 7032 9244
rect 7066 9210 7082 9244
rect 7016 9171 7082 9210
rect 7016 9137 7032 9171
rect 7066 9137 7082 9171
rect 7016 9098 7082 9137
rect 7016 9064 7032 9098
rect 7066 9064 7082 9098
rect 7016 9025 7082 9064
rect 7016 8991 7032 9025
rect 7066 8991 7082 9025
rect 7016 8952 7082 8991
rect 7016 8918 7032 8952
rect 7066 8918 7082 8952
rect 7016 8879 7082 8918
rect 7016 8845 7032 8879
rect 7066 8845 7082 8879
rect 7016 8805 7082 8845
rect 7016 8771 7032 8805
rect 7066 8771 7082 8805
rect 7016 8731 7082 8771
rect 7016 8697 7032 8731
rect 7066 8697 7082 8731
rect 7016 8657 7082 8697
rect 7016 8623 7032 8657
rect 7066 8623 7082 8657
rect 7016 8583 7082 8623
rect 7016 8549 7032 8583
rect 7066 8549 7082 8583
rect 7016 8533 7082 8549
rect 5906 8461 5972 8477
rect 5906 8427 5922 8461
rect 5956 8427 5972 8461
rect 5906 8388 5972 8427
rect 5906 8354 5922 8388
rect 5956 8354 5972 8388
rect 5906 8315 5972 8354
rect 5906 8281 5922 8315
rect 5956 8281 5972 8315
rect 5906 8242 5972 8281
rect 5906 8208 5922 8242
rect 5956 8208 5972 8242
rect 5906 8169 5972 8208
rect 5906 8135 5922 8169
rect 5956 8135 5972 8169
rect 5906 8096 5972 8135
rect 5906 8062 5922 8096
rect 5956 8062 5972 8096
rect 5906 8023 5972 8062
rect 5906 7989 5922 8023
rect 5956 7989 5972 8023
rect 5906 7949 5972 7989
rect 5906 7915 5922 7949
rect 5956 7915 5972 7949
rect 5906 7875 5972 7915
rect 5906 7841 5922 7875
rect 5956 7841 5972 7875
rect 5906 7801 5972 7841
rect 5906 7767 5922 7801
rect 5956 7767 5972 7801
rect 5906 7727 5972 7767
rect 5906 7693 5922 7727
rect 5956 7693 5972 7727
rect 5906 7677 5972 7693
rect 7016 8461 7082 8477
rect 7016 8427 7032 8461
rect 7066 8427 7082 8461
rect 7016 8388 7082 8427
rect 7016 8354 7032 8388
rect 7066 8354 7082 8388
rect 7016 8315 7082 8354
rect 7016 8281 7032 8315
rect 7066 8281 7082 8315
rect 7016 8242 7082 8281
rect 7016 8208 7032 8242
rect 7066 8208 7082 8242
rect 7016 8169 7082 8208
rect 7016 8135 7032 8169
rect 7066 8135 7082 8169
rect 7016 8096 7082 8135
rect 7016 8062 7032 8096
rect 7066 8062 7082 8096
rect 7016 8023 7082 8062
rect 7016 7989 7032 8023
rect 7066 7989 7082 8023
rect 7016 7949 7082 7989
rect 7016 7915 7032 7949
rect 7066 7915 7082 7949
rect 7016 7875 7082 7915
rect 7016 7841 7032 7875
rect 7066 7841 7082 7875
rect 7016 7801 7082 7841
rect 7016 7767 7032 7801
rect 7066 7767 7082 7801
rect 7016 7727 7082 7767
rect 7016 7693 7032 7727
rect 7066 7693 7082 7727
rect 7016 7677 7082 7693
rect 5906 7605 5972 7621
rect 5906 7571 5922 7605
rect 5956 7571 5972 7605
rect 5906 7532 5972 7571
rect 5906 7498 5922 7532
rect 5956 7498 5972 7532
rect 5906 7459 5972 7498
rect 5906 7425 5922 7459
rect 5956 7425 5972 7459
rect 5906 7386 5972 7425
rect 5906 7352 5922 7386
rect 5956 7352 5972 7386
rect 5906 7313 5972 7352
rect 5906 7279 5922 7313
rect 5956 7279 5972 7313
rect 5906 7240 5972 7279
rect 5906 7206 5922 7240
rect 5956 7206 5972 7240
rect 5906 7167 5972 7206
rect 5906 7133 5922 7167
rect 5956 7133 5972 7167
rect 5906 7093 5972 7133
rect 5906 7059 5922 7093
rect 5956 7059 5972 7093
rect 5906 7019 5972 7059
rect 5906 6985 5922 7019
rect 5956 6985 5972 7019
rect 5906 6945 5972 6985
rect 5906 6911 5922 6945
rect 5956 6911 5972 6945
rect 5906 6871 5972 6911
rect 5906 6837 5922 6871
rect 5956 6837 5972 6871
rect 5906 6821 5972 6837
rect 7016 7605 7082 7621
rect 7016 7571 7032 7605
rect 7066 7571 7082 7605
rect 7016 7532 7082 7571
rect 7016 7498 7032 7532
rect 7066 7498 7082 7532
rect 7016 7459 7082 7498
rect 7016 7425 7032 7459
rect 7066 7425 7082 7459
rect 7016 7386 7082 7425
rect 7016 7352 7032 7386
rect 7066 7352 7082 7386
rect 7016 7313 7082 7352
rect 7016 7279 7032 7313
rect 7066 7279 7082 7313
rect 7016 7240 7082 7279
rect 7016 7206 7032 7240
rect 7066 7206 7082 7240
rect 7016 7167 7082 7206
rect 7016 7133 7032 7167
rect 7066 7133 7082 7167
rect 7016 7093 7082 7133
rect 7016 7059 7032 7093
rect 7066 7059 7082 7093
rect 7016 7019 7082 7059
rect 7016 6985 7032 7019
rect 7066 6985 7082 7019
rect 7016 6945 7082 6985
rect 7016 6911 7032 6945
rect 7066 6911 7082 6945
rect 7016 6871 7082 6911
rect 7016 6837 7032 6871
rect 7066 6837 7082 6871
rect 7016 6821 7082 6837
rect 5906 6749 5972 6765
rect 5906 6715 5922 6749
rect 5956 6715 5972 6749
rect 5906 6676 5972 6715
rect 5906 6642 5922 6676
rect 5956 6642 5972 6676
rect 5906 6603 5972 6642
rect 5906 6569 5922 6603
rect 5956 6569 5972 6603
rect 5906 6530 5972 6569
rect 5906 6496 5922 6530
rect 5956 6496 5972 6530
rect 5906 6457 5972 6496
rect 5906 6423 5922 6457
rect 5956 6423 5972 6457
rect 5906 6384 5972 6423
rect 5906 6350 5922 6384
rect 5956 6350 5972 6384
rect 5906 6311 5972 6350
rect 5906 6277 5922 6311
rect 5956 6277 5972 6311
rect 5906 6237 5972 6277
rect 5906 6203 5922 6237
rect 5956 6203 5972 6237
rect 5906 6163 5972 6203
rect 5906 6129 5922 6163
rect 5956 6129 5972 6163
rect 5906 6089 5972 6129
rect 5906 6055 5922 6089
rect 5956 6055 5972 6089
rect 5906 6015 5972 6055
rect 5906 5981 5922 6015
rect 5956 5981 5972 6015
rect 5906 5965 5972 5981
rect 7016 6749 7082 6765
rect 7016 6715 7032 6749
rect 7066 6715 7082 6749
rect 7016 6676 7082 6715
rect 7016 6642 7032 6676
rect 7066 6642 7082 6676
rect 7016 6603 7082 6642
rect 7016 6569 7032 6603
rect 7066 6569 7082 6603
rect 7016 6530 7082 6569
rect 7016 6496 7032 6530
rect 7066 6496 7082 6530
rect 7016 6457 7082 6496
rect 7016 6423 7032 6457
rect 7066 6423 7082 6457
rect 7016 6384 7082 6423
rect 7016 6350 7032 6384
rect 7066 6350 7082 6384
rect 7016 6311 7082 6350
rect 7016 6277 7032 6311
rect 7066 6277 7082 6311
rect 7016 6237 7082 6277
rect 7016 6203 7032 6237
rect 7066 6203 7082 6237
rect 7016 6163 7082 6203
rect 7016 6129 7032 6163
rect 7066 6129 7082 6163
rect 7016 6089 7082 6129
rect 7016 6055 7032 6089
rect 7066 6055 7082 6089
rect 7016 6015 7082 6055
rect 7016 5981 7032 6015
rect 7066 5981 7082 6015
rect 7016 5965 7082 5981
rect 5906 5893 5972 5909
rect 5906 5859 5922 5893
rect 5956 5859 5972 5893
rect 5906 5820 5972 5859
rect 5906 5786 5922 5820
rect 5956 5786 5972 5820
rect 5906 5747 5972 5786
rect 5906 5713 5922 5747
rect 5956 5713 5972 5747
rect 5906 5674 5972 5713
rect 5906 5640 5922 5674
rect 5956 5640 5972 5674
rect 5906 5601 5972 5640
rect 5906 5567 5922 5601
rect 5956 5567 5972 5601
rect 5906 5528 5972 5567
rect 5906 5494 5922 5528
rect 5956 5494 5972 5528
rect 5906 5455 5972 5494
rect 5906 5421 5922 5455
rect 5956 5421 5972 5455
rect 5906 5381 5972 5421
rect 5906 5347 5922 5381
rect 5956 5347 5972 5381
rect 5906 5307 5972 5347
rect 5906 5273 5922 5307
rect 5956 5273 5972 5307
rect 5906 5233 5972 5273
rect 5906 5199 5922 5233
rect 5956 5199 5972 5233
rect 5906 5159 5972 5199
rect 5906 5125 5922 5159
rect 5956 5125 5972 5159
rect 5906 5109 5972 5125
rect 7016 5893 7082 5909
rect 7016 5859 7032 5893
rect 7066 5859 7082 5893
rect 7016 5820 7082 5859
rect 7016 5786 7032 5820
rect 7066 5786 7082 5820
rect 7016 5747 7082 5786
rect 7016 5713 7032 5747
rect 7066 5713 7082 5747
rect 7016 5674 7082 5713
rect 7016 5640 7032 5674
rect 7066 5640 7082 5674
rect 7016 5601 7082 5640
rect 7016 5567 7032 5601
rect 7066 5567 7082 5601
rect 7016 5528 7082 5567
rect 7016 5494 7032 5528
rect 7066 5494 7082 5528
rect 7016 5455 7082 5494
rect 7016 5421 7032 5455
rect 7066 5421 7082 5455
rect 7016 5381 7082 5421
rect 7016 5347 7032 5381
rect 7066 5347 7082 5381
rect 7016 5307 7082 5347
rect 7016 5273 7032 5307
rect 7066 5273 7082 5307
rect 7016 5233 7082 5273
rect 7016 5199 7032 5233
rect 7066 5199 7082 5233
rect 7016 5159 7082 5199
rect 7016 5125 7032 5159
rect 7066 5125 7082 5159
rect 7016 5109 7082 5125
rect 5906 5037 5972 5053
rect 5906 5003 5922 5037
rect 5956 5003 5972 5037
rect 5906 4964 5972 5003
rect 5906 4930 5922 4964
rect 5956 4930 5972 4964
rect 5906 4891 5972 4930
rect 5906 4857 5922 4891
rect 5956 4857 5972 4891
rect 5906 4818 5972 4857
rect 5906 4784 5922 4818
rect 5956 4784 5972 4818
rect 5906 4745 5972 4784
rect 5906 4711 5922 4745
rect 5956 4711 5972 4745
rect 5906 4672 5972 4711
rect 5906 4638 5922 4672
rect 5956 4638 5972 4672
rect 5906 4599 5972 4638
rect 5906 4565 5922 4599
rect 5956 4565 5972 4599
rect 5906 4525 5972 4565
rect 5906 4491 5922 4525
rect 5956 4491 5972 4525
rect 5906 4451 5972 4491
rect 5906 4417 5922 4451
rect 5956 4417 5972 4451
rect 5906 4377 5972 4417
rect 5906 4343 5922 4377
rect 5956 4343 5972 4377
rect 5906 4303 5972 4343
rect 5906 4269 5922 4303
rect 5956 4269 5972 4303
rect 5906 4253 5972 4269
rect 7016 5037 7082 5053
rect 7016 5003 7032 5037
rect 7066 5003 7082 5037
rect 7016 4964 7082 5003
rect 7016 4930 7032 4964
rect 7066 4930 7082 4964
rect 7016 4891 7082 4930
rect 7016 4857 7032 4891
rect 7066 4857 7082 4891
rect 7016 4818 7082 4857
rect 7016 4784 7032 4818
rect 7066 4784 7082 4818
rect 7016 4745 7082 4784
rect 7016 4711 7032 4745
rect 7066 4711 7082 4745
rect 7016 4672 7082 4711
rect 7016 4638 7032 4672
rect 7066 4638 7082 4672
rect 7016 4599 7082 4638
rect 7016 4565 7032 4599
rect 7066 4565 7082 4599
rect 7016 4525 7082 4565
rect 7016 4491 7032 4525
rect 7066 4491 7082 4525
rect 7016 4451 7082 4491
rect 7016 4417 7032 4451
rect 7066 4417 7082 4451
rect 7016 4377 7082 4417
rect 7016 4343 7032 4377
rect 7066 4343 7082 4377
rect 7016 4303 7082 4343
rect 7016 4269 7032 4303
rect 7066 4269 7082 4303
rect 7016 4253 7082 4269
rect 5906 4166 7082 4197
rect 5906 4132 5922 4166
rect 5956 4132 7032 4166
rect 7066 4132 7082 4166
rect 5906 4097 7082 4132
rect 7592 11224 7658 11240
rect 7592 11190 7608 11224
rect 7642 11190 7658 11224
rect 7592 11151 7658 11190
rect 7592 11117 7608 11151
rect 7642 11117 7658 11151
rect 7592 11078 7658 11117
rect 7592 11044 7608 11078
rect 7642 11044 7658 11078
rect 7592 11005 7658 11044
rect 7592 10971 7608 11005
rect 7642 10971 7658 11005
rect 7592 10932 7658 10971
rect 7592 10898 7608 10932
rect 7642 10898 7658 10932
rect 7592 10859 7658 10898
rect 7592 10825 7608 10859
rect 7642 10825 7658 10859
rect 7592 10786 7658 10825
rect 7592 10752 7608 10786
rect 7642 10752 7658 10786
rect 7592 10712 7658 10752
rect 7592 10678 7608 10712
rect 7642 10678 7658 10712
rect 7592 10638 7658 10678
rect 7592 10604 7608 10638
rect 7642 10604 7658 10638
rect 7592 10564 7658 10604
rect 7592 10530 7608 10564
rect 7642 10530 7658 10564
rect 7592 10490 7658 10530
rect 7592 10456 7608 10490
rect 7642 10456 7658 10490
rect 7592 10440 7658 10456
rect 9702 11224 9768 11240
rect 9702 11190 9718 11224
rect 9752 11190 9768 11224
rect 9702 11151 9768 11190
rect 9702 11117 9718 11151
rect 9752 11117 9768 11151
rect 9702 11078 9768 11117
rect 9702 11044 9718 11078
rect 9752 11044 9768 11078
rect 9702 11005 9768 11044
rect 9702 10971 9718 11005
rect 9752 10971 9768 11005
rect 9702 10932 9768 10971
rect 9702 10898 9718 10932
rect 9752 10898 9768 10932
rect 9702 10859 9768 10898
rect 9702 10825 9718 10859
rect 9752 10825 9768 10859
rect 9702 10786 9768 10825
rect 9702 10752 9718 10786
rect 9752 10752 9768 10786
rect 9702 10712 9768 10752
rect 9702 10678 9718 10712
rect 9752 10678 9768 10712
rect 9702 10638 9768 10678
rect 9702 10604 9718 10638
rect 9752 10604 9768 10638
rect 9702 10564 9768 10604
rect 9702 10530 9718 10564
rect 9752 10530 9768 10564
rect 9702 10490 9768 10530
rect 9702 10456 9718 10490
rect 9752 10456 9768 10490
rect 9702 10440 9768 10456
rect 7592 10138 7658 10154
rect 7592 10104 7608 10138
rect 7642 10104 7658 10138
rect 7592 10065 7658 10104
rect 7592 10031 7608 10065
rect 7642 10031 7658 10065
rect 7592 9992 7658 10031
rect 7592 9958 7608 9992
rect 7642 9958 7658 9992
rect 7592 9919 7658 9958
rect 7592 9885 7608 9919
rect 7642 9885 7658 9919
rect 7592 9846 7658 9885
rect 7592 9812 7608 9846
rect 7642 9812 7658 9846
rect 7592 9773 7658 9812
rect 7592 9739 7608 9773
rect 7642 9739 7658 9773
rect 7592 9700 7658 9739
rect 7592 9666 7608 9700
rect 7642 9666 7658 9700
rect 7592 9626 7658 9666
rect 7592 9592 7608 9626
rect 7642 9592 7658 9626
rect 7592 9552 7658 9592
rect 7592 9518 7608 9552
rect 7642 9518 7658 9552
rect 7592 9478 7658 9518
rect 7592 9444 7608 9478
rect 7642 9444 7658 9478
rect 7592 9404 7658 9444
rect 7592 9370 7608 9404
rect 7642 9370 7658 9404
rect 7592 9354 7658 9370
rect 9702 10138 9768 10154
rect 9702 10104 9718 10138
rect 9752 10104 9768 10138
rect 9702 10065 9768 10104
rect 9702 10031 9718 10065
rect 9752 10031 9768 10065
rect 9702 9992 9768 10031
rect 9702 9958 9718 9992
rect 9752 9958 9768 9992
rect 9702 9919 9768 9958
rect 9702 9885 9718 9919
rect 9752 9885 9768 9919
rect 9702 9846 9768 9885
rect 9702 9812 9718 9846
rect 9752 9812 9768 9846
rect 9702 9773 9768 9812
rect 9702 9739 9718 9773
rect 9752 9739 9768 9773
rect 9702 9700 9768 9739
rect 9702 9666 9718 9700
rect 9752 9666 9768 9700
rect 9702 9626 9768 9666
rect 9702 9592 9718 9626
rect 9752 9592 9768 9626
rect 9702 9552 9768 9592
rect 9702 9518 9718 9552
rect 9752 9518 9768 9552
rect 9702 9478 9768 9518
rect 9702 9444 9718 9478
rect 9752 9444 9768 9478
rect 9702 9404 9768 9444
rect 9702 9370 9718 9404
rect 9752 9370 9768 9404
rect 9702 9354 9768 9370
rect 7592 9282 7658 9298
rect 7592 9248 7608 9282
rect 7642 9248 7658 9282
rect 7592 9209 7658 9248
rect 7592 9175 7608 9209
rect 7642 9175 7658 9209
rect 7592 9136 7658 9175
rect 7592 9102 7608 9136
rect 7642 9102 7658 9136
rect 7592 9063 7658 9102
rect 7592 9029 7608 9063
rect 7642 9029 7658 9063
rect 7592 8990 7658 9029
rect 7592 8956 7608 8990
rect 7642 8956 7658 8990
rect 7592 8917 7658 8956
rect 7592 8883 7608 8917
rect 7642 8883 7658 8917
rect 7592 8844 7658 8883
rect 7592 8810 7608 8844
rect 7642 8810 7658 8844
rect 7592 8770 7658 8810
rect 7592 8736 7608 8770
rect 7642 8736 7658 8770
rect 7592 8696 7658 8736
rect 7592 8662 7608 8696
rect 7642 8662 7658 8696
rect 7592 8622 7658 8662
rect 7592 8588 7608 8622
rect 7642 8588 7658 8622
rect 7592 8548 7658 8588
rect 7592 8514 7608 8548
rect 7642 8514 7658 8548
rect 7592 8498 7658 8514
rect 9702 9282 9768 9298
rect 9702 9248 9718 9282
rect 9752 9248 9768 9282
rect 9702 9209 9768 9248
rect 9702 9175 9718 9209
rect 9752 9175 9768 9209
rect 9702 9136 9768 9175
rect 9702 9102 9718 9136
rect 9752 9102 9768 9136
rect 9702 9063 9768 9102
rect 9702 9029 9718 9063
rect 9752 9029 9768 9063
rect 9702 8990 9768 9029
rect 9702 8956 9718 8990
rect 9752 8956 9768 8990
rect 9702 8917 9768 8956
rect 9702 8883 9718 8917
rect 9752 8883 9768 8917
rect 9702 8844 9768 8883
rect 9702 8810 9718 8844
rect 9752 8810 9768 8844
rect 9702 8770 9768 8810
rect 9702 8736 9718 8770
rect 9752 8736 9768 8770
rect 9702 8696 9768 8736
rect 9702 8662 9718 8696
rect 9752 8662 9768 8696
rect 9702 8622 9768 8662
rect 9702 8588 9718 8622
rect 9752 8588 9768 8622
rect 9702 8548 9768 8588
rect 9702 8514 9718 8548
rect 9752 8514 9768 8548
rect 9702 8498 9768 8514
rect 7592 8196 7658 8212
rect 7592 8162 7608 8196
rect 7642 8162 7658 8196
rect 7592 8123 7658 8162
rect 7592 8089 7608 8123
rect 7642 8089 7658 8123
rect 7592 8050 7658 8089
rect 7592 8016 7608 8050
rect 7642 8016 7658 8050
rect 7592 7977 7658 8016
rect 7592 7943 7608 7977
rect 7642 7943 7658 7977
rect 7592 7904 7658 7943
rect 7592 7870 7608 7904
rect 7642 7870 7658 7904
rect 7592 7831 7658 7870
rect 7592 7797 7608 7831
rect 7642 7797 7658 7831
rect 7592 7758 7658 7797
rect 7592 7724 7608 7758
rect 7642 7724 7658 7758
rect 7592 7684 7658 7724
rect 7592 7650 7608 7684
rect 7642 7650 7658 7684
rect 7592 7610 7658 7650
rect 7592 7576 7608 7610
rect 7642 7576 7658 7610
rect 7592 7536 7658 7576
rect 7592 7502 7608 7536
rect 7642 7502 7658 7536
rect 7592 7462 7658 7502
rect 7592 7428 7608 7462
rect 7642 7428 7658 7462
rect 7592 7412 7658 7428
rect 9702 8196 9768 8212
rect 9702 8162 9718 8196
rect 9752 8162 9768 8196
rect 9702 8123 9768 8162
rect 9702 8089 9718 8123
rect 9752 8089 9768 8123
rect 9702 8050 9768 8089
rect 9702 8016 9718 8050
rect 9752 8016 9768 8050
rect 9702 7977 9768 8016
rect 9702 7943 9718 7977
rect 9752 7943 9768 7977
rect 9702 7904 9768 7943
rect 9702 7870 9718 7904
rect 9752 7870 9768 7904
rect 9702 7831 9768 7870
rect 9702 7797 9718 7831
rect 9752 7797 9768 7831
rect 9702 7758 9768 7797
rect 9702 7724 9718 7758
rect 9752 7724 9768 7758
rect 9702 7684 9768 7724
rect 9702 7650 9718 7684
rect 9752 7650 9768 7684
rect 9702 7610 9768 7650
rect 9702 7576 9718 7610
rect 9752 7576 9768 7610
rect 9702 7536 9768 7576
rect 9702 7502 9718 7536
rect 9752 7502 9768 7536
rect 9702 7462 9768 7502
rect 9702 7428 9718 7462
rect 9752 7428 9768 7462
rect 9702 7412 9768 7428
rect 7592 6464 7658 6480
rect 7592 6430 7608 6464
rect 7642 6430 7658 6464
rect 7592 6395 7658 6430
rect 7592 6361 7608 6395
rect 7642 6361 7658 6395
rect 7592 6326 7658 6361
rect 7592 6292 7608 6326
rect 7642 6292 7658 6326
rect 7592 6257 7658 6292
rect 7592 6223 7608 6257
rect 7642 6223 7658 6257
rect 7592 6188 7658 6223
rect 7592 6154 7608 6188
rect 7642 6154 7658 6188
rect 7592 6119 7658 6154
rect 7592 6085 7608 6119
rect 7642 6085 7658 6119
rect 7592 6050 7658 6085
rect 7592 6016 7608 6050
rect 7642 6016 7658 6050
rect 7592 5981 7658 6016
rect 7592 5947 7608 5981
rect 7642 5947 7658 5981
rect 7592 5912 7658 5947
rect 7592 5878 7608 5912
rect 7642 5878 7658 5912
rect 7592 5843 7658 5878
rect 7592 5809 7608 5843
rect 7642 5809 7658 5843
rect 7592 5774 7658 5809
rect 7592 5740 7608 5774
rect 7642 5740 7658 5774
rect 7592 5704 7658 5740
rect 7592 5670 7608 5704
rect 7642 5670 7658 5704
rect 7592 5654 7658 5670
rect 9702 6464 9768 6480
rect 9702 6430 9718 6464
rect 9752 6430 9768 6464
rect 9702 6395 9768 6430
rect 9702 6361 9718 6395
rect 9752 6361 9768 6395
rect 9702 6326 9768 6361
rect 9702 6292 9718 6326
rect 9752 6292 9768 6326
rect 9702 6257 9768 6292
rect 9702 6223 9718 6257
rect 9752 6223 9768 6257
rect 9702 6188 9768 6223
rect 9702 6154 9718 6188
rect 9752 6154 9768 6188
rect 9702 6119 9768 6154
rect 9702 6085 9718 6119
rect 9752 6085 9768 6119
rect 9702 6050 9768 6085
rect 9702 6016 9718 6050
rect 9752 6016 9768 6050
rect 9702 5981 9768 6016
rect 9702 5947 9718 5981
rect 9752 5947 9768 5981
rect 9702 5912 9768 5947
rect 9702 5878 9718 5912
rect 9752 5878 9768 5912
rect 9702 5843 9768 5878
rect 9702 5809 9718 5843
rect 9752 5809 9768 5843
rect 9702 5774 9768 5809
rect 9702 5740 9718 5774
rect 9752 5740 9768 5774
rect 9702 5704 9768 5740
rect 9702 5670 9718 5704
rect 9752 5670 9768 5704
rect 9702 5654 9768 5670
rect 7592 5378 7658 5394
rect 7592 5344 7608 5378
rect 7642 5344 7658 5378
rect 7592 5305 7658 5344
rect 7592 5271 7608 5305
rect 7642 5271 7658 5305
rect 7592 5232 7658 5271
rect 7592 5198 7608 5232
rect 7642 5198 7658 5232
rect 7592 5159 7658 5198
rect 7592 5125 7608 5159
rect 7642 5125 7658 5159
rect 7592 5086 7658 5125
rect 7592 5052 7608 5086
rect 7642 5052 7658 5086
rect 7592 5013 7658 5052
rect 7592 4979 7608 5013
rect 7642 4979 7658 5013
rect 7592 4940 7658 4979
rect 7592 4906 7608 4940
rect 7642 4906 7658 4940
rect 7592 4866 7658 4906
rect 7592 4832 7608 4866
rect 7642 4832 7658 4866
rect 7592 4792 7658 4832
rect 7592 4758 7608 4792
rect 7642 4758 7658 4792
rect 7592 4718 7658 4758
rect 7592 4684 7608 4718
rect 7642 4684 7658 4718
rect 7592 4644 7658 4684
rect 7592 4610 7608 4644
rect 7642 4610 7658 4644
rect 7592 4594 7658 4610
rect 9702 5378 9768 5394
rect 9702 5344 9718 5378
rect 9752 5344 9768 5378
rect 9702 5305 9768 5344
rect 9702 5271 9718 5305
rect 9752 5271 9768 5305
rect 9702 5232 9768 5271
rect 9702 5198 9718 5232
rect 9752 5198 9768 5232
rect 9702 5159 9768 5198
rect 9702 5125 9718 5159
rect 9752 5125 9768 5159
rect 9702 5086 9768 5125
rect 9702 5052 9718 5086
rect 9752 5052 9768 5086
rect 9702 5013 9768 5052
rect 9702 4979 9718 5013
rect 9752 4979 9768 5013
rect 9702 4940 9768 4979
rect 9702 4906 9718 4940
rect 9752 4906 9768 4940
rect 9702 4866 9768 4906
rect 9702 4832 9718 4866
rect 9752 4832 9768 4866
rect 9702 4792 9768 4832
rect 9702 4758 9718 4792
rect 9752 4758 9768 4792
rect 9702 4718 9768 4758
rect 9702 4684 9718 4718
rect 9752 4684 9768 4718
rect 9702 4644 9768 4684
rect 9702 4610 9718 4644
rect 9752 4610 9768 4644
rect 9702 4594 9768 4610
rect 7592 4522 7658 4538
rect 7592 4488 7608 4522
rect 7642 4488 7658 4522
rect 7592 4449 7658 4488
rect 7592 4415 7608 4449
rect 7642 4415 7658 4449
rect 7592 4376 7658 4415
rect 7592 4342 7608 4376
rect 7642 4342 7658 4376
rect 7592 4303 7658 4342
rect 7592 4269 7608 4303
rect 7642 4269 7658 4303
rect 7592 4230 7658 4269
rect 7592 4196 7608 4230
rect 7642 4196 7658 4230
rect 7592 4157 7658 4196
rect 7592 4123 7608 4157
rect 7642 4123 7658 4157
rect 7592 4084 7658 4123
rect 7592 4050 7608 4084
rect 7642 4050 7658 4084
rect 7592 4010 7658 4050
rect 7592 3976 7608 4010
rect 7642 3976 7658 4010
rect 7592 3936 7658 3976
rect 7592 3902 7608 3936
rect 7642 3902 7658 3936
rect 7592 3862 7658 3902
rect 7592 3828 7608 3862
rect 7642 3828 7658 3862
rect 7592 3788 7658 3828
rect 7592 3754 7608 3788
rect 7642 3754 7658 3788
rect 7592 3738 7658 3754
rect 9702 4522 9768 4538
rect 9702 4488 9718 4522
rect 9752 4488 9768 4522
rect 9702 4449 9768 4488
rect 9702 4415 9718 4449
rect 9752 4415 9768 4449
rect 9702 4376 9768 4415
rect 9702 4342 9718 4376
rect 9752 4342 9768 4376
rect 9702 4303 9768 4342
rect 9702 4269 9718 4303
rect 9752 4269 9768 4303
rect 9702 4230 9768 4269
rect 9702 4196 9718 4230
rect 9752 4196 9768 4230
rect 9702 4157 9768 4196
rect 9702 4123 9718 4157
rect 9752 4123 9768 4157
rect 9702 4084 9768 4123
rect 9702 4050 9718 4084
rect 9752 4050 9768 4084
rect 9702 4010 9768 4050
rect 9702 3976 9718 4010
rect 9752 3976 9768 4010
rect 9702 3936 9768 3976
rect 9702 3902 9718 3936
rect 9752 3902 9768 3936
rect 9702 3862 9768 3902
rect 9702 3828 9718 3862
rect 9752 3828 9768 3862
rect 9702 3788 9768 3828
rect 9702 3754 9718 3788
rect 9752 3754 9768 3788
rect 9702 3738 9768 3754
rect 1380 3436 1446 3452
rect 1380 3402 1396 3436
rect 1430 3402 1446 3436
rect 1380 3363 1446 3402
rect 1380 3329 1396 3363
rect 1430 3329 1446 3363
rect 1380 3290 1446 3329
rect 1380 3256 1396 3290
rect 1430 3256 1446 3290
rect 1380 3217 1446 3256
rect 1380 3183 1396 3217
rect 1430 3183 1446 3217
rect 1380 3144 1446 3183
rect 1380 3110 1396 3144
rect 1430 3110 1446 3144
rect 1380 3071 1446 3110
rect 1380 3037 1396 3071
rect 1430 3037 1446 3071
rect 1380 2998 1446 3037
rect 1380 2964 1396 2998
rect 1430 2964 1446 2998
rect 1380 2924 1446 2964
rect 1380 2890 1396 2924
rect 1430 2890 1446 2924
rect 1380 2850 1446 2890
rect 1380 2816 1396 2850
rect 1430 2816 1446 2850
rect 1380 2776 1446 2816
rect 1380 2742 1396 2776
rect 1430 2742 1446 2776
rect 1380 2702 1446 2742
rect 1380 2668 1396 2702
rect 1430 2668 1446 2702
rect 1380 2652 1446 2668
rect 3490 3436 3556 3452
rect 3490 3402 3506 3436
rect 3540 3402 3556 3436
rect 3490 3363 3556 3402
rect 3490 3329 3506 3363
rect 3540 3329 3556 3363
rect 3490 3290 3556 3329
rect 3490 3256 3506 3290
rect 3540 3256 3556 3290
rect 3490 3217 3556 3256
rect 3490 3183 3506 3217
rect 3540 3183 3556 3217
rect 3490 3144 3556 3183
rect 3490 3110 3506 3144
rect 3540 3110 3556 3144
rect 3490 3071 3556 3110
rect 3490 3037 3506 3071
rect 3540 3037 3556 3071
rect 3490 2998 3556 3037
rect 3490 2964 3506 2998
rect 3540 2964 3556 2998
rect 3490 2924 3556 2964
rect 3490 2890 3506 2924
rect 3540 2890 3556 2924
rect 3490 2850 3556 2890
rect 3490 2816 3506 2850
rect 3540 2816 3556 2850
rect 3490 2776 3556 2816
rect 3490 2742 3506 2776
rect 3540 2742 3556 2776
rect 3490 2702 3556 2742
rect 3490 2668 3506 2702
rect 3540 2668 3556 2702
rect 3490 2652 3556 2668
rect 5178 3311 5244 3327
rect 5178 3277 5194 3311
rect 5228 3277 5244 3311
rect 5178 3243 5244 3277
rect 5178 3209 5194 3243
rect 5228 3209 5244 3243
rect 5178 3175 5244 3209
rect 5178 3141 5194 3175
rect 5228 3141 5244 3175
rect 5178 3125 5244 3141
rect 7016 3311 7082 3327
rect 7016 3277 7032 3311
rect 7066 3277 7082 3311
rect 7016 3243 7082 3277
rect 7016 3209 7032 3243
rect 7066 3209 7082 3243
rect 7016 3175 7082 3209
rect 7016 3141 7032 3175
rect 7066 3141 7082 3175
rect 7016 3125 7082 3141
rect 5178 3020 5244 3069
rect 5178 2986 5194 3020
rect 5228 2986 5244 3020
rect 5178 2952 5244 2986
rect 5178 2918 5194 2952
rect 5228 2918 5244 2952
rect 5178 2869 5244 2918
rect 5178 2764 5244 2813
rect 5178 2730 5194 2764
rect 5228 2730 5244 2764
rect 5178 2696 5244 2730
rect 5178 2662 5194 2696
rect 5228 2662 5244 2696
rect 5178 2613 5244 2662
rect 5696 3048 5762 3087
rect 5696 3014 5712 3048
rect 5746 3014 5762 3048
rect 5696 2980 5762 3014
rect 5696 2946 5712 2980
rect 5746 2946 5762 2980
rect 5696 2671 5762 2946
rect 7016 3020 7082 3069
rect 7016 2986 7032 3020
rect 7066 2986 7082 3020
rect 7016 2952 7082 2986
rect 7016 2918 7032 2952
rect 7066 2918 7082 2952
rect 7016 2869 7082 2918
rect 5178 2508 5244 2557
rect 5178 2474 5194 2508
rect 5228 2474 5244 2508
rect 5178 2440 5244 2474
rect 5178 2406 5194 2440
rect 5228 2406 5244 2440
rect 5178 2357 5244 2406
rect 7016 2764 7082 2813
rect 7016 2730 7032 2764
rect 7066 2730 7082 2764
rect 7016 2696 7082 2730
rect 7016 2662 7032 2696
rect 7066 2662 7082 2696
rect 7016 2613 7082 2662
rect 7016 2508 7082 2557
rect 7016 2474 7032 2508
rect 7066 2474 7082 2508
rect 7016 2440 7082 2474
rect 7016 2406 7032 2440
rect 7066 2406 7082 2440
rect 7016 2357 7082 2406
rect 5178 2252 5244 2301
rect 5178 2218 5194 2252
rect 5228 2218 5244 2252
rect 5178 2184 5244 2218
rect 5178 2150 5194 2184
rect 5228 2150 5244 2184
rect 5178 2101 5244 2150
rect 7016 2252 7082 2301
rect 7016 2218 7032 2252
rect 7066 2218 7082 2252
rect 7016 2184 7082 2218
rect 7016 2150 7032 2184
rect 7066 2150 7082 2184
rect 7016 2101 7082 2150
rect 7592 3436 7658 3452
rect 7592 3402 7608 3436
rect 7642 3402 7658 3436
rect 7592 3363 7658 3402
rect 7592 3329 7608 3363
rect 7642 3329 7658 3363
rect 7592 3290 7658 3329
rect 7592 3256 7608 3290
rect 7642 3256 7658 3290
rect 7592 3217 7658 3256
rect 7592 3183 7608 3217
rect 7642 3183 7658 3217
rect 7592 3144 7658 3183
rect 7592 3110 7608 3144
rect 7642 3110 7658 3144
rect 7592 3071 7658 3110
rect 7592 3037 7608 3071
rect 7642 3037 7658 3071
rect 7592 2998 7658 3037
rect 7592 2964 7608 2998
rect 7642 2964 7658 2998
rect 7592 2924 7658 2964
rect 7592 2890 7608 2924
rect 7642 2890 7658 2924
rect 7592 2850 7658 2890
rect 7592 2816 7608 2850
rect 7642 2816 7658 2850
rect 7592 2776 7658 2816
rect 7592 2742 7608 2776
rect 7642 2742 7658 2776
rect 7592 2702 7658 2742
rect 7592 2668 7608 2702
rect 7642 2668 7658 2702
rect 7592 2652 7658 2668
rect 9702 3436 9768 3452
rect 9702 3402 9718 3436
rect 9752 3402 9768 3436
rect 9702 3363 9768 3402
rect 9702 3329 9718 3363
rect 9752 3329 9768 3363
rect 9702 3290 9768 3329
rect 9702 3256 9718 3290
rect 9752 3256 9768 3290
rect 9702 3217 9768 3256
rect 9702 3183 9718 3217
rect 9752 3183 9768 3217
rect 9702 3144 9768 3183
rect 9702 3110 9718 3144
rect 9752 3110 9768 3144
rect 9702 3071 9768 3110
rect 9702 3037 9718 3071
rect 9752 3037 9768 3071
rect 9702 2998 9768 3037
rect 9702 2964 9718 2998
rect 9752 2964 9768 2998
rect 9702 2924 9768 2964
rect 9702 2890 9718 2924
rect 9752 2890 9768 2924
rect 9702 2850 9768 2890
rect 9702 2816 9718 2850
rect 9752 2816 9768 2850
rect 9702 2776 9768 2816
rect 9702 2742 9718 2776
rect 9752 2742 9768 2776
rect 9702 2702 9768 2742
rect 9702 2668 9718 2702
rect 9752 2668 9768 2702
rect 9702 2652 9768 2668
rect 5178 1996 5244 2045
rect 5178 1962 5194 1996
rect 5228 1962 5244 1996
rect 5178 1928 5244 1962
rect 5178 1894 5194 1928
rect 5228 1894 5244 1928
rect 5178 1845 5244 1894
rect 7016 1996 7082 2045
rect 7016 1962 7032 1996
rect 7066 1962 7082 1996
rect 7016 1928 7082 1962
rect 7016 1894 7032 1928
rect 7066 1894 7082 1928
rect 7016 1845 7082 1894
rect 1380 1743 1446 1759
rect 1380 1709 1396 1743
rect 1430 1709 1446 1743
rect 1380 1670 1446 1709
rect 1380 1636 1396 1670
rect 1430 1636 1446 1670
rect 1380 1597 1446 1636
rect 1380 1563 1396 1597
rect 1430 1563 1446 1597
rect 1380 1524 1446 1563
rect 1380 1490 1396 1524
rect 1430 1490 1446 1524
rect 1380 1451 1446 1490
rect 1380 1417 1396 1451
rect 1430 1417 1446 1451
rect 1380 1378 1446 1417
rect 1380 1344 1396 1378
rect 1430 1344 1446 1378
rect 1380 1305 1446 1344
rect 1380 1271 1396 1305
rect 1430 1271 1446 1305
rect 1380 1231 1446 1271
rect 1380 1197 1396 1231
rect 1430 1197 1446 1231
rect 1380 1157 1446 1197
rect 1380 1123 1396 1157
rect 1430 1123 1446 1157
rect 1380 1083 1446 1123
rect 1380 1049 1396 1083
rect 1430 1049 1446 1083
rect 1380 1009 1446 1049
rect 1380 975 1396 1009
rect 1430 975 1446 1009
rect 1380 959 1446 975
rect 3490 1743 3556 1759
rect 3490 1709 3506 1743
rect 3540 1709 3556 1743
rect 3490 1670 3556 1709
rect 3490 1636 3506 1670
rect 3540 1636 3556 1670
rect 3490 1597 3556 1636
rect 3490 1563 3506 1597
rect 3540 1563 3556 1597
rect 3490 1524 3556 1563
rect 3490 1490 3506 1524
rect 3540 1490 3556 1524
rect 3490 1451 3556 1490
rect 3490 1417 3506 1451
rect 3540 1417 3556 1451
rect 3490 1378 3556 1417
rect 3490 1344 3506 1378
rect 3540 1344 3556 1378
rect 3490 1305 3556 1344
rect 3490 1271 3506 1305
rect 3540 1271 3556 1305
rect 3490 1231 3556 1271
rect 3490 1197 3506 1231
rect 3540 1197 3556 1231
rect 3490 1157 3556 1197
rect 3490 1123 3506 1157
rect 3540 1123 3556 1157
rect 3490 1083 3556 1123
rect 3490 1049 3506 1083
rect 3540 1049 3556 1083
rect 3490 1009 3556 1049
rect 3490 975 3506 1009
rect 3540 975 3556 1009
rect 3490 959 3556 975
rect 5178 1740 5244 1789
rect 5178 1706 5194 1740
rect 5228 1706 5244 1740
rect 5178 1672 5244 1706
rect 5178 1638 5194 1672
rect 5228 1638 5244 1672
rect 5178 1589 5244 1638
rect 7016 1740 7082 1789
rect 7016 1706 7032 1740
rect 7066 1706 7082 1740
rect 7016 1672 7082 1706
rect 7016 1638 7032 1672
rect 7066 1638 7082 1672
rect 7016 1589 7082 1638
rect 5178 1484 5244 1533
rect 5178 1450 5194 1484
rect 5228 1450 5244 1484
rect 5178 1416 5244 1450
rect 5178 1382 5194 1416
rect 5228 1382 5244 1416
rect 5178 1333 5244 1382
rect 7016 1484 7082 1533
rect 7016 1450 7032 1484
rect 7066 1450 7082 1484
rect 7016 1416 7082 1450
rect 7016 1382 7032 1416
rect 7066 1382 7082 1416
rect 7016 1333 7082 1382
rect 5178 1228 5244 1277
rect 5178 1194 5194 1228
rect 5228 1194 5244 1228
rect 5178 1160 5244 1194
rect 5178 1126 5194 1160
rect 5228 1126 5244 1160
rect 5178 1077 5244 1126
rect 7016 1228 7082 1277
rect 7016 1194 7032 1228
rect 7066 1194 7082 1228
rect 7016 1160 7082 1194
rect 7016 1126 7032 1160
rect 7066 1126 7082 1160
rect 7016 1077 7082 1126
rect 5178 1005 5244 1021
rect 5178 971 5194 1005
rect 5228 971 5244 1005
rect 5178 937 5244 971
rect 5178 903 5194 937
rect 5228 903 5244 937
rect 5178 887 5244 903
rect 1583 826 1783 842
rect 1583 792 1599 826
rect 1633 792 1733 826
rect 1767 792 1783 826
rect 1583 776 1783 792
rect 1892 800 2049 816
rect 1892 766 1908 800
rect 1942 766 1976 800
rect 2010 766 2049 800
rect 1892 750 2049 766
rect 2105 800 2305 816
rect 2105 766 2154 800
rect 2188 766 2222 800
rect 2256 766 2305 800
rect 2105 754 2305 766
rect 2361 800 2561 816
rect 2361 766 2410 800
rect 2444 766 2478 800
rect 2512 766 2561 800
rect 2361 754 2561 766
rect 2617 800 2817 816
rect 2617 766 2666 800
rect 2700 766 2734 800
rect 2768 766 2817 800
rect 2617 754 2817 766
rect 2873 800 3073 816
rect 2873 766 2922 800
rect 2956 766 2990 800
rect 3024 766 3073 800
rect 2873 754 3073 766
rect 3129 800 3329 816
rect 3129 766 3178 800
rect 3212 766 3246 800
rect 3280 766 3329 800
rect 3129 754 3329 766
rect 3385 800 3542 816
rect 3385 766 3424 800
rect 3458 766 3492 800
rect 3526 766 3542 800
rect 2138 750 2272 754
rect 2394 750 2528 754
rect 2650 750 2784 754
rect 2906 750 3040 754
rect 3162 750 3296 754
rect 3385 750 3542 766
rect 1949 582 2049 750
rect 3385 582 3485 750
rect 7016 1005 7082 1021
rect 7016 971 7032 1005
rect 7066 971 7082 1005
rect 7016 937 7082 971
rect 7016 903 7032 937
rect 7066 903 7082 937
rect 7016 887 7082 903
rect 7592 1743 7658 1759
rect 7592 1709 7608 1743
rect 7642 1709 7658 1743
rect 7592 1670 7658 1709
rect 7592 1636 7608 1670
rect 7642 1636 7658 1670
rect 7592 1597 7658 1636
rect 7592 1563 7608 1597
rect 7642 1563 7658 1597
rect 7592 1524 7658 1563
rect 7592 1490 7608 1524
rect 7642 1490 7658 1524
rect 7592 1451 7658 1490
rect 7592 1417 7608 1451
rect 7642 1417 7658 1451
rect 7592 1378 7658 1417
rect 7592 1344 7608 1378
rect 7642 1344 7658 1378
rect 7592 1305 7658 1344
rect 7592 1271 7608 1305
rect 7642 1271 7658 1305
rect 7592 1231 7658 1271
rect 7592 1197 7608 1231
rect 7642 1197 7658 1231
rect 7592 1157 7658 1197
rect 7592 1123 7608 1157
rect 7642 1123 7658 1157
rect 7592 1083 7658 1123
rect 7592 1049 7608 1083
rect 7642 1049 7658 1083
rect 7592 1009 7658 1049
rect 7592 975 7608 1009
rect 7642 975 7658 1009
rect 7592 959 7658 975
rect 9702 1743 9768 1759
rect 9702 1709 9718 1743
rect 9752 1709 9768 1743
rect 9702 1670 9768 1709
rect 9702 1636 9718 1670
rect 9752 1636 9768 1670
rect 9702 1597 9768 1636
rect 9702 1563 9718 1597
rect 9752 1563 9768 1597
rect 9702 1524 9768 1563
rect 9702 1490 9718 1524
rect 9752 1490 9768 1524
rect 9702 1451 9768 1490
rect 9702 1417 9718 1451
rect 9752 1417 9768 1451
rect 9702 1378 9768 1417
rect 9702 1344 9718 1378
rect 9752 1344 9768 1378
rect 9702 1305 9768 1344
rect 9702 1271 9718 1305
rect 9752 1271 9768 1305
rect 9702 1231 9768 1271
rect 9702 1197 9718 1231
rect 9752 1197 9768 1231
rect 9702 1157 9768 1197
rect 9702 1123 9718 1157
rect 9752 1123 9768 1157
rect 9702 1083 9768 1123
rect 9702 1049 9718 1083
rect 9752 1049 9768 1083
rect 9702 1009 9768 1049
rect 9702 975 9718 1009
rect 9752 975 9768 1009
rect 9702 959 9768 975
rect 5176 712 5242 755
rect 5176 678 5192 712
rect 5226 678 5242 712
rect 5176 644 5242 678
rect 5176 610 5192 644
rect 5226 610 5242 644
rect 5176 576 5242 610
rect 5176 542 5192 576
rect 5226 542 5242 576
rect 5176 499 5242 542
rect 6644 712 7082 755
rect 6644 678 7032 712
rect 7066 678 7082 712
rect 6644 655 7082 678
rect 7016 644 7082 655
rect 7016 610 7032 644
rect 7066 610 7082 644
rect 7016 599 7082 610
rect 6644 576 7082 599
rect 6644 542 7032 576
rect 7066 542 7082 576
rect 6644 499 7082 542
rect 7606 800 7763 816
rect 7606 766 7622 800
rect 7656 766 7690 800
rect 7724 766 7763 800
rect 7606 750 7763 766
rect 7819 800 8019 816
rect 7819 766 7868 800
rect 7902 766 7936 800
rect 7970 766 8019 800
rect 7819 754 8019 766
rect 8075 800 8275 816
rect 8075 766 8124 800
rect 8158 766 8192 800
rect 8226 766 8275 800
rect 8075 754 8275 766
rect 8331 800 8531 816
rect 8331 766 8380 800
rect 8414 766 8448 800
rect 8482 766 8531 800
rect 8331 754 8531 766
rect 8587 800 8787 816
rect 8587 766 8636 800
rect 8670 766 8704 800
rect 8738 766 8787 800
rect 8587 754 8787 766
rect 8843 800 9043 816
rect 8843 766 8892 800
rect 8926 766 8960 800
rect 8994 766 9043 800
rect 8843 754 9043 766
rect 9099 800 9256 816
rect 9099 766 9138 800
rect 9172 766 9206 800
rect 9240 766 9256 800
rect 7852 750 7986 754
rect 8108 750 8242 754
rect 8364 750 8498 754
rect 8620 750 8754 754
rect 8876 750 9010 754
rect 9099 750 9256 766
rect 7663 582 7763 750
rect 9099 582 9199 750
<< polycont >>
rect 1757 14043 1791 14077
rect 1757 13973 1791 14007
rect 1757 13903 1791 13937
rect 1757 13833 1791 13867
rect 1757 13763 1791 13797
rect 1757 13693 1791 13727
rect 1757 13623 1791 13657
rect 1757 13553 1791 13587
rect 1757 13483 1791 13517
rect 1757 13413 1791 13447
rect 1757 13343 1791 13377
rect 1757 13273 1791 13307
rect 1757 13203 1791 13237
rect 1757 13133 1791 13167
rect 1757 13063 1791 13097
rect 1757 12993 1791 13027
rect 1757 12923 1791 12957
rect 1757 12854 1791 12888
rect 1757 12785 1791 12819
rect 1757 12716 1791 12750
rect 1757 12647 1791 12681
rect 1757 12578 1791 12612
rect 1757 12509 1791 12543
rect 3287 14043 3321 14077
rect 3287 13973 3321 14007
rect 4245 14013 4279 14047
rect 3287 13903 3321 13937
rect 3287 13833 3321 13867
rect 3407 13919 3441 13953
rect 3407 13851 3441 13885
rect 4137 13919 4171 13953
rect 4245 13945 4279 13979
rect 4975 14013 5009 14047
rect 4975 13945 5009 13979
rect 6085 14013 6119 14047
rect 7761 14043 7795 14077
rect 6085 13945 6119 13979
rect 4137 13851 4171 13885
rect 7761 13973 7795 14007
rect 5284 13887 5318 13921
rect 5356 13887 5390 13921
rect 5428 13887 5462 13921
rect 5500 13887 5534 13921
rect 5572 13887 5606 13921
rect 5644 13887 5678 13921
rect 5715 13887 5749 13921
rect 5786 13887 5820 13921
rect 6923 13919 6957 13953
rect 3287 13763 3321 13797
rect 4245 13800 4279 13834
rect 3287 13693 3321 13727
rect 3287 13623 3321 13657
rect 3287 13553 3321 13587
rect 3407 13706 3441 13740
rect 3407 13618 3441 13652
rect 4137 13706 4171 13740
rect 4245 13712 4279 13746
rect 4975 13800 5009 13834
rect 4975 13712 5009 13746
rect 4137 13618 4171 13652
rect 4245 13544 4279 13578
rect 3287 13483 3321 13517
rect 3287 13413 3321 13447
rect 3287 13343 3321 13377
rect 3407 13450 3441 13484
rect 3407 13362 3441 13396
rect 4137 13450 4171 13484
rect 4245 13456 4279 13490
rect 4975 13544 5009 13578
rect 4975 13456 5009 13490
rect 4137 13362 4171 13396
rect 3287 13273 3321 13307
rect 4245 13288 4279 13322
rect 3287 13203 3321 13237
rect 3287 13133 3321 13167
rect 3287 13063 3321 13097
rect 3407 13194 3441 13228
rect 3407 13106 3441 13140
rect 4137 13194 4171 13228
rect 4245 13200 4279 13234
rect 4975 13288 5009 13322
rect 4975 13200 5009 13234
rect 4137 13106 4171 13140
rect 3287 12993 3321 13027
rect 4245 13032 4279 13066
rect 3287 12923 3321 12957
rect 3287 12854 3321 12888
rect 3287 12785 3321 12819
rect 3407 12938 3441 12972
rect 3407 12850 3441 12884
rect 4137 12938 4171 12972
rect 4245 12944 4279 12978
rect 4975 13031 5009 13065
rect 4975 12943 5009 12977
rect 4137 12850 4171 12884
rect 6085 13800 6119 13834
rect 6085 13712 6119 13746
rect 6923 13851 6957 13885
rect 7653 13919 7687 13953
rect 7653 13851 7687 13885
rect 7761 13903 7795 13937
rect 6815 13800 6849 13834
rect 7761 13833 7795 13867
rect 6815 13712 6849 13746
rect 6923 13706 6957 13740
rect 6923 13618 6957 13652
rect 6085 13544 6119 13578
rect 6085 13456 6119 13490
rect 7653 13706 7687 13740
rect 7653 13618 7687 13652
rect 7761 13763 7795 13797
rect 7761 13693 7795 13727
rect 7761 13623 7795 13657
rect 6815 13544 6849 13578
rect 7761 13553 7795 13587
rect 6815 13456 6849 13490
rect 6923 13450 6957 13484
rect 6923 13362 6957 13396
rect 6085 13288 6119 13322
rect 6085 13200 6119 13234
rect 7653 13450 7687 13484
rect 7653 13362 7687 13396
rect 7761 13483 7795 13517
rect 7761 13413 7795 13447
rect 7761 13343 7795 13377
rect 6815 13288 6849 13322
rect 7761 13273 7795 13307
rect 6815 13200 6849 13234
rect 6923 13194 6957 13228
rect 6923 13106 6957 13140
rect 6085 13032 6119 13066
rect 6085 12944 6119 12978
rect 7653 13194 7687 13228
rect 7653 13106 7687 13140
rect 7761 13203 7795 13237
rect 7761 13133 7795 13167
rect 6815 13031 6849 13065
rect 7761 13063 7795 13097
rect 6815 12943 6849 12977
rect 6923 12938 6957 12972
rect 6923 12850 6957 12884
rect 4245 12776 4279 12810
rect 3287 12716 3321 12750
rect 3287 12647 3321 12681
rect 3407 12705 3441 12739
rect 3407 12637 3441 12671
rect 4137 12705 4171 12739
rect 4137 12637 4171 12671
rect 4245 12688 4279 12722
rect 4975 12776 5009 12810
rect 5273 12757 5307 12791
rect 5347 12757 5381 12791
rect 5421 12757 5455 12791
rect 5495 12757 5529 12791
rect 5568 12757 5602 12791
rect 5641 12757 5675 12791
rect 5714 12757 5748 12791
rect 5787 12757 5821 12791
rect 6085 12776 6119 12810
rect 4975 12688 5009 12722
rect 3287 12578 3321 12612
rect 3287 12509 3321 12543
rect 4245 12543 4279 12577
rect 4245 12475 4279 12509
rect 4975 12543 5009 12577
rect 4975 12475 5009 12509
rect 6085 12688 6119 12722
rect 7653 12938 7687 12972
rect 7653 12850 7687 12884
rect 7761 12993 7795 13027
rect 7761 12923 7795 12957
rect 7761 12854 7795 12888
rect 6815 12776 6849 12810
rect 7761 12785 7795 12819
rect 6815 12688 6849 12722
rect 6923 12705 6957 12739
rect 6923 12637 6957 12671
rect 7653 12705 7687 12739
rect 7653 12637 7687 12671
rect 7761 12716 7795 12750
rect 7761 12647 7795 12681
rect 1422 12424 1456 12458
rect 1552 12424 1586 12458
rect 5502 12424 5536 12458
rect 5570 12424 5604 12458
rect 6815 12543 6849 12577
rect 6815 12475 6849 12509
rect 7761 12578 7795 12612
rect 7761 12509 7795 12543
rect 9291 14043 9325 14077
rect 9291 13973 9325 14007
rect 9291 13903 9325 13937
rect 9291 13833 9325 13867
rect 9291 13763 9325 13797
rect 9291 13693 9325 13727
rect 9291 13623 9325 13657
rect 9291 13553 9325 13587
rect 9291 13483 9325 13517
rect 9291 13413 9325 13447
rect 9291 13343 9325 13377
rect 9291 13273 9325 13307
rect 9291 13203 9325 13237
rect 9291 13133 9325 13167
rect 9291 13063 9325 13097
rect 9291 12993 9325 13027
rect 9291 12923 9325 12957
rect 9291 12854 9325 12888
rect 9291 12785 9325 12819
rect 9291 12716 9325 12750
rect 9291 12647 9325 12681
rect 9291 12578 9325 12612
rect 9291 12509 9325 12543
rect 9522 13887 9556 13921
rect 9617 13887 9651 13921
rect 9712 13887 9746 13921
rect 1396 11190 1430 11224
rect 1396 11117 1430 11151
rect 1396 11044 1430 11078
rect 1396 10971 1430 11005
rect 1396 10898 1430 10932
rect 1396 10825 1430 10859
rect 1396 10752 1430 10786
rect 1396 10678 1430 10712
rect 1396 10604 1430 10638
rect 1396 10530 1430 10564
rect 1396 10456 1430 10490
rect 3506 11190 3540 11224
rect 3506 11117 3540 11151
rect 3506 11044 3540 11078
rect 3506 10971 3540 11005
rect 3506 10898 3540 10932
rect 3506 10825 3540 10859
rect 3506 10752 3540 10786
rect 3506 10678 3540 10712
rect 3506 10604 3540 10638
rect 3506 10530 3540 10564
rect 3506 10456 3540 10490
rect 1396 10104 1430 10138
rect 1396 10031 1430 10065
rect 1396 9958 1430 9992
rect 1396 9885 1430 9919
rect 1396 9812 1430 9846
rect 1396 9739 1430 9773
rect 1396 9666 1430 9700
rect 1396 9592 1430 9626
rect 1396 9518 1430 9552
rect 1396 9444 1430 9478
rect 1396 9370 1430 9404
rect 3506 10104 3540 10138
rect 3506 10031 3540 10065
rect 3506 9958 3540 9992
rect 3506 9885 3540 9919
rect 3506 9812 3540 9846
rect 3506 9739 3540 9773
rect 3506 9666 3540 9700
rect 3506 9592 3540 9626
rect 3506 9518 3540 9552
rect 3506 9444 3540 9478
rect 3506 9370 3540 9404
rect 1396 9248 1430 9282
rect 1396 9175 1430 9209
rect 1396 9102 1430 9136
rect 1396 9029 1430 9063
rect 1396 8956 1430 8990
rect 1396 8883 1430 8917
rect 1396 8810 1430 8844
rect 1396 8736 1430 8770
rect 1396 8662 1430 8696
rect 1396 8588 1430 8622
rect 1396 8514 1430 8548
rect 3506 9248 3540 9282
rect 3506 9175 3540 9209
rect 3506 9102 3540 9136
rect 3506 9029 3540 9063
rect 3506 8956 3540 8990
rect 3506 8883 3540 8917
rect 3506 8810 3540 8844
rect 3506 8736 3540 8770
rect 3506 8662 3540 8696
rect 3506 8588 3540 8622
rect 3506 8514 3540 8548
rect 1396 8188 1430 8222
rect 1396 8119 1430 8153
rect 1396 8050 1430 8084
rect 1396 7981 1430 8015
rect 1396 7912 1430 7946
rect 1396 7843 1430 7877
rect 1396 7774 1430 7808
rect 1396 7705 1430 7739
rect 1396 7636 1430 7670
rect 1396 7567 1430 7601
rect 1396 7498 1430 7532
rect 1396 7428 1430 7462
rect 3506 8188 3540 8222
rect 3506 8119 3540 8153
rect 3506 8050 3540 8084
rect 3506 7981 3540 8015
rect 3506 7912 3540 7946
rect 3506 7843 3540 7877
rect 3506 7774 3540 7808
rect 3506 7705 3540 7739
rect 3506 7636 3540 7670
rect 3506 7567 3540 7601
rect 3506 7498 3540 7532
rect 3506 7428 3540 7462
rect 1396 6430 1430 6464
rect 1396 6357 1430 6391
rect 1396 6284 1430 6318
rect 1396 6211 1430 6245
rect 1396 6138 1430 6172
rect 1396 6065 1430 6099
rect 1396 5992 1430 6026
rect 1396 5918 1430 5952
rect 1396 5844 1430 5878
rect 1396 5770 1430 5804
rect 1396 5696 1430 5730
rect 3506 6430 3540 6464
rect 3506 6357 3540 6391
rect 3506 6284 3540 6318
rect 3506 6211 3540 6245
rect 3506 6138 3540 6172
rect 3506 6065 3540 6099
rect 3506 5992 3540 6026
rect 3506 5918 3540 5952
rect 3506 5844 3540 5878
rect 3506 5770 3540 5804
rect 3506 5696 3540 5730
rect 1396 5344 1430 5378
rect 1396 5271 1430 5305
rect 1396 5198 1430 5232
rect 1396 5125 1430 5159
rect 1396 5052 1430 5086
rect 1396 4979 1430 5013
rect 1396 4906 1430 4940
rect 1396 4832 1430 4866
rect 1396 4758 1430 4792
rect 1396 4684 1430 4718
rect 1396 4610 1430 4644
rect 3506 5344 3540 5378
rect 3506 5271 3540 5305
rect 3506 5198 3540 5232
rect 3506 5125 3540 5159
rect 3506 5052 3540 5086
rect 3506 4979 3540 5013
rect 3506 4906 3540 4940
rect 3506 4832 3540 4866
rect 3506 4758 3540 4792
rect 3506 4684 3540 4718
rect 3506 4610 3540 4644
rect 1396 4488 1430 4522
rect 1396 4415 1430 4449
rect 1396 4342 1430 4376
rect 1396 4269 1430 4303
rect 1396 4196 1430 4230
rect 1396 4123 1430 4157
rect 1396 4050 1430 4084
rect 1396 3976 1430 4010
rect 1396 3902 1430 3936
rect 1396 3828 1430 3862
rect 1396 3754 1430 3788
rect 3506 4488 3540 4522
rect 3506 4415 3540 4449
rect 3506 4342 3540 4376
rect 3506 4269 3540 4303
rect 3506 4196 3540 4230
rect 3506 4123 3540 4157
rect 3506 4050 3540 4084
rect 3506 3976 3540 4010
rect 3506 3902 3540 3936
rect 3506 3828 3540 3862
rect 3506 3754 3540 3788
rect 4082 11136 4116 11170
rect 5192 11136 5226 11170
rect 4082 10995 4116 11029
rect 4082 10922 4116 10956
rect 4082 10849 4116 10883
rect 4082 10776 4116 10810
rect 4082 10703 4116 10737
rect 4082 10630 4116 10664
rect 4082 10557 4116 10591
rect 4082 10483 4116 10517
rect 4082 10409 4116 10443
rect 4082 10335 4116 10369
rect 4082 10261 4116 10295
rect 5192 10995 5226 11029
rect 5192 10922 5226 10956
rect 5192 10849 5226 10883
rect 5192 10776 5226 10810
rect 5192 10703 5226 10737
rect 5192 10630 5226 10664
rect 5192 10557 5226 10591
rect 5192 10483 5226 10517
rect 5192 10409 5226 10443
rect 5192 10335 5226 10369
rect 5192 10261 5226 10295
rect 4082 10139 4116 10173
rect 4082 10066 4116 10100
rect 4082 9993 4116 10027
rect 4082 9920 4116 9954
rect 4082 9847 4116 9881
rect 4082 9774 4116 9808
rect 4082 9701 4116 9735
rect 4082 9627 4116 9661
rect 4082 9553 4116 9587
rect 4082 9479 4116 9513
rect 4082 9405 4116 9439
rect 5192 10139 5226 10173
rect 5192 10066 5226 10100
rect 5192 9993 5226 10027
rect 5192 9920 5226 9954
rect 5192 9847 5226 9881
rect 5192 9774 5226 9808
rect 5192 9701 5226 9735
rect 5192 9627 5226 9661
rect 5192 9553 5226 9587
rect 5192 9479 5226 9513
rect 5192 9405 5226 9439
rect 4082 9283 4116 9317
rect 4082 9210 4116 9244
rect 4082 9137 4116 9171
rect 4082 9064 4116 9098
rect 4082 8991 4116 9025
rect 4082 8918 4116 8952
rect 4082 8845 4116 8879
rect 4082 8771 4116 8805
rect 4082 8697 4116 8731
rect 4082 8623 4116 8657
rect 4082 8549 4116 8583
rect 5192 9283 5226 9317
rect 5192 9210 5226 9244
rect 5192 9137 5226 9171
rect 5192 9064 5226 9098
rect 5192 8991 5226 9025
rect 5192 8918 5226 8952
rect 5192 8845 5226 8879
rect 5192 8771 5226 8805
rect 5192 8697 5226 8731
rect 5192 8623 5226 8657
rect 5192 8549 5226 8583
rect 4082 8427 4116 8461
rect 4082 8354 4116 8388
rect 4082 8281 4116 8315
rect 4082 8208 4116 8242
rect 4082 8135 4116 8169
rect 4082 8062 4116 8096
rect 4082 7989 4116 8023
rect 4082 7915 4116 7949
rect 4082 7841 4116 7875
rect 4082 7767 4116 7801
rect 4082 7693 4116 7727
rect 5192 8427 5226 8461
rect 5192 8354 5226 8388
rect 5192 8281 5226 8315
rect 5192 8208 5226 8242
rect 5192 8135 5226 8169
rect 5192 8062 5226 8096
rect 5192 7989 5226 8023
rect 5192 7915 5226 7949
rect 5192 7841 5226 7875
rect 5192 7767 5226 7801
rect 5192 7693 5226 7727
rect 4082 7571 4116 7605
rect 4082 7498 4116 7532
rect 4082 7425 4116 7459
rect 4082 7352 4116 7386
rect 4082 7279 4116 7313
rect 4082 7206 4116 7240
rect 4082 7133 4116 7167
rect 4082 7059 4116 7093
rect 4082 6985 4116 7019
rect 4082 6911 4116 6945
rect 4082 6837 4116 6871
rect 5192 7571 5226 7605
rect 5192 7498 5226 7532
rect 5192 7425 5226 7459
rect 5192 7352 5226 7386
rect 5192 7279 5226 7313
rect 5192 7206 5226 7240
rect 5192 7133 5226 7167
rect 5192 7059 5226 7093
rect 5192 6985 5226 7019
rect 5192 6911 5226 6945
rect 5192 6837 5226 6871
rect 4082 6715 4116 6749
rect 4082 6642 4116 6676
rect 4082 6569 4116 6603
rect 4082 6496 4116 6530
rect 4082 6423 4116 6457
rect 4082 6350 4116 6384
rect 4082 6277 4116 6311
rect 4082 6203 4116 6237
rect 4082 6129 4116 6163
rect 4082 6055 4116 6089
rect 4082 5981 4116 6015
rect 5192 6715 5226 6749
rect 5192 6642 5226 6676
rect 5192 6569 5226 6603
rect 5192 6496 5226 6530
rect 5192 6423 5226 6457
rect 5192 6350 5226 6384
rect 5192 6277 5226 6311
rect 5192 6203 5226 6237
rect 5192 6129 5226 6163
rect 5192 6055 5226 6089
rect 5192 5981 5226 6015
rect 4082 5859 4116 5893
rect 4082 5786 4116 5820
rect 4082 5713 4116 5747
rect 4082 5640 4116 5674
rect 4082 5567 4116 5601
rect 4082 5494 4116 5528
rect 4082 5421 4116 5455
rect 4082 5347 4116 5381
rect 4082 5273 4116 5307
rect 4082 5199 4116 5233
rect 4082 5125 4116 5159
rect 5192 5859 5226 5893
rect 5192 5786 5226 5820
rect 5192 5713 5226 5747
rect 5192 5640 5226 5674
rect 5192 5567 5226 5601
rect 5192 5494 5226 5528
rect 5192 5421 5226 5455
rect 5192 5347 5226 5381
rect 5192 5273 5226 5307
rect 5192 5199 5226 5233
rect 5192 5125 5226 5159
rect 4082 5003 4116 5037
rect 4082 4930 4116 4964
rect 4082 4857 4116 4891
rect 4082 4784 4116 4818
rect 4082 4711 4116 4745
rect 4082 4638 4116 4672
rect 4082 4565 4116 4599
rect 4082 4491 4116 4525
rect 4082 4417 4116 4451
rect 4082 4343 4116 4377
rect 4082 4269 4116 4303
rect 5192 5003 5226 5037
rect 5192 4930 5226 4964
rect 5192 4857 5226 4891
rect 5192 4784 5226 4818
rect 5192 4711 5226 4745
rect 5192 4638 5226 4672
rect 5192 4565 5226 4599
rect 5192 4491 5226 4525
rect 5192 4417 5226 4451
rect 5192 4343 5226 4377
rect 5192 4269 5226 4303
rect 4082 4132 4116 4166
rect 5192 4132 5226 4166
rect 5922 11136 5956 11170
rect 7032 11136 7066 11170
rect 5922 10995 5956 11029
rect 5922 10922 5956 10956
rect 5922 10849 5956 10883
rect 5922 10776 5956 10810
rect 5922 10703 5956 10737
rect 5922 10630 5956 10664
rect 5922 10557 5956 10591
rect 5922 10483 5956 10517
rect 5922 10409 5956 10443
rect 5922 10335 5956 10369
rect 5922 10261 5956 10295
rect 7032 10995 7066 11029
rect 7032 10922 7066 10956
rect 7032 10849 7066 10883
rect 7032 10776 7066 10810
rect 7032 10703 7066 10737
rect 7032 10630 7066 10664
rect 7032 10557 7066 10591
rect 7032 10483 7066 10517
rect 7032 10409 7066 10443
rect 7032 10335 7066 10369
rect 7032 10261 7066 10295
rect 5922 10139 5956 10173
rect 5922 10066 5956 10100
rect 5922 9993 5956 10027
rect 5922 9920 5956 9954
rect 5922 9847 5956 9881
rect 5922 9774 5956 9808
rect 5922 9701 5956 9735
rect 5922 9627 5956 9661
rect 5922 9553 5956 9587
rect 5922 9479 5956 9513
rect 5922 9405 5956 9439
rect 7032 10139 7066 10173
rect 7032 10066 7066 10100
rect 7032 9993 7066 10027
rect 7032 9920 7066 9954
rect 7032 9847 7066 9881
rect 7032 9774 7066 9808
rect 7032 9701 7066 9735
rect 7032 9627 7066 9661
rect 7032 9553 7066 9587
rect 7032 9479 7066 9513
rect 7032 9405 7066 9439
rect 5922 9283 5956 9317
rect 5922 9210 5956 9244
rect 5922 9137 5956 9171
rect 5922 9064 5956 9098
rect 5922 8991 5956 9025
rect 5922 8918 5956 8952
rect 5922 8845 5956 8879
rect 5922 8771 5956 8805
rect 5922 8697 5956 8731
rect 5922 8623 5956 8657
rect 5922 8549 5956 8583
rect 7032 9283 7066 9317
rect 7032 9210 7066 9244
rect 7032 9137 7066 9171
rect 7032 9064 7066 9098
rect 7032 8991 7066 9025
rect 7032 8918 7066 8952
rect 7032 8845 7066 8879
rect 7032 8771 7066 8805
rect 7032 8697 7066 8731
rect 7032 8623 7066 8657
rect 7032 8549 7066 8583
rect 5922 8427 5956 8461
rect 5922 8354 5956 8388
rect 5922 8281 5956 8315
rect 5922 8208 5956 8242
rect 5922 8135 5956 8169
rect 5922 8062 5956 8096
rect 5922 7989 5956 8023
rect 5922 7915 5956 7949
rect 5922 7841 5956 7875
rect 5922 7767 5956 7801
rect 5922 7693 5956 7727
rect 7032 8427 7066 8461
rect 7032 8354 7066 8388
rect 7032 8281 7066 8315
rect 7032 8208 7066 8242
rect 7032 8135 7066 8169
rect 7032 8062 7066 8096
rect 7032 7989 7066 8023
rect 7032 7915 7066 7949
rect 7032 7841 7066 7875
rect 7032 7767 7066 7801
rect 7032 7693 7066 7727
rect 5922 7571 5956 7605
rect 5922 7498 5956 7532
rect 5922 7425 5956 7459
rect 5922 7352 5956 7386
rect 5922 7279 5956 7313
rect 5922 7206 5956 7240
rect 5922 7133 5956 7167
rect 5922 7059 5956 7093
rect 5922 6985 5956 7019
rect 5922 6911 5956 6945
rect 5922 6837 5956 6871
rect 7032 7571 7066 7605
rect 7032 7498 7066 7532
rect 7032 7425 7066 7459
rect 7032 7352 7066 7386
rect 7032 7279 7066 7313
rect 7032 7206 7066 7240
rect 7032 7133 7066 7167
rect 7032 7059 7066 7093
rect 7032 6985 7066 7019
rect 7032 6911 7066 6945
rect 7032 6837 7066 6871
rect 5922 6715 5956 6749
rect 5922 6642 5956 6676
rect 5922 6569 5956 6603
rect 5922 6496 5956 6530
rect 5922 6423 5956 6457
rect 5922 6350 5956 6384
rect 5922 6277 5956 6311
rect 5922 6203 5956 6237
rect 5922 6129 5956 6163
rect 5922 6055 5956 6089
rect 5922 5981 5956 6015
rect 7032 6715 7066 6749
rect 7032 6642 7066 6676
rect 7032 6569 7066 6603
rect 7032 6496 7066 6530
rect 7032 6423 7066 6457
rect 7032 6350 7066 6384
rect 7032 6277 7066 6311
rect 7032 6203 7066 6237
rect 7032 6129 7066 6163
rect 7032 6055 7066 6089
rect 7032 5981 7066 6015
rect 5922 5859 5956 5893
rect 5922 5786 5956 5820
rect 5922 5713 5956 5747
rect 5922 5640 5956 5674
rect 5922 5567 5956 5601
rect 5922 5494 5956 5528
rect 5922 5421 5956 5455
rect 5922 5347 5956 5381
rect 5922 5273 5956 5307
rect 5922 5199 5956 5233
rect 5922 5125 5956 5159
rect 7032 5859 7066 5893
rect 7032 5786 7066 5820
rect 7032 5713 7066 5747
rect 7032 5640 7066 5674
rect 7032 5567 7066 5601
rect 7032 5494 7066 5528
rect 7032 5421 7066 5455
rect 7032 5347 7066 5381
rect 7032 5273 7066 5307
rect 7032 5199 7066 5233
rect 7032 5125 7066 5159
rect 5922 5003 5956 5037
rect 5922 4930 5956 4964
rect 5922 4857 5956 4891
rect 5922 4784 5956 4818
rect 5922 4711 5956 4745
rect 5922 4638 5956 4672
rect 5922 4565 5956 4599
rect 5922 4491 5956 4525
rect 5922 4417 5956 4451
rect 5922 4343 5956 4377
rect 5922 4269 5956 4303
rect 7032 5003 7066 5037
rect 7032 4930 7066 4964
rect 7032 4857 7066 4891
rect 7032 4784 7066 4818
rect 7032 4711 7066 4745
rect 7032 4638 7066 4672
rect 7032 4565 7066 4599
rect 7032 4491 7066 4525
rect 7032 4417 7066 4451
rect 7032 4343 7066 4377
rect 7032 4269 7066 4303
rect 5922 4132 5956 4166
rect 7032 4132 7066 4166
rect 7608 11190 7642 11224
rect 7608 11117 7642 11151
rect 7608 11044 7642 11078
rect 7608 10971 7642 11005
rect 7608 10898 7642 10932
rect 7608 10825 7642 10859
rect 7608 10752 7642 10786
rect 7608 10678 7642 10712
rect 7608 10604 7642 10638
rect 7608 10530 7642 10564
rect 7608 10456 7642 10490
rect 9718 11190 9752 11224
rect 9718 11117 9752 11151
rect 9718 11044 9752 11078
rect 9718 10971 9752 11005
rect 9718 10898 9752 10932
rect 9718 10825 9752 10859
rect 9718 10752 9752 10786
rect 9718 10678 9752 10712
rect 9718 10604 9752 10638
rect 9718 10530 9752 10564
rect 9718 10456 9752 10490
rect 7608 10104 7642 10138
rect 7608 10031 7642 10065
rect 7608 9958 7642 9992
rect 7608 9885 7642 9919
rect 7608 9812 7642 9846
rect 7608 9739 7642 9773
rect 7608 9666 7642 9700
rect 7608 9592 7642 9626
rect 7608 9518 7642 9552
rect 7608 9444 7642 9478
rect 7608 9370 7642 9404
rect 9718 10104 9752 10138
rect 9718 10031 9752 10065
rect 9718 9958 9752 9992
rect 9718 9885 9752 9919
rect 9718 9812 9752 9846
rect 9718 9739 9752 9773
rect 9718 9666 9752 9700
rect 9718 9592 9752 9626
rect 9718 9518 9752 9552
rect 9718 9444 9752 9478
rect 9718 9370 9752 9404
rect 7608 9248 7642 9282
rect 7608 9175 7642 9209
rect 7608 9102 7642 9136
rect 7608 9029 7642 9063
rect 7608 8956 7642 8990
rect 7608 8883 7642 8917
rect 7608 8810 7642 8844
rect 7608 8736 7642 8770
rect 7608 8662 7642 8696
rect 7608 8588 7642 8622
rect 7608 8514 7642 8548
rect 9718 9248 9752 9282
rect 9718 9175 9752 9209
rect 9718 9102 9752 9136
rect 9718 9029 9752 9063
rect 9718 8956 9752 8990
rect 9718 8883 9752 8917
rect 9718 8810 9752 8844
rect 9718 8736 9752 8770
rect 9718 8662 9752 8696
rect 9718 8588 9752 8622
rect 9718 8514 9752 8548
rect 7608 8162 7642 8196
rect 7608 8089 7642 8123
rect 7608 8016 7642 8050
rect 7608 7943 7642 7977
rect 7608 7870 7642 7904
rect 7608 7797 7642 7831
rect 7608 7724 7642 7758
rect 7608 7650 7642 7684
rect 7608 7576 7642 7610
rect 7608 7502 7642 7536
rect 7608 7428 7642 7462
rect 9718 8162 9752 8196
rect 9718 8089 9752 8123
rect 9718 8016 9752 8050
rect 9718 7943 9752 7977
rect 9718 7870 9752 7904
rect 9718 7797 9752 7831
rect 9718 7724 9752 7758
rect 9718 7650 9752 7684
rect 9718 7576 9752 7610
rect 9718 7502 9752 7536
rect 9718 7428 9752 7462
rect 7608 6430 7642 6464
rect 7608 6361 7642 6395
rect 7608 6292 7642 6326
rect 7608 6223 7642 6257
rect 7608 6154 7642 6188
rect 7608 6085 7642 6119
rect 7608 6016 7642 6050
rect 7608 5947 7642 5981
rect 7608 5878 7642 5912
rect 7608 5809 7642 5843
rect 7608 5740 7642 5774
rect 7608 5670 7642 5704
rect 9718 6430 9752 6464
rect 9718 6361 9752 6395
rect 9718 6292 9752 6326
rect 9718 6223 9752 6257
rect 9718 6154 9752 6188
rect 9718 6085 9752 6119
rect 9718 6016 9752 6050
rect 9718 5947 9752 5981
rect 9718 5878 9752 5912
rect 9718 5809 9752 5843
rect 9718 5740 9752 5774
rect 9718 5670 9752 5704
rect 7608 5344 7642 5378
rect 7608 5271 7642 5305
rect 7608 5198 7642 5232
rect 7608 5125 7642 5159
rect 7608 5052 7642 5086
rect 7608 4979 7642 5013
rect 7608 4906 7642 4940
rect 7608 4832 7642 4866
rect 7608 4758 7642 4792
rect 7608 4684 7642 4718
rect 7608 4610 7642 4644
rect 9718 5344 9752 5378
rect 9718 5271 9752 5305
rect 9718 5198 9752 5232
rect 9718 5125 9752 5159
rect 9718 5052 9752 5086
rect 9718 4979 9752 5013
rect 9718 4906 9752 4940
rect 9718 4832 9752 4866
rect 9718 4758 9752 4792
rect 9718 4684 9752 4718
rect 9718 4610 9752 4644
rect 7608 4488 7642 4522
rect 7608 4415 7642 4449
rect 7608 4342 7642 4376
rect 7608 4269 7642 4303
rect 7608 4196 7642 4230
rect 7608 4123 7642 4157
rect 7608 4050 7642 4084
rect 7608 3976 7642 4010
rect 7608 3902 7642 3936
rect 7608 3828 7642 3862
rect 7608 3754 7642 3788
rect 9718 4488 9752 4522
rect 9718 4415 9752 4449
rect 9718 4342 9752 4376
rect 9718 4269 9752 4303
rect 9718 4196 9752 4230
rect 9718 4123 9752 4157
rect 9718 4050 9752 4084
rect 9718 3976 9752 4010
rect 9718 3902 9752 3936
rect 9718 3828 9752 3862
rect 9718 3754 9752 3788
rect 1396 3402 1430 3436
rect 1396 3329 1430 3363
rect 1396 3256 1430 3290
rect 1396 3183 1430 3217
rect 1396 3110 1430 3144
rect 1396 3037 1430 3071
rect 1396 2964 1430 2998
rect 1396 2890 1430 2924
rect 1396 2816 1430 2850
rect 1396 2742 1430 2776
rect 1396 2668 1430 2702
rect 3506 3402 3540 3436
rect 3506 3329 3540 3363
rect 3506 3256 3540 3290
rect 3506 3183 3540 3217
rect 3506 3110 3540 3144
rect 3506 3037 3540 3071
rect 3506 2964 3540 2998
rect 3506 2890 3540 2924
rect 3506 2816 3540 2850
rect 3506 2742 3540 2776
rect 3506 2668 3540 2702
rect 5194 3277 5228 3311
rect 5194 3209 5228 3243
rect 5194 3141 5228 3175
rect 7032 3277 7066 3311
rect 7032 3209 7066 3243
rect 7032 3141 7066 3175
rect 5194 2986 5228 3020
rect 5194 2918 5228 2952
rect 5194 2730 5228 2764
rect 5194 2662 5228 2696
rect 5712 3014 5746 3048
rect 5712 2946 5746 2980
rect 7032 2986 7066 3020
rect 7032 2918 7066 2952
rect 5194 2474 5228 2508
rect 5194 2406 5228 2440
rect 7032 2730 7066 2764
rect 7032 2662 7066 2696
rect 7032 2474 7066 2508
rect 7032 2406 7066 2440
rect 5194 2218 5228 2252
rect 5194 2150 5228 2184
rect 7032 2218 7066 2252
rect 7032 2150 7066 2184
rect 7608 3402 7642 3436
rect 7608 3329 7642 3363
rect 7608 3256 7642 3290
rect 7608 3183 7642 3217
rect 7608 3110 7642 3144
rect 7608 3037 7642 3071
rect 7608 2964 7642 2998
rect 7608 2890 7642 2924
rect 7608 2816 7642 2850
rect 7608 2742 7642 2776
rect 7608 2668 7642 2702
rect 9718 3402 9752 3436
rect 9718 3329 9752 3363
rect 9718 3256 9752 3290
rect 9718 3183 9752 3217
rect 9718 3110 9752 3144
rect 9718 3037 9752 3071
rect 9718 2964 9752 2998
rect 9718 2890 9752 2924
rect 9718 2816 9752 2850
rect 9718 2742 9752 2776
rect 9718 2668 9752 2702
rect 5194 1962 5228 1996
rect 5194 1894 5228 1928
rect 7032 1962 7066 1996
rect 7032 1894 7066 1928
rect 1396 1709 1430 1743
rect 1396 1636 1430 1670
rect 1396 1563 1430 1597
rect 1396 1490 1430 1524
rect 1396 1417 1430 1451
rect 1396 1344 1430 1378
rect 1396 1271 1430 1305
rect 1396 1197 1430 1231
rect 1396 1123 1430 1157
rect 1396 1049 1430 1083
rect 1396 975 1430 1009
rect 3506 1709 3540 1743
rect 3506 1636 3540 1670
rect 3506 1563 3540 1597
rect 3506 1490 3540 1524
rect 3506 1417 3540 1451
rect 3506 1344 3540 1378
rect 3506 1271 3540 1305
rect 3506 1197 3540 1231
rect 3506 1123 3540 1157
rect 3506 1049 3540 1083
rect 3506 975 3540 1009
rect 5194 1706 5228 1740
rect 5194 1638 5228 1672
rect 7032 1706 7066 1740
rect 7032 1638 7066 1672
rect 5194 1450 5228 1484
rect 5194 1382 5228 1416
rect 7032 1450 7066 1484
rect 7032 1382 7066 1416
rect 5194 1194 5228 1228
rect 5194 1126 5228 1160
rect 7032 1194 7066 1228
rect 7032 1126 7066 1160
rect 5194 971 5228 1005
rect 5194 903 5228 937
rect 1599 792 1633 826
rect 1733 792 1767 826
rect 1908 766 1942 800
rect 1976 766 2010 800
rect 2154 766 2188 800
rect 2222 766 2256 800
rect 2410 766 2444 800
rect 2478 766 2512 800
rect 2666 766 2700 800
rect 2734 766 2768 800
rect 2922 766 2956 800
rect 2990 766 3024 800
rect 3178 766 3212 800
rect 3246 766 3280 800
rect 3424 766 3458 800
rect 3492 766 3526 800
rect 7032 971 7066 1005
rect 7032 903 7066 937
rect 7608 1709 7642 1743
rect 7608 1636 7642 1670
rect 7608 1563 7642 1597
rect 7608 1490 7642 1524
rect 7608 1417 7642 1451
rect 7608 1344 7642 1378
rect 7608 1271 7642 1305
rect 7608 1197 7642 1231
rect 7608 1123 7642 1157
rect 7608 1049 7642 1083
rect 7608 975 7642 1009
rect 9718 1709 9752 1743
rect 9718 1636 9752 1670
rect 9718 1563 9752 1597
rect 9718 1490 9752 1524
rect 9718 1417 9752 1451
rect 9718 1344 9752 1378
rect 9718 1271 9752 1305
rect 9718 1197 9752 1231
rect 9718 1123 9752 1157
rect 9718 1049 9752 1083
rect 9718 975 9752 1009
rect 5192 678 5226 712
rect 5192 610 5226 644
rect 5192 542 5226 576
rect 7032 678 7066 712
rect 7032 610 7066 644
rect 7032 542 7066 576
rect 7622 766 7656 800
rect 7690 766 7724 800
rect 7868 766 7902 800
rect 7936 766 7970 800
rect 8124 766 8158 800
rect 8192 766 8226 800
rect 8380 766 8414 800
rect 8448 766 8482 800
rect 8636 766 8670 800
rect 8704 766 8738 800
rect 8892 766 8926 800
rect 8960 766 8994 800
rect 9138 766 9172 800
rect 9206 766 9240 800
<< locali >>
rect 1197 14200 1231 14234
rect 1269 14200 1299 14234
rect 1342 14200 1367 14234
rect 1415 14200 1435 14234
rect 1488 14200 1503 14234
rect 1561 14200 1571 14234
rect 1634 14200 1639 14234
rect 1741 14200 1746 14234
rect 1809 14200 1819 14234
rect 1877 14200 1892 14234
rect 1945 14200 1965 14234
rect 2013 14200 2038 14234
rect 2081 14200 2111 14234
rect 2149 14200 2183 14234
rect 2217 14200 2251 14234
rect 2289 14200 2319 14234
rect 2361 14200 2387 14234
rect 2433 14200 2455 14234
rect 2505 14200 2523 14234
rect 2577 14200 2591 14234
rect 2649 14200 2659 14234
rect 2721 14200 2727 14234
rect 2793 14200 2795 14234
rect 2829 14200 2831 14234
rect 2897 14200 2903 14234
rect 2965 14200 2975 14234
rect 3033 14200 3047 14234
rect 3101 14200 3119 14234
rect 3169 14200 3191 14234
rect 3237 14200 3263 14234
rect 3305 14200 3335 14234
rect 3373 14200 3407 14234
rect 3441 14200 3475 14234
rect 3513 14200 3543 14234
rect 3585 14200 3611 14234
rect 3657 14200 3679 14234
rect 3729 14200 3747 14234
rect 3801 14200 3815 14234
rect 3873 14200 3883 14234
rect 3945 14200 3951 14234
rect 4017 14200 4019 14234
rect 4053 14200 4055 14234
rect 4121 14200 4127 14234
rect 4189 14200 4199 14234
rect 4257 14200 4271 14234
rect 4325 14200 4343 14234
rect 4393 14200 4415 14234
rect 4461 14200 4487 14234
rect 4529 14200 4559 14234
rect 4597 14200 4631 14234
rect 4665 14200 4699 14234
rect 4737 14200 4767 14234
rect 4809 14200 4835 14234
rect 4881 14200 4903 14234
rect 4953 14200 4971 14234
rect 5025 14200 5039 14234
rect 5097 14200 5107 14234
rect 5169 14200 5175 14234
rect 5241 14200 5243 14234
rect 5277 14200 5279 14234
rect 5345 14200 5351 14234
rect 5413 14200 5423 14234
rect 5481 14200 5495 14234
rect 5549 14200 5567 14234
rect 5617 14200 5639 14234
rect 5685 14200 5711 14234
rect 5753 14200 5783 14234
rect 5821 14200 5855 14234
rect 5889 14200 5923 14234
rect 5961 14200 5991 14234
rect 6033 14200 6059 14234
rect 6105 14200 6127 14234
rect 6177 14200 6195 14234
rect 6249 14200 6263 14234
rect 6321 14200 6331 14234
rect 6393 14200 6399 14234
rect 6465 14200 6467 14234
rect 6501 14200 6503 14234
rect 6569 14200 6575 14234
rect 6637 14200 6647 14234
rect 6705 14200 6719 14234
rect 6773 14200 6791 14234
rect 6841 14200 6863 14234
rect 6909 14200 6935 14234
rect 6977 14200 7007 14234
rect 7045 14200 7079 14234
rect 7113 14200 7147 14234
rect 7185 14200 7215 14234
rect 7257 14200 7283 14234
rect 7329 14200 7351 14234
rect 7401 14200 7419 14234
rect 7473 14200 7487 14234
rect 7545 14200 7555 14234
rect 7617 14200 7623 14234
rect 7689 14200 7691 14234
rect 7725 14200 7727 14234
rect 7793 14200 7799 14234
rect 7861 14200 7871 14234
rect 7929 14200 7943 14234
rect 7997 14200 8015 14234
rect 8065 14200 8087 14234
rect 8133 14200 8159 14234
rect 8201 14200 8231 14234
rect 8269 14200 8303 14234
rect 8337 14200 8371 14234
rect 8409 14200 8439 14234
rect 8481 14200 8507 14234
rect 8553 14200 8575 14234
rect 8625 14200 8643 14234
rect 8697 14200 8711 14234
rect 8769 14200 8779 14234
rect 8841 14200 8847 14234
rect 8913 14200 8915 14234
rect 8949 14200 8951 14234
rect 9017 14200 9023 14234
rect 9085 14200 9095 14234
rect 9153 14200 9167 14234
rect 9221 14200 9239 14234
rect 9289 14200 9311 14234
rect 9357 14200 9383 14234
rect 9425 14200 9455 14234
rect 9493 14200 9527 14234
rect 9561 14200 9595 14234
rect 9633 14200 9663 14234
rect 9705 14200 9731 14234
rect 9777 14200 9799 14234
rect 9849 14200 9867 14234
rect 9921 14200 9935 14234
rect 9993 14200 10003 14234
rect 10065 14200 10071 14234
rect 10137 14200 10139 14234
rect 10173 14200 10175 14234
rect 10241 14200 10247 14234
rect 10309 14200 10319 14234
rect 10377 14200 10391 14234
rect 10445 14200 10463 14234
rect 10513 14200 10535 14234
rect 10581 14200 10607 14234
rect 10649 14200 10679 14234
rect 10717 14200 10751 14234
rect 10785 14200 10819 14234
rect 10857 14200 10887 14234
rect 10929 14200 10955 14234
rect 11001 14200 11111 14234
rect 1197 14166 1560 14200
rect 1197 14132 1371 14166
rect 1405 14132 1443 14166
rect 1477 14132 1515 14166
rect 1549 14132 1560 14166
rect 5173 14155 5921 14200
rect 1197 14124 1560 14132
rect 1231 14094 1560 14124
rect 2018 14098 2059 14132
rect 2093 14098 2134 14132
rect 2168 14098 2209 14132
rect 2243 14098 2284 14132
rect 2318 14098 2359 14132
rect 2393 14098 2434 14132
rect 2468 14098 2509 14132
rect 2543 14098 2584 14132
rect 2618 14098 2659 14132
rect 2693 14098 2734 14132
rect 2768 14098 2809 14132
rect 2843 14098 2884 14132
rect 2918 14098 2959 14132
rect 2993 14098 3033 14132
rect 5173 14121 5189 14155
rect 5223 14121 5265 14155
rect 5299 14121 5341 14155
rect 5375 14121 5417 14155
rect 5451 14121 5493 14155
rect 5527 14121 5569 14155
rect 5603 14121 5645 14155
rect 5679 14121 5721 14155
rect 5755 14121 5796 14155
rect 5830 14121 5871 14155
rect 5905 14121 5921 14155
rect 9365 14153 9903 14200
rect 1231 14066 1371 14094
rect 1197 14060 1371 14066
rect 1405 14060 1443 14094
rect 1477 14060 1515 14094
rect 1549 14060 1560 14094
rect 1197 14052 1560 14060
rect 1231 14021 1560 14052
rect 1231 13998 1371 14021
rect 1197 13987 1371 13998
rect 1405 13987 1443 14021
rect 1477 13987 1515 14021
rect 1549 13987 1560 14021
rect 1197 13980 1560 13987
rect 1231 13948 1560 13980
rect 1231 13930 1371 13948
rect 1197 13914 1371 13930
rect 1405 13914 1443 13948
rect 1477 13914 1515 13948
rect 1549 13914 1560 13948
rect 1197 13908 1560 13914
rect 1231 13875 1560 13908
rect 1231 13862 1371 13875
rect 1197 13841 1371 13862
rect 1405 13841 1443 13875
rect 1477 13841 1515 13875
rect 1549 13841 1560 13875
rect 1197 13836 1560 13841
rect 1231 13802 1560 13836
rect 1231 13794 1371 13802
rect 1197 13768 1371 13794
rect 1405 13768 1443 13802
rect 1477 13768 1515 13802
rect 1549 13768 1560 13802
rect 1197 13764 1560 13768
rect 1231 13729 1560 13764
rect 1231 13726 1371 13729
rect 1197 13695 1371 13726
rect 1405 13695 1443 13729
rect 1477 13695 1515 13729
rect 1549 13695 1560 13729
rect 1197 13692 1560 13695
rect 1231 13658 1560 13692
rect 1197 13656 1560 13658
rect 1197 13624 1371 13656
rect 1231 13622 1371 13624
rect 1405 13622 1443 13656
rect 1477 13622 1515 13656
rect 1549 13622 1560 13656
rect 1231 13586 1560 13622
rect 1197 13583 1560 13586
rect 1197 13556 1371 13583
rect 1231 13549 1371 13556
rect 1405 13549 1443 13583
rect 1477 13549 1515 13583
rect 1549 13549 1560 13583
rect 1231 13514 1560 13549
rect 1197 13510 1560 13514
rect 1197 13488 1371 13510
rect 1231 13476 1371 13488
rect 1405 13476 1443 13510
rect 1477 13476 1515 13510
rect 1549 13476 1560 13510
rect 1231 13442 1560 13476
rect 1197 13437 1560 13442
rect 1197 13420 1371 13437
rect 1231 13403 1371 13420
rect 1405 13403 1443 13437
rect 1477 13403 1515 13437
rect 1549 13403 1560 13437
rect 1231 13370 1560 13403
rect 1197 13364 1560 13370
rect 1197 13352 1371 13364
rect 1231 13330 1371 13352
rect 1405 13330 1443 13364
rect 1477 13330 1515 13364
rect 1549 13330 1560 13364
rect 1231 13298 1560 13330
rect 1197 13291 1560 13298
rect 1197 13284 1371 13291
rect 1231 13257 1371 13284
rect 1405 13257 1443 13291
rect 1477 13257 1515 13291
rect 1549 13257 1560 13291
rect 1231 13226 1560 13257
rect 1197 13218 1560 13226
rect 1197 13216 1371 13218
rect 1231 13184 1371 13216
rect 1405 13184 1443 13218
rect 1477 13184 1515 13218
rect 1549 13184 1560 13218
rect 1231 13168 1560 13184
rect 1791 14043 3287 14064
rect 5173 14083 5921 14121
rect 8049 14098 8089 14132
rect 8123 14098 8164 14132
rect 8198 14098 8239 14132
rect 8273 14098 8314 14132
rect 8348 14098 8389 14132
rect 8423 14098 8464 14132
rect 8498 14098 8539 14132
rect 8573 14098 8614 14132
rect 8648 14098 8689 14132
rect 8723 14098 8764 14132
rect 8798 14098 8839 14132
rect 8873 14098 8914 14132
rect 8948 14098 8989 14132
rect 9023 14098 9064 14132
rect 9365 14126 9399 14153
rect 9433 14126 9472 14153
rect 9506 14126 9545 14153
rect 9579 14126 9618 14153
rect 1757 14018 3321 14043
rect 1791 13973 3287 14018
rect 4245 14047 4389 14074
rect 4279 14040 4389 14047
rect 4572 14040 4610 14074
rect 4644 14040 4682 14074
rect 4865 14047 5009 14074
rect 4865 14040 4975 14047
rect 1757 13943 3321 13973
rect 1791 13903 3287 13943
rect 1757 13868 3321 13903
rect 1791 13833 3287 13868
rect 1757 13797 3321 13833
rect 1791 13759 3287 13797
rect 3407 13953 3551 13980
rect 3441 13946 3551 13953
rect 3734 13946 3772 13980
rect 3806 13946 3844 13980
rect 4027 13953 4171 13980
rect 4027 13946 4137 13953
rect 3407 13885 3441 13919
rect 3407 13824 3441 13851
rect 4137 13885 4171 13919
rect 4245 13979 4279 14013
rect 4245 13918 4279 13945
rect 4975 13979 5009 14013
rect 5173 14049 5189 14083
rect 5223 14049 5265 14083
rect 5299 14049 5341 14083
rect 5375 14049 5417 14083
rect 5451 14049 5493 14083
rect 5527 14049 5569 14083
rect 5603 14049 5645 14083
rect 5679 14049 5721 14083
rect 5755 14049 5796 14083
rect 5830 14049 5871 14083
rect 5905 14049 5921 14083
rect 5173 14011 5921 14049
rect 5173 13977 5189 14011
rect 5223 13977 5265 14011
rect 5299 13977 5341 14011
rect 5375 13977 5417 14011
rect 5451 13977 5493 14011
rect 5527 13977 5569 14011
rect 5603 13977 5645 14011
rect 5679 13977 5721 14011
rect 5755 13977 5796 14011
rect 5830 13977 5871 14011
rect 5905 13977 5921 14011
rect 6085 14047 6119 14063
rect 6252 14040 6292 14074
rect 7795 14043 9291 14064
rect 6085 14000 6119 14013
rect 7761 14018 9325 14043
rect 9365 14092 9380 14126
rect 9433 14119 9459 14126
rect 9506 14119 9538 14126
rect 9579 14119 9617 14126
rect 9652 14119 9691 14153
rect 9725 14126 9763 14153
rect 9797 14126 9835 14153
rect 9869 14126 9903 14153
rect 9730 14119 9763 14126
rect 9809 14119 9835 14126
rect 9414 14092 9459 14119
rect 9493 14092 9538 14119
rect 9572 14092 9617 14119
rect 9651 14092 9696 14119
rect 9730 14092 9775 14119
rect 9809 14092 9854 14119
rect 9888 14092 9903 14126
rect 9365 14085 9903 14092
rect 9365 14051 9399 14085
rect 9433 14051 9472 14085
rect 9506 14051 9545 14085
rect 9579 14051 9618 14085
rect 9652 14051 9691 14085
rect 9725 14051 9763 14085
rect 9797 14051 9835 14085
rect 9869 14051 9903 14085
rect 9365 14018 9903 14051
rect 11077 14132 11111 14162
rect 11077 14064 11111 14088
rect 5173 13966 5921 13977
rect 6063 13979 6103 14000
rect 6063 13966 6085 13979
rect 6137 13966 6957 14000
rect 4975 13918 5009 13945
rect 6085 13929 6119 13945
rect 6923 13953 6957 13966
rect 4245 13884 4389 13918
rect 4572 13884 4610 13918
rect 4644 13884 4682 13918
rect 4865 13884 5009 13918
rect 5318 13887 5342 13921
rect 5390 13887 5416 13921
rect 5462 13887 5490 13921
rect 5534 13887 5564 13921
rect 5606 13887 5638 13921
rect 5678 13887 5712 13921
rect 5749 13887 5786 13921
rect 5820 13887 5836 13921
rect 7250 13946 7288 13980
rect 7322 13946 7360 13980
rect 7795 13973 9291 14018
rect 7653 13953 7687 13969
rect 4137 13824 4171 13851
rect 3407 13790 3551 13824
rect 3734 13790 3772 13824
rect 3806 13790 3844 13824
rect 4027 13790 4171 13824
rect 4245 13834 4279 13850
rect 4975 13834 5009 13850
rect 1757 13727 3321 13759
rect 1791 13684 3287 13727
rect 1757 13657 3321 13684
rect 1791 13609 3287 13657
rect 1757 13587 3321 13609
rect 3407 13740 3441 13756
rect 4137 13740 4171 13756
rect 3407 13696 3441 13706
rect 4131 13696 4171 13706
rect 3407 13662 4171 13696
rect 3407 13652 3441 13662
rect 4131 13652 4171 13662
rect 4245 13746 4285 13800
rect 4975 13746 5009 13800
rect 4245 13662 4279 13712
rect 4975 13662 5009 13712
rect 4245 13628 4257 13662
rect 4291 13628 4329 13662
rect 4363 13628 4401 13662
rect 4865 13628 5009 13662
rect 5224 13753 5258 13795
rect 5224 13677 5258 13719
rect 3407 13602 3441 13618
rect 1791 13534 3287 13587
rect 3453 13534 3491 13568
rect 3525 13534 3563 13568
rect 1757 13517 3321 13534
rect 1791 13459 3287 13517
rect 1757 13447 3321 13459
rect 1791 13384 3287 13447
rect 1757 13377 3321 13384
rect 1791 13309 3287 13377
rect 3407 13484 3441 13500
rect 4137 13485 4171 13618
rect 5224 13602 5258 13643
rect 3407 13441 3441 13450
rect 4165 13484 4171 13485
rect 4131 13450 4137 13451
rect 4131 13441 4171 13450
rect 3407 13407 4171 13441
rect 3407 13396 3441 13407
rect 4131 13397 4171 13407
rect 4165 13396 4171 13397
rect 4245 13578 4279 13594
rect 4245 13490 4279 13544
rect 4245 13406 4279 13456
rect 4975 13578 5009 13594
rect 4975 13490 5009 13544
rect 4975 13406 5009 13456
rect 4245 13372 4323 13406
rect 4572 13372 4610 13406
rect 4644 13372 4682 13406
rect 4811 13372 5009 13406
rect 5224 13527 5258 13568
rect 5224 13452 5258 13493
rect 5224 13377 5258 13418
rect 3407 13346 3441 13362
rect 1757 13307 3321 13309
rect 1791 13273 3287 13307
rect 3734 13278 3772 13312
rect 3806 13278 3844 13312
rect 1757 13268 3321 13273
rect 1791 13203 3287 13268
rect 1757 13193 3321 13203
rect 1197 13124 1231 13154
rect 1197 13054 1231 13082
rect 1791 13133 3287 13193
rect 1757 13119 3321 13133
rect 1791 13063 3287 13119
rect 3407 13228 3441 13244
rect 4137 13228 4171 13362
rect 3407 13184 3441 13194
rect 4131 13184 4171 13194
rect 3407 13150 4171 13184
rect 3407 13140 3441 13150
rect 4131 13140 4171 13150
rect 4245 13322 4279 13338
rect 4245 13234 4279 13288
rect 4245 13150 4279 13200
rect 4975 13322 5009 13338
rect 4975 13234 5009 13288
rect 4975 13184 5009 13200
rect 5224 13302 5258 13343
rect 5224 13227 5258 13268
rect 5224 13152 5258 13193
rect 4245 13116 4323 13150
rect 4853 13115 4891 13149
rect 4925 13115 4963 13149
rect 3407 13090 3441 13106
rect 1757 13045 3321 13063
rect 1197 12984 1231 13009
rect 1197 12914 1231 12936
rect 1197 12844 1231 12863
rect 1197 12774 1231 12790
rect 1197 12704 1231 12717
rect 1197 12633 1231 12644
rect 1197 12562 1231 12571
rect 1357 12972 1391 13010
rect 1357 12900 1391 12938
rect 1357 12828 1391 12866
rect 1357 12755 1391 12794
rect 1357 12682 1391 12721
rect 1357 12609 1391 12648
rect 1357 12536 1391 12575
rect 1613 12972 1647 13010
rect 1613 12900 1647 12938
rect 1613 12828 1647 12866
rect 1613 12755 1647 12794
rect 1613 12682 1647 12721
rect 1613 12609 1647 12648
rect 1613 12536 1647 12575
rect 1791 12993 3287 13045
rect 3453 13022 3491 13056
rect 3525 13022 3563 13056
rect 1757 12971 3321 12993
rect 1791 12923 3287 12971
rect 1757 12897 3321 12923
rect 1791 12854 3287 12897
rect 1757 12823 3321 12854
rect 3407 12972 3441 12988
rect 4137 12972 4171 13106
rect 3407 12928 3441 12938
rect 4131 12928 4171 12938
rect 3407 12894 4171 12928
rect 3407 12884 3441 12894
rect 4131 12884 4171 12894
rect 4245 13066 4279 13082
rect 4245 12978 4279 13032
rect 4245 12894 4279 12944
rect 4975 13065 5009 13081
rect 4975 12977 5009 13031
rect 4975 12894 5009 12943
rect 4245 12860 4323 12894
rect 4572 12860 4610 12894
rect 4644 12860 4682 12894
rect 4811 12860 5009 12894
rect 5224 13077 5258 13118
rect 5224 13002 5258 13043
rect 5224 12927 5258 12968
rect 3407 12834 3441 12850
rect 4137 12834 4171 12850
rect 1791 12785 3287 12823
rect 4245 12810 4279 12826
rect 4975 12810 5009 12826
rect 1757 12750 3321 12785
rect 1791 12715 3287 12750
rect 1757 12681 3321 12715
rect 1791 12641 3287 12681
rect 1757 12612 3321 12641
rect 1791 12567 3287 12612
rect 3407 12766 3551 12800
rect 3734 12766 3772 12800
rect 3806 12766 3844 12800
rect 4027 12766 4171 12800
rect 3407 12739 3441 12766
rect 3407 12671 3441 12705
rect 4137 12739 4171 12766
rect 4137 12671 4171 12705
rect 4245 12722 4285 12776
rect 5292 12791 5346 13887
rect 5380 13752 5414 13793
rect 5380 13677 5414 13718
rect 5380 13602 5414 13643
rect 5380 13527 5414 13568
rect 5380 13452 5414 13493
rect 5380 13377 5414 13418
rect 5380 13302 5414 13343
rect 5380 13227 5414 13268
rect 5380 13152 5414 13193
rect 5380 13077 5414 13118
rect 5380 13002 5414 13043
rect 5380 12927 5414 12968
rect 5448 12791 5502 13887
rect 5536 13753 5570 13795
rect 5536 13677 5570 13719
rect 5536 13602 5570 13643
rect 5536 13527 5570 13568
rect 5536 13452 5570 13493
rect 5536 13377 5570 13418
rect 5536 13302 5570 13343
rect 5536 13227 5570 13268
rect 5536 13152 5570 13193
rect 5536 13077 5570 13118
rect 5536 13002 5570 13043
rect 5536 12927 5570 12968
rect 5604 12791 5658 13887
rect 5692 13752 5726 13793
rect 5692 13677 5726 13718
rect 5692 13602 5726 13643
rect 5692 13527 5726 13568
rect 5692 13452 5726 13493
rect 5692 13377 5726 13418
rect 5692 13302 5726 13343
rect 5692 13227 5726 13268
rect 5692 13152 5726 13193
rect 5692 13077 5726 13118
rect 5692 13002 5726 13043
rect 5692 12927 5726 12968
rect 5760 12791 5814 13887
rect 6412 13884 6450 13918
rect 6484 13884 6522 13918
rect 6923 13912 6957 13919
rect 7653 13912 7687 13919
rect 6923 13885 7687 13912
rect 6957 13878 7653 13885
rect 6085 13834 6119 13850
rect 6815 13834 6849 13850
rect 6923 13835 6957 13851
rect 7653 13835 7687 13851
rect 7761 13943 9325 13973
rect 7795 13903 9291 13943
rect 7761 13868 9325 13903
rect 5848 13753 5882 13795
rect 5848 13677 5882 13719
rect 5848 13602 5882 13643
rect 6085 13746 6125 13800
rect 7795 13833 9291 13868
rect 6815 13746 6849 13800
rect 7250 13790 7288 13824
rect 7322 13790 7360 13824
rect 7761 13797 9325 13833
rect 7795 13759 9291 13797
rect 6085 13662 6119 13712
rect 6815 13662 6849 13712
rect 6085 13628 6097 13662
rect 6131 13628 6169 13662
rect 6203 13628 6241 13662
rect 6705 13628 6849 13662
rect 6923 13740 6957 13756
rect 7653 13740 7687 13756
rect 6923 13696 6963 13706
rect 7653 13696 7687 13706
rect 6923 13662 7687 13696
rect 6923 13652 6963 13662
rect 7653 13652 7687 13662
rect 5848 13527 5882 13568
rect 5848 13452 5882 13493
rect 5848 13377 5882 13418
rect 6085 13578 6119 13594
rect 6085 13490 6119 13544
rect 6085 13406 6119 13456
rect 6815 13578 6849 13594
rect 6815 13490 6849 13544
rect 6815 13406 6849 13456
rect 6085 13372 6163 13406
rect 6412 13372 6450 13406
rect 6484 13372 6522 13406
rect 6651 13372 6849 13406
rect 6923 13485 6957 13618
rect 7653 13602 7687 13618
rect 7761 13727 9325 13759
rect 7795 13684 9291 13727
rect 7761 13657 9325 13684
rect 7795 13609 9291 13657
rect 7761 13587 9325 13609
rect 7531 13534 7569 13568
rect 7603 13534 7641 13568
rect 7795 13534 9291 13587
rect 7761 13517 9325 13534
rect 6923 13484 6929 13485
rect 6957 13450 6963 13451
rect 6923 13441 6963 13450
rect 7653 13484 7687 13500
rect 7653 13441 7687 13450
rect 6923 13407 7687 13441
rect 6923 13397 6963 13407
rect 6923 13396 6929 13397
rect 5848 13302 5882 13343
rect 7653 13396 7687 13407
rect 5848 13227 5882 13268
rect 5848 13152 5882 13193
rect 5848 13077 5882 13118
rect 6085 13322 6119 13338
rect 6085 13234 6119 13288
rect 6085 13150 6119 13200
rect 6815 13322 6849 13338
rect 6815 13234 6849 13288
rect 6085 13116 6163 13150
rect 6815 13149 6849 13200
rect 6693 13115 6731 13149
rect 6765 13115 6803 13149
rect 6837 13115 6849 13149
rect 6923 13228 6957 13362
rect 7653 13346 7687 13362
rect 7795 13459 9291 13517
rect 7761 13447 9325 13459
rect 7795 13384 9291 13447
rect 7761 13377 9325 13384
rect 7250 13278 7288 13312
rect 7322 13278 7360 13312
rect 7795 13309 9291 13377
rect 7761 13307 9325 13309
rect 7795 13273 9291 13307
rect 7761 13268 9325 13273
rect 7653 13228 7687 13244
rect 6923 13184 6963 13194
rect 7653 13184 7687 13194
rect 6923 13150 7687 13184
rect 6923 13140 6963 13150
rect 7653 13140 7687 13150
rect 5848 13002 5882 13043
rect 5848 12927 5882 12968
rect 6085 13066 6119 13082
rect 6085 12978 6119 13032
rect 6085 12894 6119 12944
rect 6815 13065 6849 13081
rect 6815 12977 6849 13031
rect 6815 12894 6849 12943
rect 6085 12860 6163 12894
rect 6412 12860 6450 12894
rect 6484 12860 6522 12894
rect 6651 12860 6849 12894
rect 6923 12972 6957 13106
rect 7653 13090 7687 13106
rect 7795 13203 9291 13268
rect 7761 13193 9325 13203
rect 7795 13133 9291 13193
rect 7761 13119 9325 13133
rect 7795 13063 9291 13119
rect 7531 13022 7569 13056
rect 7603 13022 7641 13056
rect 7761 13045 9325 13063
rect 7795 12993 9291 13045
rect 7653 12972 7687 12988
rect 6923 12928 6963 12938
rect 7653 12928 7687 12938
rect 6923 12894 7687 12928
rect 6923 12884 6963 12894
rect 7653 12884 7687 12894
rect 6923 12834 6957 12850
rect 7653 12834 7687 12850
rect 7761 12971 9325 12993
rect 7795 12923 9291 12971
rect 7761 12897 9325 12923
rect 7795 12854 9291 12897
rect 6085 12810 6119 12826
rect 6815 12810 6849 12826
rect 4975 12722 5009 12776
rect 5257 12757 5273 12791
rect 5307 12757 5347 12791
rect 5381 12757 5421 12791
rect 5455 12757 5495 12791
rect 5529 12757 5568 12791
rect 5602 12757 5641 12791
rect 5675 12757 5714 12791
rect 5748 12757 5787 12791
rect 5821 12757 5837 12791
rect 6085 12722 6125 12776
rect 4245 12672 4279 12688
rect 4975 12672 5009 12688
rect 3441 12637 3551 12644
rect 3407 12610 3551 12637
rect 3734 12610 3772 12644
rect 3806 12610 3844 12644
rect 4027 12637 4137 12644
rect 5195 12668 5345 12692
rect 4027 12610 4171 12637
rect 1757 12543 3321 12567
rect 1791 12516 3287 12543
rect 1197 12491 1231 12498
rect 4245 12577 4279 12593
rect 4245 12509 4279 12543
rect 4481 12550 4515 12604
rect 5195 12634 5219 12668
rect 5253 12634 5287 12668
rect 5321 12634 5345 12668
rect 5740 12668 5890 12692
rect 7761 12823 9325 12854
rect 6815 12722 6849 12776
rect 6085 12672 6119 12688
rect 6815 12672 6849 12688
rect 6923 12766 7067 12800
rect 7250 12766 7288 12800
rect 7322 12766 7360 12800
rect 7543 12766 7687 12800
rect 6923 12739 6957 12766
rect 4975 12577 5009 12593
rect 1197 12420 1231 12425
rect 1406 12424 1422 12458
rect 1474 12424 1529 12458
rect 1586 12424 1602 12458
rect 2018 12448 2059 12482
rect 2093 12448 2134 12482
rect 2168 12448 2209 12482
rect 2243 12448 2284 12482
rect 2318 12448 2359 12482
rect 2393 12448 2434 12482
rect 2468 12448 2509 12482
rect 2543 12448 2584 12482
rect 2618 12448 2659 12482
rect 2693 12448 2734 12482
rect 2768 12448 2809 12482
rect 2843 12448 2884 12482
rect 2918 12448 2959 12482
rect 2993 12448 3033 12482
rect 4975 12509 5009 12543
rect 4279 12475 4389 12482
rect 4245 12448 4389 12475
rect 4642 12448 4682 12482
rect 4865 12475 4975 12482
rect 4865 12448 5009 12475
rect 5195 12569 5345 12634
rect 5195 12535 5219 12569
rect 5253 12535 5287 12569
rect 5321 12535 5345 12569
rect 5195 12469 5345 12535
rect 5457 12560 5491 12626
rect 5614 12560 5648 12626
rect 5740 12634 5764 12668
rect 5798 12634 5832 12668
rect 5866 12634 5890 12668
rect 6923 12671 6957 12705
rect 5740 12569 5890 12634
rect 5740 12535 5764 12569
rect 5798 12535 5832 12569
rect 5866 12535 5890 12569
rect 5195 12435 5219 12469
rect 5253 12435 5287 12469
rect 5321 12435 5345 12469
rect 5740 12469 5890 12535
rect 7653 12739 7687 12766
rect 7653 12671 7687 12705
rect 6957 12637 7067 12644
rect 6923 12610 7067 12637
rect 7250 12610 7288 12644
rect 7322 12610 7360 12644
rect 7543 12637 7653 12644
rect 7543 12610 7687 12637
rect 7795 12785 9291 12823
rect 7761 12750 9325 12785
rect 7795 12715 9291 12750
rect 9359 14012 9909 14018
rect 9359 13978 9397 14012
rect 9431 13978 9471 14012
rect 9529 13978 9544 14012
rect 9597 13978 9617 14012
rect 9665 13978 9690 14012
rect 9733 13978 9763 14012
rect 9801 13978 9835 14012
rect 9869 13980 9909 14012
rect 9359 13944 9365 13978
rect 9399 13972 9869 13978
rect 9399 13944 9405 13972
rect 9359 13910 9405 13944
rect 9863 13946 9869 13972
rect 9903 13946 9909 13980
rect 9359 13874 9365 13910
rect 9399 13874 9405 13910
rect 9506 13887 9522 13921
rect 9556 13887 9617 13921
rect 9651 13887 9712 13921
rect 9746 13887 9762 13921
rect 9863 13907 9909 13946
rect 9359 13842 9405 13874
rect 9359 13802 9365 13842
rect 9399 13802 9405 13842
rect 9863 13873 9869 13907
rect 9903 13873 9909 13907
rect 9863 13839 9909 13873
rect 9359 13774 9405 13802
rect 9359 13730 9365 13774
rect 9399 13730 9405 13774
rect 9359 13706 9405 13730
rect 9359 13658 9365 13706
rect 9399 13658 9405 13706
rect 9359 13638 9405 13658
rect 9359 13586 9365 13638
rect 9399 13586 9405 13638
rect 9359 13570 9405 13586
rect 9359 13513 9365 13570
rect 9399 13513 9405 13570
rect 9359 13502 9405 13513
rect 9359 13440 9365 13502
rect 9399 13440 9405 13502
rect 9359 13434 9405 13440
rect 9359 13367 9365 13434
rect 9399 13367 9405 13434
rect 9359 13366 9405 13367
rect 9359 13332 9365 13366
rect 9399 13332 9405 13366
rect 9359 13328 9405 13332
rect 9359 13264 9365 13328
rect 9399 13264 9405 13328
rect 9359 13255 9405 13264
rect 9359 13196 9365 13255
rect 9399 13196 9405 13255
rect 9359 13182 9405 13196
rect 9359 13128 9365 13182
rect 9399 13128 9405 13182
rect 9359 13109 9405 13128
rect 9359 13060 9365 13109
rect 9399 13060 9405 13109
rect 9359 13036 9405 13060
rect 9359 12992 9365 13036
rect 9399 12992 9405 13036
rect 9359 12963 9405 12992
rect 9359 12924 9365 12963
rect 9399 12924 9405 12963
rect 9359 12890 9405 12924
rect 9461 13754 9495 13793
rect 9461 13681 9495 13720
rect 9461 13608 9495 13647
rect 9461 13535 9495 13574
rect 9461 13461 9495 13501
rect 9461 13387 9495 13427
rect 9461 13313 9495 13353
rect 9461 13239 9495 13279
rect 9461 13165 9495 13205
rect 9461 13091 9495 13131
rect 9461 13017 9495 13057
rect 9461 12943 9495 12983
rect 9618 13754 9652 13793
rect 9618 13681 9652 13720
rect 9618 13608 9652 13647
rect 9618 13535 9652 13574
rect 9618 13461 9652 13501
rect 9618 13387 9652 13427
rect 9618 13313 9652 13353
rect 9618 13239 9652 13279
rect 9618 13165 9652 13205
rect 9618 13091 9652 13131
rect 9618 13017 9652 13057
rect 9618 12943 9652 12983
rect 9773 13754 9807 13793
rect 9773 13681 9807 13720
rect 9773 13608 9807 13647
rect 9773 13535 9807 13574
rect 9773 13461 9807 13501
rect 9773 13387 9807 13427
rect 9773 13313 9807 13353
rect 9773 13239 9807 13279
rect 9773 13165 9807 13205
rect 9773 13091 9807 13131
rect 9773 13017 9807 13057
rect 9773 12943 9807 12983
rect 9863 13800 9869 13839
rect 9903 13800 9909 13839
rect 9863 13771 9909 13800
rect 9863 13727 9869 13771
rect 9903 13727 9909 13771
rect 9863 13703 9909 13727
rect 9863 13654 9869 13703
rect 9903 13654 9909 13703
rect 9863 13635 9909 13654
rect 9863 13581 9869 13635
rect 9903 13581 9909 13635
rect 9863 13567 9909 13581
rect 9863 13508 9869 13567
rect 9903 13508 9909 13567
rect 9863 13499 9909 13508
rect 9863 13435 9869 13499
rect 9903 13435 9909 13499
rect 9863 13431 9909 13435
rect 9863 13397 9869 13431
rect 9903 13397 9909 13431
rect 9863 13396 9909 13397
rect 9863 13329 9869 13396
rect 9903 13329 9909 13396
rect 9863 13323 9909 13329
rect 9863 13261 9869 13323
rect 9903 13261 9909 13323
rect 9863 13250 9909 13261
rect 9863 13193 9869 13250
rect 9903 13193 9909 13250
rect 9863 13177 9909 13193
rect 9863 13125 9869 13177
rect 9903 13125 9909 13177
rect 9863 13105 9909 13125
rect 9863 13057 9869 13105
rect 9903 13057 9909 13105
rect 9863 13033 9909 13057
rect 9863 12989 9869 13033
rect 9903 12989 9909 13033
rect 9863 12961 9909 12989
rect 9863 12921 9869 12961
rect 9903 12921 9909 12961
rect 9359 12856 9365 12890
rect 9399 12856 9405 12890
rect 9359 12817 9405 12856
rect 9359 12783 9365 12817
rect 9399 12791 9405 12817
rect 9863 12889 9909 12921
rect 9863 12853 9869 12889
rect 9903 12853 9909 12889
rect 9863 12819 9909 12853
rect 9863 12791 9869 12819
rect 9399 12785 9529 12791
rect 9730 12785 9869 12791
rect 9903 12785 9909 12819
rect 9359 12751 9399 12783
rect 9433 12751 9467 12785
rect 9517 12751 9535 12785
rect 9569 12751 9603 12785
rect 9637 12751 9671 12785
rect 9705 12751 9739 12785
rect 9776 12751 9837 12785
rect 9871 12751 9909 12785
rect 9359 12745 9909 12751
rect 11077 13996 11111 14014
rect 11077 13928 11111 13940
rect 11077 13860 11111 13866
rect 11077 13752 11111 13758
rect 11077 13678 11111 13690
rect 11077 13604 11111 13622
rect 11077 13530 11111 13554
rect 11077 13456 11111 13486
rect 11077 13384 11111 13418
rect 11077 13316 11111 13348
rect 11077 13248 11111 13274
rect 11077 13160 11111 13200
rect 11077 13120 11111 13126
rect 11077 13050 11111 13052
rect 11077 13012 11111 13016
rect 11077 12938 11111 12946
rect 11077 12864 11111 12876
rect 11077 12790 11111 12806
rect 7761 12681 9325 12715
rect 7795 12641 9291 12681
rect 7761 12612 9325 12641
rect 6321 12550 6355 12604
rect 6815 12577 6849 12593
rect 6815 12509 6849 12543
rect 5195 12386 5345 12435
rect 5486 12424 5500 12458
rect 5536 12424 5570 12458
rect 5606 12424 5620 12458
rect 5740 12435 5764 12469
rect 5798 12435 5832 12469
rect 5866 12435 5890 12469
rect 6085 12448 6229 12482
rect 6482 12448 6522 12482
rect 6705 12475 6815 12482
rect 7795 12567 9291 12612
rect 7761 12543 9325 12567
rect 7795 12516 9291 12543
rect 9395 12709 9873 12745
rect 9395 12690 9453 12709
rect 9395 12656 9419 12690
rect 9487 12690 9783 12709
rect 9817 12690 9873 12709
rect 9453 12656 9487 12675
rect 9521 12656 9747 12690
rect 9781 12675 9783 12690
rect 9781 12656 9815 12675
rect 9849 12656 9873 12690
rect 9395 12631 9873 12656
rect 9395 12617 9453 12631
rect 9395 12583 9419 12617
rect 9487 12617 9783 12631
rect 9817 12617 9873 12631
rect 9453 12583 9487 12597
rect 9521 12583 9747 12617
rect 9781 12597 9783 12617
rect 9781 12583 9815 12597
rect 9849 12583 9873 12617
rect 9395 12553 9873 12583
rect 9395 12543 9453 12553
rect 9395 12509 9419 12543
rect 9487 12543 9783 12553
rect 9817 12543 9873 12553
rect 9453 12509 9487 12519
rect 9521 12509 9747 12543
rect 9781 12519 9783 12543
rect 9781 12509 9815 12519
rect 9849 12509 9873 12543
rect 6705 12448 6849 12475
rect 8049 12448 8089 12482
rect 8123 12448 8164 12482
rect 8198 12448 8239 12482
rect 8273 12448 8314 12482
rect 8348 12448 8389 12482
rect 8423 12448 8464 12482
rect 8498 12448 8539 12482
rect 8573 12448 8614 12482
rect 8648 12448 8689 12482
rect 8723 12448 8764 12482
rect 8798 12448 8839 12482
rect 8873 12448 8914 12482
rect 8948 12448 8989 12482
rect 9023 12448 9064 12482
rect 9395 12475 9873 12509
rect 9395 12469 9453 12475
rect 5740 12386 5890 12435
rect 9395 12435 9419 12469
rect 9487 12469 9783 12475
rect 9817 12469 9873 12475
rect 9453 12435 9487 12441
rect 9521 12435 9747 12469
rect 9781 12441 9783 12469
rect 9781 12435 9815 12441
rect 9849 12435 9873 12469
rect 9395 12386 9873 12435
rect 11077 12716 11111 12736
rect 11077 12642 11111 12666
rect 11077 12568 11111 12596
rect 11077 12494 11111 12526
rect 11077 12420 11111 12456
rect 1231 12352 1299 12386
rect 1333 12352 1367 12386
rect 1401 12352 1435 12386
rect 1469 12352 1503 12386
rect 1537 12352 1571 12386
rect 1605 12352 1639 12386
rect 1673 12352 1707 12386
rect 1741 12352 1775 12386
rect 1809 12352 1843 12386
rect 1877 12352 1911 12386
rect 1945 12352 1979 12386
rect 2013 12352 2047 12386
rect 2081 12352 2115 12386
rect 2149 12352 2183 12386
rect 2217 12352 2251 12386
rect 2285 12352 2319 12386
rect 2353 12352 2387 12386
rect 2421 12352 2455 12386
rect 2489 12352 2523 12386
rect 2557 12352 2591 12386
rect 2625 12352 2659 12386
rect 2693 12352 2727 12386
rect 2761 12352 2795 12386
rect 2829 12352 2863 12386
rect 2897 12352 2931 12386
rect 2965 12352 2999 12386
rect 3033 12352 3067 12386
rect 3101 12352 3135 12386
rect 3169 12352 3203 12386
rect 3237 12352 3271 12386
rect 3305 12352 3339 12386
rect 3373 12352 3407 12386
rect 3441 12352 3475 12386
rect 3509 12352 3543 12386
rect 3577 12352 3611 12386
rect 3646 12352 3679 12386
rect 3727 12352 3747 12386
rect 3808 12352 3815 12386
rect 3849 12352 3855 12386
rect 3917 12352 3936 12386
rect 3985 12352 4017 12386
rect 4053 12352 4087 12386
rect 4131 12352 4155 12386
rect 4189 12352 4223 12386
rect 4257 12352 4291 12386
rect 4325 12352 4359 12386
rect 4393 12352 4427 12386
rect 4461 12352 4495 12386
rect 4529 12352 4563 12386
rect 4597 12352 4631 12386
rect 4665 12352 4699 12386
rect 4733 12352 4767 12386
rect 4801 12352 4835 12386
rect 4869 12352 4903 12386
rect 4937 12352 4971 12386
rect 5005 12352 5039 12386
rect 5073 12381 5107 12386
rect 5141 12381 5175 12386
rect 5209 12381 5243 12386
rect 5073 12352 5087 12381
rect 5141 12352 5162 12381
rect 5209 12352 5237 12381
rect 5277 12352 5311 12386
rect 5345 12381 5379 12386
rect 5413 12381 5447 12386
rect 5481 12381 5515 12386
rect 5549 12381 5583 12386
rect 5617 12381 5651 12386
rect 5685 12381 5719 12386
rect 5346 12352 5379 12381
rect 5420 12352 5447 12381
rect 5494 12352 5515 12381
rect 5568 12352 5583 12381
rect 5642 12352 5651 12381
rect 5716 12352 5719 12381
rect 5753 12381 5787 12386
rect 5821 12381 5855 12386
rect 5889 12381 5923 12386
rect 5957 12381 5991 12386
rect 5753 12352 5756 12381
rect 5821 12352 5830 12381
rect 5889 12352 5904 12381
rect 5957 12352 5978 12381
rect 6025 12352 6059 12386
rect 6093 12352 6127 12386
rect 6161 12352 6195 12386
rect 6229 12352 6263 12386
rect 6297 12352 6331 12386
rect 6365 12352 6399 12386
rect 6433 12352 6467 12386
rect 6501 12352 6535 12386
rect 6569 12352 6603 12386
rect 6637 12352 6671 12386
rect 6705 12352 6739 12386
rect 6773 12352 6807 12386
rect 6841 12352 6875 12386
rect 6933 12352 6943 12386
rect 6977 12352 6978 12386
rect 7045 12352 7058 12386
rect 7113 12352 7138 12386
rect 7181 12352 7215 12386
rect 7252 12352 7283 12386
rect 7332 12352 7351 12386
rect 7412 12352 7419 12386
rect 7453 12352 7458 12386
rect 7521 12352 7555 12386
rect 7589 12352 7623 12386
rect 7657 12352 7691 12386
rect 7725 12352 7759 12386
rect 7793 12380 7827 12386
rect 7861 12380 7895 12386
rect 7929 12380 7963 12386
rect 7997 12380 8031 12386
rect 8065 12380 8099 12386
rect 8133 12380 8167 12386
rect 8201 12380 8235 12386
rect 7793 12352 7802 12380
rect 7861 12352 7874 12380
rect 7929 12352 7946 12380
rect 7997 12352 8018 12380
rect 8065 12352 8090 12380
rect 8133 12352 8162 12380
rect 8201 12352 8234 12380
rect 8269 12352 8303 12386
rect 8337 12380 8371 12386
rect 8405 12380 8439 12386
rect 8473 12380 8507 12386
rect 8541 12380 8575 12386
rect 8609 12380 8643 12386
rect 8677 12380 8711 12386
rect 8745 12380 8779 12386
rect 8813 12380 8847 12386
rect 8340 12352 8371 12380
rect 8412 12352 8439 12380
rect 8484 12352 8507 12380
rect 8556 12352 8575 12380
rect 8628 12352 8643 12380
rect 8700 12352 8711 12380
rect 8772 12352 8779 12380
rect 8844 12352 8847 12380
rect 8881 12380 8915 12386
rect 8949 12380 8983 12386
rect 9017 12380 9052 12386
rect 9086 12380 9121 12386
rect 9155 12380 9190 12386
rect 9224 12380 9259 12386
rect 9293 12380 9328 12386
rect 9362 12380 9397 12386
rect 9431 12380 9466 12386
rect 9500 12380 9535 12386
rect 9569 12380 9604 12386
rect 8881 12352 8882 12380
rect 8949 12352 8954 12380
rect 9017 12352 9026 12380
rect 9086 12352 9098 12380
rect 9155 12352 9170 12380
rect 9224 12352 9242 12380
rect 9293 12352 9314 12380
rect 9362 12352 9386 12380
rect 9431 12352 9458 12380
rect 9500 12352 9530 12380
rect 9569 12352 9602 12380
rect 9638 12352 9673 12386
rect 9707 12380 9742 12386
rect 9776 12380 9811 12386
rect 9845 12380 9880 12386
rect 9914 12380 9949 12386
rect 9983 12380 10018 12386
rect 9708 12352 9742 12380
rect 9781 12352 9811 12380
rect 9854 12352 9880 12380
rect 9927 12352 9949 12380
rect 10000 12352 10018 12380
rect 10052 12380 10087 12386
rect 10121 12380 10156 12386
rect 10190 12380 10225 12386
rect 10259 12380 10294 12386
rect 10052 12352 10065 12380
rect 10121 12352 10141 12380
rect 10190 12352 10217 12380
rect 10259 12352 10293 12380
rect 10328 12352 10363 12386
rect 10397 12380 10432 12386
rect 10466 12380 10501 12386
rect 10535 12380 10583 12386
rect 10617 12380 10659 12386
rect 10693 12380 10735 12386
rect 10769 12380 10811 12386
rect 10845 12380 10886 12386
rect 10920 12380 10961 12386
rect 10403 12352 10432 12380
rect 10480 12352 10501 12380
rect 10557 12352 10583 12380
rect 10634 12352 10659 12380
rect 10711 12352 10735 12380
rect 10788 12352 10811 12380
rect 10865 12352 10886 12380
rect 10942 12352 10961 12380
rect 10995 12352 11111 12386
rect 5121 12347 5162 12352
rect 5196 12347 5237 12352
rect 5271 12347 5312 12352
rect 5346 12347 5386 12352
rect 5420 12347 5460 12352
rect 5494 12347 5534 12352
rect 5568 12347 5608 12352
rect 5642 12347 5682 12352
rect 5716 12347 5756 12352
rect 5790 12347 5830 12352
rect 5864 12347 5904 12352
rect 5938 12347 5978 12352
rect 7836 12346 7874 12352
rect 7908 12346 7946 12352
rect 7980 12346 8018 12352
rect 8052 12346 8090 12352
rect 8124 12346 8162 12352
rect 8196 12346 8234 12352
rect 8268 12346 8306 12352
rect 8340 12346 8378 12352
rect 8412 12346 8450 12352
rect 8484 12346 8522 12352
rect 8556 12346 8594 12352
rect 8628 12346 8666 12352
rect 8700 12346 8738 12352
rect 8772 12346 8810 12352
rect 8844 12346 8882 12352
rect 8916 12346 8954 12352
rect 8988 12346 9026 12352
rect 9060 12346 9098 12352
rect 9132 12346 9170 12352
rect 9204 12346 9242 12352
rect 9276 12346 9314 12352
rect 9348 12346 9386 12352
rect 9420 12346 9458 12352
rect 9492 12346 9530 12352
rect 9564 12346 9602 12352
rect 9636 12346 9674 12352
rect 9708 12346 9747 12352
rect 9781 12346 9820 12352
rect 9854 12346 9893 12352
rect 9927 12346 9966 12352
rect 10000 12346 10065 12352
rect 10099 12346 10141 12352
rect 10175 12346 10217 12352
rect 10251 12346 10293 12352
rect 10327 12346 10369 12352
rect 10403 12346 10446 12352
rect 10480 12346 10523 12352
rect 10557 12346 10600 12352
rect 10634 12346 10677 12352
rect 10711 12346 10754 12352
rect 10788 12346 10831 12352
rect 10865 12346 10908 12352
rect 1685 12171 1743 12175
rect 1777 12171 1836 12175
rect 1870 12171 1929 12175
rect 2321 12171 2363 12175
rect 2397 12171 2439 12175
rect 2473 12171 2515 12175
rect 2549 12171 2592 12175
rect 2626 12171 2669 12175
rect 2703 12171 2746 12175
rect 2780 12171 2823 12175
rect 2857 12171 2900 12175
rect 2934 12171 2977 12175
rect 3011 12171 3054 12175
rect 3088 12171 3131 12175
rect 3165 12171 3208 12175
rect 3242 12171 3285 12175
rect 5111 12171 5154 12175
rect 5188 12171 5231 12175
rect 5265 12171 5308 12175
rect 5342 12171 5385 12175
rect 5419 12171 5463 12175
rect 5497 12171 5541 12175
rect 5575 12171 5619 12175
rect 5653 12171 5697 12175
rect 5731 12171 5775 12175
rect 5809 12171 5853 12175
rect 5887 12171 5931 12175
rect 6923 12171 6971 12175
rect 7005 12171 7053 12175
rect 7087 12171 7135 12175
rect 7169 12171 7218 12175
rect 7252 12171 7301 12175
rect 7335 12171 7384 12175
rect 7837 12171 7876 12175
rect 7910 12171 7949 12175
rect 7983 12171 8022 12175
rect 8056 12171 8095 12175
rect 8129 12171 8168 12175
rect 8202 12171 8241 12175
rect 8275 12171 8314 12175
rect 8348 12171 8387 12175
rect 8421 12171 8460 12175
rect 8494 12171 8533 12175
rect 8567 12171 8606 12175
rect 8640 12171 8680 12175
rect 8714 12171 8754 12175
rect 8788 12171 8828 12175
rect 9456 12171 9501 12175
rect 9535 12171 9580 12175
rect 9614 12171 9659 12175
rect 9693 12171 9739 12175
rect 9773 12171 9819 12175
rect 10041 12171 10082 12175
rect 10116 12171 10157 12175
rect 10191 12171 10233 12175
rect 10517 12171 10558 12175
rect 10592 12171 10633 12175
rect 10667 12171 10709 12175
rect 10743 12171 10785 12175
rect 10819 12171 10861 12175
rect 10895 12171 10937 12175
rect 10971 12171 11013 12175
rect 11047 12171 11089 12175
rect 1204 12137 1228 12171
rect 1262 12137 1297 12171
rect 1331 12137 1366 12171
rect 1400 12137 1435 12171
rect 1469 12137 1504 12171
rect 1538 12137 1573 12171
rect 1607 12137 1642 12171
rect 1685 12141 1711 12171
rect 1777 12141 1780 12171
rect 1676 12137 1711 12141
rect 1745 12137 1780 12141
rect 1814 12141 1836 12171
rect 1814 12137 1849 12141
rect 1883 12137 1918 12171
rect 1963 12141 1987 12171
rect 1952 12137 1987 12141
rect 2021 12137 2056 12171
rect 2090 12137 2125 12171
rect 2159 12137 2194 12171
rect 2228 12137 2263 12171
rect 2321 12141 2332 12171
rect 2397 12141 2401 12171
rect 2297 12137 2332 12141
rect 2366 12137 2401 12141
rect 2435 12141 2439 12171
rect 2504 12141 2515 12171
rect 2573 12141 2592 12171
rect 2642 12141 2669 12171
rect 2435 12137 2470 12141
rect 2504 12137 2539 12141
rect 2573 12137 2608 12141
rect 2642 12137 2677 12141
rect 2711 12137 2746 12171
rect 2780 12137 2815 12171
rect 2857 12141 2884 12171
rect 2934 12141 2953 12171
rect 3011 12141 3022 12171
rect 3088 12141 3091 12171
rect 2849 12137 2884 12141
rect 2918 12137 2953 12141
rect 2987 12137 3022 12141
rect 3056 12137 3091 12141
rect 3125 12141 3131 12171
rect 3194 12141 3208 12171
rect 3263 12141 3285 12171
rect 3125 12137 3160 12141
rect 3194 12137 3229 12141
rect 3263 12137 3298 12141
rect 3332 12137 3367 12171
rect 3401 12137 3436 12171
rect 3470 12137 3505 12171
rect 3539 12137 3574 12171
rect 3608 12137 3643 12171
rect 3677 12137 3712 12171
rect 3746 12137 3781 12171
rect 3815 12137 3850 12171
rect 3884 12137 3919 12171
rect 3953 12137 3988 12171
rect 11123 12141 11165 12175
rect 1204 12103 3988 12137
rect 11094 12103 11199 12141
rect 1204 12069 1228 12103
rect 1262 12069 1297 12103
rect 1331 12069 1366 12103
rect 1400 12069 1435 12103
rect 1469 12069 1504 12103
rect 1538 12069 1573 12103
rect 1607 12069 1642 12103
rect 1685 12069 1711 12103
rect 1777 12069 1780 12103
rect 1814 12069 1836 12103
rect 1883 12069 1918 12103
rect 1963 12069 1987 12103
rect 2021 12069 2056 12103
rect 2090 12069 2125 12103
rect 2159 12069 2194 12103
rect 2228 12069 2263 12103
rect 2321 12069 2332 12103
rect 2397 12069 2401 12103
rect 2435 12069 2439 12103
rect 2504 12069 2515 12103
rect 2573 12069 2592 12103
rect 2642 12069 2669 12103
rect 2711 12069 2746 12103
rect 2780 12069 2815 12103
rect 2857 12069 2884 12103
rect 2934 12069 2953 12103
rect 3011 12069 3022 12103
rect 3088 12069 3091 12103
rect 3125 12069 3131 12103
rect 3194 12069 3208 12103
rect 3263 12069 3285 12103
rect 3332 12069 3367 12103
rect 3401 12069 3436 12103
rect 3470 12069 3505 12103
rect 3539 12069 3574 12103
rect 3608 12069 3643 12103
rect 3677 12069 3712 12103
rect 3746 12069 3781 12103
rect 3815 12069 3850 12103
rect 3884 12069 3919 12103
rect 3953 12069 3988 12103
rect 11123 12069 11165 12103
rect 1204 12035 3988 12069
rect 1204 12001 1228 12035
rect 1262 12001 1297 12035
rect 1331 12001 1366 12035
rect 1400 12001 1435 12035
rect 1469 12001 1504 12035
rect 1538 12001 1573 12035
rect 1607 12001 1642 12035
rect 1676 12031 1711 12035
rect 1745 12031 1780 12035
rect 1685 12001 1711 12031
rect 1777 12001 1780 12031
rect 1814 12031 1849 12035
rect 1814 12001 1836 12031
rect 1883 12001 1918 12035
rect 1952 12031 1987 12035
rect 1963 12001 1987 12031
rect 2021 12001 2056 12035
rect 2090 12001 2125 12035
rect 2159 12001 2194 12035
rect 2228 12001 2263 12035
rect 2297 12031 2332 12035
rect 2366 12031 2401 12035
rect 2321 12001 2332 12031
rect 2397 12001 2401 12031
rect 2435 12031 2470 12035
rect 2504 12031 2539 12035
rect 2573 12031 2608 12035
rect 2642 12031 2677 12035
rect 2435 12001 2439 12031
rect 2504 12001 2515 12031
rect 2573 12001 2592 12031
rect 2642 12001 2669 12031
rect 2711 12001 2746 12035
rect 2780 12001 2815 12035
rect 2849 12031 2884 12035
rect 2918 12031 2953 12035
rect 2987 12031 3022 12035
rect 3056 12031 3091 12035
rect 2857 12001 2884 12031
rect 2934 12001 2953 12031
rect 3011 12001 3022 12031
rect 3088 12001 3091 12031
rect 3125 12031 3160 12035
rect 3194 12031 3229 12035
rect 3263 12031 3298 12035
rect 3125 12001 3131 12031
rect 3194 12001 3208 12031
rect 3263 12001 3285 12031
rect 3332 12001 3367 12035
rect 3401 12001 3436 12035
rect 3470 12001 3505 12035
rect 3539 12001 3574 12035
rect 3608 12001 3643 12035
rect 3677 12001 3712 12035
rect 3746 12001 3781 12035
rect 3815 12001 3850 12035
rect 3884 12001 3919 12035
rect 3953 12001 3988 12035
rect 11094 12031 11199 12069
rect 1685 11997 1743 12001
rect 1777 11997 1836 12001
rect 1870 11997 1929 12001
rect 2321 11997 2363 12001
rect 2397 11997 2439 12001
rect 2473 11997 2515 12001
rect 2549 11997 2592 12001
rect 2626 11997 2669 12001
rect 2703 11997 2746 12001
rect 2780 11997 2823 12001
rect 2857 11997 2900 12001
rect 2934 11997 2977 12001
rect 3011 11997 3054 12001
rect 3088 11997 3131 12001
rect 3165 11997 3208 12001
rect 3242 11997 3285 12001
rect 5111 11997 5154 12001
rect 5188 11997 5231 12001
rect 5265 11997 5308 12001
rect 5342 11997 5385 12001
rect 5419 11997 5463 12001
rect 5497 11997 5541 12001
rect 5575 11997 5619 12001
rect 5653 11997 5697 12001
rect 5731 11997 5775 12001
rect 5809 11997 5853 12001
rect 5887 11997 5931 12001
rect 6923 11997 6971 12001
rect 7005 11997 7053 12001
rect 7087 11997 7135 12001
rect 7169 11997 7218 12001
rect 7252 11997 7301 12001
rect 7335 11997 7384 12001
rect 7837 11997 7876 12001
rect 7910 11997 7949 12001
rect 7983 11997 8022 12001
rect 8056 11997 8095 12001
rect 8129 11997 8168 12001
rect 8202 11997 8241 12001
rect 8275 11997 8314 12001
rect 8348 11997 8387 12001
rect 8421 11997 8460 12001
rect 8494 11997 8533 12001
rect 8567 11997 8606 12001
rect 8640 11997 8680 12001
rect 8714 11997 8754 12001
rect 8788 11997 8828 12001
rect 9456 11997 9501 12001
rect 9535 11997 9580 12001
rect 9614 11997 9659 12001
rect 9693 11997 9739 12001
rect 9773 11997 9819 12001
rect 10041 11997 10082 12001
rect 10116 11997 10157 12001
rect 10191 11997 10233 12001
rect 10517 11997 10558 12001
rect 10592 11997 10633 12001
rect 10667 11997 10709 12001
rect 10743 11997 10785 12001
rect 10819 11997 10861 12001
rect 10895 11997 10937 12001
rect 10971 11997 11013 12001
rect 11047 11997 11089 12001
rect 11123 11997 11165 12031
rect 1117 11699 1185 11723
rect 1151 11689 1185 11699
rect 1321 11689 1355 11723
rect 1389 11689 1423 11723
rect 1457 11689 1491 11723
rect 1525 11689 1559 11723
rect 1593 11689 1627 11723
rect 1664 11689 1695 11723
rect 1747 11689 1763 11723
rect 1830 11689 1831 11723
rect 1865 11689 1879 11723
rect 1933 11689 1962 11723
rect 2001 11689 2035 11723
rect 2069 11689 2103 11723
rect 2137 11689 2171 11723
rect 2205 11689 2230 11723
rect 2273 11689 2302 11723
rect 2341 11689 2374 11723
rect 2409 11689 2443 11723
rect 2480 11689 2511 11723
rect 2552 11689 2579 11723
rect 2625 11689 2647 11723
rect 2698 11689 2715 11723
rect 2771 11689 2810 11723
rect 2875 11689 2883 11723
rect 2943 11689 2956 11723
rect 3011 11689 3029 11723
rect 3079 11689 3102 11723
rect 3147 11689 3175 11723
rect 3215 11689 3248 11723
rect 3283 11689 3317 11723
rect 3355 11689 3385 11723
rect 3419 11689 3453 11723
rect 3487 11689 3521 11723
rect 3555 11689 3577 11723
rect 3623 11689 3657 11723
rect 3691 11689 3693 11723
rect 3759 11689 3765 11723
rect 3827 11689 3843 11723
rect 3895 11689 3921 11723
rect 3963 11689 3997 11723
rect 4034 11689 4065 11723
rect 4113 11689 4133 11723
rect 4192 11689 4201 11723
rect 4235 11689 4269 11723
rect 4303 11689 4337 11723
rect 4371 11689 4405 11723
rect 4439 11689 4473 11723
rect 4533 11689 4541 11723
rect 4607 11689 4609 11723
rect 4643 11689 4647 11723
rect 4711 11689 4721 11723
rect 4779 11689 4813 11723
rect 4847 11689 4881 11723
rect 4915 11689 4949 11723
rect 4983 11689 5017 11723
rect 5051 11689 5061 11723
rect 5119 11689 5145 11723
rect 5187 11689 5221 11723
rect 5264 11689 5289 11723
rect 5349 11689 5357 11723
rect 5391 11689 5400 11723
rect 5459 11689 5485 11723
rect 5519 11689 5557 11723
rect 5591 11689 5629 11723
rect 5663 11689 5688 11723
rect 5737 11689 5756 11723
rect 5811 11689 5824 11723
rect 5885 11689 5892 11723
rect 5959 11689 5960 11723
rect 5994 11689 5999 11723
rect 6062 11689 6096 11723
rect 6130 11689 6164 11723
rect 6198 11689 6232 11723
rect 6266 11689 6300 11723
rect 6334 11689 6339 11723
rect 6402 11689 6413 11723
rect 6470 11689 6487 11723
rect 6538 11689 6561 11723
rect 6606 11689 6640 11723
rect 6674 11689 6708 11723
rect 6742 11689 6776 11723
rect 6810 11689 6844 11723
rect 6878 11689 6901 11723
rect 6946 11689 6976 11723
rect 7014 11689 7048 11723
rect 7085 11689 7116 11723
rect 7160 11689 7184 11723
rect 7235 11689 7252 11723
rect 7310 11689 7320 11723
rect 7385 11689 7388 11723
rect 7422 11689 7423 11723
rect 7490 11689 7524 11723
rect 7558 11689 7592 11723
rect 7626 11689 7660 11723
rect 7694 11689 7728 11723
rect 7762 11689 7796 11723
rect 7860 11689 7901 11723
rect 7957 11689 7976 11723
rect 8025 11689 8051 11723
rect 8093 11689 8126 11723
rect 8161 11689 8195 11723
rect 8235 11689 8263 11723
rect 8310 11689 8331 11723
rect 8386 11689 8399 11723
rect 8462 11689 8467 11723
rect 8501 11689 8504 11723
rect 8569 11689 8580 11723
rect 8637 11689 8656 11723
rect 8705 11689 8732 11723
rect 8773 11689 8807 11723
rect 8842 11689 8875 11723
rect 8918 11689 8943 11723
rect 8977 11689 9011 11723
rect 9045 11689 9079 11723
rect 9113 11689 9147 11723
rect 9181 11689 9215 11723
rect 9249 11689 9283 11723
rect 9317 11689 9347 11723
rect 9385 11689 9419 11723
rect 9461 11689 9487 11723
rect 9541 11689 9555 11723
rect 9621 11689 9623 11723
rect 9657 11689 9667 11723
rect 9725 11689 9747 11723
rect 9793 11689 9827 11723
rect 9861 11689 9895 11723
rect 9933 11689 9963 11723
rect 1151 11665 1219 11689
rect 1117 11655 1219 11665
rect 3693 11655 3751 11689
rect 3693 11650 3717 11655
rect 3727 11616 3751 11621
rect 3693 11587 3751 11616
rect 3693 11577 3717 11587
rect 3727 11543 3751 11553
rect 3693 11519 3751 11543
rect 3693 11504 3717 11519
rect 3727 11470 3751 11485
rect 3693 11451 3751 11470
rect 3693 11431 3717 11451
rect 1464 11395 2246 11421
rect 2280 11395 2319 11429
rect 2353 11395 2392 11429
rect 2426 11395 2465 11429
rect 2499 11395 2538 11429
rect 2572 11395 2611 11429
rect 1464 11357 2611 11395
rect 1464 11353 2246 11357
rect 2280 11323 2319 11357
rect 2353 11323 2392 11357
rect 2426 11323 2465 11357
rect 2499 11323 2538 11357
rect 2572 11323 2611 11357
rect 1219 11246 1287 11281
rect 2280 11251 2319 11285
rect 2353 11251 2392 11285
rect 2426 11251 2465 11285
rect 2499 11251 2538 11285
rect 2572 11251 2611 11285
rect 3221 11387 3468 11421
rect 3727 11397 3751 11417
rect 3221 11353 3446 11387
rect 3693 11383 3751 11397
rect 3693 11359 3717 11383
rect 5554 11655 5557 11689
rect 5591 11655 5594 11689
rect 5554 11651 5594 11655
rect 5554 11587 5557 11651
rect 5591 11587 5594 11651
rect 5554 11579 5594 11587
rect 5554 11519 5557 11579
rect 5591 11519 5594 11579
rect 5554 11507 5594 11519
rect 5554 11451 5557 11507
rect 5591 11451 5594 11507
rect 5554 11435 5594 11451
rect 5554 11383 5557 11435
rect 5591 11383 5594 11435
rect 5554 11363 5594 11383
rect 3727 11325 3751 11349
rect 3693 11315 3751 11325
rect 3693 11287 3717 11315
rect 3727 11253 3751 11281
rect 1219 11212 1253 11246
rect 3693 11247 3751 11253
rect 1219 11177 1287 11212
rect 1219 11143 1253 11177
rect 1219 11108 1287 11143
rect 1219 11074 1253 11108
rect 1219 11039 1287 11074
rect 1219 11005 1253 11039
rect 1219 10970 1287 11005
rect 1219 10936 1253 10970
rect 1219 10901 1287 10936
rect 1219 10867 1253 10901
rect 1219 10832 1287 10867
rect 1219 10798 1253 10832
rect 1219 10763 1287 10798
rect 1219 10729 1253 10763
rect 1219 10694 1287 10729
rect 1219 10660 1253 10694
rect 1219 10625 1287 10660
rect 1219 10591 1253 10625
rect 1219 10556 1287 10591
rect 1219 10522 1253 10556
rect 1219 10487 1287 10522
rect 1219 10453 1253 10487
rect 1219 10418 1287 10453
rect 1396 11228 1430 11240
rect 3506 11228 3540 11240
rect 1430 11190 3506 11217
rect 1396 11154 3540 11190
rect 1430 11117 3506 11154
rect 1396 11080 3540 11117
rect 1430 11044 3506 11080
rect 1396 11006 3540 11044
rect 1430 10971 3506 11006
rect 1396 10932 3540 10971
rect 1430 10898 3506 10932
rect 1396 10859 3540 10898
rect 1430 10824 3506 10859
rect 1396 10786 3540 10824
rect 1430 10750 3506 10786
rect 1396 10712 3540 10750
rect 1430 10676 3506 10712
rect 1396 10638 3540 10676
rect 1430 10602 3506 10638
rect 1396 10564 3540 10602
rect 1430 10527 3506 10564
rect 1396 10490 3540 10527
rect 1430 10463 3506 10490
rect 1396 10440 1430 10452
rect 3506 10440 3540 10452
rect 3693 11215 3717 11247
rect 3727 11181 3751 11213
rect 3693 11179 3751 11181
rect 3693 11145 3717 11179
rect 3693 11143 3751 11145
rect 3727 11111 3751 11143
rect 3693 11077 3717 11109
rect 3693 11071 3751 11077
rect 3727 11043 3751 11071
rect 3693 11009 3717 11037
rect 3693 10999 3751 11009
rect 3727 10975 3751 10999
rect 3693 10941 3717 10965
rect 3693 10927 3751 10941
rect 3727 10907 3751 10927
rect 3693 10873 3717 10893
rect 3693 10855 3751 10873
rect 3727 10839 3751 10855
rect 3693 10805 3717 10821
rect 3693 10783 3751 10805
rect 3727 10771 3751 10783
rect 3693 10737 3717 10749
rect 3693 10711 3751 10737
rect 3727 10703 3751 10711
rect 3693 10669 3717 10677
rect 3693 10639 3751 10669
rect 3727 10635 3751 10639
rect 3693 10601 3717 10605
rect 3693 10567 3751 10601
rect 3693 10499 3751 10533
rect 3693 10495 3717 10499
rect 3727 10461 3751 10465
rect 1219 10384 1253 10418
rect 3693 10431 3751 10461
rect 3693 10423 3717 10431
rect 1219 10349 1287 10384
rect 2280 10362 2319 10396
rect 2353 10362 2392 10396
rect 2426 10362 2465 10396
rect 2499 10362 2538 10396
rect 2572 10362 2611 10396
rect 1219 10315 1253 10349
rect 1219 10280 1287 10315
rect 1219 10246 1253 10280
rect 1219 10211 1287 10246
rect 1219 10177 1253 10211
rect 1219 10142 1287 10177
rect 1464 10324 2611 10327
rect 1464 10290 2246 10324
rect 2280 10290 2319 10324
rect 2353 10290 2392 10324
rect 2426 10290 2465 10324
rect 2499 10290 2538 10324
rect 2572 10290 2611 10324
rect 1464 10252 2611 10290
rect 1464 10218 2246 10252
rect 2280 10218 2319 10252
rect 2353 10218 2392 10252
rect 2426 10218 2465 10252
rect 2499 10218 2538 10252
rect 2572 10218 2611 10252
rect 3727 10389 3751 10397
rect 3693 10363 3751 10389
rect 3693 10351 3717 10363
rect 3221 10218 3446 10327
rect 1464 10165 3446 10218
rect 3727 10317 3751 10329
rect 3693 10295 3751 10317
rect 3693 10279 3717 10295
rect 3727 10245 3751 10261
rect 3693 10227 3751 10245
rect 3693 10207 3717 10227
rect 3727 10173 3751 10193
rect 3693 10159 3751 10173
rect 1219 10108 1253 10142
rect 1219 10073 1287 10108
rect 1219 10039 1253 10073
rect 1219 10004 1287 10039
rect 1219 9970 1253 10004
rect 1219 9935 1287 9970
rect 1219 9901 1253 9935
rect 1219 9866 1287 9901
rect 1219 9832 1253 9866
rect 1219 9797 1287 9832
rect 1219 9763 1253 9797
rect 1219 9728 1287 9763
rect 1219 9694 1253 9728
rect 1219 9659 1287 9694
rect 1219 9625 1253 9659
rect 1219 9590 1287 9625
rect 1219 9556 1253 9590
rect 1219 9521 1287 9556
rect 1219 9487 1253 9521
rect 1219 9452 1287 9487
rect 1219 9418 1253 9452
rect 1219 9383 1287 9418
rect 1219 9349 1253 9383
rect 1396 10142 1430 10154
rect 3506 10142 3540 10154
rect 1430 10104 3506 10131
rect 1396 10068 3540 10104
rect 1430 10031 3506 10068
rect 1396 9994 3540 10031
rect 1430 9958 3506 9994
rect 1396 9920 3540 9958
rect 1430 9885 3506 9920
rect 1396 9846 3540 9885
rect 1430 9812 3506 9846
rect 1396 9773 3540 9812
rect 1430 9738 3506 9773
rect 1396 9700 3540 9738
rect 1430 9664 3506 9700
rect 1396 9626 3540 9664
rect 1430 9590 3506 9626
rect 1396 9552 3540 9590
rect 1430 9516 3506 9552
rect 1396 9478 3540 9516
rect 1430 9441 3506 9478
rect 1396 9404 3540 9441
rect 1430 9377 3506 9404
rect 1396 9354 1430 9366
rect 3506 9354 3540 9366
rect 3693 10135 3717 10159
rect 3727 10101 3751 10125
rect 3693 10091 3751 10101
rect 3693 10063 3717 10091
rect 3727 10029 3751 10057
rect 3693 10023 3751 10029
rect 3693 9991 3717 10023
rect 3727 9957 3751 9989
rect 3693 9955 3751 9957
rect 3693 9921 3717 9955
rect 3693 9919 3751 9921
rect 3727 9887 3751 9919
rect 3693 9853 3717 9885
rect 3693 9847 3751 9853
rect 3727 9819 3751 9847
rect 3693 9785 3717 9813
rect 3693 9775 3751 9785
rect 3727 9751 3751 9775
rect 3693 9717 3717 9741
rect 3693 9703 3751 9717
rect 3727 9683 3751 9703
rect 3693 9649 3717 9669
rect 3693 9631 3751 9649
rect 3727 9615 3751 9631
rect 3693 9581 3717 9597
rect 3693 9559 3751 9581
rect 3727 9547 3751 9559
rect 3693 9513 3717 9525
rect 3693 9487 3751 9513
rect 3727 9479 3751 9487
rect 3693 9445 3717 9453
rect 3693 9415 3751 9445
rect 3727 9411 3751 9415
rect 3693 9377 3717 9381
rect 1219 9314 1287 9349
rect 3693 9343 3751 9377
rect 1219 9280 1253 9314
rect 2280 9309 2319 9343
rect 2353 9309 2392 9343
rect 2426 9309 2465 9343
rect 2499 9309 2538 9343
rect 2572 9309 2611 9343
rect 2645 9309 2683 9343
rect 2717 9309 2755 9343
rect 2789 9309 2827 9343
rect 2861 9309 2899 9343
rect 2933 9309 2971 9343
rect 3005 9309 3043 9343
rect 3077 9309 3115 9343
rect 3149 9309 3187 9343
rect 1219 9245 1287 9280
rect 1219 9211 1253 9245
rect 1219 9176 1287 9211
rect 1219 9142 1253 9176
rect 1219 9107 1287 9142
rect 1219 9073 1253 9107
rect 1219 9038 1287 9073
rect 1219 9004 1253 9038
rect 1219 8969 1287 9004
rect 1219 8935 1253 8969
rect 1219 8900 1287 8935
rect 1219 8866 1253 8900
rect 1219 8831 1287 8866
rect 1219 8797 1253 8831
rect 1219 8762 1287 8797
rect 1219 8728 1253 8762
rect 1219 8693 1287 8728
rect 1219 8659 1253 8693
rect 1219 8624 1287 8659
rect 1219 8590 1253 8624
rect 1219 8555 1287 8590
rect 1219 8521 1253 8555
rect 1219 8486 1287 8521
rect 1396 9286 1430 9298
rect 3506 9286 3540 9298
rect 1430 9248 3506 9275
rect 1396 9212 3540 9248
rect 1430 9175 3506 9212
rect 1396 9138 3540 9175
rect 1430 9102 3506 9138
rect 1396 9064 3540 9102
rect 1430 9029 3506 9064
rect 1396 8990 3540 9029
rect 1430 8956 3506 8990
rect 1396 8917 3540 8956
rect 1430 8882 3506 8917
rect 1396 8844 3540 8882
rect 1430 8808 3506 8844
rect 1396 8770 3540 8808
rect 1430 8734 3506 8770
rect 1396 8696 3540 8734
rect 1430 8660 3506 8696
rect 1396 8622 3540 8660
rect 1430 8585 3506 8622
rect 1396 8548 3540 8585
rect 1430 8521 3506 8548
rect 1396 8498 1430 8510
rect 3506 8498 3540 8510
rect 3693 9275 3751 9309
rect 3693 9271 3717 9275
rect 3727 9237 3751 9241
rect 3693 9207 3751 9237
rect 3693 9199 3717 9207
rect 3727 9165 3751 9173
rect 3693 9139 3751 9165
rect 3693 9127 3717 9139
rect 3727 9093 3751 9105
rect 3693 9071 3751 9093
rect 3693 9055 3717 9071
rect 3727 9021 3751 9037
rect 3693 9003 3751 9021
rect 3693 8983 3717 9003
rect 3727 8949 3751 8969
rect 3693 8935 3751 8949
rect 3693 8911 3717 8935
rect 3727 8877 3751 8901
rect 3693 8867 3751 8877
rect 3693 8839 3717 8867
rect 3727 8805 3751 8833
rect 3693 8799 3751 8805
rect 3693 8767 3717 8799
rect 3727 8733 3751 8765
rect 3693 8731 3751 8733
rect 3693 8697 3717 8731
rect 3693 8695 3751 8697
rect 3727 8663 3751 8695
rect 3693 8629 3717 8661
rect 3693 8623 3751 8629
rect 3727 8595 3751 8623
rect 3693 8561 3717 8589
rect 3693 8551 3751 8561
rect 3727 8527 3751 8551
rect 1219 8452 1253 8486
rect 3693 8493 3717 8517
rect 3693 8479 3751 8493
rect 3727 8459 3751 8479
rect 1219 8417 1287 8452
rect 2280 8423 2319 8457
rect 2353 8423 2392 8457
rect 2426 8423 2465 8457
rect 2499 8423 2538 8457
rect 2572 8423 2611 8457
rect 1219 8383 1253 8417
rect 1219 8348 1287 8383
rect 1219 8314 1253 8348
rect 1219 8279 1287 8314
rect 1464 8351 2246 8385
rect 2280 8351 2319 8385
rect 2353 8351 2392 8385
rect 2426 8351 2465 8385
rect 2499 8351 2538 8385
rect 2572 8351 2611 8385
rect 1464 8313 2611 8351
rect 1464 8279 2246 8313
rect 2280 8279 2319 8313
rect 2353 8279 2392 8313
rect 2426 8279 2465 8313
rect 2499 8279 2538 8313
rect 2572 8279 2611 8313
rect 3693 8425 3717 8445
rect 3693 8407 3751 8425
rect 3727 8391 3751 8407
rect 3221 8279 3446 8385
rect 3693 8357 3717 8373
rect 3693 8335 3751 8357
rect 3727 8323 3751 8335
rect 3693 8289 3717 8301
rect 1219 8245 1253 8279
rect 3693 8263 3751 8289
rect 3727 8255 3751 8263
rect 1219 8210 1287 8245
rect 1219 8176 1253 8210
rect 1219 8141 1287 8176
rect 1219 8107 1253 8141
rect 1219 8072 1287 8107
rect 1219 8038 1253 8072
rect 1219 8003 1287 8038
rect 1219 7969 1253 8003
rect 1219 7934 1287 7969
rect 1219 7900 1253 7934
rect 1219 7865 1287 7900
rect 1219 7831 1253 7865
rect 1219 7796 1287 7831
rect 1219 7762 1253 7796
rect 1219 7727 1287 7762
rect 1219 7693 1253 7727
rect 1219 7658 1287 7693
rect 1219 7624 1253 7658
rect 1219 7589 1287 7624
rect 1219 7555 1253 7589
rect 1219 7520 1287 7555
rect 1219 7486 1253 7520
rect 1219 7451 1287 7486
rect 1219 7417 1253 7451
rect 1219 7382 1287 7417
rect 1430 8188 3506 8189
rect 1396 8180 3540 8188
rect 1430 8119 3506 8180
rect 1396 8108 3540 8119
rect 1430 8050 3506 8108
rect 1396 8036 3540 8050
rect 1430 7981 3506 8036
rect 1396 7964 3540 7981
rect 1430 7912 3506 7964
rect 1396 7892 3540 7912
rect 1430 7843 3506 7892
rect 1396 7820 3540 7843
rect 1430 7774 3506 7820
rect 1396 7748 3540 7774
rect 1430 7705 3506 7748
rect 1396 7676 3540 7705
rect 1430 7636 3506 7676
rect 1396 7604 3540 7636
rect 1430 7567 3506 7604
rect 1396 7532 3540 7567
rect 1430 7497 3506 7532
rect 1396 7462 3540 7497
rect 1430 7435 3506 7462
rect 1396 7412 1430 7424
rect 3506 7412 3540 7424
rect 3693 8221 3717 8229
rect 3693 8191 3751 8221
rect 3727 8187 3751 8191
rect 3693 8153 3717 8157
rect 3693 8119 3751 8153
rect 3693 8051 3751 8085
rect 3693 8047 3717 8051
rect 3727 8013 3751 8017
rect 3693 7983 3751 8013
rect 3693 7975 3717 7983
rect 3727 7941 3751 7949
rect 3693 7915 3751 7941
rect 3693 7903 3717 7915
rect 3727 7869 3751 7881
rect 3693 7847 3751 7869
rect 3693 7831 3717 7847
rect 3727 7797 3751 7813
rect 3693 7779 3751 7797
rect 3693 7759 3717 7779
rect 3727 7725 3751 7745
rect 3693 7711 3751 7725
rect 3693 7687 3717 7711
rect 3727 7653 3751 7677
rect 3693 7643 3751 7653
rect 3693 7615 3717 7643
rect 3727 7581 3751 7609
rect 3693 7575 3751 7581
rect 3693 7543 3717 7575
rect 3727 7509 3751 7541
rect 3693 7507 3751 7509
rect 3693 7473 3717 7507
rect 3693 7471 3751 7473
rect 3727 7439 3751 7471
rect 3693 7405 3717 7437
rect 1219 7348 1253 7382
rect 2280 7367 2319 7401
rect 2353 7367 2392 7401
rect 2426 7367 2465 7401
rect 2499 7367 2538 7401
rect 2572 7367 2611 7401
rect 1219 7313 1287 7348
rect 1219 7279 1253 7313
rect 1219 7244 1287 7279
rect 1219 7210 1253 7244
rect 1464 7295 2246 7299
rect 2280 7295 2319 7329
rect 2353 7295 2392 7329
rect 2426 7295 2465 7329
rect 2499 7295 2538 7329
rect 2572 7295 2611 7329
rect 1464 7257 2611 7295
rect 1464 7231 2246 7257
rect 2280 7223 2319 7257
rect 2353 7223 2392 7257
rect 2426 7223 2465 7257
rect 2499 7223 2538 7257
rect 2572 7223 2611 7257
rect 3693 7399 3751 7405
rect 3727 7371 3751 7399
rect 3693 7337 3717 7365
rect 3693 7327 3751 7337
rect 3727 7303 3751 7327
rect 3221 7265 3446 7299
rect 3693 7269 3717 7293
rect 3221 7231 3468 7265
rect 3693 7255 3751 7269
rect 3727 7235 3751 7255
rect 1219 7175 1287 7210
rect 1219 7141 1253 7175
rect 1219 7106 1287 7141
rect 1219 7072 1253 7106
rect 1219 7037 1287 7072
rect 1219 7003 1253 7037
rect 1219 6963 1287 7003
rect 3693 7201 3717 7221
rect 3693 7183 3751 7201
rect 3727 7167 3751 7183
rect 3693 7133 3717 7149
rect 3693 7111 3751 7133
rect 3727 7099 3751 7111
rect 3693 7065 3717 7077
rect 3693 7039 3751 7065
rect 3727 7031 3751 7039
rect 3693 6997 3717 7005
rect 3693 6967 3751 6997
rect 3727 6963 3751 6967
rect 1287 6929 1321 6963
rect 1355 6929 1389 6963
rect 1423 6929 1457 6963
rect 1491 6929 1525 6963
rect 1559 6929 1593 6963
rect 1627 6929 1661 6963
rect 1695 6929 1729 6963
rect 1763 6929 1797 6963
rect 1831 6929 1865 6963
rect 1899 6929 1933 6963
rect 1967 6929 2001 6963
rect 2035 6929 2069 6963
rect 2103 6929 2137 6963
rect 2171 6929 2205 6963
rect 2239 6929 2273 6963
rect 2307 6929 2341 6963
rect 2375 6929 2409 6963
rect 2443 6929 2477 6963
rect 2511 6929 2545 6963
rect 2579 6929 2613 6963
rect 2647 6929 2681 6963
rect 2715 6929 2749 6963
rect 2783 6929 2817 6963
rect 2851 6929 2885 6963
rect 2919 6929 2953 6963
rect 2987 6929 3021 6963
rect 3055 6929 3089 6963
rect 3123 6929 3157 6963
rect 3191 6929 3225 6963
rect 3259 6929 3293 6963
rect 3327 6929 3361 6963
rect 3395 6929 3429 6963
rect 3463 6929 3497 6963
rect 3531 6929 3565 6963
rect 3599 6929 3633 6963
rect 3667 6933 3693 6963
rect 3667 6929 3717 6933
rect 3693 6895 3751 6929
rect 3693 6827 3751 6861
rect 3693 6823 3717 6827
rect 3727 6789 3751 6793
rect 3693 6759 3751 6789
rect 3693 6751 3717 6759
rect 3727 6717 3751 6725
rect 3693 6691 3751 6717
rect 3693 6679 3717 6691
rect 1464 6635 2022 6661
rect 2056 6635 2095 6669
rect 2129 6635 2168 6669
rect 2202 6635 2241 6669
rect 2275 6635 2314 6669
rect 2348 6635 2387 6669
rect 1464 6597 2387 6635
rect 1464 6593 2022 6597
rect 2056 6563 2095 6597
rect 2129 6563 2168 6597
rect 2202 6563 2241 6597
rect 2275 6563 2314 6597
rect 2348 6563 2387 6597
rect 2056 6491 2095 6525
rect 2129 6491 2168 6525
rect 2202 6491 2241 6525
rect 2275 6491 2314 6525
rect 2348 6491 2387 6525
rect 2997 6627 3468 6661
rect 3727 6645 3751 6657
rect 2997 6593 3446 6627
rect 3693 6623 3751 6645
rect 3693 6607 3717 6623
rect 3727 6573 3751 6589
rect 3693 6555 3751 6573
rect 3693 6535 3717 6555
rect 3727 6501 3751 6521
rect 3693 6487 3751 6501
rect 1396 6468 1430 6480
rect 3506 6468 3540 6480
rect 1430 6430 3506 6457
rect 1396 6394 3540 6430
rect 1430 6357 3506 6394
rect 1396 6320 3540 6357
rect 1430 6284 3506 6320
rect 1396 6246 3540 6284
rect 1430 6211 3506 6246
rect 1396 6172 3540 6211
rect 1430 6138 3506 6172
rect 1396 6099 3540 6138
rect 1430 6064 3506 6099
rect 1396 6026 3540 6064
rect 1430 5990 3506 6026
rect 1396 5952 3540 5990
rect 1430 5916 3506 5952
rect 1396 5878 3540 5916
rect 1430 5842 3506 5878
rect 1396 5804 3540 5842
rect 1430 5767 3506 5804
rect 1396 5730 3540 5767
rect 1430 5703 3506 5730
rect 1396 5680 1430 5692
rect 3506 5680 3540 5692
rect 3693 6463 3717 6487
rect 3727 6429 3751 6453
rect 3693 6419 3751 6429
rect 3693 6391 3717 6419
rect 3727 6357 3751 6385
rect 3693 6351 3751 6357
rect 3693 6319 3717 6351
rect 3727 6285 3751 6317
rect 3693 6283 3751 6285
rect 3693 6249 3717 6283
rect 3693 6247 3751 6249
rect 3727 6215 3751 6247
rect 3693 6181 3717 6213
rect 3693 6175 3751 6181
rect 3727 6147 3751 6175
rect 3693 6113 3717 6141
rect 3693 6103 3751 6113
rect 3727 6079 3751 6103
rect 3693 6045 3717 6069
rect 3693 6031 3751 6045
rect 3727 6011 3751 6031
rect 3693 5977 3717 5997
rect 3693 5959 3751 5977
rect 3727 5943 3751 5959
rect 3693 5909 3717 5925
rect 3693 5887 3751 5909
rect 3727 5875 3751 5887
rect 3693 5841 3717 5853
rect 3693 5815 3751 5841
rect 3727 5807 3751 5815
rect 3693 5773 3717 5781
rect 3693 5743 3751 5773
rect 3727 5739 3751 5743
rect 3693 5705 3717 5709
rect 3693 5671 3751 5705
rect 1464 5576 2022 5600
rect 2056 5576 2095 5610
rect 2129 5576 2168 5610
rect 2202 5576 2241 5610
rect 2275 5576 2314 5610
rect 2348 5576 2387 5610
rect 1464 5538 2387 5576
rect 1464 5504 2022 5538
rect 2056 5504 2095 5538
rect 2129 5504 2168 5538
rect 2202 5504 2241 5538
rect 2275 5504 2314 5538
rect 2348 5504 2387 5538
rect 1464 5466 2387 5504
rect 1464 5464 2022 5466
rect 2056 5432 2095 5466
rect 2129 5432 2168 5466
rect 2202 5432 2241 5466
rect 2275 5432 2314 5466
rect 2348 5432 2387 5466
rect 3693 5603 3751 5637
rect 2997 5464 3446 5600
rect 3693 5599 3717 5603
rect 3727 5565 3751 5569
rect 3693 5535 3751 5565
rect 3693 5527 3717 5535
rect 3727 5493 3751 5501
rect 3693 5467 3751 5493
rect 3693 5455 3717 5467
rect 3727 5421 3751 5433
rect 3693 5399 3751 5421
rect 1396 5382 1430 5394
rect 3506 5382 3540 5394
rect 1430 5344 3506 5371
rect 1396 5308 3540 5344
rect 1430 5271 3506 5308
rect 1396 5234 3540 5271
rect 1430 5198 3506 5234
rect 1396 5160 3540 5198
rect 1430 5125 3506 5160
rect 1396 5086 3540 5125
rect 1430 5052 3506 5086
rect 1396 5013 3540 5052
rect 1430 4978 3506 5013
rect 1396 4940 3540 4978
rect 1430 4904 3506 4940
rect 1396 4866 3540 4904
rect 1430 4830 3506 4866
rect 1396 4792 3540 4830
rect 1430 4756 3506 4792
rect 1396 4718 3540 4756
rect 1430 4681 3506 4718
rect 1396 4644 3540 4681
rect 1430 4617 3506 4644
rect 1396 4594 1430 4606
rect 3506 4594 3540 4606
rect 3693 5383 3717 5399
rect 3727 5349 3751 5365
rect 3693 5331 3751 5349
rect 3693 5311 3717 5331
rect 3727 5277 3751 5297
rect 3693 5263 3751 5277
rect 3693 5239 3717 5263
rect 3727 5205 3751 5229
rect 3693 5195 3751 5205
rect 3693 5167 3717 5195
rect 3727 5133 3751 5161
rect 3693 5127 3751 5133
rect 3693 5095 3717 5127
rect 3727 5061 3751 5093
rect 3693 5059 3751 5061
rect 3693 5025 3717 5059
rect 3693 5023 3751 5025
rect 3727 4991 3751 5023
rect 3693 4957 3717 4989
rect 3693 4951 3751 4957
rect 3727 4923 3751 4951
rect 3693 4889 3717 4917
rect 3693 4879 3751 4889
rect 3727 4855 3751 4879
rect 3693 4821 3717 4845
rect 3693 4807 3751 4821
rect 3727 4787 3751 4807
rect 3693 4753 3717 4773
rect 3693 4735 3751 4753
rect 3727 4719 3751 4735
rect 3693 4685 3717 4701
rect 3693 4663 3751 4685
rect 3727 4651 3751 4663
rect 3693 4617 3717 4629
rect 3693 4591 3751 4617
rect 3727 4583 3751 4591
rect 2056 4549 2095 4583
rect 2129 4549 2168 4583
rect 2202 4549 2241 4583
rect 2275 4549 2314 4583
rect 2348 4549 2387 4583
rect 2421 4549 2459 4583
rect 2493 4549 2531 4583
rect 2565 4549 2603 4583
rect 2637 4549 2675 4583
rect 2709 4549 2747 4583
rect 2781 4549 2819 4583
rect 2853 4549 2891 4583
rect 2925 4549 2963 4583
rect 3693 4549 3717 4557
rect 1117 3878 1185 3913
rect 1151 3844 1185 3878
rect 1117 3809 1185 3844
rect 1151 3775 1185 3809
rect 1117 3740 1185 3775
rect 1151 3706 1185 3740
rect 1396 4526 1430 4538
rect 3506 4526 3540 4538
rect 1430 4488 3506 4515
rect 1396 4452 3540 4488
rect 1430 4415 3506 4452
rect 1396 4378 3540 4415
rect 1430 4342 3506 4378
rect 1396 4304 3540 4342
rect 1430 4269 3506 4304
rect 1396 4230 3540 4269
rect 1430 4196 3506 4230
rect 1396 4157 3540 4196
rect 1430 4122 3506 4157
rect 1396 4084 3540 4122
rect 1430 4048 3506 4084
rect 1396 4010 3540 4048
rect 1430 3974 3506 4010
rect 1396 3936 3540 3974
rect 1430 3900 3506 3936
rect 1396 3862 3540 3900
rect 1430 3825 3506 3862
rect 1396 3788 3540 3825
rect 1430 3761 3506 3788
rect 1396 3738 1430 3750
rect 3506 3738 3540 3750
rect 3693 4519 3751 4549
rect 3727 4515 3751 4519
rect 3693 4481 3717 4485
rect 3693 4447 3751 4481
rect 3693 4379 3751 4413
rect 3693 4375 3717 4379
rect 3727 4341 3751 4345
rect 3693 4311 3751 4341
rect 3693 4303 3717 4311
rect 3727 4269 3751 4277
rect 3693 4243 3751 4269
rect 3693 4231 3717 4243
rect 3727 4197 3751 4209
rect 3693 4175 3751 4197
rect 3693 4159 3717 4175
rect 3727 4125 3751 4141
rect 3693 4107 3751 4125
rect 3693 4087 3717 4107
rect 3727 4053 3751 4073
rect 3693 4039 3751 4053
rect 3693 4015 3717 4039
rect 3727 3981 3751 4005
rect 3693 3971 3751 3981
rect 3693 3943 3717 3971
rect 3727 3909 3751 3937
rect 4000 11252 4034 11362
rect 4072 11328 4102 11362
rect 4136 11328 4150 11362
rect 4204 11328 4238 11362
rect 4272 11328 4306 11362
rect 4340 11328 4374 11362
rect 4408 11328 4442 11362
rect 4476 11328 4510 11362
rect 4544 11328 4578 11362
rect 4612 11328 4646 11362
rect 4680 11328 4714 11362
rect 4748 11328 4782 11362
rect 4816 11328 4850 11362
rect 4884 11328 4918 11362
rect 4952 11328 4986 11362
rect 5020 11328 5054 11362
rect 5104 11328 5122 11362
rect 5184 11328 5190 11362
rect 5224 11328 5308 11362
rect 5274 11324 5308 11328
rect 5274 11251 5308 11290
rect 4000 11180 4034 11205
rect 4000 11108 4034 11136
rect 4082 11212 4150 11246
rect 4572 11214 4610 11248
rect 4644 11214 4682 11248
rect 5100 11212 5226 11246
rect 4082 11170 4116 11212
rect 5192 11170 5226 11212
rect 4116 11136 5192 11170
rect 4082 11120 4116 11136
rect 5192 11120 5226 11136
rect 5274 11178 5308 11205
rect 5274 11105 5308 11136
rect 4000 11036 4034 11067
rect 4572 11056 4610 11090
rect 4644 11056 4682 11090
rect 4000 10964 4034 10998
rect 4000 10894 4034 10929
rect 4000 10825 4034 10858
rect 4000 10756 4034 10786
rect 4000 10687 4034 10714
rect 4000 10618 4034 10642
rect 4000 10549 4034 10570
rect 4000 10480 4034 10498
rect 4000 10411 4034 10426
rect 4000 10342 4034 10354
rect 4000 10273 4034 10282
rect 4082 11029 4116 11045
rect 4082 10956 4116 10995
rect 4082 10883 4116 10922
rect 4082 10810 4116 10849
rect 4082 10775 4116 10776
rect 5192 11033 5226 11045
rect 5192 10959 5226 10995
rect 5192 10885 5226 10922
rect 5192 10811 5226 10849
rect 5192 10775 5226 10776
rect 4082 10737 5226 10775
rect 4116 10703 5192 10737
rect 4082 10664 5226 10703
rect 4116 10630 5192 10664
rect 4082 10629 5192 10630
rect 4082 10591 5226 10629
rect 4116 10557 5192 10591
rect 4082 10555 5192 10557
rect 4082 10517 5226 10555
rect 4116 10516 5192 10517
rect 4082 10443 4116 10483
rect 4082 10369 4116 10409
rect 4082 10295 4116 10335
rect 4082 10245 4116 10261
rect 5192 10443 5226 10481
rect 5192 10369 5226 10407
rect 5192 10295 5226 10332
rect 5192 10245 5226 10257
rect 5274 11032 5308 11067
rect 5274 10963 5308 10998
rect 5274 10894 5308 10925
rect 5274 10825 5308 10852
rect 5274 10756 5308 10779
rect 5274 10687 5308 10706
rect 5274 10618 5308 10633
rect 5274 10549 5308 10560
rect 5274 10480 5308 10487
rect 5274 10411 5308 10414
rect 5274 10375 5308 10377
rect 5274 10302 5308 10308
rect 4000 10204 4034 10210
rect 4874 10200 4912 10234
rect 4946 10200 4984 10234
rect 5274 10229 5308 10239
rect 4000 10135 4034 10138
rect 4000 10100 4034 10101
rect 4000 10028 4034 10032
rect 4000 9956 4034 9963
rect 4000 9884 4034 9894
rect 4000 9812 4034 9825
rect 4000 9740 4034 9756
rect 4000 9668 4034 9687
rect 4000 9596 4034 9618
rect 4000 9524 4034 9549
rect 4000 9452 4034 9480
rect 4000 9380 4034 9411
rect 4082 10173 4116 10189
rect 4082 10100 4116 10139
rect 4082 10027 4116 10066
rect 4082 9954 4116 9993
rect 4082 9919 4116 9920
rect 5192 10177 5226 10189
rect 5192 10103 5226 10139
rect 5192 10029 5226 10066
rect 5192 9955 5226 9993
rect 5192 9919 5226 9920
rect 4082 9881 5226 9919
rect 4116 9847 5192 9881
rect 4082 9808 5226 9847
rect 4116 9774 5192 9808
rect 4082 9773 5192 9774
rect 4082 9735 5226 9773
rect 4116 9701 5192 9735
rect 4082 9699 5192 9701
rect 4082 9661 5226 9699
rect 4116 9660 5192 9661
rect 4082 9587 4116 9627
rect 4082 9513 4116 9553
rect 4082 9439 4116 9479
rect 4082 9389 4116 9405
rect 5192 9587 5226 9625
rect 5192 9513 5226 9551
rect 5192 9439 5226 9476
rect 5192 9389 5226 9401
rect 5274 10156 5308 10170
rect 5274 10083 5308 10101
rect 5274 10010 5308 10032
rect 5274 9937 5308 9963
rect 5274 9864 5308 9894
rect 5274 9791 5308 9825
rect 5274 9721 5308 9756
rect 5274 9652 5308 9684
rect 5274 9583 5308 9611
rect 5274 9514 5308 9538
rect 5274 9445 5308 9465
rect 4572 9344 4610 9378
rect 4644 9344 4682 9378
rect 5274 9376 5308 9392
rect 4000 9308 4034 9342
rect 4000 9238 4034 9273
rect 4000 9169 4034 9202
rect 4000 9100 4034 9130
rect 4000 9031 4034 9058
rect 4000 8962 4034 8986
rect 4000 8893 4034 8914
rect 4000 8824 4034 8842
rect 4000 8755 4034 8770
rect 4000 8686 4034 8698
rect 4000 8617 4034 8626
rect 4000 8548 4034 8554
rect 4082 9321 4116 9333
rect 4082 9247 4116 9283
rect 4082 9173 4116 9210
rect 4082 9099 4116 9137
rect 4082 9063 4116 9064
rect 5192 9317 5226 9333
rect 5192 9244 5226 9283
rect 5192 9171 5226 9210
rect 5192 9098 5226 9137
rect 5192 9063 5226 9064
rect 4082 9025 5226 9063
rect 4116 8991 5192 9025
rect 4082 8952 5226 8991
rect 4116 8918 5192 8952
rect 4116 8917 5226 8918
rect 4082 8879 5226 8917
rect 4116 8845 5192 8879
rect 4116 8843 5226 8845
rect 4082 8805 5226 8843
rect 4116 8804 5192 8805
rect 4082 8731 4116 8769
rect 4082 8657 4116 8695
rect 4082 8583 4116 8620
rect 4082 8533 4116 8545
rect 5192 8731 5226 8771
rect 5192 8657 5226 8697
rect 5192 8583 5226 8623
rect 5192 8533 5226 8549
rect 5274 9307 5308 9319
rect 5274 9238 5308 9246
rect 5274 9169 5308 9173
rect 5274 9134 5308 9135
rect 5274 9061 5308 9066
rect 5274 8988 5308 8997
rect 5274 8915 5308 8928
rect 5274 8842 5308 8859
rect 5274 8769 5308 8790
rect 5274 8696 5308 8721
rect 5274 8623 5308 8652
rect 5274 8550 5308 8583
rect 4270 8488 4308 8522
rect 4342 8488 4380 8522
rect 4000 8479 4034 8482
rect 5274 8479 5308 8514
rect 4000 8444 4034 8445
rect 4000 8372 4034 8376
rect 4000 8300 4034 8307
rect 4000 8228 4034 8238
rect 4000 8156 4034 8169
rect 4000 8084 4034 8100
rect 4000 8012 4034 8031
rect 4000 7940 4034 7962
rect 4000 7868 4034 7893
rect 4000 7796 4034 7824
rect 4000 7724 4034 7755
rect 4000 7652 4034 7686
rect 4082 8465 4116 8477
rect 4082 8391 4116 8427
rect 4082 8317 4116 8354
rect 4082 8243 4116 8281
rect 4082 8207 4116 8208
rect 5192 8461 5226 8477
rect 5192 8388 5226 8427
rect 5192 8315 5226 8354
rect 5192 8242 5226 8281
rect 5192 8207 5226 8208
rect 4082 8169 5226 8207
rect 4116 8135 5192 8169
rect 4082 8096 5226 8135
rect 4116 8062 5192 8096
rect 4116 8061 5226 8062
rect 4082 8023 5226 8061
rect 4116 7989 5192 8023
rect 4116 7987 5226 7989
rect 4082 7949 5226 7987
rect 4116 7948 5192 7949
rect 4082 7875 4116 7913
rect 4082 7801 4116 7839
rect 4082 7727 4116 7764
rect 4082 7677 4116 7689
rect 5192 7875 5226 7915
rect 5192 7801 5226 7841
rect 5192 7727 5226 7767
rect 5192 7677 5226 7693
rect 5274 8410 5308 8443
rect 5274 8341 5308 8370
rect 5274 8272 5308 8297
rect 5274 8203 5308 8224
rect 5274 8134 5308 8151
rect 5274 8065 5308 8078
rect 5274 7996 5308 8006
rect 5274 7927 5308 7934
rect 5274 7858 5308 7862
rect 5274 7789 5308 7790
rect 5274 7752 5308 7755
rect 5274 7680 5308 7686
rect 4572 7632 4610 7666
rect 4644 7632 4682 7666
rect 4000 7583 4034 7617
rect 4000 7515 4034 7546
rect 4000 7447 4034 7474
rect 4000 7379 4034 7402
rect 4000 7311 4034 7330
rect 4000 7243 4034 7258
rect 4000 7175 4034 7186
rect 4000 7107 4034 7113
rect 4000 7039 4034 7040
rect 4000 7001 4034 7005
rect 4000 6928 4034 6937
rect 4000 6855 4034 6869
rect 4082 7605 4116 7621
rect 4082 7532 4116 7571
rect 4082 7459 4116 7498
rect 4082 7386 4116 7425
rect 4082 7351 4116 7352
rect 5192 7609 5226 7621
rect 5192 7535 5226 7571
rect 5192 7461 5226 7498
rect 5192 7387 5226 7425
rect 5192 7351 5226 7352
rect 4082 7313 5226 7351
rect 4116 7279 5192 7313
rect 4082 7240 5226 7279
rect 4116 7206 5192 7240
rect 4082 7205 5192 7206
rect 4082 7167 5226 7205
rect 4116 7133 5192 7167
rect 4082 7131 5192 7133
rect 4082 7093 5226 7131
rect 4116 7092 5192 7093
rect 4082 7019 4116 7059
rect 4082 6945 4116 6985
rect 4082 6871 4116 6911
rect 4082 6821 4116 6837
rect 5192 7019 5226 7057
rect 5192 6945 5226 6983
rect 5192 6871 5226 6908
rect 5192 6821 5226 6833
rect 5274 7608 5308 7617
rect 5274 7536 5308 7549
rect 5274 7464 5308 7481
rect 5274 7392 5308 7413
rect 5274 7320 5308 7345
rect 5274 7248 5308 7277
rect 5274 7176 5308 7209
rect 5274 7107 5308 7141
rect 5274 7039 5308 7070
rect 5274 6971 5308 6998
rect 5274 6903 5308 6926
rect 5274 6835 5308 6854
rect 4000 6782 4034 6801
rect 4874 6776 4912 6810
rect 4946 6776 4984 6810
rect 5274 6767 5308 6782
rect 4000 6709 4034 6733
rect 4000 6636 4034 6665
rect 4000 6563 4034 6597
rect 4000 6495 4034 6529
rect 4000 6427 4034 6456
rect 4000 6359 4034 6383
rect 4000 6291 4034 6310
rect 4000 6223 4034 6237
rect 4000 6155 4034 6164
rect 4000 6087 4034 6091
rect 4000 6052 4034 6053
rect 4000 5979 4034 5985
rect 4082 6749 4116 6765
rect 4082 6676 4116 6715
rect 4082 6603 4116 6642
rect 4082 6530 4116 6569
rect 4082 6495 4116 6496
rect 5192 6753 5226 6765
rect 5192 6679 5226 6715
rect 5192 6605 5226 6642
rect 5192 6531 5226 6569
rect 5192 6495 5226 6496
rect 4082 6457 5226 6495
rect 4116 6423 5192 6457
rect 4082 6384 5226 6423
rect 4116 6350 5192 6384
rect 4082 6349 5192 6350
rect 4082 6311 5226 6349
rect 4116 6277 5192 6311
rect 4082 6275 5192 6277
rect 4082 6237 5226 6275
rect 4116 6236 5192 6237
rect 4082 6163 4116 6203
rect 4082 6089 4116 6129
rect 4082 6015 4116 6055
rect 4082 5965 4116 5981
rect 5192 6163 5226 6201
rect 5192 6089 5226 6127
rect 5192 6015 5226 6052
rect 5192 5965 5226 5977
rect 5274 6699 5308 6710
rect 5274 6631 5308 6638
rect 5274 6563 5308 6566
rect 5274 6528 5308 6529
rect 5274 6456 5308 6461
rect 5274 6384 5308 6393
rect 5274 6312 5308 6325
rect 5274 6240 5308 6257
rect 5274 6168 5308 6189
rect 5274 6096 5308 6121
rect 5274 6024 5308 6053
rect 4572 5920 4610 5954
rect 4644 5920 4682 5954
rect 5274 5952 5308 5985
rect 4000 5906 4034 5917
rect 4000 5833 4034 5849
rect 4000 5760 4034 5781
rect 4000 5687 4034 5713
rect 4000 5614 4034 5645
rect 4000 5543 4034 5577
rect 4000 5475 4034 5507
rect 4000 5407 4034 5434
rect 4000 5339 4034 5361
rect 4000 5271 4034 5288
rect 4000 5203 4034 5215
rect 4000 5135 4034 5142
rect 4082 5897 4116 5909
rect 4082 5823 4116 5859
rect 4082 5749 4116 5786
rect 4082 5675 4116 5713
rect 4082 5639 4116 5640
rect 5192 5893 5226 5909
rect 5192 5820 5226 5859
rect 5192 5747 5226 5786
rect 5192 5674 5226 5713
rect 5192 5639 5226 5640
rect 4082 5601 5226 5639
rect 4116 5567 5192 5601
rect 4082 5528 5226 5567
rect 4116 5494 5192 5528
rect 4116 5493 5226 5494
rect 4082 5455 5226 5493
rect 4116 5421 5192 5455
rect 4116 5419 5226 5421
rect 4082 5381 5226 5419
rect 4116 5380 5192 5381
rect 4082 5307 4116 5345
rect 4082 5233 4116 5271
rect 4082 5159 4116 5196
rect 4082 5109 4116 5121
rect 5192 5307 5226 5347
rect 5192 5233 5226 5273
rect 5192 5159 5226 5199
rect 5192 5109 5226 5125
rect 5274 5883 5308 5917
rect 5274 5815 5308 5846
rect 5274 5747 5308 5774
rect 5274 5679 5308 5702
rect 5274 5611 5308 5630
rect 5274 5543 5308 5558
rect 5274 5475 5308 5486
rect 5274 5407 5308 5414
rect 5274 5339 5308 5342
rect 5274 5304 5308 5305
rect 5274 5232 5308 5237
rect 5274 5160 5308 5169
rect 4000 5067 4034 5069
rect 4270 5064 4308 5098
rect 4342 5064 4380 5098
rect 5274 5088 5308 5101
rect 4000 5030 4034 5033
rect 4000 4957 4034 4965
rect 4000 4884 4034 4897
rect 4000 4811 4034 4829
rect 4000 4738 4034 4761
rect 4000 4665 4034 4693
rect 4000 4592 4034 4625
rect 4000 4523 4034 4557
rect 4000 4455 4034 4485
rect 4000 4387 4034 4412
rect 4000 4319 4034 4339
rect 4000 4251 4034 4266
rect 4082 5041 4116 5053
rect 4082 4967 4116 5003
rect 4082 4893 4116 4930
rect 4082 4819 4116 4857
rect 4082 4783 4116 4784
rect 5192 5037 5226 5053
rect 5192 4964 5226 5003
rect 5192 4891 5226 4930
rect 5192 4818 5226 4857
rect 5192 4783 5226 4784
rect 4082 4745 5226 4783
rect 4116 4711 5192 4745
rect 4082 4672 5226 4711
rect 4116 4638 5192 4672
rect 4116 4637 5226 4638
rect 4082 4599 5226 4637
rect 4116 4565 5192 4599
rect 4116 4563 5226 4565
rect 4082 4525 5226 4563
rect 4116 4524 5192 4525
rect 4082 4451 4116 4489
rect 4082 4377 4116 4415
rect 4082 4303 4116 4340
rect 4082 4253 4116 4265
rect 5192 4451 5226 4491
rect 5192 4377 5226 4417
rect 5192 4303 5226 4343
rect 5192 4253 5226 4269
rect 5274 5016 5308 5033
rect 5274 4944 5308 4965
rect 5274 4872 5308 4897
rect 5274 4800 5308 4829
rect 5274 4728 5308 4761
rect 5274 4659 5308 4693
rect 5274 4591 5308 4622
rect 5274 4523 5308 4550
rect 5274 4455 5308 4478
rect 5274 4387 5308 4406
rect 5274 4319 5308 4334
rect 5274 4251 5308 4262
rect 4572 4208 4610 4242
rect 4644 4208 4682 4242
rect 4000 4183 4034 4193
rect 5274 4183 5308 4190
rect 4000 4115 4034 4120
rect 4082 4166 4116 4182
rect 5192 4166 5226 4182
rect 4116 4132 5192 4166
rect 4082 4086 4116 4132
rect 5192 4086 5226 4132
rect 4082 4052 4150 4086
rect 4572 4050 4610 4084
rect 4644 4050 4682 4084
rect 5100 4052 5226 4086
rect 5274 4115 5308 4118
rect 5274 4080 5308 4081
rect 4000 4008 4034 4047
rect 4000 3936 4034 3974
rect 5274 4004 5308 4046
rect 4068 3936 4102 3970
rect 4136 3936 4138 3970
rect 4204 3936 4224 3970
rect 4272 3936 4306 3970
rect 4344 3936 4374 3970
rect 4431 3936 4442 3970
rect 4476 3936 4510 3970
rect 4544 3936 4578 3970
rect 4612 3936 4646 3970
rect 4680 3936 4714 3970
rect 4748 3936 4782 3970
rect 4816 3936 4843 3970
rect 4884 3936 4918 3970
rect 4955 3936 4986 3970
rect 5033 3936 5054 3970
rect 5112 3936 5122 3970
rect 5156 3936 5157 3970
rect 5224 3936 5236 3970
rect 5270 3936 5308 3970
rect 5554 11315 5557 11363
rect 5591 11315 5594 11363
rect 7397 11655 7457 11689
rect 7431 11650 7457 11655
rect 7397 11616 7423 11621
rect 7397 11587 7457 11616
rect 7431 11577 7457 11587
rect 7397 11543 7423 11553
rect 7397 11519 7457 11543
rect 7431 11504 7457 11519
rect 7397 11470 7423 11485
rect 7397 11451 7457 11470
rect 7431 11431 7457 11451
rect 9899 11655 9963 11689
rect 9899 11650 9929 11655
rect 9933 11616 9963 11621
rect 9899 11587 9963 11616
rect 9899 11577 9929 11587
rect 9933 11543 9963 11553
rect 9899 11519 9963 11543
rect 9899 11504 9929 11519
rect 9933 11470 9963 11485
rect 9899 11451 9963 11470
rect 9899 11431 9929 11451
rect 7397 11397 7423 11417
rect 7397 11383 7457 11397
rect 7680 11387 7927 11421
rect 5554 11291 5594 11315
rect 5554 11247 5557 11291
rect 5591 11247 5594 11291
rect 5554 11219 5594 11247
rect 5554 11179 5557 11219
rect 5591 11179 5594 11219
rect 5554 11147 5594 11179
rect 5554 11111 5557 11147
rect 5591 11111 5594 11147
rect 5554 11077 5594 11111
rect 5554 11041 5557 11077
rect 5591 11041 5594 11077
rect 5554 11009 5594 11041
rect 5554 10969 5557 11009
rect 5591 10969 5594 11009
rect 5554 10941 5594 10969
rect 5554 10897 5557 10941
rect 5591 10897 5594 10941
rect 5554 10873 5594 10897
rect 5554 10825 5557 10873
rect 5591 10825 5594 10873
rect 5554 10805 5594 10825
rect 5554 10753 5557 10805
rect 5591 10753 5594 10805
rect 5554 10737 5594 10753
rect 5554 10681 5557 10737
rect 5591 10681 5594 10737
rect 5554 10669 5594 10681
rect 5554 10609 5557 10669
rect 5591 10609 5594 10669
rect 5554 10601 5594 10609
rect 5554 10537 5557 10601
rect 5591 10537 5594 10601
rect 5554 10533 5594 10537
rect 5554 10431 5557 10533
rect 5591 10431 5594 10533
rect 5554 10427 5594 10431
rect 5554 10363 5557 10427
rect 5591 10363 5594 10427
rect 5554 10355 5594 10363
rect 5554 10295 5557 10355
rect 5591 10295 5594 10355
rect 5554 10283 5594 10295
rect 5554 10227 5557 10283
rect 5591 10227 5594 10283
rect 5554 10211 5594 10227
rect 5554 10159 5557 10211
rect 5591 10159 5594 10211
rect 5554 10139 5594 10159
rect 5554 10091 5557 10139
rect 5591 10091 5594 10139
rect 5554 10067 5594 10091
rect 5554 10023 5557 10067
rect 5591 10023 5594 10067
rect 5554 9995 5594 10023
rect 5554 9955 5557 9995
rect 5591 9955 5594 9995
rect 5554 9923 5594 9955
rect 5554 9887 5557 9923
rect 5591 9887 5594 9923
rect 5554 9853 5594 9887
rect 5554 9817 5557 9853
rect 5591 9817 5594 9853
rect 5554 9785 5594 9817
rect 5554 9745 5557 9785
rect 5591 9745 5594 9785
rect 5554 9717 5594 9745
rect 5554 9673 5557 9717
rect 5591 9673 5594 9717
rect 5554 9649 5594 9673
rect 5554 9601 5557 9649
rect 5591 9601 5594 9649
rect 5554 9581 5594 9601
rect 5554 9529 5557 9581
rect 5591 9529 5594 9581
rect 5554 9513 5594 9529
rect 5554 9457 5557 9513
rect 5591 9457 5594 9513
rect 5554 9445 5594 9457
rect 5554 9385 5557 9445
rect 5591 9385 5594 9445
rect 5554 9377 5594 9385
rect 5554 9313 5557 9377
rect 5591 9313 5594 9377
rect 5554 9309 5594 9313
rect 5554 9207 5557 9309
rect 5591 9207 5594 9309
rect 5554 9203 5594 9207
rect 5554 9139 5557 9203
rect 5591 9139 5594 9203
rect 5554 9131 5594 9139
rect 5554 9071 5557 9131
rect 5591 9071 5594 9131
rect 5554 9059 5594 9071
rect 5554 9003 5557 9059
rect 5591 9003 5594 9059
rect 5554 8987 5594 9003
rect 5554 8935 5557 8987
rect 5591 8935 5594 8987
rect 5554 8915 5594 8935
rect 5554 8867 5557 8915
rect 5591 8867 5594 8915
rect 5554 8843 5594 8867
rect 5554 8799 5557 8843
rect 5591 8799 5594 8843
rect 5554 8771 5594 8799
rect 5554 8731 5557 8771
rect 5591 8731 5594 8771
rect 5554 8699 5594 8731
rect 5554 8663 5557 8699
rect 5591 8663 5594 8699
rect 5554 8629 5594 8663
rect 5554 8593 5557 8629
rect 5591 8593 5594 8629
rect 5554 8561 5594 8593
rect 5554 8521 5557 8561
rect 5591 8521 5594 8561
rect 5554 8493 5594 8521
rect 5554 8449 5557 8493
rect 5591 8449 5594 8493
rect 5554 8425 5594 8449
rect 5554 8377 5557 8425
rect 5591 8377 5594 8425
rect 5554 8357 5594 8377
rect 5554 8305 5557 8357
rect 5591 8305 5594 8357
rect 5554 8289 5594 8305
rect 5554 8233 5557 8289
rect 5591 8233 5594 8289
rect 5554 8221 5594 8233
rect 5554 8161 5557 8221
rect 5591 8161 5594 8221
rect 5554 8153 5594 8161
rect 5554 8089 5557 8153
rect 5591 8089 5594 8153
rect 5554 8085 5594 8089
rect 5554 7983 5557 8085
rect 5591 7983 5594 8085
rect 5554 7979 5594 7983
rect 5554 7915 5557 7979
rect 5591 7915 5594 7979
rect 5554 7907 5594 7915
rect 5554 7847 5557 7907
rect 5591 7847 5594 7907
rect 5554 7835 5594 7847
rect 5554 7779 5557 7835
rect 5591 7779 5594 7835
rect 5554 7763 5594 7779
rect 5554 7711 5557 7763
rect 5591 7711 5594 7763
rect 5554 7691 5594 7711
rect 5554 7643 5557 7691
rect 5591 7643 5594 7691
rect 5554 7619 5594 7643
rect 5554 7575 5557 7619
rect 5591 7575 5594 7619
rect 5554 7547 5594 7575
rect 5554 7507 5557 7547
rect 5591 7507 5594 7547
rect 5554 7475 5594 7507
rect 5554 7439 5557 7475
rect 5591 7439 5594 7475
rect 5554 7405 5594 7439
rect 5554 7369 5557 7405
rect 5591 7369 5594 7405
rect 5554 7337 5594 7369
rect 5554 7297 5557 7337
rect 5591 7297 5594 7337
rect 5554 7269 5594 7297
rect 5554 7225 5557 7269
rect 5591 7225 5594 7269
rect 5554 7201 5594 7225
rect 5554 7153 5557 7201
rect 5591 7153 5594 7201
rect 5554 7133 5594 7153
rect 5554 7081 5557 7133
rect 5591 7081 5594 7133
rect 5554 7065 5594 7081
rect 5554 7009 5557 7065
rect 5591 7009 5594 7065
rect 5554 6997 5594 7009
rect 5554 6937 5557 6997
rect 5591 6937 5594 6997
rect 5554 6929 5594 6937
rect 5554 6865 5557 6929
rect 5591 6865 5594 6929
rect 5554 6861 5594 6865
rect 5554 6827 5557 6861
rect 5591 6827 5594 6861
rect 5554 6826 5594 6827
rect 5554 6759 5557 6826
rect 5591 6759 5594 6826
rect 5554 6753 5594 6759
rect 5554 6691 5557 6753
rect 5591 6691 5594 6753
rect 5554 6680 5594 6691
rect 5554 6623 5557 6680
rect 5591 6623 5594 6680
rect 5554 6607 5594 6623
rect 5554 6555 5557 6607
rect 5591 6555 5594 6607
rect 5554 6534 5594 6555
rect 5554 6487 5557 6534
rect 5591 6487 5594 6534
rect 5554 6461 5594 6487
rect 5554 6419 5557 6461
rect 5591 6419 5594 6461
rect 5554 6388 5594 6419
rect 5554 6351 5557 6388
rect 5591 6351 5594 6388
rect 5554 6317 5594 6351
rect 5554 6281 5557 6317
rect 5591 6281 5594 6317
rect 5554 6249 5594 6281
rect 5554 6208 5557 6249
rect 5591 6208 5594 6249
rect 5554 6181 5594 6208
rect 5554 6135 5557 6181
rect 5591 6135 5594 6181
rect 5554 6113 5594 6135
rect 5554 6062 5557 6113
rect 5591 6062 5594 6113
rect 5554 6045 5594 6062
rect 5554 5989 5557 6045
rect 5591 5989 5594 6045
rect 5554 5977 5594 5989
rect 5554 5916 5557 5977
rect 5591 5916 5594 5977
rect 5554 5909 5594 5916
rect 5554 5843 5557 5909
rect 5591 5843 5594 5909
rect 5554 5841 5594 5843
rect 5554 5807 5557 5841
rect 5591 5807 5594 5841
rect 5554 5804 5594 5807
rect 5554 5739 5557 5804
rect 5591 5739 5594 5804
rect 5554 5731 5594 5739
rect 5554 5671 5557 5731
rect 5591 5671 5594 5731
rect 5554 5658 5594 5671
rect 5554 5603 5557 5658
rect 5591 5603 5594 5658
rect 5554 5585 5594 5603
rect 5554 5535 5557 5585
rect 5591 5535 5594 5585
rect 5554 5512 5594 5535
rect 5554 5467 5557 5512
rect 5591 5467 5594 5512
rect 5554 5439 5594 5467
rect 5554 5399 5557 5439
rect 5591 5399 5594 5439
rect 5554 5366 5594 5399
rect 5554 5331 5557 5366
rect 5591 5331 5594 5366
rect 5554 5297 5594 5331
rect 5554 5259 5557 5297
rect 5591 5259 5594 5297
rect 5554 5229 5594 5259
rect 5554 5186 5557 5229
rect 5591 5186 5594 5229
rect 5554 5161 5594 5186
rect 5554 5113 5557 5161
rect 5591 5113 5594 5161
rect 5554 5093 5594 5113
rect 5554 5040 5557 5093
rect 5591 5040 5594 5093
rect 5554 5025 5594 5040
rect 5554 4967 5557 5025
rect 5591 4967 5594 5025
rect 5554 4957 5594 4967
rect 5554 4894 5557 4957
rect 5591 4894 5594 4957
rect 5554 4889 5594 4894
rect 5554 4787 5557 4889
rect 5591 4787 5594 4889
rect 5554 4782 5594 4787
rect 5554 4719 5557 4782
rect 5591 4719 5594 4782
rect 5554 4709 5594 4719
rect 5554 4651 5557 4709
rect 5591 4651 5594 4709
rect 5554 4636 5594 4651
rect 5554 4583 5557 4636
rect 5591 4583 5594 4636
rect 5554 4563 5594 4583
rect 5554 4515 5557 4563
rect 5591 4515 5594 4563
rect 5554 4490 5594 4515
rect 5554 4447 5557 4490
rect 5591 4447 5594 4490
rect 5554 4417 5594 4447
rect 5554 4379 5557 4417
rect 5591 4379 5594 4417
rect 5554 4345 5594 4379
rect 5554 4310 5557 4345
rect 5591 4310 5594 4345
rect 5554 4277 5594 4310
rect 5554 4237 5557 4277
rect 5591 4237 5594 4277
rect 5554 4209 5594 4237
rect 5554 4164 5557 4209
rect 5591 4164 5594 4209
rect 5554 4141 5594 4164
rect 5554 4091 5557 4141
rect 5591 4091 5594 4141
rect 5554 4073 5594 4091
rect 5554 4018 5557 4073
rect 5591 4018 5594 4073
rect 5554 4005 5594 4018
rect 5554 3945 5557 4005
rect 5591 3945 5594 4005
rect 5554 3937 5594 3945
rect 3693 3903 3751 3909
rect 3693 3871 3717 3903
rect 3727 3837 3751 3869
rect 3693 3835 3751 3837
rect 3693 3801 3717 3835
rect 3693 3799 3751 3801
rect 3727 3767 3751 3799
rect 1117 3671 1185 3706
rect 3693 3733 3717 3765
rect 3693 3727 3751 3733
rect 3727 3699 3751 3727
rect 1151 3637 1185 3671
rect 2056 3663 2095 3697
rect 2129 3663 2168 3697
rect 2202 3663 2241 3697
rect 2275 3663 2314 3697
rect 2348 3663 2387 3697
rect 1117 3602 1185 3637
rect 1151 3568 1185 3602
rect 1117 3533 1185 3568
rect 1464 3591 2022 3625
rect 2056 3591 2095 3625
rect 2129 3591 2168 3625
rect 2202 3591 2241 3625
rect 2275 3591 2314 3625
rect 2348 3591 2387 3625
rect 3693 3665 3717 3693
rect 5554 3872 5557 3937
rect 5591 3872 5594 3937
rect 5840 11252 5874 11362
rect 5912 11328 5942 11362
rect 5976 11328 5990 11362
rect 6044 11328 6078 11362
rect 6112 11328 6146 11362
rect 6180 11328 6214 11362
rect 6248 11328 6282 11362
rect 6316 11328 6350 11362
rect 6384 11328 6418 11362
rect 6452 11328 6486 11362
rect 6520 11328 6554 11362
rect 6588 11328 6622 11362
rect 6656 11328 6690 11362
rect 6724 11328 6758 11362
rect 6792 11328 6826 11362
rect 6860 11328 6894 11362
rect 6944 11328 6962 11362
rect 7024 11328 7030 11362
rect 7064 11328 7148 11362
rect 7114 11324 7148 11328
rect 7114 11251 7148 11290
rect 5840 11180 5874 11205
rect 5840 11108 5874 11136
rect 5922 11212 5990 11246
rect 6412 11214 6450 11248
rect 6484 11214 6522 11248
rect 6940 11212 7066 11246
rect 5922 11170 5956 11212
rect 7032 11170 7066 11212
rect 5956 11136 7032 11170
rect 5922 11120 5956 11136
rect 7032 11120 7066 11136
rect 7114 11178 7148 11205
rect 7114 11105 7148 11136
rect 5840 11036 5874 11067
rect 6412 11056 6450 11090
rect 6484 11056 6522 11090
rect 5840 10964 5874 10998
rect 5840 10894 5874 10929
rect 5840 10825 5874 10858
rect 5840 10756 5874 10786
rect 5840 10687 5874 10714
rect 5840 10618 5874 10642
rect 5840 10549 5874 10570
rect 5840 10480 5874 10498
rect 5840 10411 5874 10426
rect 5840 10342 5874 10354
rect 5840 10273 5874 10282
rect 5922 11029 5956 11045
rect 5922 10956 5956 10995
rect 5922 10883 5956 10922
rect 5922 10810 5956 10849
rect 5922 10775 5956 10776
rect 7032 11033 7066 11045
rect 7032 10959 7066 10995
rect 7032 10885 7066 10922
rect 7032 10811 7066 10849
rect 7032 10775 7066 10776
rect 5922 10737 7066 10775
rect 5956 10703 7032 10737
rect 5922 10664 7066 10703
rect 5956 10630 7032 10664
rect 5922 10629 7032 10630
rect 5922 10591 7066 10629
rect 5956 10557 7032 10591
rect 5922 10555 7032 10557
rect 5922 10517 7066 10555
rect 5956 10516 7032 10517
rect 5922 10443 5956 10483
rect 5922 10369 5956 10409
rect 5922 10295 5956 10335
rect 5922 10245 5956 10261
rect 7032 10443 7066 10481
rect 7032 10369 7066 10407
rect 7032 10295 7066 10332
rect 7032 10245 7066 10257
rect 7114 11032 7148 11067
rect 7114 10963 7148 10998
rect 7114 10894 7148 10925
rect 7114 10825 7148 10852
rect 7114 10756 7148 10779
rect 7114 10687 7148 10706
rect 7114 10618 7148 10633
rect 7114 10549 7148 10560
rect 7114 10480 7148 10487
rect 7114 10411 7148 10414
rect 7114 10375 7148 10377
rect 7114 10302 7148 10308
rect 5840 10204 5874 10210
rect 6714 10200 6752 10234
rect 6786 10200 6824 10234
rect 7114 10229 7148 10239
rect 5840 10135 5874 10138
rect 5840 10100 5874 10101
rect 5840 10028 5874 10032
rect 5840 9956 5874 9963
rect 5840 9884 5874 9894
rect 5840 9812 5874 9825
rect 5840 9740 5874 9756
rect 5840 9668 5874 9687
rect 5840 9596 5874 9618
rect 5840 9524 5874 9549
rect 5840 9452 5874 9480
rect 5840 9380 5874 9411
rect 5922 10173 5956 10189
rect 5922 10100 5956 10139
rect 5922 10027 5956 10066
rect 5922 9954 5956 9993
rect 5922 9919 5956 9920
rect 7032 10177 7066 10189
rect 7032 10103 7066 10139
rect 7032 10029 7066 10066
rect 7032 9955 7066 9993
rect 7032 9919 7066 9920
rect 5922 9881 7066 9919
rect 5956 9847 7032 9881
rect 5922 9808 7066 9847
rect 5956 9774 7032 9808
rect 5922 9773 7032 9774
rect 5922 9735 7066 9773
rect 5956 9701 7032 9735
rect 5922 9699 7032 9701
rect 5922 9661 7066 9699
rect 5956 9660 7032 9661
rect 5922 9587 5956 9627
rect 5922 9513 5956 9553
rect 5922 9439 5956 9479
rect 5922 9389 5956 9405
rect 7032 9587 7066 9625
rect 7032 9513 7066 9551
rect 7032 9439 7066 9476
rect 7032 9389 7066 9401
rect 7114 10156 7148 10170
rect 7114 10083 7148 10101
rect 7114 10010 7148 10032
rect 7114 9937 7148 9963
rect 7114 9864 7148 9894
rect 7114 9791 7148 9825
rect 7114 9721 7148 9756
rect 7114 9652 7148 9684
rect 7114 9583 7148 9611
rect 7114 9514 7148 9538
rect 7114 9445 7148 9465
rect 6412 9344 6450 9378
rect 6484 9344 6522 9378
rect 7114 9376 7148 9392
rect 5840 9308 5874 9342
rect 5840 9238 5874 9273
rect 5840 9169 5874 9202
rect 5840 9100 5874 9130
rect 5840 9031 5874 9058
rect 5840 8962 5874 8986
rect 5840 8893 5874 8914
rect 5840 8824 5874 8842
rect 5840 8755 5874 8770
rect 5840 8686 5874 8698
rect 5840 8617 5874 8626
rect 5840 8548 5874 8554
rect 5922 9321 5956 9333
rect 5922 9247 5956 9283
rect 5922 9173 5956 9210
rect 5922 9099 5956 9137
rect 5922 9063 5956 9064
rect 7032 9317 7066 9333
rect 7032 9244 7066 9283
rect 7032 9171 7066 9210
rect 7032 9098 7066 9137
rect 7032 9063 7066 9064
rect 5922 9025 7066 9063
rect 5956 8991 7032 9025
rect 5922 8952 7066 8991
rect 5956 8918 7032 8952
rect 5956 8917 7066 8918
rect 5922 8879 7066 8917
rect 5956 8845 7032 8879
rect 5956 8843 7066 8845
rect 5922 8805 7066 8843
rect 5956 8804 7032 8805
rect 5922 8731 5956 8769
rect 5922 8657 5956 8695
rect 5922 8583 5956 8620
rect 5922 8533 5956 8545
rect 7032 8731 7066 8771
rect 7032 8657 7066 8697
rect 7032 8583 7066 8623
rect 7032 8533 7066 8549
rect 7114 9307 7148 9319
rect 7114 9238 7148 9246
rect 7114 9169 7148 9173
rect 7114 9134 7148 9135
rect 7114 9061 7148 9066
rect 7114 8988 7148 8997
rect 7114 8915 7148 8928
rect 7114 8842 7148 8859
rect 7114 8769 7148 8790
rect 7114 8696 7148 8721
rect 7114 8623 7148 8652
rect 7114 8550 7148 8583
rect 6110 8488 6148 8522
rect 6182 8488 6220 8522
rect 5840 8479 5874 8482
rect 7114 8479 7148 8514
rect 5840 8444 5874 8445
rect 5840 8372 5874 8376
rect 5840 8300 5874 8307
rect 5840 8228 5874 8238
rect 5840 8156 5874 8169
rect 5840 8084 5874 8100
rect 5840 8012 5874 8031
rect 5840 7940 5874 7962
rect 5840 7868 5874 7893
rect 5840 7796 5874 7824
rect 5840 7724 5874 7755
rect 5840 7652 5874 7686
rect 5922 8465 5956 8477
rect 5922 8391 5956 8427
rect 5922 8317 5956 8354
rect 5922 8243 5956 8281
rect 5922 8207 5956 8208
rect 7032 8461 7066 8477
rect 7032 8388 7066 8427
rect 7032 8315 7066 8354
rect 7032 8242 7066 8281
rect 7032 8207 7066 8208
rect 5922 8169 7066 8207
rect 5956 8135 7032 8169
rect 5922 8096 7066 8135
rect 5956 8062 7032 8096
rect 5956 8061 7066 8062
rect 5922 8023 7066 8061
rect 5956 7989 7032 8023
rect 5956 7987 7066 7989
rect 5922 7949 7066 7987
rect 5956 7948 7032 7949
rect 5922 7875 5956 7913
rect 5922 7801 5956 7839
rect 5922 7727 5956 7764
rect 5922 7677 5956 7689
rect 7032 7875 7066 7915
rect 7032 7801 7066 7841
rect 7032 7727 7066 7767
rect 7032 7677 7066 7693
rect 7114 8410 7148 8443
rect 7114 8341 7148 8370
rect 7114 8272 7148 8297
rect 7114 8203 7148 8224
rect 7114 8134 7148 8151
rect 7114 8065 7148 8078
rect 7114 7996 7148 8006
rect 7114 7927 7148 7934
rect 7114 7858 7148 7862
rect 7114 7789 7148 7790
rect 7114 7752 7148 7755
rect 7114 7680 7148 7686
rect 6412 7632 6450 7666
rect 6484 7632 6522 7666
rect 5840 7583 5874 7617
rect 5840 7515 5874 7546
rect 5840 7447 5874 7474
rect 5840 7379 5874 7402
rect 5840 7311 5874 7330
rect 5840 7243 5874 7258
rect 5840 7175 5874 7186
rect 5840 7107 5874 7113
rect 5840 7039 5874 7040
rect 5840 7001 5874 7005
rect 5840 6928 5874 6937
rect 5840 6855 5874 6869
rect 5922 7605 5956 7621
rect 5922 7532 5956 7571
rect 5922 7459 5956 7498
rect 5922 7386 5956 7425
rect 5922 7351 5956 7352
rect 7032 7609 7066 7621
rect 7032 7535 7066 7571
rect 7032 7461 7066 7498
rect 7032 7387 7066 7425
rect 7032 7351 7066 7352
rect 5922 7313 7066 7351
rect 5956 7279 7032 7313
rect 5922 7240 7066 7279
rect 5956 7206 7032 7240
rect 5922 7205 7032 7206
rect 5922 7167 7066 7205
rect 5956 7133 7032 7167
rect 5922 7131 7032 7133
rect 5922 7093 7066 7131
rect 5956 7092 7032 7093
rect 5922 7019 5956 7059
rect 5922 6945 5956 6985
rect 5922 6871 5956 6911
rect 5922 6821 5956 6837
rect 7032 7019 7066 7057
rect 7032 6945 7066 6983
rect 7032 6871 7066 6908
rect 7032 6821 7066 6833
rect 7114 7608 7148 7617
rect 7114 7536 7148 7549
rect 7114 7464 7148 7481
rect 7114 7392 7148 7413
rect 7114 7320 7148 7345
rect 7114 7248 7148 7277
rect 7114 7176 7148 7209
rect 7114 7107 7148 7141
rect 7114 7039 7148 7070
rect 7114 6971 7148 6998
rect 7114 6903 7148 6926
rect 7114 6835 7148 6854
rect 5840 6782 5874 6801
rect 6714 6776 6752 6810
rect 6786 6776 6824 6810
rect 7114 6767 7148 6782
rect 5840 6709 5874 6733
rect 5840 6636 5874 6665
rect 5840 6563 5874 6597
rect 5840 6495 5874 6529
rect 5840 6427 5874 6456
rect 5840 6359 5874 6383
rect 5840 6291 5874 6310
rect 5840 6223 5874 6237
rect 5840 6155 5874 6164
rect 5840 6087 5874 6091
rect 5840 6052 5874 6053
rect 5840 5979 5874 5985
rect 5922 6749 5956 6765
rect 5922 6676 5956 6715
rect 5922 6603 5956 6642
rect 5922 6530 5956 6569
rect 5922 6495 5956 6496
rect 7032 6753 7066 6765
rect 7032 6679 7066 6715
rect 7032 6605 7066 6642
rect 7032 6531 7066 6569
rect 7032 6495 7066 6496
rect 5922 6457 7066 6495
rect 5956 6423 7032 6457
rect 5922 6384 7066 6423
rect 5956 6350 7032 6384
rect 5922 6349 7032 6350
rect 5922 6311 7066 6349
rect 5956 6277 7032 6311
rect 5922 6275 7032 6277
rect 5922 6237 7066 6275
rect 5956 6236 7032 6237
rect 5922 6163 5956 6203
rect 5922 6089 5956 6129
rect 5922 6015 5956 6055
rect 5922 5965 5956 5981
rect 7032 6163 7066 6201
rect 7032 6089 7066 6127
rect 7032 6015 7066 6052
rect 7032 5965 7066 5977
rect 7114 6699 7148 6710
rect 7114 6631 7148 6638
rect 7114 6563 7148 6566
rect 7114 6528 7148 6529
rect 7114 6456 7148 6461
rect 7114 6384 7148 6393
rect 7114 6312 7148 6325
rect 7114 6240 7148 6257
rect 7114 6168 7148 6189
rect 7114 6096 7148 6121
rect 7114 6024 7148 6053
rect 6412 5920 6450 5954
rect 6484 5920 6522 5954
rect 7114 5952 7148 5985
rect 5840 5906 5874 5917
rect 5840 5833 5874 5849
rect 5840 5760 5874 5781
rect 5840 5687 5874 5713
rect 5840 5614 5874 5645
rect 5840 5543 5874 5577
rect 5840 5475 5874 5507
rect 5840 5407 5874 5434
rect 5840 5339 5874 5361
rect 5840 5271 5874 5288
rect 5840 5203 5874 5215
rect 5840 5135 5874 5142
rect 5922 5897 5956 5909
rect 5922 5823 5956 5859
rect 5922 5749 5956 5786
rect 5922 5675 5956 5713
rect 5922 5639 5956 5640
rect 7032 5893 7066 5909
rect 7032 5820 7066 5859
rect 7032 5747 7066 5786
rect 7032 5674 7066 5713
rect 7032 5639 7066 5640
rect 5922 5601 7066 5639
rect 5956 5567 7032 5601
rect 5922 5528 7066 5567
rect 5956 5494 7032 5528
rect 5956 5493 7066 5494
rect 5922 5455 7066 5493
rect 5956 5421 7032 5455
rect 5956 5419 7066 5421
rect 5922 5381 7066 5419
rect 5956 5380 7032 5381
rect 5922 5307 5956 5345
rect 5922 5233 5956 5271
rect 5922 5159 5956 5196
rect 5922 5109 5956 5121
rect 7032 5307 7066 5347
rect 7032 5233 7066 5273
rect 7032 5159 7066 5199
rect 7032 5109 7066 5125
rect 7114 5883 7148 5917
rect 7114 5815 7148 5846
rect 7114 5747 7148 5774
rect 7114 5679 7148 5702
rect 7114 5611 7148 5630
rect 7114 5543 7148 5558
rect 7114 5475 7148 5486
rect 7114 5407 7148 5414
rect 7114 5339 7148 5342
rect 7114 5304 7148 5305
rect 7114 5232 7148 5237
rect 7114 5160 7148 5169
rect 5840 5067 5874 5069
rect 6110 5064 6148 5098
rect 6182 5064 6220 5098
rect 7114 5088 7148 5101
rect 5840 5030 5874 5033
rect 5840 4957 5874 4965
rect 5840 4884 5874 4897
rect 5840 4811 5874 4829
rect 5840 4738 5874 4761
rect 5840 4665 5874 4693
rect 5840 4592 5874 4625
rect 5840 4523 5874 4557
rect 5840 4455 5874 4485
rect 5840 4387 5874 4412
rect 5840 4319 5874 4339
rect 5840 4251 5874 4266
rect 5922 5041 5956 5053
rect 5922 4967 5956 5003
rect 5922 4893 5956 4930
rect 5922 4819 5956 4857
rect 5922 4783 5956 4784
rect 7032 5037 7066 5053
rect 7032 4964 7066 5003
rect 7032 4891 7066 4930
rect 7032 4818 7066 4857
rect 7032 4783 7066 4784
rect 5922 4745 7066 4783
rect 5956 4711 7032 4745
rect 5922 4672 7066 4711
rect 5956 4638 7032 4672
rect 5956 4637 7066 4638
rect 5922 4599 7066 4637
rect 5956 4565 7032 4599
rect 5956 4563 7066 4565
rect 5922 4525 7066 4563
rect 5956 4524 7032 4525
rect 5922 4451 5956 4489
rect 5922 4377 5956 4415
rect 5922 4303 5956 4340
rect 5922 4253 5956 4265
rect 7032 4451 7066 4491
rect 7032 4377 7066 4417
rect 7032 4303 7066 4343
rect 7032 4253 7066 4269
rect 7114 5016 7148 5033
rect 7114 4944 7148 4965
rect 7114 4872 7148 4897
rect 7114 4800 7148 4829
rect 7114 4728 7148 4761
rect 7114 4659 7148 4693
rect 7114 4591 7148 4622
rect 7114 4523 7148 4550
rect 7114 4455 7148 4478
rect 7114 4387 7148 4406
rect 7114 4319 7148 4334
rect 7114 4251 7148 4262
rect 6412 4208 6450 4242
rect 6484 4208 6522 4242
rect 5840 4183 5874 4193
rect 7114 4183 7148 4190
rect 5840 4115 5874 4120
rect 5922 4166 5956 4182
rect 7032 4166 7066 4182
rect 5956 4132 7032 4166
rect 5922 4086 5956 4132
rect 7032 4086 7066 4132
rect 5922 4052 5990 4086
rect 6412 4050 6450 4084
rect 6484 4050 6522 4084
rect 6940 4052 7066 4086
rect 7114 4115 7148 4118
rect 7114 4080 7148 4081
rect 5840 4008 5874 4047
rect 5840 3936 5874 3974
rect 7114 4004 7148 4046
rect 5908 3936 5942 3970
rect 5976 3936 5978 3970
rect 6044 3936 6064 3970
rect 6112 3936 6146 3970
rect 6184 3936 6214 3970
rect 6271 3936 6282 3970
rect 6316 3936 6350 3970
rect 6384 3936 6418 3970
rect 6452 3936 6486 3970
rect 6520 3936 6554 3970
rect 6588 3936 6622 3970
rect 6656 3936 6671 3970
rect 6724 3936 6752 3970
rect 6792 3936 6826 3970
rect 6867 3936 6894 3970
rect 6948 3936 6962 3970
rect 7029 3936 7030 3970
rect 7064 3936 7076 3970
rect 7110 3936 7148 3970
rect 7431 11359 7457 11383
rect 7702 11353 7927 11387
rect 7397 11325 7423 11349
rect 7397 11315 7457 11325
rect 7431 11287 7457 11315
rect 7397 11253 7423 11281
rect 7397 11247 7457 11253
rect 8537 11395 8576 11429
rect 8610 11395 8649 11429
rect 8683 11395 8722 11429
rect 8756 11395 8795 11429
rect 8829 11395 8868 11429
rect 8902 11395 9684 11421
rect 8537 11357 9684 11395
rect 8537 11323 8576 11357
rect 8610 11323 8649 11357
rect 8683 11323 8722 11357
rect 8756 11323 8795 11357
rect 8829 11323 8868 11357
rect 8902 11353 9684 11357
rect 9933 11397 9963 11417
rect 9899 11383 9963 11397
rect 9899 11358 9929 11383
rect 9933 11324 9963 11349
rect 9899 11315 9963 11324
rect 9899 11285 9929 11315
rect 8537 11251 8576 11285
rect 8610 11251 8649 11285
rect 8683 11251 8722 11285
rect 8756 11251 8795 11285
rect 8829 11251 8868 11285
rect 9933 11251 9963 11281
rect 7431 11215 7457 11247
rect 9899 11247 9963 11251
rect 7397 11181 7423 11213
rect 7397 11179 7457 11181
rect 7431 11145 7457 11179
rect 7397 11143 7457 11145
rect 7397 11111 7423 11143
rect 7431 11077 7457 11109
rect 7397 11071 7457 11077
rect 7397 11043 7423 11071
rect 7431 11009 7457 11037
rect 7397 10999 7457 11009
rect 7397 10975 7423 10999
rect 7431 10941 7457 10965
rect 7397 10927 7457 10941
rect 7397 10907 7423 10927
rect 7431 10873 7457 10893
rect 7397 10855 7457 10873
rect 7397 10839 7423 10855
rect 7431 10805 7457 10821
rect 7397 10783 7457 10805
rect 7397 10771 7423 10783
rect 7431 10737 7457 10749
rect 7397 10711 7457 10737
rect 7397 10703 7423 10711
rect 7431 10669 7457 10677
rect 7397 10639 7457 10669
rect 7397 10635 7423 10639
rect 7431 10601 7457 10605
rect 7397 10567 7457 10601
rect 7397 10499 7457 10533
rect 7431 10495 7457 10499
rect 7397 10461 7423 10465
rect 7397 10431 7457 10461
rect 7608 11228 7642 11240
rect 9718 11228 9752 11240
rect 7642 11190 9718 11217
rect 7608 11154 9752 11190
rect 7642 11117 9718 11154
rect 7608 11080 9752 11117
rect 7642 11044 9718 11080
rect 7608 11006 9752 11044
rect 7642 10971 9718 11006
rect 7608 10932 9752 10971
rect 7642 10898 9718 10932
rect 7608 10859 9752 10898
rect 7642 10824 9718 10859
rect 7608 10786 9752 10824
rect 7642 10750 9718 10786
rect 7608 10712 9752 10750
rect 7642 10676 9718 10712
rect 7608 10638 9752 10676
rect 7642 10602 9718 10638
rect 7608 10564 9752 10602
rect 7642 10527 9718 10564
rect 7608 10490 9752 10527
rect 7642 10463 9718 10490
rect 7608 10440 7642 10452
rect 9718 10440 9752 10452
rect 9899 11213 9929 11247
rect 9899 11212 9963 11213
rect 9933 11179 9963 11212
rect 9899 11145 9929 11178
rect 9899 11139 9963 11145
rect 9933 11111 9963 11139
rect 9899 11077 9929 11105
rect 9899 11066 9963 11077
rect 9933 11043 9963 11066
rect 9899 11009 9929 11032
rect 9899 10993 9963 11009
rect 9933 10975 9963 10993
rect 9899 10941 9929 10959
rect 9899 10920 9963 10941
rect 9933 10907 9963 10920
rect 9899 10873 9929 10886
rect 9899 10847 9963 10873
rect 9933 10839 9963 10847
rect 9899 10805 9929 10813
rect 9899 10774 9963 10805
rect 9933 10771 9963 10774
rect 9899 10737 9929 10740
rect 9899 10703 9963 10737
rect 9899 10701 9929 10703
rect 9933 10667 9963 10669
rect 9899 10635 9963 10667
rect 9899 10628 9929 10635
rect 9933 10594 9963 10601
rect 9899 10567 9963 10594
rect 9899 10555 9929 10567
rect 9933 10521 9963 10533
rect 9899 10499 9963 10521
rect 9899 10482 9929 10499
rect 9933 10448 9963 10465
rect 7431 10423 7457 10431
rect 7397 10389 7423 10397
rect 9899 10431 9963 10448
rect 9899 10409 9929 10431
rect 7397 10363 7457 10389
rect 7431 10351 7457 10363
rect 7397 10317 7423 10329
rect 7397 10295 7457 10317
rect 7431 10279 7457 10295
rect 7397 10245 7423 10261
rect 7397 10227 7457 10245
rect 7702 10239 7927 10375
rect 7431 10207 7457 10227
rect 8537 10362 8576 10396
rect 8610 10362 8649 10396
rect 8683 10362 8722 10396
rect 8756 10362 8795 10396
rect 8829 10362 8868 10396
rect 9933 10375 9963 10397
rect 8902 10362 9684 10375
rect 8537 10324 9684 10362
rect 8537 10290 8576 10324
rect 8610 10290 8649 10324
rect 8683 10290 8722 10324
rect 8756 10290 8795 10324
rect 8829 10290 8868 10324
rect 8902 10290 9684 10324
rect 8537 10252 9684 10290
rect 8537 10218 8576 10252
rect 8610 10218 8649 10252
rect 8683 10218 8722 10252
rect 8756 10218 8795 10252
rect 8829 10218 8868 10252
rect 8902 10239 9684 10252
rect 9899 10363 9963 10375
rect 9899 10336 9929 10363
rect 9933 10302 9963 10329
rect 9899 10295 9963 10302
rect 9899 10263 9929 10295
rect 9933 10229 9963 10261
rect 9899 10227 9963 10229
rect 7397 10173 7423 10193
rect 7397 10159 7457 10173
rect 7431 10135 7457 10159
rect 9899 10193 9929 10227
rect 9899 10190 9963 10193
rect 9933 10159 9963 10190
rect 7397 10101 7423 10125
rect 7397 10091 7457 10101
rect 7431 10063 7457 10091
rect 7397 10029 7423 10057
rect 7397 10023 7457 10029
rect 7431 9991 7457 10023
rect 7397 9957 7423 9989
rect 7397 9955 7457 9957
rect 7431 9921 7457 9955
rect 7397 9919 7457 9921
rect 7397 9887 7423 9919
rect 7431 9853 7457 9885
rect 7397 9847 7457 9853
rect 7397 9819 7423 9847
rect 7431 9785 7457 9813
rect 7397 9775 7457 9785
rect 7397 9751 7423 9775
rect 7431 9717 7457 9741
rect 7397 9703 7457 9717
rect 7397 9683 7423 9703
rect 7431 9649 7457 9669
rect 7397 9631 7457 9649
rect 7397 9615 7423 9631
rect 7431 9581 7457 9597
rect 7397 9559 7457 9581
rect 7397 9547 7423 9559
rect 7431 9513 7457 9525
rect 7397 9487 7457 9513
rect 7397 9479 7423 9487
rect 7431 9445 7457 9453
rect 7397 9415 7457 9445
rect 7397 9411 7423 9415
rect 7431 9377 7457 9381
rect 7397 9343 7457 9377
rect 7608 10142 7642 10154
rect 9718 10142 9752 10154
rect 7642 10104 9718 10131
rect 7608 10068 9752 10104
rect 7642 10031 9718 10068
rect 7608 9994 9752 10031
rect 7642 9958 9718 9994
rect 7608 9920 9752 9958
rect 7642 9885 9718 9920
rect 7608 9846 9752 9885
rect 7642 9812 9718 9846
rect 7608 9773 9752 9812
rect 7642 9738 9718 9773
rect 7608 9700 9752 9738
rect 7642 9664 9718 9700
rect 7608 9626 9752 9664
rect 7642 9590 9718 9626
rect 7608 9552 9752 9590
rect 7642 9516 9718 9552
rect 7608 9478 9752 9516
rect 7642 9441 9718 9478
rect 7608 9404 9752 9441
rect 7642 9403 9718 9404
rect 7608 9354 7642 9366
rect 9718 9354 9752 9366
rect 9899 10125 9929 10156
rect 9899 10117 9963 10125
rect 9933 10091 9963 10117
rect 9899 10057 9929 10083
rect 9899 10044 9963 10057
rect 9933 10023 9963 10044
rect 9899 9989 9929 10010
rect 9899 9971 9963 9989
rect 9933 9955 9963 9971
rect 9899 9921 9929 9937
rect 9899 9898 9963 9921
rect 9933 9887 9963 9898
rect 9899 9853 9929 9864
rect 9899 9825 9963 9853
rect 9933 9819 9963 9825
rect 9899 9785 9929 9791
rect 9899 9752 9963 9785
rect 9933 9751 9963 9752
rect 9899 9717 9929 9718
rect 9899 9683 9963 9717
rect 9899 9679 9929 9683
rect 9933 9645 9963 9649
rect 9899 9615 9963 9645
rect 9899 9606 9929 9615
rect 9933 9572 9963 9581
rect 9899 9547 9963 9572
rect 9899 9533 9929 9547
rect 9933 9499 9963 9513
rect 9899 9479 9963 9499
rect 9899 9460 9929 9479
rect 9933 9426 9963 9445
rect 9899 9411 9963 9426
rect 9899 9387 9929 9411
rect 9933 9353 9963 9377
rect 9899 9343 9963 9353
rect 7961 9309 7999 9343
rect 8033 9309 8071 9343
rect 8105 9309 8143 9343
rect 8177 9309 8215 9343
rect 8249 9309 8287 9343
rect 8321 9309 8359 9343
rect 8393 9309 8431 9343
rect 8465 9309 8503 9343
rect 8537 9309 8576 9343
rect 8610 9309 8649 9343
rect 8683 9309 8722 9343
rect 8756 9309 8795 9343
rect 8829 9309 8868 9343
rect 9899 9314 9929 9343
rect 7397 9275 7457 9309
rect 7431 9271 7457 9275
rect 7397 9237 7423 9241
rect 7397 9207 7457 9237
rect 7431 9199 7457 9207
rect 7397 9165 7423 9173
rect 7397 9139 7457 9165
rect 7431 9127 7457 9139
rect 7397 9093 7423 9105
rect 7397 9071 7457 9093
rect 7431 9055 7457 9071
rect 7397 9021 7423 9037
rect 7397 9003 7457 9021
rect 7431 8983 7457 9003
rect 7397 8949 7423 8969
rect 7397 8935 7457 8949
rect 7431 8911 7457 8935
rect 7397 8877 7423 8901
rect 7397 8867 7457 8877
rect 7431 8839 7457 8867
rect 7397 8805 7423 8833
rect 7397 8799 7457 8805
rect 7431 8767 7457 8799
rect 7397 8733 7423 8765
rect 7397 8731 7457 8733
rect 7431 8697 7457 8731
rect 7397 8695 7457 8697
rect 7397 8663 7423 8695
rect 7431 8629 7457 8661
rect 7397 8623 7457 8629
rect 7397 8595 7423 8623
rect 7431 8561 7457 8589
rect 7397 8551 7457 8561
rect 7397 8527 7423 8551
rect 7431 8493 7457 8517
rect 7608 9286 7642 9298
rect 9718 9286 9752 9298
rect 7642 9248 9718 9275
rect 7608 9212 9752 9248
rect 7642 9175 9718 9212
rect 7608 9138 9752 9175
rect 7642 9102 9718 9138
rect 7608 9064 9752 9102
rect 7642 9029 9718 9064
rect 7608 8990 9752 9029
rect 7642 8956 9718 8990
rect 7608 8917 9752 8956
rect 7642 8882 9718 8917
rect 7608 8844 9752 8882
rect 7642 8808 9718 8844
rect 7608 8770 9752 8808
rect 7642 8734 9718 8770
rect 7608 8696 9752 8734
rect 7642 8660 9718 8696
rect 7608 8622 9752 8660
rect 7642 8585 9718 8622
rect 7608 8548 9752 8585
rect 7642 8547 9718 8548
rect 7608 8498 7642 8510
rect 9718 8498 9752 8510
rect 9933 9280 9963 9309
rect 9899 9275 9963 9280
rect 9899 9241 9929 9275
rect 9933 9207 9963 9241
rect 9899 9173 9929 9207
rect 9899 9168 9963 9173
rect 9933 9139 9963 9168
rect 9899 9105 9929 9134
rect 9899 9095 9963 9105
rect 9933 9071 9963 9095
rect 9899 9037 9929 9061
rect 9899 9022 9963 9037
rect 9933 9003 9963 9022
rect 9899 8969 9929 8988
rect 9899 8949 9963 8969
rect 9933 8935 9963 8949
rect 9899 8901 9929 8915
rect 9899 8876 9963 8901
rect 9933 8867 9963 8876
rect 9899 8833 9929 8842
rect 9899 8803 9963 8833
rect 9933 8799 9963 8803
rect 9899 8765 9929 8769
rect 9899 8731 9963 8765
rect 9899 8730 9929 8731
rect 9933 8696 9963 8697
rect 9899 8663 9963 8696
rect 9899 8657 9929 8663
rect 9933 8623 9963 8629
rect 9899 8595 9963 8623
rect 9899 8584 9929 8595
rect 9933 8550 9963 8561
rect 9899 8527 9963 8550
rect 9899 8511 9929 8527
rect 7397 8479 7457 8493
rect 7397 8459 7423 8479
rect 7961 8449 7999 8483
rect 8033 8449 8071 8483
rect 8105 8449 8143 8483
rect 8177 8449 8215 8483
rect 8249 8449 8287 8483
rect 8321 8449 8359 8483
rect 8393 8449 8431 8483
rect 8465 8449 8503 8483
rect 8537 8449 8576 8483
rect 8610 8449 8649 8483
rect 8683 8449 8722 8483
rect 8756 8449 8795 8483
rect 8829 8449 8868 8483
rect 9933 8477 9963 8493
rect 9899 8459 9963 8477
rect 7431 8425 7457 8445
rect 7397 8407 7457 8425
rect 9899 8438 9929 8459
rect 7397 8391 7423 8407
rect 7431 8357 7457 8373
rect 7397 8335 7457 8357
rect 7397 8323 7423 8335
rect 7702 8359 9684 8411
rect 7702 8325 7927 8359
rect 7431 8289 7457 8301
rect 7397 8263 7457 8289
rect 7397 8255 7423 8263
rect 8537 8325 8576 8359
rect 8610 8325 8649 8359
rect 8683 8325 8722 8359
rect 8756 8325 8795 8359
rect 8829 8325 8868 8359
rect 8902 8325 9684 8359
rect 9933 8404 9963 8425
rect 9899 8391 9963 8404
rect 9899 8365 9929 8391
rect 9933 8331 9963 8357
rect 9899 8323 9963 8331
rect 9899 8292 9929 8323
rect 8537 8253 8576 8287
rect 8610 8253 8649 8287
rect 8683 8253 8722 8287
rect 8756 8253 8795 8287
rect 8829 8253 8868 8287
rect 9933 8258 9963 8289
rect 9899 8255 9963 8258
rect 7431 8221 7457 8229
rect 7397 8191 7457 8221
rect 9899 8221 9929 8255
rect 9899 8219 9963 8221
rect 7397 8187 7423 8191
rect 7431 8153 7457 8157
rect 7397 8119 7457 8153
rect 7397 8051 7457 8085
rect 7431 8047 7457 8051
rect 7397 8013 7423 8017
rect 7397 7983 7457 8013
rect 7431 7975 7457 7983
rect 7397 7941 7423 7949
rect 7397 7915 7457 7941
rect 7431 7903 7457 7915
rect 7397 7869 7423 7881
rect 7397 7847 7457 7869
rect 7431 7831 7457 7847
rect 7397 7797 7423 7813
rect 7397 7779 7457 7797
rect 7431 7759 7457 7779
rect 7397 7725 7423 7745
rect 7397 7711 7457 7725
rect 7431 7687 7457 7711
rect 7397 7653 7423 7677
rect 7397 7643 7457 7653
rect 7431 7615 7457 7643
rect 7397 7581 7423 7609
rect 7397 7575 7457 7581
rect 7431 7543 7457 7575
rect 7397 7509 7423 7541
rect 7397 7507 7457 7509
rect 7431 7473 7457 7507
rect 7397 7471 7457 7473
rect 7397 7439 7423 7471
rect 7431 7405 7457 7437
rect 7608 8200 7642 8212
rect 9718 8200 9752 8212
rect 7642 8162 9718 8189
rect 7608 8126 9752 8162
rect 7642 8089 9718 8126
rect 7608 8052 9752 8089
rect 7642 8016 9718 8052
rect 7608 7978 9752 8016
rect 7642 7943 9718 7978
rect 7608 7904 9752 7943
rect 7642 7870 9718 7904
rect 7608 7831 9752 7870
rect 7642 7796 9718 7831
rect 7608 7758 9752 7796
rect 7642 7722 9718 7758
rect 7608 7684 9752 7722
rect 7642 7648 9718 7684
rect 7608 7610 9752 7648
rect 7642 7574 9718 7610
rect 7608 7536 9752 7574
rect 7642 7499 9718 7536
rect 7608 7462 9752 7499
rect 7642 7435 9718 7462
rect 7608 7412 7642 7424
rect 9718 7412 9752 7424
rect 9933 8187 9963 8219
rect 9899 8153 9929 8185
rect 9899 8146 9963 8153
rect 9933 8119 9963 8146
rect 9899 8085 9929 8112
rect 9899 8073 9963 8085
rect 9933 8051 9963 8073
rect 9899 8017 9929 8039
rect 9963 8017 9997 8040
rect 9899 8006 9997 8017
rect 10031 8006 10065 8040
rect 10099 8006 10133 8040
rect 10167 8006 10201 8040
rect 10235 8006 10269 8040
rect 10303 8006 10317 8040
rect 10371 8006 10389 8040
rect 10439 8006 10461 8040
rect 10507 8006 10533 8040
rect 10575 8006 10605 8040
rect 10643 8006 10677 8040
rect 10711 8006 10745 8040
rect 10783 8006 10813 8040
rect 10855 8006 10881 8040
rect 10927 8006 10949 8040
rect 10999 8006 11017 8040
rect 11071 8006 11085 8040
rect 11143 8006 11153 8040
rect 11215 8006 11221 8040
rect 11287 8006 11289 8040
rect 11323 8006 11325 8040
rect 11391 8006 11397 8040
rect 11459 8006 11469 8040
rect 11527 8006 11541 8040
rect 11595 8006 11613 8040
rect 11663 8006 11685 8040
rect 11731 8006 11757 8040
rect 11799 8006 11829 8040
rect 11867 8006 11901 8040
rect 11935 8006 11969 8040
rect 12007 8006 12037 8040
rect 12079 8006 12105 8040
rect 12151 8006 12173 8040
rect 12223 8006 12241 8040
rect 12295 8006 12309 8040
rect 12367 8006 12377 8040
rect 12439 8006 12445 8040
rect 12512 8006 12513 8040
rect 12547 8006 12551 8040
rect 12615 8006 12624 8040
rect 12683 8006 12697 8040
rect 12751 8006 12770 8040
rect 12819 8006 12853 8040
rect 12887 8006 12921 8040
rect 12955 8006 12989 8040
rect 13023 8006 13103 8040
rect 9899 8000 9963 8006
rect 9933 7983 9963 8000
rect 9899 7949 9929 7966
rect 9899 7927 9963 7949
rect 9933 7915 9963 7927
rect 9899 7881 9929 7893
rect 9899 7854 9963 7881
rect 9933 7847 9963 7854
rect 9899 7813 9929 7820
rect 9899 7782 9963 7813
rect 9933 7779 9963 7782
rect 9899 7745 9929 7748
rect 9899 7711 9963 7745
rect 9899 7710 9929 7711
rect 13069 7938 13103 7972
rect 13069 7870 13103 7904
rect 13069 7802 13103 7836
rect 13069 7734 13103 7768
rect 10212 7699 10277 7705
rect 9933 7676 9963 7677
rect 9899 7643 9963 7676
rect 9899 7638 9929 7643
rect 9933 7604 9963 7609
rect 9899 7575 9963 7604
rect 9899 7566 9929 7575
rect 9933 7532 9963 7541
rect 9899 7507 9963 7532
rect 9899 7494 9929 7507
rect 9933 7460 9963 7473
rect 9899 7439 9963 7460
rect 9899 7422 9929 7439
rect 7397 7399 7457 7405
rect 7397 7371 7423 7399
rect 7431 7337 7457 7365
rect 7397 7327 7457 7337
rect 7397 7303 7423 7327
rect 7431 7269 7457 7293
rect 7397 7255 7457 7269
rect 7702 7265 7927 7299
rect 7397 7235 7423 7255
rect 7680 7231 7927 7265
rect 8537 7367 8576 7401
rect 8610 7367 8649 7401
rect 8683 7367 8722 7401
rect 8756 7367 8795 7401
rect 8829 7367 8868 7401
rect 9933 7388 9963 7405
rect 9899 7371 9963 7388
rect 9899 7350 9929 7371
rect 8537 7295 8576 7329
rect 8610 7295 8649 7329
rect 8683 7295 8722 7329
rect 8756 7295 8795 7329
rect 8829 7295 8868 7329
rect 9933 7316 9963 7337
rect 9899 7303 9963 7316
rect 8902 7295 9684 7299
rect 8537 7257 9684 7295
rect 8537 7223 8576 7257
rect 8610 7223 8649 7257
rect 8683 7223 8722 7257
rect 8756 7223 8795 7257
rect 8829 7223 8868 7257
rect 8902 7231 9684 7257
rect 9899 7278 9929 7303
rect 9933 7244 9963 7269
rect 9899 7235 9963 7244
rect 7431 7201 7457 7221
rect 7397 7183 7457 7201
rect 7397 7167 7423 7183
rect 7431 7133 7457 7149
rect 7397 7111 7457 7133
rect 7397 7099 7423 7111
rect 7431 7065 7457 7077
rect 7397 7039 7457 7065
rect 7397 7031 7423 7039
rect 7431 6997 7457 7005
rect 7397 6967 7457 6997
rect 7397 6963 7423 6967
rect 9899 7206 9929 7235
rect 9933 7172 9963 7201
rect 9899 7167 9963 7172
rect 9899 7134 9929 7167
rect 9933 7100 9963 7133
rect 9899 7099 9963 7100
rect 9899 7065 9929 7099
rect 9899 7062 9963 7065
rect 9933 7031 9963 7062
rect 9899 6997 9929 7028
rect 9899 6990 9963 6997
rect 9933 6963 9963 6990
rect 7457 6933 7481 6963
rect 7431 6929 7481 6933
rect 7515 6929 7549 6963
rect 7583 6929 7617 6963
rect 7651 6929 7685 6963
rect 7719 6929 7753 6963
rect 7787 6929 7821 6963
rect 7855 6929 7889 6963
rect 7923 6929 7957 6963
rect 7991 6929 8025 6963
rect 8059 6929 8093 6963
rect 8127 6929 8161 6963
rect 8195 6929 8229 6963
rect 8263 6929 8297 6963
rect 8331 6929 8365 6963
rect 8399 6929 8433 6963
rect 8467 6929 8501 6963
rect 8535 6929 8569 6963
rect 8603 6929 8637 6963
rect 8671 6929 8705 6963
rect 8739 6929 8773 6963
rect 8807 6929 8841 6963
rect 8875 6929 8909 6963
rect 8943 6929 8977 6963
rect 9011 6929 9045 6963
rect 9079 6929 9113 6963
rect 9147 6929 9181 6963
rect 9215 6929 9249 6963
rect 9283 6929 9317 6963
rect 9351 6929 9385 6963
rect 9419 6929 9453 6963
rect 9487 6929 9521 6963
rect 9555 6929 9589 6963
rect 9623 6929 9657 6963
rect 9691 6929 9725 6963
rect 9759 6929 9793 6963
rect 9827 6929 9861 6963
rect 9895 6956 9899 6963
rect 9895 6929 9929 6956
rect 7397 6895 7457 6929
rect 7397 6827 7457 6861
rect 7431 6823 7457 6827
rect 7397 6789 7423 6793
rect 7397 6759 7457 6789
rect 7431 6751 7457 6759
rect 7397 6717 7423 6725
rect 7397 6691 7457 6717
rect 7431 6679 7457 6691
rect 9899 6918 9963 6929
rect 9933 6895 9963 6918
rect 9899 6861 9929 6884
rect 9899 6846 9963 6861
rect 9933 6827 9963 6846
rect 9899 6793 9929 6812
rect 9899 6774 9963 6793
rect 9933 6759 9963 6774
rect 9899 6725 9929 6740
rect 9899 6702 9963 6725
rect 9933 6691 9963 6702
rect 7397 6645 7423 6657
rect 7397 6623 7457 6645
rect 7680 6627 8151 6661
rect 7431 6607 7457 6623
rect 7702 6593 8151 6627
rect 7397 6573 7423 6589
rect 7397 6555 7457 6573
rect 7431 6535 7457 6555
rect 7397 6501 7423 6521
rect 7397 6487 7457 6501
rect 8761 6635 8800 6669
rect 8834 6635 8873 6669
rect 8907 6635 8946 6669
rect 8980 6635 9019 6669
rect 9053 6635 9092 6669
rect 9126 6635 9684 6661
rect 8761 6597 9684 6635
rect 8761 6563 8800 6597
rect 8834 6563 8873 6597
rect 8907 6563 8946 6597
rect 8980 6563 9019 6597
rect 9053 6563 9092 6597
rect 9126 6593 9684 6597
rect 9899 6657 9929 6668
rect 9899 6630 9963 6657
rect 9933 6623 9963 6630
rect 9899 6589 9929 6596
rect 9899 6558 9963 6589
rect 9933 6555 9963 6558
rect 8761 6491 8800 6525
rect 8834 6491 8873 6525
rect 8907 6491 8946 6525
rect 8980 6491 9019 6525
rect 9053 6491 9092 6525
rect 9899 6521 9929 6524
rect 7431 6463 7457 6487
rect 9899 6487 9963 6521
rect 9899 6486 9929 6487
rect 7397 6429 7423 6453
rect 7397 6419 7457 6429
rect 7431 6391 7457 6419
rect 7397 6357 7423 6385
rect 7397 6351 7457 6357
rect 7431 6319 7457 6351
rect 7397 6285 7423 6317
rect 7397 6283 7457 6285
rect 7431 6249 7457 6283
rect 7397 6247 7457 6249
rect 7397 6215 7423 6247
rect 7431 6181 7457 6213
rect 7397 6175 7457 6181
rect 7397 6147 7423 6175
rect 7431 6113 7457 6141
rect 7397 6103 7457 6113
rect 7397 6079 7423 6103
rect 7431 6045 7457 6069
rect 7397 6031 7457 6045
rect 7397 6011 7423 6031
rect 7431 5977 7457 5997
rect 7397 5959 7457 5977
rect 7397 5943 7423 5959
rect 7431 5909 7457 5925
rect 7397 5887 7457 5909
rect 7397 5875 7423 5887
rect 7431 5841 7457 5853
rect 7397 5815 7457 5841
rect 7397 5807 7423 5815
rect 7431 5773 7457 5781
rect 7397 5743 7457 5773
rect 7397 5739 7423 5743
rect 7431 5705 7457 5709
rect 7397 5671 7457 5705
rect 7608 6468 7642 6480
rect 9718 6468 9752 6480
rect 7642 6430 9718 6457
rect 7608 6395 9752 6430
rect 7642 6358 9718 6395
rect 7608 6326 9752 6358
rect 7642 6282 9718 6326
rect 7608 6257 9752 6282
rect 7642 6205 9718 6257
rect 7608 6188 9752 6205
rect 7642 6128 9718 6188
rect 7608 6119 9752 6128
rect 7642 6051 9718 6119
rect 7608 6050 9752 6051
rect 7642 6016 9718 6050
rect 7608 6008 9752 6016
rect 7642 5947 9718 6008
rect 7608 5931 9752 5947
rect 7642 5878 9718 5931
rect 7608 5854 9752 5878
rect 7642 5809 9718 5854
rect 7608 5777 9752 5809
rect 7642 5740 9718 5777
rect 7608 5704 9752 5740
rect 7642 5703 9718 5704
rect 7608 5654 7642 5666
rect 9718 5654 9752 5666
rect 9933 6452 9963 6453
rect 9899 6419 9963 6452
rect 9899 6414 9929 6419
rect 9933 6380 9963 6385
rect 9899 6351 9963 6380
rect 9899 6342 9929 6351
rect 9933 6308 9963 6317
rect 9899 6283 9963 6308
rect 9899 6270 9929 6283
rect 9933 6236 9963 6249
rect 9899 6215 9963 6236
rect 9899 6198 9929 6215
rect 9933 6164 9963 6181
rect 9899 6147 9963 6164
rect 9899 6126 9929 6147
rect 9933 6092 9963 6113
rect 9899 6079 9963 6092
rect 9899 6054 9929 6079
rect 9933 6020 9963 6045
rect 9899 6011 9963 6020
rect 9899 5982 9929 6011
rect 9933 5948 9963 5977
rect 9899 5943 9963 5948
rect 9899 5910 9929 5943
rect 9933 5876 9963 5909
rect 9899 5875 9963 5876
rect 9899 5841 9929 5875
rect 9899 5838 9963 5841
rect 9933 5807 9963 5838
rect 9899 5773 9929 5804
rect 9899 5766 9963 5773
rect 9933 5739 9963 5766
rect 9899 5705 9929 5732
rect 9899 5694 9963 5705
rect 9933 5671 9963 5694
rect 7397 5603 7457 5637
rect 9899 5637 9929 5660
rect 9899 5622 9963 5637
rect 7431 5599 7457 5603
rect 7397 5565 7423 5569
rect 7397 5535 7457 5565
rect 7431 5527 7457 5535
rect 7397 5493 7423 5501
rect 7397 5467 7457 5493
rect 7431 5455 7457 5467
rect 7702 5439 8151 5575
rect 7397 5421 7423 5433
rect 8761 5576 8800 5610
rect 8834 5576 8873 5610
rect 8907 5576 8946 5610
rect 8980 5576 9019 5610
rect 9053 5576 9092 5610
rect 9933 5603 9963 5622
rect 8761 5538 9684 5575
rect 8761 5504 8800 5538
rect 8834 5504 8873 5538
rect 8907 5504 8946 5538
rect 8980 5504 9019 5538
rect 9053 5504 9092 5538
rect 9126 5504 9684 5538
rect 8761 5466 9684 5504
rect 8761 5432 8800 5466
rect 8834 5432 8873 5466
rect 8907 5432 8946 5466
rect 8980 5432 9019 5466
rect 9053 5432 9092 5466
rect 9126 5439 9684 5466
rect 9899 5569 9929 5588
rect 9899 5550 9963 5569
rect 9933 5535 9963 5550
rect 9899 5501 9929 5516
rect 9899 5478 9963 5501
rect 9933 5467 9963 5478
rect 9899 5433 9929 5444
rect 7397 5399 7457 5421
rect 7431 5383 7457 5399
rect 9899 5406 9963 5433
rect 9933 5399 9963 5406
rect 7397 5349 7423 5365
rect 7397 5331 7457 5349
rect 7431 5311 7457 5331
rect 7397 5277 7423 5297
rect 7397 5263 7457 5277
rect 7431 5239 7457 5263
rect 7397 5205 7423 5229
rect 7397 5195 7457 5205
rect 7431 5167 7457 5195
rect 7397 5133 7423 5161
rect 7397 5127 7457 5133
rect 7431 5095 7457 5127
rect 7397 5061 7423 5093
rect 7397 5059 7457 5061
rect 7431 5025 7457 5059
rect 7397 5023 7457 5025
rect 7397 4991 7423 5023
rect 7431 4957 7457 4989
rect 7397 4951 7457 4957
rect 7397 4923 7423 4951
rect 7431 4889 7457 4917
rect 7397 4879 7457 4889
rect 7397 4855 7423 4879
rect 7431 4821 7457 4845
rect 7397 4807 7457 4821
rect 7397 4787 7423 4807
rect 7431 4753 7457 4773
rect 7397 4735 7457 4753
rect 7397 4719 7423 4735
rect 7431 4685 7457 4701
rect 7397 4663 7457 4685
rect 7397 4651 7423 4663
rect 7431 4617 7457 4629
rect 7397 4591 7457 4617
rect 7608 5382 7642 5394
rect 9718 5382 9752 5394
rect 7642 5344 9718 5371
rect 7608 5308 9752 5344
rect 7642 5271 9718 5308
rect 7608 5234 9752 5271
rect 7642 5198 9718 5234
rect 7608 5160 9752 5198
rect 7642 5125 9718 5160
rect 7608 5086 9752 5125
rect 7642 5052 9718 5086
rect 7608 5013 9752 5052
rect 7642 4978 9718 5013
rect 7608 4940 9752 4978
rect 7642 4904 9718 4940
rect 7608 4866 9752 4904
rect 7642 4830 9718 4866
rect 7608 4792 9752 4830
rect 7642 4756 9718 4792
rect 7608 4718 9752 4756
rect 7642 4681 9718 4718
rect 7608 4644 9752 4681
rect 7642 4617 9718 4644
rect 7608 4594 7642 4606
rect 9718 4594 9752 4606
rect 9899 5365 9929 5372
rect 9899 5334 9963 5365
rect 9933 5331 9963 5334
rect 9899 5297 9929 5300
rect 9899 5263 9963 5297
rect 9899 5262 9929 5263
rect 9933 5228 9963 5229
rect 9899 5195 9963 5228
rect 9899 5190 9929 5195
rect 9933 5156 9963 5161
rect 9899 5127 9963 5156
rect 9899 5118 9929 5127
rect 9933 5084 9963 5093
rect 9899 5059 9963 5084
rect 9899 5046 9929 5059
rect 9933 5012 9963 5025
rect 9899 4991 9963 5012
rect 9899 4974 9929 4991
rect 9933 4940 9963 4957
rect 9899 4923 9963 4940
rect 9899 4902 9929 4923
rect 9933 4868 9963 4889
rect 9899 4855 9963 4868
rect 9899 4830 9929 4855
rect 9933 4796 9963 4821
rect 9899 4787 9963 4796
rect 9899 4758 9929 4787
rect 9933 4724 9963 4753
rect 9899 4719 9963 4724
rect 9899 4686 9929 4719
rect 9933 4652 9963 4685
rect 9899 4651 9963 4652
rect 9899 4617 9929 4651
rect 9899 4614 9963 4617
rect 7397 4583 7423 4591
rect 9933 4583 9963 4614
rect 7431 4549 7457 4557
rect 8185 4549 8223 4583
rect 8257 4549 8295 4583
rect 8329 4549 8367 4583
rect 8401 4549 8439 4583
rect 8473 4549 8511 4583
rect 8545 4549 8583 4583
rect 8617 4549 8655 4583
rect 8689 4549 8727 4583
rect 8761 4549 8800 4583
rect 8834 4549 8873 4583
rect 8907 4549 8946 4583
rect 8980 4549 9019 4583
rect 9053 4549 9092 4583
rect 9899 4549 9929 4580
rect 7397 4519 7457 4549
rect 9899 4542 9963 4549
rect 7397 4515 7423 4519
rect 7431 4481 7457 4485
rect 7397 4447 7457 4481
rect 7397 4379 7457 4413
rect 7431 4375 7457 4379
rect 7397 4341 7423 4345
rect 7397 4311 7457 4341
rect 7431 4303 7457 4311
rect 7397 4269 7423 4277
rect 7397 4243 7457 4269
rect 7431 4231 7457 4243
rect 7397 4197 7423 4209
rect 7397 4175 7457 4197
rect 7431 4159 7457 4175
rect 7397 4125 7423 4141
rect 7397 4107 7457 4125
rect 7431 4087 7457 4107
rect 7397 4053 7423 4073
rect 7397 4039 7457 4053
rect 7431 4015 7457 4039
rect 7397 3981 7423 4005
rect 7397 3971 7457 3981
rect 7431 3943 7457 3971
rect 5554 3869 5594 3872
rect 5554 3835 5557 3869
rect 5591 3835 5594 3869
rect 5554 3833 5594 3835
rect 5554 3767 5557 3833
rect 5591 3767 5594 3833
rect 5554 3760 5594 3767
rect 5554 3726 5557 3760
rect 5591 3726 5594 3760
rect 5554 3687 5594 3726
rect 7397 3909 7423 3937
rect 7397 3903 7457 3909
rect 7431 3871 7457 3903
rect 7397 3837 7423 3869
rect 7397 3835 7457 3837
rect 7431 3801 7457 3835
rect 7397 3799 7457 3801
rect 7397 3767 7423 3799
rect 7431 3733 7457 3765
rect 7608 4526 7642 4538
rect 9718 4526 9752 4538
rect 7642 4488 9718 4515
rect 7608 4452 9752 4488
rect 7642 4415 9718 4452
rect 7608 4378 9752 4415
rect 7642 4342 9718 4378
rect 7608 4304 9752 4342
rect 7642 4269 9718 4304
rect 7608 4230 9752 4269
rect 7642 4196 9718 4230
rect 7608 4157 9752 4196
rect 7642 4122 9718 4157
rect 7608 4084 9752 4122
rect 7642 4048 9718 4084
rect 7608 4010 9752 4048
rect 7642 3974 9718 4010
rect 7608 3936 9752 3974
rect 7642 3900 9718 3936
rect 7608 3862 9752 3900
rect 7642 3825 9718 3862
rect 7608 3788 9752 3825
rect 7642 3761 9718 3788
rect 7608 3738 7642 3750
rect 9718 3738 9752 3750
rect 9933 4515 9963 4542
rect 9899 4481 9929 4508
rect 9899 4470 9963 4481
rect 9933 4447 9963 4470
rect 9899 4413 9929 4436
rect 9899 4398 9963 4413
rect 9933 4379 9963 4398
rect 9899 4345 9929 4364
rect 9899 4326 9963 4345
rect 9933 4311 9963 4326
rect 9899 4277 9929 4292
rect 9899 4254 9963 4277
rect 9933 4243 9963 4254
rect 9899 4209 9929 4220
rect 9899 4182 9963 4209
rect 9933 4175 9963 4182
rect 9899 4141 9929 4148
rect 9899 4110 9963 4141
rect 9933 4107 9963 4110
rect 9899 4073 9929 4076
rect 9899 4039 9963 4073
rect 9899 4038 9929 4039
rect 9933 4004 9963 4005
rect 9899 3971 9963 4004
rect 9899 3966 9929 3971
rect 9933 3932 9963 3937
rect 9899 3903 9963 3932
rect 9899 3894 9929 3903
rect 9933 3860 9963 3869
rect 9899 3835 9963 3860
rect 9899 3822 9929 3835
rect 9933 3788 9963 3801
rect 9899 3767 9963 3788
rect 9899 3750 9929 3767
rect 7397 3727 7457 3733
rect 7397 3699 7423 3727
rect 9933 3716 9963 3733
rect 9899 3699 9963 3716
rect 3751 3665 3785 3687
rect 3693 3655 3785 3665
rect 3727 3653 3785 3655
rect 3819 3653 3853 3687
rect 3887 3653 3921 3687
rect 3955 3653 3989 3687
rect 4023 3653 4057 3687
rect 4091 3653 4125 3687
rect 4159 3653 4193 3687
rect 4227 3653 4261 3687
rect 4295 3653 4329 3687
rect 4363 3653 4397 3687
rect 4431 3653 4465 3687
rect 4499 3653 4533 3687
rect 4567 3653 4601 3687
rect 4635 3653 4669 3687
rect 4703 3653 4737 3687
rect 4771 3653 4805 3687
rect 4839 3653 4873 3687
rect 4907 3653 4941 3687
rect 4975 3653 5009 3687
rect 5043 3653 5077 3687
rect 5111 3653 5145 3687
rect 5179 3653 5213 3687
rect 5247 3653 5281 3687
rect 5315 3653 5349 3687
rect 5383 3653 5417 3687
rect 5451 3653 5485 3687
rect 5519 3653 5557 3687
rect 5591 3653 5625 3687
rect 5659 3653 5693 3687
rect 5727 3653 5761 3687
rect 5795 3653 5829 3687
rect 5863 3653 5897 3687
rect 5931 3653 5965 3687
rect 5999 3653 6033 3687
rect 6067 3653 6101 3687
rect 6135 3653 6169 3687
rect 6203 3653 6237 3687
rect 6271 3653 6305 3687
rect 6339 3653 6373 3687
rect 6407 3653 6441 3687
rect 6475 3653 6509 3687
rect 6543 3653 6577 3687
rect 6611 3653 6645 3687
rect 6679 3653 6713 3687
rect 6747 3653 6781 3687
rect 6815 3653 6849 3687
rect 6883 3653 6917 3687
rect 6951 3653 6985 3687
rect 7019 3653 7053 3687
rect 7087 3653 7121 3687
rect 7155 3653 7189 3687
rect 7223 3653 7257 3687
rect 7291 3653 7325 3687
rect 7359 3665 7397 3687
rect 7431 3665 7457 3693
rect 7359 3655 7457 3665
rect 7359 3653 7423 3655
rect 3727 3631 3751 3653
rect 2997 3591 3446 3625
rect 1464 3565 3446 3591
rect 3693 3597 3717 3621
rect 3693 3583 3751 3597
rect 1151 3499 1185 3533
rect 3727 3563 3751 3583
rect 3693 3529 3717 3549
rect 1117 3464 1185 3499
rect 2056 3493 2095 3527
rect 2129 3493 2168 3527
rect 2202 3493 2241 3527
rect 2275 3493 2314 3527
rect 2348 3493 2387 3527
rect 2421 3493 2459 3527
rect 2493 3493 2531 3527
rect 2565 3493 2603 3527
rect 2637 3493 2675 3527
rect 2709 3493 2747 3527
rect 2781 3493 2819 3527
rect 2853 3493 2891 3527
rect 2925 3493 2963 3527
rect 3693 3511 3751 3529
rect 3727 3495 3751 3511
rect 1151 3430 1185 3464
rect 3693 3461 3717 3477
rect 1117 3395 1185 3430
rect 1151 3361 1185 3395
rect 1117 3326 1185 3361
rect 1151 3292 1185 3326
rect 1117 3257 1185 3292
rect 1151 3223 1185 3257
rect 1117 3188 1185 3223
rect 1151 3154 1185 3188
rect 1117 3119 1185 3154
rect 1151 3085 1185 3119
rect 1117 3050 1185 3085
rect 1151 3016 1185 3050
rect 1117 2981 1185 3016
rect 1151 2947 1185 2981
rect 1117 2912 1185 2947
rect 1151 2878 1185 2912
rect 1117 2843 1185 2878
rect 1151 2809 1185 2843
rect 1117 2774 1185 2809
rect 1151 2740 1185 2774
rect 1117 2705 1185 2740
rect 1151 2671 1185 2705
rect 1117 2636 1185 2671
rect 1396 3440 1430 3452
rect 3506 3440 3540 3452
rect 1430 3402 3506 3429
rect 1396 3366 3540 3402
rect 1430 3329 3506 3366
rect 1396 3292 3540 3329
rect 1430 3256 3506 3292
rect 1396 3218 3540 3256
rect 1430 3183 3506 3218
rect 1396 3144 3540 3183
rect 1430 3110 3506 3144
rect 1396 3071 3540 3110
rect 1430 3036 3506 3071
rect 1396 2998 3540 3036
rect 1430 2962 3506 2998
rect 1396 2924 3540 2962
rect 1430 2888 3506 2924
rect 1396 2850 3540 2888
rect 1430 2814 3506 2850
rect 1396 2776 3540 2814
rect 1430 2739 3506 2776
rect 1396 2702 3540 2739
rect 1430 2675 3506 2702
rect 1396 2652 1430 2664
rect 3506 2652 3540 2664
rect 3693 3439 3751 3461
rect 3727 3427 3751 3439
rect 3693 3393 3717 3405
rect 3693 3367 3751 3393
rect 7397 3631 7423 3653
rect 7431 3597 7457 3621
rect 7397 3583 7457 3597
rect 7397 3563 7423 3583
rect 7702 3591 8151 3625
rect 8761 3663 8800 3697
rect 8834 3663 8873 3697
rect 8907 3663 8946 3697
rect 8980 3663 9019 3697
rect 9053 3663 9092 3697
rect 9899 3678 9929 3699
rect 9933 3644 9963 3665
rect 9899 3631 9963 3644
rect 8761 3591 8800 3625
rect 8834 3591 8873 3625
rect 8907 3591 8946 3625
rect 8980 3591 9019 3625
rect 9053 3591 9092 3625
rect 9126 3591 9684 3625
rect 7702 3565 9684 3591
rect 9899 3606 9929 3631
rect 9933 3572 9963 3597
rect 7431 3529 7457 3549
rect 7397 3511 7457 3529
rect 9899 3563 9963 3572
rect 9899 3534 9929 3563
rect 7397 3495 7423 3511
rect 8185 3493 8223 3527
rect 8257 3493 8295 3527
rect 8329 3493 8367 3527
rect 8401 3493 8439 3527
rect 8473 3493 8511 3527
rect 8545 3493 8583 3527
rect 8617 3493 8655 3527
rect 8689 3493 8727 3527
rect 8761 3493 8800 3527
rect 8834 3493 8873 3527
rect 8907 3493 8946 3527
rect 8980 3493 9019 3527
rect 9053 3493 9092 3527
rect 9933 3500 9963 3529
rect 9899 3495 9963 3500
rect 7431 3461 7457 3477
rect 7397 3439 7457 3461
rect 9899 3462 9929 3495
rect 7397 3427 7423 3439
rect 7431 3393 7457 3405
rect 3727 3359 3751 3367
rect 3693 3325 3717 3333
rect 3693 3295 3751 3325
rect 3727 3291 3751 3295
rect 3693 3257 3717 3261
rect 3693 3223 3751 3257
rect 3693 3155 3751 3189
rect 3693 3151 3717 3155
rect 3727 3117 3751 3121
rect 3693 3087 3751 3117
rect 3693 3079 3717 3087
rect 3727 3045 3751 3053
rect 3693 3019 3751 3045
rect 3693 3007 3717 3019
rect 3727 2973 3751 2985
rect 3693 2951 3751 2973
rect 3693 2935 3717 2951
rect 3727 2901 3751 2917
rect 3693 2883 3751 2901
rect 3693 2863 3717 2883
rect 3727 2829 3751 2849
rect 3693 2815 3751 2829
rect 3693 2791 3717 2815
rect 3727 2757 3751 2781
rect 3693 2747 3751 2757
rect 3693 2719 3717 2747
rect 3727 2685 3751 2713
rect 3693 2679 3751 2685
rect 1151 2602 1185 2636
rect 3693 2647 3717 2679
rect 1117 2577 1185 2602
rect 2056 2607 2095 2641
rect 2129 2607 2168 2641
rect 2202 2607 2241 2641
rect 2275 2607 2314 2641
rect 2348 2607 2387 2641
rect 1117 2573 1287 2577
rect 1117 2567 1185 2573
rect 1151 2533 1185 2567
rect 1219 2542 1287 2573
rect 1117 2509 1185 2533
rect 1219 2509 1253 2542
rect 1117 2508 1253 2509
rect 1117 2501 1287 2508
rect 1117 2498 1185 2501
rect 1151 2464 1185 2498
rect 1219 2473 1287 2501
rect 1117 2441 1185 2464
rect 1219 2441 1253 2473
rect 1117 2439 1253 2441
rect 1464 2535 2022 2539
rect 2056 2535 2095 2569
rect 2129 2535 2168 2569
rect 2202 2535 2241 2569
rect 2275 2535 2314 2569
rect 2348 2535 2387 2569
rect 1464 2497 2387 2535
rect 1464 2471 2022 2497
rect 2056 2463 2095 2497
rect 2129 2463 2168 2497
rect 2202 2463 2241 2497
rect 2275 2463 2314 2497
rect 2348 2463 2387 2497
rect 3727 2613 3751 2645
rect 3693 2611 3751 2613
rect 3693 2577 3717 2611
rect 3693 2575 3751 2577
rect 3727 2543 3751 2575
rect 2997 2505 3446 2539
rect 3693 2509 3717 2541
rect 2997 2471 3468 2505
rect 3693 2503 3751 2509
rect 3727 2475 3751 2503
rect 1117 2429 1287 2439
rect 1151 2395 1185 2429
rect 1219 2404 1287 2429
rect 1117 2373 1185 2395
rect 1219 2373 1253 2404
rect 1117 2370 1253 2373
rect 1117 2360 1287 2370
rect 1151 2357 1287 2360
rect 1151 2326 1185 2357
rect 1117 2305 1185 2326
rect 1219 2335 1287 2357
rect 1219 2305 1253 2335
rect 1117 2301 1253 2305
rect 1117 2291 1287 2301
rect 1151 2285 1287 2291
rect 1151 2257 1185 2285
rect 1117 2237 1185 2257
rect 1219 2266 1287 2285
rect 1219 2237 1253 2266
rect 1117 2232 1253 2237
rect 1117 2222 1287 2232
rect 1151 2213 1287 2222
rect 1151 2188 1185 2213
rect 1219 2203 1287 2213
rect 3693 2441 3717 2469
rect 3693 2431 3751 2441
rect 3727 2407 3751 2431
rect 3693 2373 3717 2397
rect 3693 2359 3751 2373
rect 3727 2339 3751 2359
rect 3693 2305 3717 2325
rect 3693 2287 3751 2305
rect 3727 2271 3751 2287
rect 3693 2237 3717 2253
rect 3693 2215 3751 2237
rect 1117 2169 1185 2188
rect 1219 2197 1371 2203
rect 1219 2169 1253 2197
rect 1117 2163 1253 2169
rect 1287 2169 1371 2197
rect 1405 2169 1439 2203
rect 1473 2169 1507 2203
rect 1541 2169 1575 2203
rect 1609 2169 1643 2203
rect 1677 2169 1711 2203
rect 1745 2169 1779 2203
rect 1813 2169 1847 2203
rect 1881 2169 1915 2203
rect 1949 2169 1983 2203
rect 2017 2169 2051 2203
rect 2085 2169 2119 2203
rect 2153 2169 2187 2203
rect 2221 2169 2255 2203
rect 2289 2169 2323 2203
rect 2357 2169 2391 2203
rect 2425 2169 2459 2203
rect 2493 2169 2527 2203
rect 2561 2169 2595 2203
rect 2629 2169 2663 2203
rect 2697 2169 2731 2203
rect 2765 2169 2799 2203
rect 2833 2169 2867 2203
rect 2901 2169 2935 2203
rect 2969 2169 3003 2203
rect 3037 2169 3071 2203
rect 3105 2169 3139 2203
rect 3173 2169 3207 2203
rect 3241 2169 3275 2203
rect 3309 2169 3343 2203
rect 3377 2169 3411 2203
rect 3445 2169 3479 2203
rect 3513 2169 3547 2203
rect 3581 2169 3615 2203
rect 3649 2169 3683 2203
rect 3727 2181 3751 2215
rect 3717 2169 3751 2181
rect 4000 3354 4034 3378
rect 5100 3336 5228 3370
rect 4000 3285 4034 3320
rect 4000 3216 4034 3251
rect 4000 3147 4034 3182
rect 5194 3311 5228 3336
rect 5194 3243 5228 3277
rect 5194 3175 5228 3209
rect 5194 3125 5228 3141
rect 5276 3354 5310 3378
rect 5276 3285 5310 3320
rect 5276 3248 5310 3251
rect 5838 3354 5872 3378
rect 6940 3336 7066 3370
rect 5838 3285 5872 3320
rect 5838 3248 5872 3251
rect 5276 3216 5344 3248
rect 5310 3214 5344 3216
rect 5378 3214 5415 3248
rect 5449 3214 5486 3248
rect 5520 3214 5557 3248
rect 5591 3214 5628 3248
rect 5662 3214 5699 3248
rect 5733 3214 5770 3248
rect 5804 3216 5872 3248
rect 5804 3214 5838 3216
rect 5276 3147 5310 3182
rect 4000 3078 4034 3113
rect 4000 3009 4034 3044
rect 5838 3147 5872 3182
rect 5276 3078 5310 3113
rect 5447 3098 5493 3132
rect 5527 3098 5573 3132
rect 7032 3311 7066 3336
rect 7032 3243 7066 3277
rect 7032 3175 7066 3209
rect 7032 3125 7066 3141
rect 7114 3354 7148 3378
rect 7114 3285 7148 3320
rect 7114 3216 7148 3251
rect 7114 3147 7148 3182
rect 5838 3078 5872 3113
rect 4000 2940 4034 2975
rect 4000 2871 4034 2906
rect 4000 2802 4034 2837
rect 4000 2733 4034 2768
rect 4000 2664 4034 2699
rect 4000 2595 4034 2630
rect 4000 2526 4034 2561
rect 4000 2457 4034 2492
rect 4000 2388 4034 2423
rect 4000 2319 4034 2354
rect 4000 2250 4034 2285
rect 4000 2181 4034 2216
rect 1117 2153 1287 2163
rect 1151 2141 1287 2153
rect 1151 2119 1185 2141
rect 1117 2101 1185 2119
rect 1219 2128 1287 2141
rect 1219 2101 1253 2128
rect 1117 2094 1253 2101
rect 1117 2084 1287 2094
rect 1151 2069 1287 2084
rect 1151 2050 1185 2069
rect 1117 2033 1185 2050
rect 1219 2059 1287 2069
rect 4000 2112 4034 2147
rect 1219 2033 1253 2059
rect 1117 2025 1253 2033
rect 1117 2015 1287 2025
rect 1151 1999 1287 2015
rect 1151 1981 1185 1999
rect 1117 1963 1185 1981
rect 1219 1990 1287 1999
rect 1219 1963 1253 1990
rect 1117 1956 1253 1963
rect 1117 1946 1287 1956
rect 1151 1931 1287 1946
rect 1151 1912 1185 1931
rect 1117 1891 1185 1912
rect 1219 1921 1287 1931
rect 1219 1891 1253 1921
rect 1117 1887 1253 1891
rect 3767 2026 3773 2060
rect 3807 2026 3845 2060
rect 3879 2026 3885 2060
rect 3767 1985 3885 2026
rect 3767 1951 3773 1985
rect 3807 1951 3845 1985
rect 3879 1951 3885 1985
rect 3767 1920 3885 1951
rect 4000 2043 4034 2078
rect 4000 1974 4034 2009
rect 4000 1920 4034 1940
rect 1117 1877 1287 1887
rect 1468 1886 1492 1920
rect 1526 1886 1562 1920
rect 1596 1886 1632 1920
rect 1666 1886 1702 1920
rect 1736 1886 1772 1920
rect 1806 1886 1842 1920
rect 1876 1886 1912 1920
rect 1946 1886 1982 1920
rect 2016 1886 2052 1920
rect 2086 1886 2122 1920
rect 2156 1886 2192 1920
rect 2226 1886 2262 1920
rect 2296 1886 2332 1920
rect 2366 1886 2402 1920
rect 2436 1886 2472 1920
rect 2506 1886 2542 1920
rect 2576 1886 2611 1920
rect 2645 1886 2680 1920
rect 2714 1886 2749 1920
rect 2783 1886 2818 1920
rect 2852 1886 2887 1920
rect 2921 1886 2956 1920
rect 2990 1886 3025 1920
rect 3059 1886 3094 1920
rect 3128 1886 3163 1920
rect 3197 1886 3232 1920
rect 3266 1886 3301 1920
rect 3335 1886 3370 1920
rect 3404 1886 3439 1920
rect 3473 1886 3508 1920
rect 3542 1910 4034 1920
rect 3542 1896 3773 1910
rect 3807 1896 3845 1910
rect 3879 1904 4034 1910
rect 3879 1896 4000 1904
rect 3542 1886 3709 1896
rect 1151 1863 1287 1877
rect 1151 1843 1185 1863
rect 1117 1819 1185 1843
rect 1219 1852 1287 1863
rect 1219 1819 1253 1852
rect 1117 1818 1253 1819
rect 1117 1808 1287 1818
rect 1151 1795 1287 1808
rect 1151 1774 1185 1795
rect 1219 1783 1287 1795
rect 1117 1747 1185 1774
rect 1219 1749 1253 1783
rect 3646 1862 3709 1886
rect 3743 1876 3773 1896
rect 3743 1862 3777 1876
rect 3811 1862 3845 1896
rect 3879 1862 3913 1896
rect 3947 1870 4000 1896
rect 3947 1862 4034 1870
rect 3646 1852 4034 1862
rect 3612 1835 4034 1852
rect 3612 1827 3773 1835
rect 3807 1827 3845 1835
rect 3879 1834 4034 1835
rect 3879 1827 4000 1834
rect 3612 1816 3709 1827
rect 3646 1793 3709 1816
rect 3743 1801 3773 1827
rect 3743 1793 3777 1801
rect 3811 1793 3845 1827
rect 3879 1793 3913 1827
rect 3947 1800 4000 1827
rect 3947 1793 4034 1800
rect 3646 1782 4034 1793
rect 3612 1764 4034 1782
rect 3612 1760 4000 1764
rect 1219 1747 1287 1749
rect 1117 1739 1287 1747
rect 1151 1727 1287 1739
rect 1151 1705 1185 1727
rect 1219 1714 1287 1727
rect 1117 1675 1185 1705
rect 1219 1680 1253 1714
rect 1219 1675 1287 1680
rect 1117 1670 1287 1675
rect 1151 1659 1287 1670
rect 1151 1636 1185 1659
rect 1219 1645 1287 1659
rect 1117 1603 1185 1636
rect 1219 1611 1253 1645
rect 1219 1603 1287 1611
rect 1117 1601 1287 1603
rect 1151 1591 1287 1601
rect 1151 1567 1185 1591
rect 1117 1532 1185 1567
rect 1219 1576 1287 1591
rect 1151 1531 1185 1532
rect 1219 1542 1253 1576
rect 1219 1531 1287 1542
rect 1151 1523 1287 1531
rect 1151 1498 1185 1523
rect 1117 1463 1185 1498
rect 1219 1507 1287 1523
rect 1151 1459 1185 1463
rect 1219 1473 1253 1507
rect 1219 1459 1287 1473
rect 1151 1455 1287 1459
rect 1151 1429 1185 1455
rect 1117 1394 1185 1429
rect 1219 1438 1287 1455
rect 1151 1360 1185 1394
rect 1219 1404 1253 1438
rect 1117 1353 1185 1360
rect 1219 1369 1287 1404
rect 1219 1353 1253 1369
rect 1117 1349 1253 1353
rect 1117 1325 1185 1349
rect 1151 1291 1185 1325
rect 1219 1335 1253 1349
rect 1117 1285 1185 1291
rect 1219 1300 1287 1335
rect 1219 1285 1253 1300
rect 1117 1277 1253 1285
rect 1117 1256 1185 1277
rect 1151 1222 1185 1256
rect 1219 1266 1253 1277
rect 1117 1217 1185 1222
rect 1219 1231 1287 1266
rect 1219 1217 1253 1231
rect 1117 1205 1253 1217
rect 1117 1187 1185 1205
rect 1151 1153 1185 1187
rect 1219 1197 1253 1205
rect 1117 1149 1185 1153
rect 1219 1162 1287 1197
rect 1219 1149 1253 1162
rect 1117 1133 1253 1149
rect 1117 1118 1185 1133
rect 1151 1084 1185 1118
rect 1219 1128 1253 1133
rect 1117 1081 1185 1084
rect 1219 1093 1287 1128
rect 1219 1081 1253 1093
rect 1117 1061 1253 1081
rect 1117 1049 1185 1061
rect 1151 1015 1185 1049
rect 1219 1059 1253 1061
rect 1117 1013 1185 1015
rect 1219 1024 1287 1059
rect 1219 1013 1253 1024
rect 1117 990 1253 1013
rect 1117 989 1287 990
rect 1117 980 1185 989
rect 1151 946 1185 980
rect 1219 955 1287 989
rect 1396 1747 1430 1759
rect 3506 1747 3540 1759
rect 1430 1709 3506 1736
rect 1396 1673 3540 1709
rect 1430 1636 3506 1673
rect 1396 1599 3540 1636
rect 1430 1563 3506 1599
rect 1396 1525 3540 1563
rect 1430 1490 3506 1525
rect 1396 1451 3540 1490
rect 1430 1417 3506 1451
rect 1396 1378 3540 1417
rect 1430 1343 3506 1378
rect 1396 1305 3540 1343
rect 1430 1269 3506 1305
rect 1396 1231 3540 1269
rect 1430 1195 3506 1231
rect 1396 1157 3540 1195
rect 1430 1121 3506 1157
rect 1396 1083 3540 1121
rect 1430 1046 3506 1083
rect 1396 1009 3540 1046
rect 1430 982 3506 1009
rect 1396 959 1430 971
rect 3506 959 3540 971
rect 3612 1758 3773 1760
rect 3807 1758 3845 1760
rect 3879 1758 4000 1760
rect 3612 1746 3709 1758
rect 3646 1724 3709 1746
rect 3743 1726 3773 1758
rect 3743 1724 3777 1726
rect 3811 1724 3845 1758
rect 3879 1724 3913 1758
rect 3947 1730 4000 1758
rect 3947 1724 4034 1730
rect 3646 1712 4034 1724
rect 3612 1694 4034 1712
rect 3612 1689 4000 1694
rect 3612 1676 3709 1689
rect 3646 1655 3709 1676
rect 3743 1685 3777 1689
rect 3743 1655 3773 1685
rect 3811 1655 3845 1689
rect 3879 1655 3913 1689
rect 3947 1660 4000 1689
rect 3947 1655 4034 1660
rect 3646 1651 3773 1655
rect 3807 1651 3845 1655
rect 3879 1651 4034 1655
rect 3646 1642 4034 1651
rect 3612 1624 4034 1642
rect 3612 1620 4000 1624
rect 3612 1606 3709 1620
rect 3646 1586 3709 1606
rect 3743 1610 3777 1620
rect 3743 1586 3773 1610
rect 3811 1586 3845 1620
rect 3879 1586 3913 1620
rect 3947 1590 4000 1620
rect 3947 1586 4034 1590
rect 3646 1576 3773 1586
rect 3807 1576 3845 1586
rect 3879 1576 4034 1586
rect 3646 1572 4034 1576
rect 3612 1554 4034 1572
rect 3612 1551 4000 1554
rect 3612 1536 3709 1551
rect 3646 1517 3709 1536
rect 3743 1535 3777 1551
rect 3743 1517 3773 1535
rect 3811 1517 3845 1551
rect 3879 1517 3913 1551
rect 3947 1520 4000 1551
rect 3947 1517 4034 1520
rect 3646 1502 3773 1517
rect 3612 1501 3773 1502
rect 3807 1501 3845 1517
rect 3879 1501 4034 1517
rect 3612 1484 4034 1501
rect 3612 1482 4000 1484
rect 3612 1466 3709 1482
rect 3646 1448 3709 1466
rect 3743 1460 3777 1482
rect 3743 1448 3773 1460
rect 3811 1448 3845 1482
rect 3879 1448 3913 1482
rect 3947 1450 4000 1482
rect 3947 1448 4034 1450
rect 3646 1432 3773 1448
rect 3612 1426 3773 1432
rect 3807 1426 3845 1448
rect 3879 1426 4034 1448
rect 3612 1414 4034 1426
rect 3612 1413 4000 1414
rect 3612 1396 3709 1413
rect 3646 1379 3709 1396
rect 3743 1385 3777 1413
rect 3743 1379 3773 1385
rect 3811 1379 3845 1413
rect 3879 1379 3913 1413
rect 3947 1380 4000 1413
rect 3947 1379 4034 1380
rect 3646 1362 3773 1379
rect 3612 1351 3773 1362
rect 3807 1351 3845 1379
rect 3879 1351 4034 1379
rect 3612 1344 4034 1351
rect 3612 1326 3709 1344
rect 3646 1310 3709 1326
rect 3743 1310 3777 1344
rect 3811 1310 3845 1344
rect 3879 1310 3913 1344
rect 3947 1310 4000 1344
rect 3646 1292 3773 1310
rect 3612 1276 3773 1292
rect 3807 1276 3845 1310
rect 3879 1276 4034 1310
rect 3612 1274 4034 1276
rect 3612 1257 3709 1274
rect 3646 1240 3709 1257
rect 3743 1240 3777 1274
rect 3811 1240 3845 1274
rect 3879 1240 3913 1274
rect 3947 1240 4000 1274
rect 3646 1235 4034 1240
rect 3646 1223 3773 1235
rect 3612 1204 3773 1223
rect 3807 1204 3845 1235
rect 3879 1204 4034 1235
rect 3612 1188 3709 1204
rect 3646 1170 3709 1188
rect 3743 1201 3773 1204
rect 3743 1170 3777 1201
rect 3811 1170 3845 1204
rect 3879 1170 3913 1204
rect 3947 1170 4000 1204
rect 3646 1160 4034 1170
rect 3646 1154 3773 1160
rect 3612 1134 3773 1154
rect 3807 1134 3845 1160
rect 3879 1134 4034 1160
rect 3612 1119 3709 1134
rect 3646 1100 3709 1119
rect 3743 1126 3773 1134
rect 3743 1100 3777 1126
rect 3811 1100 3845 1134
rect 3879 1100 3913 1134
rect 3947 1100 4000 1134
rect 5194 2964 5228 2986
rect 5194 2892 5228 2918
rect 5194 2820 5228 2858
rect 5194 2764 5228 2786
rect 5194 2696 5228 2714
rect 5194 2604 5228 2642
rect 5194 2532 5228 2570
rect 5194 2459 5228 2474
rect 5194 2386 5228 2406
rect 5194 2313 5228 2352
rect 5194 2252 5228 2279
rect 5194 2184 5228 2206
rect 5194 2094 5228 2133
rect 5194 2021 5228 2060
rect 5194 1948 5228 1962
rect 5194 1875 5228 1894
rect 5194 1802 5228 1841
rect 5194 1740 5228 1768
rect 5194 1672 5228 1695
rect 5194 1583 5228 1622
rect 5194 1510 5228 1549
rect 5194 1437 5228 1450
rect 5194 1364 5228 1382
rect 5194 1291 5228 1330
rect 5194 1228 5228 1257
rect 5194 1160 5228 1184
rect 5194 1110 5228 1111
rect 5276 3009 5310 3044
rect 5276 2940 5310 2975
rect 5712 3048 5746 3064
rect 5712 2980 5746 3014
rect 5712 2930 5746 2942
rect 5838 3009 5872 3044
rect 7114 3078 7148 3113
rect 5838 2940 5872 2975
rect 5276 2871 5310 2906
rect 5587 2862 5627 2896
rect 5661 2862 5701 2896
rect 5838 2871 5872 2906
rect 5276 2802 5310 2837
rect 5276 2733 5310 2768
rect 5276 2664 5310 2699
rect 5838 2802 5872 2837
rect 5838 2733 5872 2768
rect 5838 2664 5872 2699
rect 5276 2595 5310 2630
rect 5447 2627 5493 2661
rect 5527 2627 5573 2661
rect 5276 2544 5310 2561
rect 5838 2595 5872 2630
rect 5838 2544 5872 2561
rect 5276 2526 5563 2544
rect 5310 2520 5563 2526
rect 5597 2526 5872 2544
rect 5597 2520 5838 2526
rect 5310 2492 5359 2520
rect 5276 2486 5359 2492
rect 5393 2486 5427 2520
rect 5461 2486 5495 2520
rect 5529 2486 5563 2520
rect 5597 2486 5631 2520
rect 5665 2486 5699 2520
rect 5733 2486 5767 2520
rect 5801 2492 5838 2520
rect 5801 2486 5872 2492
rect 5276 2471 5872 2486
rect 5276 2457 5563 2471
rect 5310 2451 5563 2457
rect 5597 2457 5872 2471
rect 5597 2451 5838 2457
rect 5310 2423 5359 2451
rect 5276 2417 5359 2423
rect 5393 2417 5427 2451
rect 5461 2417 5495 2451
rect 5529 2417 5563 2451
rect 5597 2417 5631 2451
rect 5665 2417 5699 2451
rect 5733 2417 5767 2451
rect 5801 2423 5838 2451
rect 5801 2417 5872 2423
rect 5276 2398 5872 2417
rect 5276 2388 5563 2398
rect 5310 2382 5563 2388
rect 5597 2388 5872 2398
rect 5597 2382 5838 2388
rect 5310 2354 5359 2382
rect 5276 2348 5359 2354
rect 5393 2348 5427 2382
rect 5461 2348 5495 2382
rect 5529 2348 5563 2382
rect 5597 2348 5631 2382
rect 5665 2348 5699 2382
rect 5733 2348 5767 2382
rect 5801 2354 5838 2382
rect 5801 2348 5872 2354
rect 5276 2325 5872 2348
rect 5276 2319 5563 2325
rect 5310 2313 5563 2319
rect 5597 2319 5872 2325
rect 5597 2313 5838 2319
rect 5310 2285 5359 2313
rect 5276 2279 5359 2285
rect 5393 2279 5427 2313
rect 5461 2279 5495 2313
rect 5529 2279 5563 2313
rect 5597 2279 5631 2313
rect 5665 2279 5699 2313
rect 5733 2279 5767 2313
rect 5801 2285 5838 2313
rect 5801 2279 5872 2285
rect 5276 2252 5872 2279
rect 5276 2250 5563 2252
rect 5310 2244 5563 2250
rect 5597 2250 5872 2252
rect 5597 2244 5838 2250
rect 5310 2216 5359 2244
rect 5276 2210 5359 2216
rect 5393 2210 5427 2244
rect 5461 2210 5495 2244
rect 5529 2210 5563 2244
rect 5597 2210 5631 2244
rect 5665 2210 5699 2244
rect 5733 2210 5767 2244
rect 5801 2216 5838 2244
rect 5801 2210 5872 2216
rect 5276 2181 5872 2210
rect 5310 2179 5838 2181
rect 5310 2175 5563 2179
rect 5597 2175 5838 2179
rect 5310 2147 5359 2175
rect 5276 2141 5359 2147
rect 5393 2141 5427 2175
rect 5461 2141 5495 2175
rect 5529 2141 5563 2175
rect 5597 2141 5631 2175
rect 5665 2141 5699 2175
rect 5733 2141 5767 2175
rect 5801 2147 5838 2175
rect 5801 2141 5872 2147
rect 5276 2112 5872 2141
rect 5310 2106 5838 2112
rect 5310 2078 5359 2106
rect 5276 2072 5359 2078
rect 5393 2072 5427 2106
rect 5461 2072 5495 2106
rect 5529 2072 5563 2106
rect 5597 2072 5631 2106
rect 5665 2072 5699 2106
rect 5733 2072 5767 2106
rect 5801 2078 5838 2106
rect 5801 2072 5872 2078
rect 5276 2043 5872 2072
rect 5310 2037 5838 2043
rect 5310 2009 5359 2037
rect 5276 2003 5359 2009
rect 5393 2003 5427 2037
rect 5461 2003 5495 2037
rect 5529 2003 5563 2037
rect 5597 2003 5631 2037
rect 5665 2003 5699 2037
rect 5733 2003 5767 2037
rect 5801 2009 5838 2037
rect 5801 2003 5872 2009
rect 5276 1999 5563 2003
rect 5597 1999 5872 2003
rect 5276 1974 5872 1999
rect 5310 1968 5838 1974
rect 5310 1940 5359 1968
rect 5276 1934 5359 1940
rect 5393 1934 5427 1968
rect 5461 1934 5495 1968
rect 5529 1934 5563 1968
rect 5597 1934 5631 1968
rect 5665 1934 5699 1968
rect 5733 1934 5767 1968
rect 5801 1940 5838 1968
rect 5801 1934 5872 1940
rect 5276 1926 5563 1934
rect 5597 1926 5872 1934
rect 5276 1905 5872 1926
rect 5310 1899 5838 1905
rect 5310 1871 5359 1899
rect 5276 1865 5359 1871
rect 5393 1865 5427 1899
rect 5461 1865 5495 1899
rect 5529 1865 5563 1899
rect 5597 1865 5631 1899
rect 5665 1865 5699 1899
rect 5733 1865 5767 1899
rect 5801 1871 5838 1899
rect 5801 1865 5872 1871
rect 5276 1853 5563 1865
rect 5597 1853 5872 1865
rect 5276 1836 5872 1853
rect 5310 1830 5838 1836
rect 5310 1802 5359 1830
rect 5276 1796 5359 1802
rect 5393 1796 5427 1830
rect 5461 1796 5495 1830
rect 5529 1796 5563 1830
rect 5597 1796 5631 1830
rect 5665 1796 5699 1830
rect 5733 1796 5767 1830
rect 5801 1802 5838 1830
rect 5801 1796 5872 1802
rect 5276 1780 5563 1796
rect 5597 1780 5872 1796
rect 5276 1766 5872 1780
rect 5310 1761 5838 1766
rect 5310 1732 5359 1761
rect 5276 1727 5359 1732
rect 5393 1727 5427 1761
rect 5461 1727 5495 1761
rect 5529 1727 5563 1761
rect 5597 1727 5631 1761
rect 5665 1727 5699 1761
rect 5733 1727 5767 1761
rect 5801 1732 5838 1761
rect 5801 1727 5872 1732
rect 5276 1706 5563 1727
rect 5597 1706 5872 1727
rect 5276 1696 5872 1706
rect 5310 1692 5838 1696
rect 5310 1662 5359 1692
rect 5276 1658 5359 1662
rect 5393 1658 5427 1692
rect 5461 1658 5495 1692
rect 5529 1658 5563 1692
rect 5597 1658 5631 1692
rect 5665 1658 5699 1692
rect 5733 1658 5767 1692
rect 5801 1662 5838 1692
rect 5801 1658 5872 1662
rect 5276 1632 5563 1658
rect 5597 1632 5872 1658
rect 5276 1626 5872 1632
rect 5310 1623 5838 1626
rect 5310 1592 5359 1623
rect 5276 1589 5359 1592
rect 5393 1589 5427 1623
rect 5461 1589 5495 1623
rect 5529 1589 5563 1623
rect 5597 1589 5631 1623
rect 5665 1589 5699 1623
rect 5733 1589 5767 1623
rect 5801 1592 5838 1623
rect 5801 1589 5872 1592
rect 5276 1558 5563 1589
rect 5597 1558 5872 1589
rect 5276 1556 5872 1558
rect 5310 1554 5838 1556
rect 5310 1522 5359 1554
rect 5276 1520 5359 1522
rect 5393 1520 5427 1554
rect 5461 1520 5495 1554
rect 5529 1520 5563 1554
rect 5597 1520 5631 1554
rect 5665 1520 5699 1554
rect 5733 1520 5767 1554
rect 5801 1522 5838 1554
rect 5801 1520 5872 1522
rect 5276 1518 5872 1520
rect 5276 1486 5563 1518
rect 5310 1485 5563 1486
rect 5597 1486 5872 1518
rect 5597 1485 5838 1486
rect 5310 1452 5359 1485
rect 5276 1451 5359 1452
rect 5393 1451 5427 1485
rect 5461 1451 5495 1485
rect 5529 1451 5563 1485
rect 5597 1451 5631 1485
rect 5665 1451 5699 1485
rect 5733 1451 5767 1485
rect 5801 1452 5838 1485
rect 5801 1451 5872 1452
rect 5276 1444 5872 1451
rect 5276 1416 5563 1444
rect 5597 1416 5872 1444
rect 5310 1382 5359 1416
rect 5393 1382 5427 1416
rect 5461 1382 5495 1416
rect 5529 1382 5563 1416
rect 5597 1382 5631 1416
rect 5665 1382 5699 1416
rect 5733 1382 5767 1416
rect 5801 1382 5838 1416
rect 5276 1370 5872 1382
rect 5276 1346 5563 1370
rect 5597 1346 5872 1370
rect 5310 1312 5359 1346
rect 5393 1312 5427 1346
rect 5461 1312 5495 1346
rect 5529 1312 5563 1346
rect 5597 1312 5631 1346
rect 5665 1312 5699 1346
rect 5733 1312 5767 1346
rect 5801 1312 5838 1346
rect 5276 1296 5872 1312
rect 5276 1276 5563 1296
rect 5597 1276 5872 1296
rect 5310 1242 5359 1276
rect 5393 1242 5427 1276
rect 5461 1242 5495 1276
rect 5529 1242 5563 1276
rect 5597 1242 5631 1276
rect 5665 1242 5699 1276
rect 5733 1242 5767 1276
rect 5801 1242 5838 1276
rect 5276 1222 5872 1242
rect 5276 1206 5563 1222
rect 5597 1206 5872 1222
rect 5310 1172 5359 1206
rect 5393 1172 5427 1206
rect 5461 1172 5495 1206
rect 5529 1172 5563 1206
rect 5597 1172 5631 1206
rect 5665 1172 5699 1206
rect 5733 1172 5767 1206
rect 5801 1172 5838 1206
rect 5276 1148 5872 1172
rect 5276 1136 5563 1148
rect 5597 1136 5872 1148
rect 3646 1085 4034 1100
rect 3612 1064 3773 1085
rect 3807 1064 3845 1085
rect 3879 1064 4034 1085
rect 3612 1050 3709 1064
rect 3646 1030 3709 1050
rect 3743 1051 3773 1064
rect 3743 1030 3777 1051
rect 3811 1030 3845 1064
rect 3879 1030 3913 1064
rect 3947 1030 4000 1064
rect 3646 1016 4034 1030
rect 5310 1102 5359 1136
rect 5393 1102 5427 1136
rect 5461 1102 5495 1136
rect 5529 1102 5563 1136
rect 5597 1102 5631 1136
rect 5665 1102 5699 1136
rect 5733 1102 5767 1136
rect 5801 1102 5838 1136
rect 7032 2964 7066 2986
rect 7032 2892 7066 2918
rect 7032 2820 7066 2858
rect 7032 2764 7066 2786
rect 7032 2696 7066 2714
rect 7032 2604 7066 2642
rect 7032 2532 7066 2570
rect 7032 2459 7066 2474
rect 7032 2386 7066 2406
rect 7032 2313 7066 2352
rect 7032 2252 7066 2279
rect 7032 2184 7066 2206
rect 7032 2094 7066 2133
rect 7032 2021 7066 2060
rect 7032 1948 7066 1962
rect 7032 1875 7066 1894
rect 7032 1802 7066 1841
rect 7032 1740 7066 1768
rect 7032 1672 7066 1695
rect 7032 1583 7066 1622
rect 7032 1510 7066 1549
rect 7032 1437 7066 1450
rect 7032 1364 7066 1382
rect 7032 1291 7066 1330
rect 7032 1228 7066 1257
rect 7032 1160 7066 1184
rect 7032 1110 7066 1111
rect 7114 3009 7148 3044
rect 7114 2940 7148 2975
rect 7114 2871 7148 2906
rect 7114 2802 7148 2837
rect 7114 2733 7148 2768
rect 7114 2664 7148 2699
rect 7114 2595 7148 2630
rect 7114 2526 7148 2561
rect 7114 2457 7148 2492
rect 7114 2388 7148 2423
rect 7114 2319 7148 2354
rect 7114 2250 7148 2285
rect 7114 2181 7148 2216
rect 7397 3367 7457 3393
rect 7397 3359 7423 3367
rect 7431 3325 7457 3333
rect 7397 3295 7457 3325
rect 7397 3291 7423 3295
rect 7431 3257 7457 3261
rect 7397 3223 7457 3257
rect 7397 3155 7457 3189
rect 7431 3151 7457 3155
rect 7397 3117 7423 3121
rect 7397 3087 7457 3117
rect 7431 3079 7457 3087
rect 7397 3045 7423 3053
rect 7397 3019 7457 3045
rect 7431 3007 7457 3019
rect 7397 2973 7423 2985
rect 7397 2951 7457 2973
rect 7431 2935 7457 2951
rect 7397 2901 7423 2917
rect 7397 2883 7457 2901
rect 7431 2863 7457 2883
rect 7397 2829 7423 2849
rect 7397 2815 7457 2829
rect 7431 2791 7457 2815
rect 7397 2757 7423 2781
rect 7397 2747 7457 2757
rect 7431 2719 7457 2747
rect 7397 2685 7423 2713
rect 7397 2679 7457 2685
rect 7431 2647 7457 2679
rect 7608 3440 7642 3452
rect 9718 3440 9752 3452
rect 7642 3402 9718 3429
rect 7608 3366 9752 3402
rect 7642 3329 9718 3366
rect 7608 3292 9752 3329
rect 7642 3256 9718 3292
rect 7608 3218 9752 3256
rect 7642 3183 9718 3218
rect 7608 3144 9752 3183
rect 7642 3110 9718 3144
rect 7608 3071 9752 3110
rect 7642 3036 9718 3071
rect 7608 2998 9752 3036
rect 7642 2962 9718 2998
rect 7608 2924 9752 2962
rect 7642 2888 9718 2924
rect 7608 2850 9752 2888
rect 7642 2814 9718 2850
rect 7608 2776 9752 2814
rect 7642 2739 9718 2776
rect 7608 2702 9752 2739
rect 7642 2675 9718 2702
rect 7608 2652 7642 2664
rect 9718 2652 9752 2664
rect 9933 3428 9963 3461
rect 9899 3427 9963 3428
rect 9899 3393 9929 3427
rect 9899 3390 9963 3393
rect 9933 3359 9963 3390
rect 9899 3325 9929 3356
rect 9899 3318 9963 3325
rect 9933 3291 9963 3318
rect 9899 3257 9929 3284
rect 9899 3246 9963 3257
rect 9933 3223 9963 3246
rect 9899 3189 9929 3212
rect 9899 3174 9963 3189
rect 9933 3155 9963 3174
rect 9899 3121 9929 3140
rect 9899 3102 9963 3121
rect 9933 3087 9963 3102
rect 9899 3053 9929 3068
rect 9899 3030 9963 3053
rect 9933 3019 9963 3030
rect 9899 2985 9929 2996
rect 9899 2958 9963 2985
rect 9933 2951 9963 2958
rect 9899 2917 9929 2924
rect 9899 2886 9963 2917
rect 9933 2883 9963 2886
rect 9899 2849 9929 2852
rect 9899 2815 9963 2849
rect 9899 2814 9929 2815
rect 9933 2780 9963 2781
rect 9899 2747 9963 2780
rect 9899 2742 9929 2747
rect 9933 2708 9963 2713
rect 9899 2679 9963 2708
rect 9899 2670 9929 2679
rect 7397 2613 7423 2645
rect 7397 2611 7457 2613
rect 7431 2577 7457 2611
rect 7397 2575 7457 2577
rect 7397 2543 7423 2575
rect 7431 2509 7457 2541
rect 7397 2503 7457 2509
rect 7702 2505 8151 2539
rect 7397 2475 7423 2503
rect 7680 2471 8151 2505
rect 7431 2441 7457 2469
rect 8761 2607 8800 2641
rect 8834 2607 8873 2641
rect 8907 2607 8946 2641
rect 8980 2607 9019 2641
rect 9053 2607 9092 2641
rect 9933 2636 9963 2645
rect 9899 2611 9963 2636
rect 9899 2598 9929 2611
rect 8761 2535 8800 2569
rect 8834 2535 8873 2569
rect 8907 2535 8946 2569
rect 8980 2535 9019 2569
rect 9053 2535 9092 2569
rect 9933 2564 9963 2577
rect 9899 2543 9963 2564
rect 9126 2535 9684 2539
rect 8761 2497 9684 2535
rect 8761 2463 8800 2497
rect 8834 2463 8873 2497
rect 8907 2463 8946 2497
rect 8980 2463 9019 2497
rect 9053 2463 9092 2497
rect 9126 2471 9684 2497
rect 9899 2526 9929 2543
rect 9933 2492 9963 2509
rect 9899 2475 9963 2492
rect 7397 2431 7457 2441
rect 7397 2407 7423 2431
rect 7431 2373 7457 2397
rect 7397 2359 7457 2373
rect 7397 2339 7423 2359
rect 7431 2305 7457 2325
rect 7397 2287 7457 2305
rect 7397 2271 7423 2287
rect 7431 2237 7457 2253
rect 7397 2215 7457 2237
rect 7397 2181 7423 2215
rect 9899 2454 9929 2475
rect 9933 2420 9963 2441
rect 9899 2407 9963 2420
rect 9899 2382 9929 2407
rect 9933 2348 9963 2373
rect 9899 2339 9963 2348
rect 9899 2310 9929 2339
rect 9933 2276 9963 2305
rect 9899 2271 9963 2276
rect 9899 2238 9929 2271
rect 9933 2204 9963 2237
rect 9899 2203 9963 2204
rect 7397 2169 7431 2181
rect 7465 2169 7499 2203
rect 7533 2169 7567 2203
rect 7601 2169 7635 2203
rect 7669 2169 7703 2203
rect 7737 2169 7771 2203
rect 7805 2169 7839 2203
rect 7873 2169 7907 2203
rect 7941 2169 7975 2203
rect 8009 2169 8043 2203
rect 8077 2169 8111 2203
rect 8145 2169 8179 2203
rect 8213 2169 8247 2203
rect 8281 2169 8315 2203
rect 8349 2169 8383 2203
rect 8417 2169 8451 2203
rect 8485 2169 8519 2203
rect 8553 2169 8587 2203
rect 8621 2169 8655 2203
rect 8689 2169 8723 2203
rect 8757 2169 8791 2203
rect 8825 2169 8859 2203
rect 8893 2169 8927 2203
rect 8961 2169 8995 2203
rect 9029 2169 9063 2203
rect 9097 2169 9131 2203
rect 9165 2169 9199 2203
rect 9233 2169 9267 2203
rect 9301 2169 9335 2203
rect 9369 2169 9403 2203
rect 9437 2169 9471 2203
rect 9505 2169 9539 2203
rect 9573 2169 9607 2203
rect 9641 2169 9675 2203
rect 9709 2169 9743 2203
rect 9777 2169 9811 2203
rect 9845 2169 9929 2203
rect 7114 2112 7148 2147
rect 7114 2043 7148 2078
rect 9899 2166 9963 2169
rect 9933 2135 9963 2166
rect 9899 2101 9929 2132
rect 9899 2094 9963 2101
rect 9933 2067 9963 2094
rect 7114 1974 7148 2009
rect 7114 1920 7148 1940
rect 7265 2026 7271 2060
rect 7305 2026 7343 2060
rect 7377 2026 7383 2060
rect 7265 1985 7383 2026
rect 7265 1951 7271 1985
rect 7305 1951 7343 1985
rect 7377 1951 7383 1985
rect 7265 1920 7383 1951
rect 9899 2033 9929 2060
rect 9899 2022 9963 2033
rect 9933 1999 9963 2022
rect 9899 1965 9929 1988
rect 9899 1950 9963 1965
rect 9933 1931 9963 1950
rect 7114 1910 7606 1920
rect 7114 1904 7271 1910
rect 7148 1896 7271 1904
rect 7305 1896 7343 1910
rect 7377 1896 7606 1910
rect 7148 1870 7207 1896
rect 7114 1862 7207 1870
rect 7241 1876 7271 1896
rect 7241 1862 7275 1876
rect 7309 1862 7343 1896
rect 7377 1862 7411 1896
rect 7445 1886 7606 1896
rect 7640 1886 7675 1920
rect 7709 1886 7744 1920
rect 7778 1886 7813 1920
rect 7847 1886 7882 1920
rect 7916 1886 7951 1920
rect 7985 1886 8020 1920
rect 8054 1886 8089 1920
rect 8123 1886 8158 1920
rect 8192 1886 8227 1920
rect 8261 1886 8296 1920
rect 8330 1886 8365 1920
rect 8399 1886 8434 1920
rect 8468 1886 8503 1920
rect 8537 1886 8572 1920
rect 8606 1886 8642 1920
rect 8676 1886 8712 1920
rect 8746 1886 8782 1920
rect 8816 1886 8852 1920
rect 8886 1886 8922 1920
rect 8956 1886 8992 1920
rect 9026 1886 9062 1920
rect 9096 1886 9132 1920
rect 9166 1886 9202 1920
rect 9236 1886 9272 1920
rect 9306 1886 9342 1920
rect 9376 1886 9412 1920
rect 9446 1886 9482 1920
rect 9516 1886 9552 1920
rect 9586 1886 9622 1920
rect 9656 1886 9680 1920
rect 9899 1897 9929 1916
rect 7445 1862 7502 1886
rect 7114 1852 7502 1862
rect 7114 1835 7536 1852
rect 7114 1834 7271 1835
rect 7148 1827 7271 1834
rect 7305 1827 7343 1835
rect 7377 1827 7536 1835
rect 7148 1800 7207 1827
rect 7114 1793 7207 1800
rect 7241 1801 7271 1827
rect 7241 1793 7275 1801
rect 7309 1793 7343 1827
rect 7377 1793 7411 1827
rect 7445 1816 7536 1827
rect 7445 1793 7502 1816
rect 7114 1782 7502 1793
rect 7114 1764 7536 1782
rect 7148 1760 7536 1764
rect 7148 1758 7271 1760
rect 7305 1758 7343 1760
rect 7377 1758 7536 1760
rect 9899 1878 9963 1897
rect 9933 1863 9963 1878
rect 9899 1829 9929 1844
rect 9899 1806 9963 1829
rect 9933 1795 9963 1806
rect 9899 1761 9929 1772
rect 7148 1730 7207 1758
rect 7114 1724 7207 1730
rect 7241 1726 7271 1758
rect 7241 1724 7275 1726
rect 7309 1724 7343 1758
rect 7377 1724 7411 1758
rect 7445 1746 7536 1758
rect 7445 1724 7502 1746
rect 7114 1712 7502 1724
rect 7114 1694 7536 1712
rect 7148 1689 7536 1694
rect 7148 1660 7207 1689
rect 7114 1655 7207 1660
rect 7241 1685 7275 1689
rect 7241 1655 7271 1685
rect 7309 1655 7343 1689
rect 7377 1655 7411 1689
rect 7445 1676 7536 1689
rect 7445 1655 7502 1676
rect 7114 1651 7271 1655
rect 7305 1651 7343 1655
rect 7377 1651 7502 1655
rect 7114 1642 7502 1651
rect 7114 1624 7536 1642
rect 7148 1620 7536 1624
rect 7148 1590 7207 1620
rect 7114 1586 7207 1590
rect 7241 1610 7275 1620
rect 7241 1586 7271 1610
rect 7309 1586 7343 1620
rect 7377 1586 7411 1620
rect 7445 1606 7536 1620
rect 7445 1586 7502 1606
rect 7114 1576 7271 1586
rect 7305 1576 7343 1586
rect 7377 1576 7502 1586
rect 7114 1572 7502 1576
rect 7114 1554 7536 1572
rect 7148 1551 7536 1554
rect 7148 1520 7207 1551
rect 7114 1517 7207 1520
rect 7241 1535 7275 1551
rect 7241 1517 7271 1535
rect 7309 1517 7343 1551
rect 7377 1517 7411 1551
rect 7445 1536 7536 1551
rect 7445 1517 7502 1536
rect 7114 1501 7271 1517
rect 7305 1501 7343 1517
rect 7377 1502 7502 1517
rect 7377 1501 7536 1502
rect 7114 1484 7536 1501
rect 7148 1482 7536 1484
rect 7148 1450 7207 1482
rect 7114 1448 7207 1450
rect 7241 1460 7275 1482
rect 7241 1448 7271 1460
rect 7309 1448 7343 1482
rect 7377 1448 7411 1482
rect 7445 1466 7536 1482
rect 7445 1448 7502 1466
rect 7114 1426 7271 1448
rect 7305 1426 7343 1448
rect 7377 1432 7502 1448
rect 7377 1426 7536 1432
rect 7114 1414 7536 1426
rect 7148 1413 7536 1414
rect 7148 1380 7207 1413
rect 7114 1379 7207 1380
rect 7241 1385 7275 1413
rect 7241 1379 7271 1385
rect 7309 1379 7343 1413
rect 7377 1379 7411 1413
rect 7445 1396 7536 1413
rect 7445 1379 7502 1396
rect 7114 1351 7271 1379
rect 7305 1351 7343 1379
rect 7377 1362 7502 1379
rect 7377 1351 7536 1362
rect 7114 1344 7536 1351
rect 7148 1310 7207 1344
rect 7241 1310 7275 1344
rect 7309 1310 7343 1344
rect 7377 1310 7411 1344
rect 7445 1326 7536 1344
rect 7445 1310 7502 1326
rect 7114 1276 7271 1310
rect 7305 1276 7343 1310
rect 7377 1292 7502 1310
rect 7377 1276 7536 1292
rect 7114 1274 7536 1276
rect 7148 1240 7207 1274
rect 7241 1240 7275 1274
rect 7309 1240 7343 1274
rect 7377 1240 7411 1274
rect 7445 1257 7536 1274
rect 7445 1240 7502 1257
rect 7114 1235 7502 1240
rect 7114 1204 7271 1235
rect 7305 1204 7343 1235
rect 7377 1223 7502 1235
rect 7377 1204 7536 1223
rect 7148 1170 7207 1204
rect 7241 1201 7271 1204
rect 7241 1170 7275 1201
rect 7309 1170 7343 1204
rect 7377 1170 7411 1204
rect 7445 1188 7536 1204
rect 7445 1170 7502 1188
rect 7114 1160 7502 1170
rect 7114 1134 7271 1160
rect 7305 1134 7343 1160
rect 7377 1154 7502 1160
rect 7377 1134 7536 1154
rect 5276 1074 5872 1102
rect 5276 1066 5563 1074
rect 5597 1066 5872 1074
rect 5310 1032 5359 1066
rect 5393 1032 5427 1066
rect 5461 1032 5495 1066
rect 5529 1032 5563 1066
rect 5597 1032 5631 1066
rect 5665 1032 5699 1066
rect 5733 1032 5767 1066
rect 5801 1032 5838 1066
rect 3612 1010 4034 1016
rect 3612 994 3773 1010
rect 3807 994 3845 1010
rect 3879 994 4034 1010
rect 3612 981 3709 994
rect 1117 945 1185 946
rect 1219 945 1253 955
rect 1117 921 1253 945
rect 1117 917 1287 921
rect 1117 911 1185 917
rect 1151 877 1185 911
rect 1219 886 1287 917
rect 1219 877 1253 886
rect 1117 852 1253 877
rect 3646 960 3709 981
rect 3743 976 3773 994
rect 3743 960 3777 976
rect 3811 960 3845 994
rect 3879 960 3913 994
rect 3947 960 4000 994
rect 3646 947 4034 960
rect 3612 935 4034 947
rect 3612 924 3773 935
rect 3807 924 3845 935
rect 3879 924 4034 935
rect 3612 912 3709 924
rect 3646 890 3709 912
rect 3743 901 3773 924
rect 3743 890 3777 901
rect 3811 890 3845 924
rect 3879 890 3913 924
rect 3947 890 4000 924
rect 5194 1005 5228 1021
rect 5194 937 5228 971
rect 3646 878 4034 890
rect 1117 845 1287 852
rect 1117 842 1185 845
rect 1151 809 1185 842
rect 1219 817 1287 845
rect 1219 809 1253 817
rect 1151 808 1253 809
rect 1117 783 1253 808
rect 1583 792 1599 826
rect 1658 792 1716 826
rect 1767 792 1783 826
rect 3506 800 3540 829
rect 3612 860 4034 878
rect 5100 903 5194 910
rect 5100 876 5228 903
rect 5276 1000 5872 1032
rect 7148 1100 7207 1134
rect 7241 1126 7271 1134
rect 7241 1100 7275 1126
rect 7309 1100 7343 1134
rect 7377 1100 7411 1134
rect 7445 1119 7536 1134
rect 7445 1100 7502 1119
rect 7114 1085 7502 1100
rect 7114 1064 7271 1085
rect 7305 1064 7343 1085
rect 7377 1064 7536 1085
rect 7148 1030 7207 1064
rect 7241 1051 7271 1064
rect 7241 1030 7275 1051
rect 7309 1030 7343 1064
rect 7377 1030 7411 1064
rect 7445 1050 7536 1064
rect 7445 1030 7502 1050
rect 5276 996 5563 1000
rect 5597 996 5872 1000
rect 5310 962 5359 996
rect 5393 962 5427 996
rect 5461 962 5495 996
rect 5529 962 5563 996
rect 5597 962 5631 996
rect 5665 962 5699 996
rect 5733 962 5767 996
rect 5801 962 5838 996
rect 5276 926 5872 962
rect 5310 892 5359 926
rect 5393 892 5427 926
rect 5461 892 5495 926
rect 5529 892 5563 926
rect 5597 892 5631 926
rect 5665 892 5699 926
rect 5733 892 5767 926
rect 5801 892 5838 926
rect 7032 1005 7066 1021
rect 7032 937 7066 971
rect 3612 854 3773 860
rect 3807 854 3845 860
rect 3879 854 4034 860
rect 3612 843 3709 854
rect 3646 820 3709 843
rect 3743 826 3773 854
rect 3743 820 3777 826
rect 3811 820 3845 854
rect 3879 820 3913 854
rect 3947 820 4000 854
rect 3646 809 4034 820
rect 1117 775 1287 783
rect 1117 773 1185 775
rect 1151 739 1185 773
rect 1219 748 1287 775
rect 1892 766 1908 800
rect 1942 766 1976 800
rect 2010 766 2026 800
rect 2094 766 2154 800
rect 2188 766 2222 800
rect 2256 766 2410 800
rect 2444 766 2478 800
rect 2512 766 2666 800
rect 2700 766 2734 800
rect 2768 766 2922 800
rect 2956 766 2990 800
rect 3024 766 3175 800
rect 3212 766 3246 800
rect 3281 766 3296 800
rect 3408 766 3424 800
rect 3458 766 3492 800
rect 3526 791 3542 800
rect 3540 766 3542 791
rect 3612 785 4034 809
rect 3612 784 3773 785
rect 3807 784 3845 785
rect 3879 784 4034 785
rect 3612 774 3709 784
rect 1219 739 1253 748
rect 1117 714 1253 739
rect 1117 707 1287 714
rect 1117 704 1185 707
rect 1151 670 1185 704
rect 1219 679 1287 707
rect 1117 667 1185 670
rect 1219 667 1253 679
rect 1117 645 1253 667
rect 1117 639 1287 645
rect 1117 635 1185 639
rect 1151 601 1185 635
rect 1219 610 1287 639
rect 1117 595 1185 601
rect 1219 595 1253 610
rect 1117 576 1253 595
rect 1117 571 1287 576
rect 1117 566 1185 571
rect 1151 532 1185 566
rect 1219 541 1287 571
rect 1904 708 1938 766
rect 1538 654 1572 692
rect 1538 582 1572 620
rect 1794 636 1828 674
rect 1794 564 1828 602
rect 1117 523 1185 532
rect 1219 523 1253 541
rect 1117 507 1253 523
rect 1904 636 1938 674
rect 2060 728 2094 766
rect 3646 750 3709 774
rect 3743 751 3773 784
rect 3743 750 3777 751
rect 3811 750 3845 784
rect 3879 750 3913 784
rect 3947 750 4000 784
rect 3646 740 4034 750
rect 2060 656 2094 694
rect 2316 636 2350 674
rect 1904 564 1938 602
rect 2316 564 2350 602
rect 2572 658 2606 696
rect 2572 586 2606 624
rect 2828 636 2862 674
rect 2828 564 2862 602
rect 3612 714 4034 740
rect 5276 856 5872 892
rect 6940 903 7032 910
rect 6940 876 7066 903
rect 7114 1016 7502 1030
rect 7114 1010 7536 1016
rect 7114 994 7271 1010
rect 7305 994 7343 1010
rect 7377 994 7536 1010
rect 7148 960 7207 994
rect 7241 976 7271 994
rect 7241 960 7275 976
rect 7309 960 7343 994
rect 7377 960 7411 994
rect 7445 981 7536 994
rect 7445 960 7502 981
rect 7114 947 7502 960
rect 7608 1747 7642 1759
rect 9718 1747 9752 1759
rect 7642 1709 9718 1736
rect 7608 1673 9752 1709
rect 7642 1636 9718 1673
rect 7608 1599 9752 1636
rect 7642 1563 9718 1599
rect 7608 1525 9752 1563
rect 7642 1490 9718 1525
rect 7608 1451 9752 1490
rect 7642 1417 9718 1451
rect 7608 1378 9752 1417
rect 7642 1343 9718 1378
rect 7608 1305 9752 1343
rect 7642 1269 9718 1305
rect 7608 1231 9752 1269
rect 7642 1195 9718 1231
rect 7608 1157 9752 1195
rect 7642 1121 9718 1157
rect 7608 1083 9752 1121
rect 7642 1046 9718 1083
rect 7608 1009 9752 1046
rect 7642 982 9718 1009
rect 7608 959 7642 971
rect 9718 959 9752 971
rect 9899 1734 9963 1761
rect 9933 1727 9963 1734
rect 9899 1693 9929 1700
rect 9899 1662 9963 1693
rect 9933 1659 9963 1662
rect 9899 1625 9929 1628
rect 9899 1591 9963 1625
rect 9899 1590 9929 1591
rect 9933 1556 9963 1557
rect 9899 1523 9963 1556
rect 9899 1518 9929 1523
rect 9933 1484 9963 1489
rect 9899 1455 9963 1484
rect 9899 1446 9929 1455
rect 9933 1412 9963 1421
rect 9899 1387 9963 1412
rect 9899 1374 9929 1387
rect 9933 1340 9963 1353
rect 9899 1319 9963 1340
rect 9899 1302 9929 1319
rect 9933 1268 9963 1285
rect 9899 1251 9963 1268
rect 9899 1230 9929 1251
rect 9933 1196 9963 1217
rect 9899 1183 9963 1196
rect 9899 1158 9929 1183
rect 9933 1124 9963 1149
rect 9899 1115 9963 1124
rect 9899 1086 9929 1115
rect 9933 1052 9963 1081
rect 9899 1047 9963 1052
rect 9899 1014 9929 1047
rect 9933 980 9963 1013
rect 9899 979 9963 980
rect 7114 935 7536 947
rect 7114 924 7271 935
rect 7305 924 7343 935
rect 7377 924 7536 935
rect 7148 890 7207 924
rect 7241 901 7271 924
rect 7241 890 7275 901
rect 7309 890 7343 924
rect 7377 890 7411 924
rect 7445 912 7536 924
rect 7445 890 7502 912
rect 7114 878 7502 890
rect 5310 822 5359 856
rect 5393 822 5427 856
rect 5461 822 5495 856
rect 5529 822 5563 856
rect 5597 822 5631 856
rect 5665 822 5699 856
rect 5733 822 5767 856
rect 5801 822 5838 856
rect 5276 818 5563 822
rect 5597 818 5872 822
rect 5276 786 5872 818
rect 5310 752 5359 786
rect 5393 752 5427 786
rect 5461 752 5495 786
rect 5529 752 5563 786
rect 5597 752 5631 786
rect 5665 752 5699 786
rect 5733 752 5767 786
rect 5801 752 5838 786
rect 5276 744 5563 752
rect 5597 744 5872 752
rect 3612 705 3709 714
rect 3084 658 3118 696
rect 3084 586 3118 624
rect 3506 633 3540 671
rect 3646 680 3709 705
rect 3743 710 3777 714
rect 3743 680 3773 710
rect 3811 680 3845 714
rect 3879 680 3913 714
rect 3947 680 4000 714
rect 3646 676 3773 680
rect 3807 676 3845 680
rect 3879 676 4034 680
rect 3646 671 4034 676
rect 3612 644 4034 671
rect 3612 636 3709 644
rect 3646 610 3709 636
rect 3743 634 3777 644
rect 3743 610 3773 634
rect 3811 610 3845 644
rect 3879 610 3913 644
rect 3947 610 4000 644
rect 3646 602 3773 610
rect 3612 600 3773 602
rect 3807 600 3845 610
rect 3879 600 4034 610
rect 3612 574 4034 600
rect 3340 553 3374 574
rect 3302 519 3340 553
rect 3612 540 3709 574
rect 3743 558 3777 574
rect 3743 540 3773 558
rect 3811 540 3845 574
rect 3879 540 3913 574
rect 3947 540 4000 574
rect 3612 524 3773 540
rect 3807 524 3845 540
rect 3879 524 4034 540
rect 5192 712 5226 728
rect 5192 644 5226 658
rect 5192 600 5226 610
rect 5192 526 5226 542
rect 5276 716 5872 744
rect 7114 860 7536 878
rect 9899 945 9929 979
rect 9899 942 9963 945
rect 9933 911 9963 942
rect 9899 877 9929 908
rect 9899 870 9963 877
rect 7114 854 7271 860
rect 7305 854 7343 860
rect 7377 854 7536 860
rect 7148 820 7207 854
rect 7241 826 7271 854
rect 7241 820 7275 826
rect 7309 820 7343 854
rect 7377 820 7411 854
rect 7445 843 7536 854
rect 7445 820 7502 843
rect 7114 809 7502 820
rect 7114 785 7536 809
rect 7114 784 7271 785
rect 7305 784 7343 785
rect 7377 784 7536 785
rect 7148 750 7207 784
rect 7241 751 7271 784
rect 7241 750 7275 751
rect 7309 750 7343 784
rect 7377 750 7411 784
rect 7445 774 7536 784
rect 7445 750 7502 774
rect 7114 740 7502 750
rect 7587 800 7621 826
rect 9933 843 9963 870
rect 9899 809 9929 836
rect 7587 788 7622 800
rect 7621 766 7622 788
rect 7656 766 7690 800
rect 7724 766 7740 800
rect 7852 766 7868 800
rect 7902 766 7936 800
rect 7970 766 8124 800
rect 8158 766 8192 800
rect 8226 766 8380 800
rect 8414 766 8448 800
rect 8482 766 8636 800
rect 8670 766 8704 800
rect 8738 766 8892 800
rect 8926 766 8960 800
rect 8994 766 9054 800
rect 9122 766 9138 800
rect 9172 766 9206 800
rect 9240 766 9256 800
rect 9899 798 9963 809
rect 9933 775 9963 798
rect 5310 682 5359 716
rect 5393 682 5427 716
rect 5461 682 5495 716
rect 5529 682 5563 716
rect 5597 682 5631 716
rect 5665 682 5699 716
rect 5733 682 5767 716
rect 5801 682 5838 716
rect 5276 670 5563 682
rect 5597 670 5872 682
rect 5276 646 5872 670
rect 5310 612 5359 646
rect 5393 612 5427 646
rect 5461 612 5495 646
rect 5529 612 5563 646
rect 5597 612 5631 646
rect 5665 612 5699 646
rect 5733 612 5767 646
rect 5801 612 5838 646
rect 5276 596 5563 612
rect 5597 596 5872 612
rect 5276 576 5872 596
rect 5310 542 5359 576
rect 5393 542 5427 576
rect 5461 542 5495 576
rect 5529 542 5563 576
rect 5597 542 5631 576
rect 5665 542 5699 576
rect 5733 542 5767 576
rect 5801 542 5838 576
rect 1117 503 1287 507
rect 1117 497 1185 503
rect 1151 463 1185 497
rect 1219 472 1287 503
rect 3612 504 4034 524
rect 1117 451 1185 463
rect 1219 451 1253 472
rect 1117 438 1253 451
rect 1530 446 1554 480
rect 1588 446 1623 480
rect 1657 446 1692 480
rect 1726 446 1761 480
rect 1795 446 1830 480
rect 1864 446 1899 480
rect 1933 446 1968 480
rect 2002 446 2038 480
rect 2072 446 2108 480
rect 2142 446 2178 480
rect 2212 446 2248 480
rect 2282 446 2318 480
rect 2352 446 2388 480
rect 2422 446 2458 480
rect 2492 446 2528 480
rect 2562 446 2598 480
rect 2632 446 2668 480
rect 2702 446 2738 480
rect 2772 446 2808 480
rect 2842 446 2878 480
rect 2912 446 2948 480
rect 2982 446 3018 480
rect 3052 446 3088 480
rect 3122 446 3158 480
rect 3192 446 3228 480
rect 3262 446 3298 480
rect 3332 446 3368 480
rect 3402 446 3438 480
rect 3472 446 3508 480
rect 3542 446 3578 480
rect 3612 470 3709 504
rect 3743 482 3777 504
rect 3743 470 3773 482
rect 3811 470 3845 504
rect 3879 470 3913 504
rect 3947 470 4000 504
rect 3612 448 3773 470
rect 3807 448 3845 470
rect 3879 448 4034 470
rect 5276 522 5563 542
rect 5597 522 5872 542
rect 5276 506 5872 522
rect 7032 712 7066 728
rect 7032 644 7066 658
rect 7032 576 7066 586
rect 7114 714 7536 740
rect 7148 680 7207 714
rect 7241 710 7275 714
rect 7241 680 7271 710
rect 7309 680 7343 714
rect 7377 680 7411 714
rect 7445 705 7536 714
rect 7445 680 7502 705
rect 7114 676 7271 680
rect 7305 676 7343 680
rect 7377 676 7502 680
rect 7114 671 7502 676
rect 7114 644 7536 671
rect 7148 610 7207 644
rect 7241 634 7275 644
rect 7241 610 7271 634
rect 7309 610 7343 644
rect 7377 610 7411 644
rect 7445 636 7536 644
rect 7445 610 7502 636
rect 7114 600 7271 610
rect 7305 600 7343 610
rect 7377 602 7502 610
rect 7618 636 7652 674
rect 8030 658 8064 696
rect 7377 600 7536 602
rect 7114 574 7536 600
rect 8030 586 8064 624
rect 7148 540 7207 574
rect 7241 558 7275 574
rect 7241 540 7271 558
rect 7309 540 7343 574
rect 7377 540 7411 574
rect 7445 540 7536 574
rect 7808 544 7846 578
rect 8286 636 8320 674
rect 8286 564 8320 602
rect 7114 524 7271 540
rect 7305 524 7343 540
rect 7377 524 7536 540
rect 9054 728 9088 766
rect 8542 658 8576 696
rect 8542 586 8576 624
rect 8798 636 8832 674
rect 9054 656 9088 694
rect 9210 708 9244 766
rect 9210 636 9244 674
rect 8798 564 8832 602
rect 9210 564 9244 602
rect 9899 741 9929 764
rect 9899 726 9963 741
rect 9933 707 9963 726
rect 9899 673 9929 692
rect 9899 654 9963 673
rect 9933 639 9963 654
rect 9899 605 9929 620
rect 9899 582 9963 605
rect 9933 571 9963 582
rect 9899 537 9929 548
rect 5310 472 5359 506
rect 5393 472 5427 506
rect 5461 472 5495 506
rect 5529 472 5563 506
rect 5597 472 5631 506
rect 5665 472 5699 506
rect 5733 472 5767 506
rect 5801 472 5838 506
rect 5276 448 5563 472
rect 5597 448 5872 472
rect 7114 504 7536 524
rect 7148 470 7207 504
rect 7241 482 7275 504
rect 7241 470 7271 482
rect 7309 470 7343 504
rect 7377 470 7411 504
rect 7445 470 7536 504
rect 9899 510 9963 537
rect 9933 503 9963 510
rect 7114 448 7271 470
rect 7305 448 7343 470
rect 7377 448 7536 470
rect 3612 446 4034 448
rect 7114 446 7536 448
rect 7570 446 7606 480
rect 7640 446 7676 480
rect 7710 446 7746 480
rect 7780 446 7816 480
rect 7850 446 7886 480
rect 7920 446 7956 480
rect 7990 446 8026 480
rect 8060 446 8096 480
rect 8130 446 8166 480
rect 8200 446 8236 480
rect 8270 446 8306 480
rect 8340 446 8376 480
rect 8410 446 8446 480
rect 8480 446 8516 480
rect 8550 446 8586 480
rect 8620 446 8656 480
rect 8690 446 8726 480
rect 8760 446 8796 480
rect 8830 446 8866 480
rect 8900 446 8936 480
rect 8970 446 9006 480
rect 9040 446 9076 480
rect 9110 446 9146 480
rect 9180 446 9215 480
rect 9249 446 9284 480
rect 9318 446 9353 480
rect 9387 446 9422 480
rect 9456 446 9491 480
rect 9525 446 9560 480
rect 9594 446 9618 480
rect 9899 469 9929 476
rect 1117 435 1287 438
rect 1117 428 1185 435
rect 1151 394 1185 428
rect 1219 403 1287 435
rect 1117 379 1185 394
rect 1219 379 1253 403
rect 1117 369 1253 379
rect 1117 367 1287 369
rect 1117 359 1185 367
rect 1151 325 1185 359
rect 1219 334 1287 367
rect 1117 307 1185 325
rect 1219 307 1253 334
rect 1117 300 1253 307
rect 1117 299 1287 300
rect 1117 290 1185 299
rect 1151 256 1185 290
rect 1219 265 1287 299
rect 1117 235 1185 256
rect 1219 235 1253 265
rect 1117 231 1253 235
rect 1117 221 1185 231
rect 1151 187 1185 221
rect 1219 197 1287 231
rect 9899 438 9963 469
rect 10239 7671 10277 7699
rect 10317 7671 10349 7705
rect 10385 7671 10419 7705
rect 10455 7671 10487 7705
rect 10527 7671 10555 7705
rect 10599 7671 10623 7705
rect 10671 7671 10691 7705
rect 10743 7671 10759 7705
rect 10816 7671 10827 7705
rect 10889 7671 10895 7705
rect 10962 7671 10963 7705
rect 10997 7671 11001 7705
rect 11065 7671 11074 7705
rect 11133 7671 11147 7705
rect 11201 7671 11220 7705
rect 11269 7671 11293 7705
rect 11337 7671 11366 7705
rect 11405 7671 11439 7705
rect 11473 7671 11507 7705
rect 11546 7671 11575 7705
rect 11619 7671 11643 7705
rect 11692 7671 11711 7705
rect 11765 7671 11779 7705
rect 11838 7671 11847 7705
rect 11911 7671 11915 7705
rect 11949 7671 11950 7705
rect 12017 7671 12023 7705
rect 12085 7671 12096 7705
rect 12153 7671 12169 7705
rect 12221 7671 12242 7705
rect 12289 7671 12315 7705
rect 12357 7671 12388 7705
rect 12425 7671 12459 7705
rect 12495 7671 12527 7705
rect 12568 7671 12595 7705
rect 12641 7671 12663 7705
rect 12714 7671 12731 7705
rect 12787 7671 12799 7705
rect 10205 7637 10212 7665
rect 10205 7627 10246 7637
rect 10239 7603 10246 7627
rect 10205 7569 10212 7593
rect 10205 7555 10246 7569
rect 10239 7535 10246 7555
rect 10205 7501 10212 7521
rect 10205 7483 10246 7501
rect 10239 7467 10246 7483
rect 10205 7433 10212 7449
rect 10205 7411 10246 7433
rect 10239 7399 10246 7411
rect 10205 7365 10212 7377
rect 10205 7339 10246 7365
rect 10239 7331 10246 7339
rect 10205 7297 10212 7305
rect 10205 7267 10246 7297
rect 10239 7263 10246 7267
rect 10205 7229 10212 7233
rect 10205 7195 10246 7229
rect 10205 7127 10246 7161
rect 10205 7123 10212 7127
rect 10239 7089 10246 7093
rect 10205 7059 10246 7089
rect 10205 7051 10212 7059
rect 10239 7017 10246 7025
rect 10205 6991 10246 7017
rect 10205 6979 10212 6991
rect 10239 6945 10246 6957
rect 10205 6923 10246 6945
rect 10205 6907 10212 6923
rect 10239 6873 10246 6889
rect 10205 6855 10246 6873
rect 10205 6835 10212 6855
rect 10239 6801 10246 6821
rect 10205 6787 10246 6801
rect 10205 6763 10212 6787
rect 10239 6729 10246 6753
rect 10205 6719 10246 6729
rect 10205 6691 10212 6719
rect 10239 6657 10246 6685
rect 10205 6651 10246 6657
rect 10205 6619 10212 6651
rect 10239 6585 10246 6617
rect 10205 6583 10246 6585
rect 10205 6549 10212 6583
rect 10205 6547 10246 6549
rect 10239 6515 10246 6547
rect 10205 6481 10212 6513
rect 10205 6475 10246 6481
rect 10239 6447 10246 6475
rect 10205 6413 10212 6441
rect 10205 6403 10246 6413
rect 10239 6379 10246 6403
rect 10205 6345 10212 6369
rect 10205 6331 10246 6345
rect 10239 6311 10246 6331
rect 10205 6277 10212 6297
rect 10205 6259 10246 6277
rect 10239 6243 10246 6259
rect 10205 6209 10212 6225
rect 10205 6187 10246 6209
rect 10239 6175 10246 6187
rect 10205 6141 10212 6153
rect 10205 6115 10246 6141
rect 10239 6107 10246 6115
rect 10205 6073 10212 6081
rect 10205 6043 10246 6073
rect 10239 6039 10246 6043
rect 10205 6005 10212 6009
rect 10205 5971 10246 6005
rect 10205 5903 10246 5937
rect 10205 5899 10212 5903
rect 10239 5865 10246 5869
rect 10205 5835 10246 5865
rect 10205 5827 10212 5835
rect 10239 5793 10246 5801
rect 10205 5767 10246 5793
rect 10205 5755 10212 5767
rect 10239 5721 10246 5733
rect 10205 5699 10246 5721
rect 10205 5683 10212 5699
rect 10239 5649 10246 5665
rect 10205 5631 10246 5649
rect 10205 5611 10212 5631
rect 10239 5577 10246 5597
rect 10205 5563 10246 5577
rect 10205 5539 10212 5563
rect 10239 5505 10246 5529
rect 10205 5495 10246 5505
rect 10205 5467 10212 5495
rect 10239 5433 10246 5461
rect 10205 5427 10246 5433
rect 10205 5395 10212 5427
rect 10239 5361 10246 5393
rect 10205 5359 10246 5361
rect 10205 5325 10212 5359
rect 10205 5323 10246 5325
rect 10239 5291 10246 5323
rect 10205 5257 10212 5289
rect 10205 5251 10246 5257
rect 10239 5223 10246 5251
rect 10205 5189 10212 5217
rect 10205 5179 10246 5189
rect 10239 5155 10246 5179
rect 10205 5121 10212 5145
rect 10205 5107 10246 5121
rect 10239 5087 10246 5107
rect 10205 5053 10212 5073
rect 10205 5035 10246 5053
rect 10239 5019 10246 5035
rect 10205 4985 10212 5001
rect 10205 4963 10246 4985
rect 10239 4951 10246 4963
rect 10205 4917 10212 4929
rect 10205 4891 10246 4917
rect 10239 4883 10246 4891
rect 10205 4849 10212 4857
rect 10205 4819 10246 4849
rect 10239 4815 10246 4819
rect 10205 4781 10212 4785
rect 10205 4747 10246 4781
rect 10205 4679 10246 4713
rect 10205 4675 10212 4679
rect 10239 4641 10246 4645
rect 10205 4611 10246 4641
rect 10205 4603 10212 4611
rect 10239 4569 10246 4577
rect 10205 4543 10246 4569
rect 10205 4531 10212 4543
rect 10239 4497 10246 4509
rect 10205 4475 10246 4497
rect 10205 4459 10212 4475
rect 10239 4425 10246 4441
rect 10205 4407 10246 4425
rect 10205 4387 10212 4407
rect 10239 4353 10246 4373
rect 10205 4339 10246 4353
rect 10205 4315 10212 4339
rect 10239 4281 10246 4305
rect 10205 4271 10246 4281
rect 10205 4243 10212 4271
rect 10239 4209 10246 4237
rect 10205 4203 10246 4209
rect 10205 4171 10212 4203
rect 10239 4137 10246 4169
rect 10205 4135 10246 4137
rect 10205 4101 10212 4135
rect 10205 4099 10246 4101
rect 10239 4067 10246 4099
rect 10205 4033 10212 4065
rect 10205 4027 10246 4033
rect 10239 3999 10246 4027
rect 10205 3965 10212 3993
rect 10205 3955 10246 3965
rect 10239 3931 10246 3955
rect 10205 3897 10212 3921
rect 10205 3883 10246 3897
rect 10239 3863 10246 3883
rect 10205 3829 10212 3849
rect 10205 3811 10246 3829
rect 10239 3795 10246 3811
rect 10205 3761 10212 3777
rect 10205 3739 10246 3761
rect 10239 3727 10246 3739
rect 10205 3693 10212 3705
rect 10205 3667 10246 3693
rect 10239 3659 10246 3667
rect 10205 3625 10212 3633
rect 10205 3595 10246 3625
rect 10239 3591 10246 3595
rect 10205 3557 10212 3561
rect 10205 3523 10246 3557
rect 10205 3455 10246 3489
rect 10205 3451 10212 3455
rect 10239 3417 10246 3421
rect 10205 3387 10246 3417
rect 10205 3379 10212 3387
rect 10239 3345 10246 3353
rect 10205 3319 10246 3345
rect 10205 3307 10212 3319
rect 10239 3273 10246 3285
rect 10205 3251 10246 3273
rect 10205 3235 10212 3251
rect 10239 3201 10246 3217
rect 10205 3183 10246 3201
rect 10205 3163 10212 3183
rect 10239 3129 10246 3149
rect 10205 3115 10246 3129
rect 10205 3091 10212 3115
rect 10239 3057 10246 3081
rect 10205 3047 10246 3057
rect 10205 3019 10212 3047
rect 10239 2985 10246 3013
rect 10205 2979 10246 2985
rect 10205 2947 10212 2979
rect 10239 2913 10246 2945
rect 10205 2911 10246 2913
rect 10205 2877 10212 2911
rect 10205 2875 10246 2877
rect 10239 2843 10246 2875
rect 10205 2809 10212 2841
rect 10205 2803 10246 2809
rect 10239 2775 10246 2803
rect 10205 2741 10212 2769
rect 10205 2731 10246 2741
rect 10239 2707 10246 2731
rect 10205 2673 10212 2697
rect 10205 2659 10246 2673
rect 10239 2639 10246 2659
rect 10205 2605 10212 2625
rect 10205 2587 10246 2605
rect 10239 2571 10246 2587
rect 10205 2537 10212 2553
rect 10205 2515 10246 2537
rect 10239 2503 10246 2515
rect 10205 2469 10212 2481
rect 10205 2443 10246 2469
rect 10239 2435 10246 2443
rect 10205 2401 10212 2409
rect 10205 2371 10246 2401
rect 10239 2367 10246 2371
rect 10205 2333 10212 2337
rect 10205 2299 10246 2333
rect 10205 2231 10246 2265
rect 10205 2227 10212 2231
rect 10239 2193 10246 2197
rect 10205 2163 10246 2193
rect 10205 2155 10212 2163
rect 10239 2121 10246 2129
rect 10205 2095 10246 2121
rect 10205 2083 10212 2095
rect 10239 2049 10246 2061
rect 10205 2027 10246 2049
rect 10205 2011 10212 2027
rect 10239 1977 10246 1993
rect 10205 1959 10246 1977
rect 10205 1939 10212 1959
rect 10239 1905 10246 1925
rect 10205 1891 10246 1905
rect 10205 1867 10212 1891
rect 10239 1833 10246 1857
rect 10205 1823 10246 1833
rect 10205 1795 10212 1823
rect 10239 1761 10246 1789
rect 10205 1755 10246 1761
rect 10205 1723 10212 1755
rect 10239 1689 10246 1721
rect 10205 1687 10246 1689
rect 10205 1653 10212 1687
rect 10205 1651 10246 1653
rect 10239 1619 10246 1651
rect 10205 1585 10212 1617
rect 10205 1579 10246 1585
rect 10239 1551 10246 1579
rect 10205 1517 10212 1545
rect 10205 1507 10246 1517
rect 10239 1483 10246 1507
rect 10205 1449 10212 1473
rect 10205 1435 10246 1449
rect 10239 1415 10246 1435
rect 10205 1381 10212 1401
rect 10205 1363 10246 1381
rect 10239 1347 10246 1363
rect 10205 1313 10212 1329
rect 10205 1291 10246 1313
rect 10239 1279 10246 1291
rect 10205 1245 10212 1257
rect 10205 1219 10246 1245
rect 10239 1211 10246 1219
rect 10205 1177 10212 1185
rect 10205 1147 10246 1177
rect 10239 1143 10246 1147
rect 10205 1109 10212 1113
rect 10205 1075 10246 1109
rect 10205 1007 10246 1041
rect 10205 1003 10212 1007
rect 10239 969 10246 973
rect 10205 939 10246 969
rect 10205 930 10212 939
rect 10239 896 10246 905
rect 10205 871 10246 896
rect 10205 857 10212 871
rect 10239 823 10246 837
rect 10205 803 10246 823
rect 10205 784 10212 803
rect 10239 750 10246 769
rect 10205 735 10246 750
rect 10205 711 10212 735
rect 10239 677 10246 701
rect 10205 667 10246 677
rect 10205 638 10212 667
rect 10239 604 10246 633
rect 10205 599 10246 604
rect 10205 565 10212 599
rect 10239 531 10246 565
rect 10205 492 10246 531
rect 10239 458 10246 492
rect 13069 7666 13103 7700
rect 13069 7598 13103 7632
rect 13069 7530 13103 7564
rect 13069 7462 13103 7496
rect 13069 7394 13103 7428
rect 13069 7326 13103 7360
rect 13069 7258 13103 7292
rect 13069 7190 13103 7224
rect 13069 7122 13103 7126
rect 13069 7016 13103 7020
rect 13069 6944 13103 6952
rect 13069 6872 13103 6884
rect 13069 6800 13103 6816
rect 13069 6728 13103 6748
rect 13069 6656 13103 6680
rect 13069 6584 13103 6612
rect 13069 6512 13103 6544
rect 13069 6442 13103 6476
rect 13069 6374 13103 6406
rect 13069 6306 13103 6334
rect 13069 6238 13103 6262
rect 13069 6170 13103 6190
rect 13069 6102 13103 6118
rect 13069 6034 13103 6046
rect 13069 5966 13103 5974
rect 13069 5898 13103 5902
rect 13069 5792 13103 5796
rect 13069 5720 13103 5728
rect 13069 5648 13103 5660
rect 13069 5576 13103 5592
rect 13069 5504 13103 5524
rect 13069 5432 13103 5456
rect 13069 5360 13103 5388
rect 13069 5288 13103 5320
rect 13069 5218 13103 5252
rect 13069 5150 13103 5182
rect 13069 5082 13103 5110
rect 13069 5014 13103 5038
rect 13069 4946 13103 4966
rect 13069 4878 13103 4894
rect 13069 4810 13103 4822
rect 13069 4742 13103 4750
rect 13069 4674 13103 4678
rect 13069 4568 13103 4572
rect 13069 4496 13103 4504
rect 13069 4424 13103 4436
rect 13069 4352 13103 4368
rect 13069 4280 13103 4300
rect 13069 4208 13103 4232
rect 13069 4136 13103 4164
rect 13069 4064 13103 4096
rect 13069 3994 13103 4028
rect 13069 3926 13103 3958
rect 13069 3858 13103 3886
rect 13069 3790 13103 3814
rect 13069 3722 13103 3742
rect 13069 3654 13103 3670
rect 13069 3586 13103 3598
rect 13069 3518 13103 3526
rect 13069 3450 13103 3454
rect 13069 3344 13103 3348
rect 13069 3272 13103 3280
rect 13069 3200 13103 3212
rect 13069 3128 13103 3144
rect 13069 3056 13103 3076
rect 13069 2984 13103 3008
rect 13069 2912 13103 2940
rect 13069 2840 13103 2872
rect 13069 2770 13103 2804
rect 13069 2702 13103 2734
rect 13069 2634 13103 2662
rect 13069 2566 13103 2589
rect 13069 2498 13103 2516
rect 13069 2430 13103 2443
rect 13069 2362 13103 2370
rect 13069 2294 13103 2297
rect 13069 2258 13103 2260
rect 13069 2185 13103 2192
rect 13069 2112 13103 2124
rect 13069 2039 13103 2056
rect 13069 1966 13103 1988
rect 13069 1893 13103 1920
rect 13069 1820 13103 1852
rect 13069 1750 13103 1784
rect 13069 1682 13103 1713
rect 13069 1614 13103 1640
rect 13069 1546 13103 1567
rect 13069 1478 13103 1494
rect 13069 1410 13103 1421
rect 13069 1342 13103 1348
rect 13069 1274 13103 1275
rect 13069 1236 13103 1240
rect 13069 1163 13103 1172
rect 13069 1090 13103 1104
rect 13069 1017 13103 1036
rect 13069 944 13103 968
rect 13069 871 13103 900
rect 13069 798 13103 832
rect 13069 730 13103 764
rect 13069 662 13103 691
rect 13069 594 13103 618
rect 13069 526 13103 545
rect 10212 446 10246 458
rect 10311 446 10314 480
rect 10348 446 10350 480
rect 10416 446 10423 480
rect 10484 446 10496 480
rect 10552 446 10569 480
rect 10620 446 10642 480
rect 10676 446 10690 480
rect 10749 446 10758 480
rect 10822 446 10826 480
rect 10860 446 10861 480
rect 10928 446 10934 480
rect 10996 446 11007 480
rect 11064 446 11080 480
rect 11132 446 11153 480
rect 11200 446 11226 480
rect 11268 446 11299 480
rect 11336 446 11370 480
rect 11406 446 11438 480
rect 11479 446 11506 480
rect 11552 446 11574 480
rect 11625 446 11642 480
rect 11698 446 11710 480
rect 11771 446 11778 480
rect 11844 446 11846 480
rect 11880 446 11883 480
rect 11948 446 11956 480
rect 12016 446 12029 480
rect 12084 446 12102 480
rect 12152 446 12175 480
rect 12220 446 12248 480
rect 12288 446 12321 480
rect 12356 446 12390 480
rect 12427 446 12458 480
rect 12499 446 12526 480
rect 12571 446 12594 480
rect 12643 446 12662 480
rect 12715 446 12730 480
rect 12787 446 12799 480
rect 13069 458 13103 472
rect 9933 435 9963 438
rect 9899 401 9929 404
rect 9899 367 9963 401
rect 9899 366 9929 367
rect 9933 332 9963 333
rect 9899 299 9963 332
rect 9899 294 9929 299
rect 9933 260 9963 265
rect 9899 231 9963 260
rect 9899 222 9929 231
rect 13069 390 13103 399
rect 13069 322 13103 326
rect 13069 287 13103 288
rect 13069 214 13103 253
rect 1117 163 1185 187
rect 1219 163 1257 197
rect 1316 163 1329 197
rect 1384 163 1401 197
rect 1452 163 1473 197
rect 1520 163 1545 197
rect 1588 163 1617 197
rect 1656 163 1689 197
rect 1724 163 1758 197
rect 1795 163 1826 197
rect 1867 163 1894 197
rect 1939 163 1962 197
rect 2011 163 2030 197
rect 2083 163 2098 197
rect 2155 163 2166 197
rect 2227 163 2234 197
rect 2299 163 2302 197
rect 2336 163 2337 197
rect 2404 163 2409 197
rect 2472 163 2481 197
rect 2540 163 2553 197
rect 2608 163 2625 197
rect 2676 163 2697 197
rect 2744 163 2769 197
rect 2812 163 2841 197
rect 2880 163 2913 197
rect 2948 163 2982 197
rect 3019 163 3050 197
rect 3091 163 3118 197
rect 3163 163 3186 197
rect 3235 163 3254 197
rect 3307 163 3322 197
rect 3379 163 3390 197
rect 3451 163 3458 197
rect 3523 163 3526 197
rect 3560 163 3561 197
rect 3628 163 3633 197
rect 3696 163 3705 197
rect 3764 163 3777 197
rect 3832 163 3849 197
rect 3900 163 3921 197
rect 3968 163 3993 197
rect 4036 163 4065 197
rect 4104 163 4137 197
rect 4172 163 4206 197
rect 4243 163 4274 197
rect 4315 163 4342 197
rect 4387 163 4410 197
rect 4459 163 4478 197
rect 4531 163 4546 197
rect 4603 163 4614 197
rect 4675 163 4682 197
rect 4747 163 4750 197
rect 4784 163 4785 197
rect 4852 163 4857 197
rect 4920 163 4929 197
rect 4988 163 5001 197
rect 5056 163 5073 197
rect 5124 163 5145 197
rect 5192 163 5217 197
rect 5260 163 5289 197
rect 5328 163 5361 197
rect 5396 163 5430 197
rect 5467 163 5498 197
rect 5539 163 5566 197
rect 5611 163 5649 197
rect 5702 163 5721 197
rect 5770 163 5793 197
rect 5838 163 5865 197
rect 5906 163 5937 197
rect 5974 163 6008 197
rect 6043 163 6076 197
rect 6115 163 6144 197
rect 6187 163 6212 197
rect 6259 163 6280 197
rect 6331 163 6348 197
rect 6403 163 6416 197
rect 6475 163 6484 197
rect 6547 163 6552 197
rect 6619 163 6620 197
rect 6654 163 6657 197
rect 6722 163 6729 197
rect 6790 163 6801 197
rect 6858 163 6873 197
rect 6926 163 6945 197
rect 6994 163 7017 197
rect 7062 163 7089 197
rect 7130 163 7161 197
rect 7198 163 7232 197
rect 7267 163 7300 197
rect 7339 163 7368 197
rect 7411 163 7436 197
rect 7483 163 7504 197
rect 7555 163 7572 197
rect 7627 163 7640 197
rect 7699 163 7708 197
rect 7771 163 7776 197
rect 7843 163 7844 197
rect 7878 163 7881 197
rect 7946 163 7953 197
rect 8014 163 8025 197
rect 8082 163 8097 197
rect 8150 163 8169 197
rect 8218 163 8241 197
rect 8286 163 8313 197
rect 8354 163 8385 197
rect 8422 163 8456 197
rect 8491 163 8524 197
rect 8563 163 8592 197
rect 8635 163 8660 197
rect 8707 163 8728 197
rect 8779 163 8796 197
rect 8851 163 8864 197
rect 8923 163 8932 197
rect 8995 163 9000 197
rect 9067 163 9068 197
rect 9102 163 9105 197
rect 9170 163 9177 197
rect 9238 163 9249 197
rect 9306 163 9321 197
rect 9374 163 9393 197
rect 9442 163 9465 197
rect 9510 163 9537 197
rect 9578 163 9609 197
rect 9646 163 9680 197
rect 9715 163 9748 197
rect 9788 163 9816 197
rect 9861 188 9899 197
rect 9933 188 9971 197
rect 9861 163 9971 188
rect 10005 163 10043 197
rect 10078 163 10111 197
rect 10151 163 10179 197
rect 10223 163 10247 197
rect 10295 163 10315 197
rect 10367 163 10383 197
rect 10439 163 10451 197
rect 10511 163 10519 197
rect 10583 163 10587 197
rect 10689 163 10693 197
rect 10757 163 10765 197
rect 10825 163 10837 197
rect 10893 163 10909 197
rect 10961 163 10981 197
rect 11029 163 11053 197
rect 11097 163 11125 197
rect 11165 163 11197 197
rect 11233 163 11267 197
rect 11303 163 11335 197
rect 11375 163 11403 197
rect 11447 163 11471 197
rect 11519 163 11539 197
rect 11591 163 11607 197
rect 11663 163 11675 197
rect 11735 163 11743 197
rect 11807 163 11811 197
rect 11913 163 11917 197
rect 11981 163 11989 197
rect 12049 163 12061 197
rect 12117 163 12133 197
rect 12185 163 12205 197
rect 12253 163 12277 197
rect 12321 163 12349 197
rect 12389 163 12421 197
rect 12457 163 12491 197
rect 12527 163 12559 197
rect 12599 163 12627 197
rect 12671 163 12695 197
rect 12743 163 12763 197
rect 12815 163 12831 197
rect 12887 163 12899 197
rect 12959 163 12967 197
rect 13031 163 13035 197
rect 13069 163 13103 180
<< viali >>
rect 1235 14200 1265 14234
rect 1265 14200 1269 14234
rect 1308 14200 1333 14234
rect 1333 14200 1342 14234
rect 1381 14200 1401 14234
rect 1401 14200 1415 14234
rect 1454 14200 1469 14234
rect 1469 14200 1488 14234
rect 1527 14200 1537 14234
rect 1537 14200 1561 14234
rect 1600 14200 1605 14234
rect 1605 14200 1634 14234
rect 1673 14200 1707 14234
rect 1746 14200 1775 14234
rect 1775 14200 1780 14234
rect 1819 14200 1843 14234
rect 1843 14200 1853 14234
rect 1892 14200 1911 14234
rect 1911 14200 1926 14234
rect 1965 14200 1979 14234
rect 1979 14200 1999 14234
rect 2038 14200 2047 14234
rect 2047 14200 2072 14234
rect 2111 14200 2115 14234
rect 2115 14200 2145 14234
rect 2183 14200 2217 14234
rect 2255 14200 2285 14234
rect 2285 14200 2289 14234
rect 2327 14200 2353 14234
rect 2353 14200 2361 14234
rect 2399 14200 2421 14234
rect 2421 14200 2433 14234
rect 2471 14200 2489 14234
rect 2489 14200 2505 14234
rect 2543 14200 2557 14234
rect 2557 14200 2577 14234
rect 2615 14200 2625 14234
rect 2625 14200 2649 14234
rect 2687 14200 2693 14234
rect 2693 14200 2721 14234
rect 2759 14200 2761 14234
rect 2761 14200 2793 14234
rect 2831 14200 2863 14234
rect 2863 14200 2865 14234
rect 2903 14200 2931 14234
rect 2931 14200 2937 14234
rect 2975 14200 2999 14234
rect 2999 14200 3009 14234
rect 3047 14200 3067 14234
rect 3067 14200 3081 14234
rect 3119 14200 3135 14234
rect 3135 14200 3153 14234
rect 3191 14200 3203 14234
rect 3203 14200 3225 14234
rect 3263 14200 3271 14234
rect 3271 14200 3297 14234
rect 3335 14200 3339 14234
rect 3339 14200 3369 14234
rect 3407 14200 3441 14234
rect 3479 14200 3509 14234
rect 3509 14200 3513 14234
rect 3551 14200 3577 14234
rect 3577 14200 3585 14234
rect 3623 14200 3645 14234
rect 3645 14200 3657 14234
rect 3695 14200 3713 14234
rect 3713 14200 3729 14234
rect 3767 14200 3781 14234
rect 3781 14200 3801 14234
rect 3839 14200 3849 14234
rect 3849 14200 3873 14234
rect 3911 14200 3917 14234
rect 3917 14200 3945 14234
rect 3983 14200 3985 14234
rect 3985 14200 4017 14234
rect 4055 14200 4087 14234
rect 4087 14200 4089 14234
rect 4127 14200 4155 14234
rect 4155 14200 4161 14234
rect 4199 14200 4223 14234
rect 4223 14200 4233 14234
rect 4271 14200 4291 14234
rect 4291 14200 4305 14234
rect 4343 14200 4359 14234
rect 4359 14200 4377 14234
rect 4415 14200 4427 14234
rect 4427 14200 4449 14234
rect 4487 14200 4495 14234
rect 4495 14200 4521 14234
rect 4559 14200 4563 14234
rect 4563 14200 4593 14234
rect 4631 14200 4665 14234
rect 4703 14200 4733 14234
rect 4733 14200 4737 14234
rect 4775 14200 4801 14234
rect 4801 14200 4809 14234
rect 4847 14200 4869 14234
rect 4869 14200 4881 14234
rect 4919 14200 4937 14234
rect 4937 14200 4953 14234
rect 4991 14200 5005 14234
rect 5005 14200 5025 14234
rect 5063 14200 5073 14234
rect 5073 14200 5097 14234
rect 5135 14200 5141 14234
rect 5141 14200 5169 14234
rect 5207 14200 5209 14234
rect 5209 14200 5241 14234
rect 5279 14200 5311 14234
rect 5311 14200 5313 14234
rect 5351 14200 5379 14234
rect 5379 14200 5385 14234
rect 5423 14200 5447 14234
rect 5447 14200 5457 14234
rect 5495 14200 5515 14234
rect 5515 14200 5529 14234
rect 5567 14200 5583 14234
rect 5583 14200 5601 14234
rect 5639 14200 5651 14234
rect 5651 14200 5673 14234
rect 5711 14200 5719 14234
rect 5719 14200 5745 14234
rect 5783 14200 5787 14234
rect 5787 14200 5817 14234
rect 5855 14200 5889 14234
rect 5927 14200 5957 14234
rect 5957 14200 5961 14234
rect 5999 14200 6025 14234
rect 6025 14200 6033 14234
rect 6071 14200 6093 14234
rect 6093 14200 6105 14234
rect 6143 14200 6161 14234
rect 6161 14200 6177 14234
rect 6215 14200 6229 14234
rect 6229 14200 6249 14234
rect 6287 14200 6297 14234
rect 6297 14200 6321 14234
rect 6359 14200 6365 14234
rect 6365 14200 6393 14234
rect 6431 14200 6433 14234
rect 6433 14200 6465 14234
rect 6503 14200 6535 14234
rect 6535 14200 6537 14234
rect 6575 14200 6603 14234
rect 6603 14200 6609 14234
rect 6647 14200 6671 14234
rect 6671 14200 6681 14234
rect 6719 14200 6739 14234
rect 6739 14200 6753 14234
rect 6791 14200 6807 14234
rect 6807 14200 6825 14234
rect 6863 14200 6875 14234
rect 6875 14200 6897 14234
rect 6935 14200 6943 14234
rect 6943 14200 6969 14234
rect 7007 14200 7011 14234
rect 7011 14200 7041 14234
rect 7079 14200 7113 14234
rect 7151 14200 7181 14234
rect 7181 14200 7185 14234
rect 7223 14200 7249 14234
rect 7249 14200 7257 14234
rect 7295 14200 7317 14234
rect 7317 14200 7329 14234
rect 7367 14200 7385 14234
rect 7385 14200 7401 14234
rect 7439 14200 7453 14234
rect 7453 14200 7473 14234
rect 7511 14200 7521 14234
rect 7521 14200 7545 14234
rect 7583 14200 7589 14234
rect 7589 14200 7617 14234
rect 7655 14200 7657 14234
rect 7657 14200 7689 14234
rect 7727 14200 7759 14234
rect 7759 14200 7761 14234
rect 7799 14200 7827 14234
rect 7827 14200 7833 14234
rect 7871 14200 7895 14234
rect 7895 14200 7905 14234
rect 7943 14200 7963 14234
rect 7963 14200 7977 14234
rect 8015 14200 8031 14234
rect 8031 14200 8049 14234
rect 8087 14200 8099 14234
rect 8099 14200 8121 14234
rect 8159 14200 8167 14234
rect 8167 14200 8193 14234
rect 8231 14200 8235 14234
rect 8235 14200 8265 14234
rect 8303 14200 8337 14234
rect 8375 14200 8405 14234
rect 8405 14200 8409 14234
rect 8447 14200 8473 14234
rect 8473 14200 8481 14234
rect 8519 14200 8541 14234
rect 8541 14200 8553 14234
rect 8591 14200 8609 14234
rect 8609 14200 8625 14234
rect 8663 14200 8677 14234
rect 8677 14200 8697 14234
rect 8735 14200 8745 14234
rect 8745 14200 8769 14234
rect 8807 14200 8813 14234
rect 8813 14200 8841 14234
rect 8879 14200 8881 14234
rect 8881 14200 8913 14234
rect 8951 14200 8983 14234
rect 8983 14200 8985 14234
rect 9023 14200 9051 14234
rect 9051 14200 9057 14234
rect 9095 14200 9119 14234
rect 9119 14200 9129 14234
rect 9167 14200 9187 14234
rect 9187 14200 9201 14234
rect 9239 14200 9255 14234
rect 9255 14200 9273 14234
rect 9311 14200 9323 14234
rect 9323 14200 9345 14234
rect 9383 14200 9391 14234
rect 9391 14200 9417 14234
rect 9455 14200 9459 14234
rect 9459 14200 9489 14234
rect 9527 14200 9561 14234
rect 9599 14200 9629 14234
rect 9629 14200 9633 14234
rect 9671 14200 9697 14234
rect 9697 14200 9705 14234
rect 9743 14200 9765 14234
rect 9765 14200 9777 14234
rect 9815 14200 9833 14234
rect 9833 14200 9849 14234
rect 9887 14200 9901 14234
rect 9901 14200 9921 14234
rect 9959 14200 9969 14234
rect 9969 14200 9993 14234
rect 10031 14200 10037 14234
rect 10037 14200 10065 14234
rect 10103 14200 10105 14234
rect 10105 14200 10137 14234
rect 10175 14200 10207 14234
rect 10207 14200 10209 14234
rect 10247 14200 10275 14234
rect 10275 14200 10281 14234
rect 10319 14200 10343 14234
rect 10343 14200 10353 14234
rect 10391 14200 10411 14234
rect 10411 14200 10425 14234
rect 10463 14200 10479 14234
rect 10479 14200 10497 14234
rect 10535 14200 10547 14234
rect 10547 14200 10569 14234
rect 10607 14200 10615 14234
rect 10615 14200 10641 14234
rect 10679 14200 10683 14234
rect 10683 14200 10713 14234
rect 10751 14200 10785 14234
rect 10823 14200 10853 14234
rect 10853 14200 10857 14234
rect 10895 14200 10921 14234
rect 10921 14200 10929 14234
rect 10967 14200 10989 14234
rect 10989 14200 11001 14234
rect 1197 14100 1231 14124
rect 1197 14090 1231 14100
rect 1984 14098 2018 14132
rect 2059 14098 2093 14132
rect 2134 14098 2168 14132
rect 2209 14098 2243 14132
rect 2284 14098 2318 14132
rect 2359 14098 2393 14132
rect 2434 14098 2468 14132
rect 2509 14098 2543 14132
rect 2584 14098 2618 14132
rect 2659 14098 2693 14132
rect 2734 14098 2768 14132
rect 2809 14098 2843 14132
rect 2884 14098 2918 14132
rect 2959 14098 2993 14132
rect 3033 14098 3067 14132
rect 1197 14032 1231 14052
rect 1197 14018 1231 14032
rect 1197 13964 1231 13980
rect 1197 13946 1231 13964
rect 1197 13896 1231 13908
rect 1197 13874 1231 13896
rect 1197 13828 1231 13836
rect 1197 13802 1231 13828
rect 1197 13760 1231 13764
rect 1197 13730 1231 13760
rect 1197 13658 1231 13692
rect 1197 13590 1231 13620
rect 1197 13586 1231 13590
rect 1197 13522 1231 13548
rect 1197 13514 1231 13522
rect 1197 13454 1231 13476
rect 1197 13442 1231 13454
rect 1197 13386 1231 13404
rect 1197 13370 1231 13386
rect 1197 13318 1231 13332
rect 1197 13298 1231 13318
rect 1197 13250 1231 13260
rect 1197 13226 1231 13250
rect 1197 13182 1231 13188
rect 1197 13154 1231 13182
rect 1757 14077 1791 14093
rect 1757 14059 1791 14077
rect 3287 14077 3321 14093
rect 3287 14059 3321 14077
rect 8015 14098 8049 14132
rect 8089 14098 8123 14132
rect 8164 14098 8198 14132
rect 8239 14098 8273 14132
rect 8314 14098 8348 14132
rect 8389 14098 8423 14132
rect 8464 14098 8498 14132
rect 8539 14098 8573 14132
rect 8614 14098 8648 14132
rect 8689 14098 8723 14132
rect 8764 14098 8798 14132
rect 8839 14098 8873 14132
rect 8914 14098 8948 14132
rect 8989 14098 9023 14132
rect 9064 14098 9098 14132
rect 1757 14007 1791 14018
rect 1757 13984 1791 14007
rect 3287 14007 3321 14018
rect 3287 13984 3321 14007
rect 4538 14040 4572 14074
rect 4610 14040 4644 14074
rect 4682 14040 4716 14074
rect 1757 13937 1791 13943
rect 1757 13909 1791 13937
rect 3287 13937 3321 13943
rect 3287 13909 3321 13937
rect 1757 13867 1791 13868
rect 1757 13834 1791 13867
rect 3287 13867 3321 13868
rect 3287 13834 3321 13867
rect 1757 13763 1791 13793
rect 1757 13759 1791 13763
rect 3287 13763 3321 13793
rect 3700 13946 3734 13980
rect 3772 13946 3806 13980
rect 3844 13946 3878 13980
rect 7761 14077 7795 14093
rect 6218 14040 6252 14074
rect 6292 14040 6326 14074
rect 7761 14059 7795 14077
rect 9291 14077 9325 14093
rect 9291 14059 9325 14077
rect 9380 14119 9399 14126
rect 9399 14119 9414 14126
rect 9459 14119 9472 14126
rect 9472 14119 9493 14126
rect 9538 14119 9545 14126
rect 9545 14119 9572 14126
rect 9617 14119 9618 14126
rect 9618 14119 9651 14126
rect 9696 14119 9725 14126
rect 9725 14119 9730 14126
rect 9775 14119 9797 14126
rect 9797 14119 9809 14126
rect 9854 14119 9869 14126
rect 9869 14119 9888 14126
rect 9380 14092 9414 14119
rect 9459 14092 9493 14119
rect 9538 14092 9572 14119
rect 9617 14092 9651 14119
rect 9696 14092 9730 14119
rect 9775 14092 9809 14119
rect 9854 14092 9888 14119
rect 11077 14166 11111 14196
rect 11077 14162 11111 14166
rect 11077 14098 11111 14122
rect 11077 14088 11111 14098
rect 11077 14030 11111 14048
rect 7761 14007 7795 14018
rect 6029 13966 6063 14000
rect 6103 13979 6137 14000
rect 6103 13966 6119 13979
rect 6119 13966 6137 13979
rect 7761 13984 7795 14007
rect 4538 13884 4572 13918
rect 4610 13884 4644 13918
rect 4682 13884 4716 13918
rect 5268 13887 5284 13921
rect 5284 13887 5302 13921
rect 5342 13887 5356 13921
rect 5356 13887 5376 13921
rect 5416 13887 5428 13921
rect 5428 13887 5450 13921
rect 5490 13887 5500 13921
rect 5500 13887 5524 13921
rect 5564 13887 5572 13921
rect 5572 13887 5598 13921
rect 5638 13887 5644 13921
rect 5644 13887 5672 13921
rect 5712 13887 5715 13921
rect 5715 13887 5746 13921
rect 5786 13887 5820 13921
rect 7216 13946 7250 13980
rect 7288 13946 7322 13980
rect 7360 13946 7394 13980
rect 9291 14007 9325 14018
rect 9291 13984 9325 14007
rect 3700 13790 3734 13824
rect 3772 13790 3806 13824
rect 3844 13790 3878 13824
rect 4251 13800 4279 13834
rect 4279 13800 4285 13834
rect 3287 13759 3321 13763
rect 1757 13693 1791 13718
rect 1757 13684 1791 13693
rect 3287 13693 3321 13718
rect 3287 13684 3321 13693
rect 1757 13623 1791 13643
rect 1757 13609 1791 13623
rect 3287 13623 3321 13643
rect 3287 13609 3321 13623
rect 4131 13706 4137 13740
rect 4137 13706 4165 13740
rect 4131 13618 4137 13652
rect 4137 13618 4165 13652
rect 4251 13712 4279 13746
rect 4279 13712 4285 13746
rect 4257 13628 4291 13662
rect 4329 13628 4363 13662
rect 4401 13628 4435 13662
rect 5224 13795 5258 13829
rect 5224 13719 5258 13753
rect 5224 13643 5258 13677
rect 1757 13553 1791 13568
rect 1757 13534 1791 13553
rect 3287 13553 3321 13568
rect 3287 13534 3321 13553
rect 3419 13534 3453 13568
rect 3491 13534 3525 13568
rect 3563 13534 3597 13568
rect 1757 13483 1791 13493
rect 1757 13459 1791 13483
rect 3287 13483 3321 13493
rect 3287 13459 3321 13483
rect 1757 13413 1791 13418
rect 1757 13384 1791 13413
rect 3287 13413 3321 13418
rect 3287 13384 3321 13413
rect 1757 13309 1791 13343
rect 4131 13484 4165 13485
rect 4131 13451 4137 13484
rect 4137 13451 4165 13484
rect 4131 13396 4165 13397
rect 4131 13363 4137 13396
rect 4137 13363 4165 13396
rect 4538 13372 4572 13406
rect 4610 13372 4644 13406
rect 4682 13372 4716 13406
rect 5224 13568 5258 13602
rect 5224 13493 5258 13527
rect 5224 13418 5258 13452
rect 3287 13309 3321 13343
rect 3700 13278 3734 13312
rect 3772 13278 3806 13312
rect 3844 13278 3878 13312
rect 1757 13237 1791 13268
rect 1757 13234 1791 13237
rect 3287 13237 3321 13268
rect 3287 13234 3321 13237
rect 1197 13090 1231 13116
rect 1197 13082 1231 13090
rect 1757 13167 1791 13193
rect 1757 13159 1791 13167
rect 3287 13167 3321 13193
rect 3287 13159 3321 13167
rect 1757 13097 1791 13119
rect 1757 13085 1791 13097
rect 3287 13097 3321 13119
rect 3287 13085 3321 13097
rect 5224 13343 5258 13377
rect 4131 13194 4137 13228
rect 4137 13194 4165 13228
rect 4131 13106 4137 13140
rect 4137 13106 4165 13140
rect 5224 13268 5258 13302
rect 5224 13193 5258 13227
rect 4819 13115 4853 13149
rect 4891 13115 4925 13149
rect 4963 13115 4997 13149
rect 5224 13118 5258 13152
rect 1197 13020 1231 13043
rect 1197 13009 1231 13020
rect 1197 12950 1231 12970
rect 1197 12936 1231 12950
rect 1197 12880 1231 12897
rect 1197 12863 1231 12880
rect 1197 12810 1231 12824
rect 1197 12790 1231 12810
rect 1197 12740 1231 12751
rect 1197 12717 1231 12740
rect 1197 12670 1231 12678
rect 1197 12644 1231 12670
rect 1197 12599 1231 12605
rect 1197 12571 1231 12599
rect 1197 12528 1231 12532
rect 1197 12498 1231 12528
rect 1357 13010 1391 13044
rect 1357 12938 1391 12972
rect 1357 12866 1391 12900
rect 1357 12794 1391 12828
rect 1357 12721 1391 12755
rect 1357 12648 1391 12682
rect 1357 12575 1391 12609
rect 1357 12502 1391 12536
rect 1613 13010 1647 13044
rect 1613 12938 1647 12972
rect 1613 12866 1647 12900
rect 1613 12794 1647 12828
rect 1613 12721 1647 12755
rect 1613 12648 1647 12682
rect 1613 12575 1647 12609
rect 1613 12502 1647 12536
rect 1757 13027 1791 13045
rect 1757 13011 1791 13027
rect 3287 13027 3321 13045
rect 3287 13011 3321 13027
rect 3419 13022 3453 13056
rect 3491 13022 3525 13056
rect 3563 13022 3597 13056
rect 1757 12957 1791 12971
rect 1757 12937 1791 12957
rect 3287 12957 3321 12971
rect 3287 12937 3321 12957
rect 1757 12888 1791 12897
rect 1757 12863 1791 12888
rect 3287 12888 3321 12897
rect 3287 12863 3321 12888
rect 4131 12938 4137 12972
rect 4137 12938 4165 12972
rect 4131 12850 4137 12884
rect 4137 12850 4165 12884
rect 4538 12860 4572 12894
rect 4610 12860 4644 12894
rect 4682 12860 4716 12894
rect 5224 13043 5258 13077
rect 5224 12968 5258 13002
rect 5224 12893 5258 12927
rect 1757 12819 1791 12823
rect 1757 12789 1791 12819
rect 3287 12819 3321 12823
rect 3287 12789 3321 12819
rect 1757 12716 1791 12749
rect 1757 12715 1791 12716
rect 3287 12716 3321 12749
rect 3287 12715 3321 12716
rect 1757 12647 1791 12675
rect 1757 12641 1791 12647
rect 3287 12647 3321 12675
rect 3287 12641 3321 12647
rect 1757 12578 1791 12601
rect 1757 12567 1791 12578
rect 3700 12766 3734 12800
rect 3772 12766 3806 12800
rect 3844 12766 3878 12800
rect 4251 12776 4279 12810
rect 4279 12776 4285 12810
rect 4251 12688 4279 12722
rect 4279 12688 4285 12722
rect 5380 13793 5414 13827
rect 5380 13718 5414 13752
rect 5380 13643 5414 13677
rect 5380 13568 5414 13602
rect 5380 13493 5414 13527
rect 5380 13418 5414 13452
rect 5380 13343 5414 13377
rect 5380 13268 5414 13302
rect 5380 13193 5414 13227
rect 5380 13118 5414 13152
rect 5380 13043 5414 13077
rect 5380 12968 5414 13002
rect 5380 12893 5414 12927
rect 5536 13795 5570 13829
rect 5536 13719 5570 13753
rect 5536 13643 5570 13677
rect 5536 13568 5570 13602
rect 5536 13493 5570 13527
rect 5536 13418 5570 13452
rect 5536 13343 5570 13377
rect 5536 13268 5570 13302
rect 5536 13193 5570 13227
rect 5536 13118 5570 13152
rect 5536 13043 5570 13077
rect 5536 12968 5570 13002
rect 5536 12893 5570 12927
rect 5692 13793 5726 13827
rect 5692 13718 5726 13752
rect 5692 13643 5726 13677
rect 5692 13568 5726 13602
rect 5692 13493 5726 13527
rect 5692 13418 5726 13452
rect 5692 13343 5726 13377
rect 5692 13268 5726 13302
rect 5692 13193 5726 13227
rect 5692 13118 5726 13152
rect 5692 13043 5726 13077
rect 5692 12968 5726 13002
rect 5692 12893 5726 12927
rect 6378 13884 6412 13918
rect 6450 13884 6484 13918
rect 6522 13884 6556 13918
rect 7761 13937 7795 13943
rect 7761 13909 7795 13937
rect 9291 13937 9325 13943
rect 9291 13909 9325 13937
rect 7761 13867 7795 13868
rect 5848 13795 5882 13829
rect 5848 13719 5882 13753
rect 5848 13643 5882 13677
rect 6091 13800 6119 13834
rect 6119 13800 6125 13834
rect 6091 13712 6119 13746
rect 6119 13712 6125 13746
rect 7761 13834 7795 13867
rect 9291 13867 9325 13868
rect 9291 13834 9325 13867
rect 7216 13790 7250 13824
rect 7288 13790 7322 13824
rect 7360 13790 7394 13824
rect 7761 13763 7795 13793
rect 7761 13759 7795 13763
rect 9291 13763 9325 13793
rect 9291 13759 9325 13763
rect 6097 13628 6131 13662
rect 6169 13628 6203 13662
rect 6241 13628 6275 13662
rect 6929 13706 6957 13740
rect 6957 13706 6963 13740
rect 5848 13568 5882 13602
rect 6929 13618 6957 13652
rect 6957 13618 6963 13652
rect 5848 13493 5882 13527
rect 5848 13418 5882 13452
rect 5848 13343 5882 13377
rect 6378 13372 6412 13406
rect 6450 13372 6484 13406
rect 6522 13372 6556 13406
rect 7761 13693 7795 13718
rect 7761 13684 7795 13693
rect 9291 13693 9325 13718
rect 9291 13684 9325 13693
rect 7761 13623 7795 13643
rect 7761 13609 7795 13623
rect 9291 13623 9325 13643
rect 9291 13609 9325 13623
rect 7497 13534 7531 13568
rect 7569 13534 7603 13568
rect 7641 13534 7675 13568
rect 7761 13553 7795 13568
rect 7761 13534 7795 13553
rect 9291 13553 9325 13568
rect 9291 13534 9325 13553
rect 6929 13484 6963 13485
rect 6929 13451 6957 13484
rect 6957 13451 6963 13484
rect 6929 13396 6963 13397
rect 6929 13363 6957 13396
rect 6957 13363 6963 13396
rect 5848 13268 5882 13302
rect 5848 13193 5882 13227
rect 5848 13118 5882 13152
rect 6659 13115 6693 13149
rect 6731 13115 6765 13149
rect 6803 13115 6837 13149
rect 7761 13483 7795 13493
rect 7761 13459 7795 13483
rect 9291 13483 9325 13493
rect 9291 13459 9325 13483
rect 7761 13413 7795 13418
rect 7761 13384 7795 13413
rect 9291 13413 9325 13418
rect 9291 13384 9325 13413
rect 7216 13278 7250 13312
rect 7288 13278 7322 13312
rect 7360 13278 7394 13312
rect 7761 13309 7795 13343
rect 9291 13309 9325 13343
rect 6929 13194 6957 13228
rect 6957 13194 6963 13228
rect 6929 13106 6957 13140
rect 6957 13106 6963 13140
rect 5848 13043 5882 13077
rect 5848 12968 5882 13002
rect 5848 12893 5882 12927
rect 6378 12860 6412 12894
rect 6450 12860 6484 12894
rect 6522 12860 6556 12894
rect 7761 13237 7795 13268
rect 7761 13234 7795 13237
rect 9291 13237 9325 13268
rect 9291 13234 9325 13237
rect 7761 13167 7795 13193
rect 7761 13159 7795 13167
rect 9291 13167 9325 13193
rect 9291 13159 9325 13167
rect 7761 13097 7795 13119
rect 7761 13085 7795 13097
rect 9291 13097 9325 13119
rect 9291 13085 9325 13097
rect 7497 13022 7531 13056
rect 7569 13022 7603 13056
rect 7641 13022 7675 13056
rect 7761 13027 7795 13045
rect 7761 13011 7795 13027
rect 9291 13027 9325 13045
rect 9291 13011 9325 13027
rect 6929 12938 6957 12972
rect 6957 12938 6963 12972
rect 6929 12850 6957 12884
rect 6957 12850 6963 12884
rect 7761 12957 7795 12971
rect 7761 12937 7795 12957
rect 9291 12957 9325 12971
rect 9291 12937 9325 12957
rect 7761 12888 7795 12897
rect 7761 12863 7795 12888
rect 9291 12888 9325 12897
rect 9291 12863 9325 12888
rect 6091 12776 6119 12810
rect 6119 12776 6125 12810
rect 3700 12610 3734 12644
rect 3772 12610 3806 12644
rect 3844 12610 3878 12644
rect 3287 12578 3321 12601
rect 4481 12604 4515 12638
rect 3287 12567 3321 12578
rect 1757 12509 1791 12527
rect 1757 12493 1791 12509
rect 3287 12509 3321 12527
rect 3287 12493 3321 12509
rect 6091 12688 6119 12722
rect 6119 12688 6125 12722
rect 7761 12819 7795 12823
rect 7216 12766 7250 12800
rect 7288 12766 7322 12800
rect 7360 12766 7394 12800
rect 4481 12516 4515 12550
rect 1197 12457 1231 12459
rect 1197 12425 1231 12457
rect 1440 12424 1456 12458
rect 1456 12424 1474 12458
rect 1529 12424 1552 12458
rect 1552 12424 1563 12458
rect 1984 12448 2018 12482
rect 2059 12448 2093 12482
rect 2134 12448 2168 12482
rect 2209 12448 2243 12482
rect 2284 12448 2318 12482
rect 2359 12448 2393 12482
rect 2434 12448 2468 12482
rect 2509 12448 2543 12482
rect 2584 12448 2618 12482
rect 2659 12448 2693 12482
rect 2734 12448 2768 12482
rect 2809 12448 2843 12482
rect 2884 12448 2918 12482
rect 2959 12448 2993 12482
rect 3033 12448 3067 12482
rect 4608 12448 4642 12482
rect 4682 12448 4716 12482
rect 5457 12626 5491 12660
rect 5457 12526 5491 12560
rect 5614 12626 5648 12660
rect 5614 12526 5648 12560
rect 6321 12604 6355 12638
rect 7216 12610 7250 12644
rect 7288 12610 7322 12644
rect 7360 12610 7394 12644
rect 7761 12789 7795 12819
rect 9291 12819 9325 12823
rect 9291 12789 9325 12819
rect 7761 12716 7795 12749
rect 7761 12715 7795 12716
rect 9291 12716 9325 12749
rect 9397 13978 9431 14012
rect 9471 13978 9495 14012
rect 9495 13978 9505 14012
rect 9544 13978 9563 14012
rect 9563 13978 9578 14012
rect 9617 13978 9631 14012
rect 9631 13978 9651 14012
rect 9690 13978 9699 14012
rect 9699 13978 9724 14012
rect 9763 13978 9767 14012
rect 9767 13978 9797 14012
rect 9869 13946 9903 13980
rect 9365 13876 9399 13908
rect 9365 13874 9399 13876
rect 9522 13887 9556 13921
rect 9617 13887 9651 13921
rect 9712 13887 9746 13921
rect 9365 13808 9399 13836
rect 9365 13802 9399 13808
rect 9869 13873 9903 13907
rect 9365 13740 9399 13764
rect 9365 13730 9399 13740
rect 9365 13672 9399 13692
rect 9365 13658 9399 13672
rect 9365 13604 9399 13620
rect 9365 13586 9399 13604
rect 9365 13536 9399 13547
rect 9365 13513 9399 13536
rect 9365 13468 9399 13474
rect 9365 13440 9399 13468
rect 9365 13400 9399 13401
rect 9365 13367 9399 13400
rect 9365 13298 9399 13328
rect 9365 13294 9399 13298
rect 9365 13230 9399 13255
rect 9365 13221 9399 13230
rect 9365 13162 9399 13182
rect 9365 13148 9399 13162
rect 9365 13094 9399 13109
rect 9365 13075 9399 13094
rect 9365 13026 9399 13036
rect 9365 13002 9399 13026
rect 9365 12958 9399 12963
rect 9365 12929 9399 12958
rect 9461 13793 9495 13827
rect 9461 13720 9495 13754
rect 9461 13647 9495 13681
rect 9461 13574 9495 13608
rect 9461 13501 9495 13535
rect 9461 13427 9495 13461
rect 9461 13353 9495 13387
rect 9461 13279 9495 13313
rect 9461 13205 9495 13239
rect 9461 13131 9495 13165
rect 9461 13057 9495 13091
rect 9461 12983 9495 13017
rect 9461 12909 9495 12943
rect 9618 13793 9652 13827
rect 9618 13720 9652 13754
rect 9618 13647 9652 13681
rect 9618 13574 9652 13608
rect 9618 13501 9652 13535
rect 9618 13427 9652 13461
rect 9618 13353 9652 13387
rect 9618 13279 9652 13313
rect 9618 13205 9652 13239
rect 9618 13131 9652 13165
rect 9618 13057 9652 13091
rect 9618 12983 9652 13017
rect 9618 12909 9652 12943
rect 9773 13793 9807 13827
rect 9773 13720 9807 13754
rect 9773 13647 9807 13681
rect 9773 13574 9807 13608
rect 9773 13501 9807 13535
rect 9773 13427 9807 13461
rect 9773 13353 9807 13387
rect 9773 13279 9807 13313
rect 9773 13205 9807 13239
rect 9773 13131 9807 13165
rect 9773 13057 9807 13091
rect 9773 12983 9807 13017
rect 9773 12909 9807 12943
rect 9869 13805 9903 13834
rect 9869 13800 9903 13805
rect 9869 13737 9903 13761
rect 9869 13727 9903 13737
rect 9869 13669 9903 13688
rect 9869 13654 9903 13669
rect 9869 13601 9903 13615
rect 9869 13581 9903 13601
rect 9869 13533 9903 13542
rect 9869 13508 9903 13533
rect 9869 13465 9903 13469
rect 9869 13435 9903 13465
rect 9869 13363 9903 13396
rect 9869 13362 9903 13363
rect 9869 13295 9903 13323
rect 9869 13289 9903 13295
rect 9869 13227 9903 13250
rect 9869 13216 9903 13227
rect 9869 13159 9903 13177
rect 9869 13143 9903 13159
rect 9869 13091 9903 13105
rect 9869 13071 9903 13091
rect 9869 13023 9903 13033
rect 9869 12999 9903 13023
rect 9869 12955 9903 12961
rect 9869 12927 9903 12955
rect 9365 12856 9399 12890
rect 9365 12783 9399 12817
rect 9869 12887 9903 12889
rect 9869 12855 9903 12887
rect 9483 12751 9501 12785
rect 9501 12751 9517 12785
rect 9742 12751 9773 12785
rect 9773 12751 9776 12785
rect 9837 12751 9871 12785
rect 11077 14014 11111 14030
rect 11077 13962 11111 13974
rect 11077 13940 11111 13962
rect 11077 13894 11111 13900
rect 11077 13866 11111 13894
rect 11077 13792 11111 13826
rect 11077 13724 11111 13752
rect 11077 13718 11111 13724
rect 11077 13656 11111 13678
rect 11077 13644 11111 13656
rect 11077 13588 11111 13604
rect 11077 13570 11111 13588
rect 11077 13520 11111 13530
rect 11077 13496 11111 13520
rect 11077 13452 11111 13456
rect 11077 13422 11111 13452
rect 11077 13350 11111 13382
rect 11077 13348 11111 13350
rect 11077 13282 11111 13308
rect 11077 13274 11111 13282
rect 11077 13214 11111 13234
rect 11077 13200 11111 13214
rect 11077 13126 11111 13160
rect 11077 13052 11111 13086
rect 11077 12980 11111 13012
rect 11077 12978 11111 12980
rect 11077 12910 11111 12938
rect 11077 12904 11111 12910
rect 11077 12840 11111 12864
rect 11077 12830 11111 12840
rect 11077 12770 11111 12790
rect 11077 12756 11111 12770
rect 9291 12715 9325 12716
rect 7761 12647 7795 12675
rect 7761 12641 7795 12647
rect 9291 12647 9325 12675
rect 9291 12641 9325 12647
rect 6321 12516 6355 12550
rect 5500 12424 5502 12458
rect 5502 12424 5534 12458
rect 5572 12424 5604 12458
rect 5604 12424 5606 12458
rect 6448 12448 6482 12482
rect 6522 12448 6556 12482
rect 7761 12578 7795 12601
rect 7761 12567 7795 12578
rect 9291 12578 9325 12601
rect 9291 12567 9325 12578
rect 7761 12509 7795 12527
rect 7761 12493 7795 12509
rect 9291 12509 9325 12527
rect 9291 12493 9325 12509
rect 9453 12675 9487 12709
rect 9783 12690 9817 12709
rect 9783 12675 9815 12690
rect 9815 12675 9817 12690
rect 9453 12597 9487 12631
rect 9783 12617 9817 12631
rect 9783 12597 9815 12617
rect 9815 12597 9817 12617
rect 9453 12519 9487 12553
rect 9783 12543 9817 12553
rect 9783 12519 9815 12543
rect 9815 12519 9817 12543
rect 8015 12448 8049 12482
rect 8089 12448 8123 12482
rect 8164 12448 8198 12482
rect 8239 12448 8273 12482
rect 8314 12448 8348 12482
rect 8389 12448 8423 12482
rect 8464 12448 8498 12482
rect 8539 12448 8573 12482
rect 8614 12448 8648 12482
rect 8689 12448 8723 12482
rect 8764 12448 8798 12482
rect 8839 12448 8873 12482
rect 8914 12448 8948 12482
rect 8989 12448 9023 12482
rect 9064 12448 9098 12482
rect 9453 12441 9487 12475
rect 9783 12469 9817 12475
rect 9783 12441 9815 12469
rect 9815 12441 9817 12469
rect 11077 12700 11111 12716
rect 11077 12682 11111 12700
rect 11077 12630 11111 12642
rect 11077 12608 11111 12630
rect 11077 12560 11111 12568
rect 11077 12534 11111 12560
rect 11077 12490 11111 12494
rect 11077 12460 11111 12490
rect 11077 12386 11111 12420
rect 1197 12352 1231 12386
rect 3612 12352 3645 12386
rect 3645 12352 3646 12386
rect 3693 12352 3713 12386
rect 3713 12352 3727 12386
rect 3774 12352 3781 12386
rect 3781 12352 3808 12386
rect 3855 12352 3883 12386
rect 3883 12352 3889 12386
rect 3936 12352 3951 12386
rect 3951 12352 3970 12386
rect 4017 12352 4019 12386
rect 4019 12352 4051 12386
rect 4097 12352 4121 12386
rect 4121 12352 4131 12386
rect 5087 12352 5107 12381
rect 5107 12352 5121 12381
rect 5162 12352 5175 12381
rect 5175 12352 5196 12381
rect 5237 12352 5243 12381
rect 5243 12352 5271 12381
rect 5312 12352 5345 12381
rect 5345 12352 5346 12381
rect 5386 12352 5413 12381
rect 5413 12352 5420 12381
rect 5460 12352 5481 12381
rect 5481 12352 5494 12381
rect 5534 12352 5549 12381
rect 5549 12352 5568 12381
rect 5608 12352 5617 12381
rect 5617 12352 5642 12381
rect 5682 12352 5685 12381
rect 5685 12352 5716 12381
rect 5756 12352 5787 12381
rect 5787 12352 5790 12381
rect 5830 12352 5855 12381
rect 5855 12352 5864 12381
rect 5904 12352 5923 12381
rect 5923 12352 5938 12381
rect 5978 12352 5991 12381
rect 5991 12352 6012 12381
rect 6899 12352 6909 12386
rect 6909 12352 6933 12386
rect 6978 12352 7011 12386
rect 7011 12352 7012 12386
rect 7058 12352 7079 12386
rect 7079 12352 7092 12386
rect 7138 12352 7147 12386
rect 7147 12352 7172 12386
rect 7218 12352 7249 12386
rect 7249 12352 7252 12386
rect 7298 12352 7317 12386
rect 7317 12352 7332 12386
rect 7378 12352 7385 12386
rect 7385 12352 7412 12386
rect 7458 12352 7487 12386
rect 7487 12352 7492 12386
rect 7802 12352 7827 12380
rect 7827 12352 7836 12380
rect 7874 12352 7895 12380
rect 7895 12352 7908 12380
rect 7946 12352 7963 12380
rect 7963 12352 7980 12380
rect 8018 12352 8031 12380
rect 8031 12352 8052 12380
rect 8090 12352 8099 12380
rect 8099 12352 8124 12380
rect 8162 12352 8167 12380
rect 8167 12352 8196 12380
rect 8234 12352 8235 12380
rect 8235 12352 8268 12380
rect 8306 12352 8337 12380
rect 8337 12352 8340 12380
rect 8378 12352 8405 12380
rect 8405 12352 8412 12380
rect 8450 12352 8473 12380
rect 8473 12352 8484 12380
rect 8522 12352 8541 12380
rect 8541 12352 8556 12380
rect 8594 12352 8609 12380
rect 8609 12352 8628 12380
rect 8666 12352 8677 12380
rect 8677 12352 8700 12380
rect 8738 12352 8745 12380
rect 8745 12352 8772 12380
rect 8810 12352 8813 12380
rect 8813 12352 8844 12380
rect 8882 12352 8915 12380
rect 8915 12352 8916 12380
rect 8954 12352 8983 12380
rect 8983 12352 8988 12380
rect 9026 12352 9052 12380
rect 9052 12352 9060 12380
rect 9098 12352 9121 12380
rect 9121 12352 9132 12380
rect 9170 12352 9190 12380
rect 9190 12352 9204 12380
rect 9242 12352 9259 12380
rect 9259 12352 9276 12380
rect 9314 12352 9328 12380
rect 9328 12352 9348 12380
rect 9386 12352 9397 12380
rect 9397 12352 9420 12380
rect 9458 12352 9466 12380
rect 9466 12352 9492 12380
rect 9530 12352 9535 12380
rect 9535 12352 9564 12380
rect 9602 12352 9604 12380
rect 9604 12352 9636 12380
rect 9674 12352 9707 12380
rect 9707 12352 9708 12380
rect 9747 12352 9776 12380
rect 9776 12352 9781 12380
rect 9820 12352 9845 12380
rect 9845 12352 9854 12380
rect 9893 12352 9914 12380
rect 9914 12352 9927 12380
rect 9966 12352 9983 12380
rect 9983 12352 10000 12380
rect 10065 12352 10087 12380
rect 10087 12352 10099 12380
rect 10141 12352 10156 12380
rect 10156 12352 10175 12380
rect 10217 12352 10225 12380
rect 10225 12352 10251 12380
rect 10293 12352 10294 12380
rect 10294 12352 10327 12380
rect 10369 12352 10397 12380
rect 10397 12352 10403 12380
rect 10446 12352 10466 12380
rect 10466 12352 10480 12380
rect 10523 12352 10535 12380
rect 10535 12352 10557 12380
rect 10600 12352 10617 12380
rect 10617 12352 10634 12380
rect 10677 12352 10693 12380
rect 10693 12352 10711 12380
rect 10754 12352 10769 12380
rect 10769 12352 10788 12380
rect 10831 12352 10845 12380
rect 10845 12352 10865 12380
rect 10908 12352 10920 12380
rect 10920 12352 10942 12380
rect 5087 12347 5121 12352
rect 5162 12347 5196 12352
rect 5237 12347 5271 12352
rect 5312 12347 5346 12352
rect 5386 12347 5420 12352
rect 5460 12347 5494 12352
rect 5534 12347 5568 12352
rect 5608 12347 5642 12352
rect 5682 12347 5716 12352
rect 5756 12347 5790 12352
rect 5830 12347 5864 12352
rect 5904 12347 5938 12352
rect 5978 12347 6012 12352
rect 7802 12346 7836 12352
rect 7874 12346 7908 12352
rect 7946 12346 7980 12352
rect 8018 12346 8052 12352
rect 8090 12346 8124 12352
rect 8162 12346 8196 12352
rect 8234 12346 8268 12352
rect 8306 12346 8340 12352
rect 8378 12346 8412 12352
rect 8450 12346 8484 12352
rect 8522 12346 8556 12352
rect 8594 12346 8628 12352
rect 8666 12346 8700 12352
rect 8738 12346 8772 12352
rect 8810 12346 8844 12352
rect 8882 12346 8916 12352
rect 8954 12346 8988 12352
rect 9026 12346 9060 12352
rect 9098 12346 9132 12352
rect 9170 12346 9204 12352
rect 9242 12346 9276 12352
rect 9314 12346 9348 12352
rect 9386 12346 9420 12352
rect 9458 12346 9492 12352
rect 9530 12346 9564 12352
rect 9602 12346 9636 12352
rect 9674 12346 9708 12352
rect 9747 12346 9781 12352
rect 9820 12346 9854 12352
rect 9893 12346 9927 12352
rect 9966 12346 10000 12352
rect 10065 12346 10099 12352
rect 10141 12346 10175 12352
rect 10217 12346 10251 12352
rect 10293 12346 10327 12352
rect 10369 12346 10403 12352
rect 10446 12346 10480 12352
rect 10523 12346 10557 12352
rect 10600 12346 10634 12352
rect 10677 12346 10711 12352
rect 10754 12346 10788 12352
rect 10831 12346 10865 12352
rect 10908 12346 10942 12352
rect 1651 12171 1685 12175
rect 1743 12171 1777 12175
rect 1836 12171 1870 12175
rect 1929 12171 1963 12175
rect 2287 12171 2321 12175
rect 2363 12171 2397 12175
rect 2439 12171 2473 12175
rect 2515 12171 2549 12175
rect 2592 12171 2626 12175
rect 2669 12171 2703 12175
rect 2746 12171 2780 12175
rect 2823 12171 2857 12175
rect 2900 12171 2934 12175
rect 2977 12171 3011 12175
rect 3054 12171 3088 12175
rect 3131 12171 3165 12175
rect 3208 12171 3242 12175
rect 3285 12171 3319 12175
rect 5077 12171 5111 12175
rect 5154 12171 5188 12175
rect 5231 12171 5265 12175
rect 5308 12171 5342 12175
rect 5385 12171 5419 12175
rect 5463 12171 5497 12175
rect 5541 12171 5575 12175
rect 5619 12171 5653 12175
rect 5697 12171 5731 12175
rect 5775 12171 5809 12175
rect 5853 12171 5887 12175
rect 5931 12171 5965 12175
rect 6889 12171 6923 12175
rect 6971 12171 7005 12175
rect 7053 12171 7087 12175
rect 7135 12171 7169 12175
rect 7218 12171 7252 12175
rect 7301 12171 7335 12175
rect 7384 12171 7418 12175
rect 7803 12171 7837 12175
rect 7876 12171 7910 12175
rect 7949 12171 7983 12175
rect 8022 12171 8056 12175
rect 8095 12171 8129 12175
rect 8168 12171 8202 12175
rect 8241 12171 8275 12175
rect 8314 12171 8348 12175
rect 8387 12171 8421 12175
rect 8460 12171 8494 12175
rect 8533 12171 8567 12175
rect 8606 12171 8640 12175
rect 8680 12171 8714 12175
rect 8754 12171 8788 12175
rect 8828 12171 8862 12175
rect 9422 12171 9456 12175
rect 9501 12171 9535 12175
rect 9580 12171 9614 12175
rect 9659 12171 9693 12175
rect 9739 12171 9773 12175
rect 9819 12171 9853 12175
rect 10007 12171 10041 12175
rect 10082 12171 10116 12175
rect 10157 12171 10191 12175
rect 10233 12171 10267 12175
rect 10483 12171 10517 12175
rect 10558 12171 10592 12175
rect 10633 12171 10667 12175
rect 10709 12171 10743 12175
rect 10785 12171 10819 12175
rect 10861 12171 10895 12175
rect 10937 12171 10971 12175
rect 11013 12171 11047 12175
rect 11089 12171 11123 12175
rect 1651 12141 1676 12171
rect 1676 12141 1685 12171
rect 1743 12141 1745 12171
rect 1745 12141 1777 12171
rect 1836 12141 1849 12171
rect 1849 12141 1870 12171
rect 1929 12141 1952 12171
rect 1952 12141 1963 12171
rect 2287 12141 2297 12171
rect 2297 12141 2321 12171
rect 2363 12141 2366 12171
rect 2366 12141 2397 12171
rect 2439 12141 2470 12171
rect 2470 12141 2473 12171
rect 2515 12141 2539 12171
rect 2539 12141 2549 12171
rect 2592 12141 2608 12171
rect 2608 12141 2626 12171
rect 2669 12141 2677 12171
rect 2677 12141 2703 12171
rect 2746 12141 2780 12171
rect 2823 12141 2849 12171
rect 2849 12141 2857 12171
rect 2900 12141 2918 12171
rect 2918 12141 2934 12171
rect 2977 12141 2987 12171
rect 2987 12141 3011 12171
rect 3054 12141 3056 12171
rect 3056 12141 3088 12171
rect 3131 12141 3160 12171
rect 3160 12141 3165 12171
rect 3208 12141 3229 12171
rect 3229 12141 3242 12171
rect 3285 12141 3298 12171
rect 3298 12141 3319 12171
rect 5077 12141 5111 12171
rect 5154 12141 5188 12171
rect 5231 12141 5265 12171
rect 5308 12141 5342 12171
rect 5385 12141 5419 12171
rect 5463 12141 5497 12171
rect 5541 12141 5575 12171
rect 5619 12141 5653 12171
rect 5697 12141 5731 12171
rect 5775 12141 5809 12171
rect 5853 12141 5887 12171
rect 5931 12141 5965 12171
rect 6889 12141 6923 12171
rect 6971 12141 7005 12171
rect 7053 12141 7087 12171
rect 7135 12141 7169 12171
rect 7218 12141 7252 12171
rect 7301 12141 7335 12171
rect 7384 12141 7418 12171
rect 7803 12141 7837 12171
rect 7876 12141 7910 12171
rect 7949 12141 7983 12171
rect 8022 12141 8056 12171
rect 8095 12141 8129 12171
rect 8168 12141 8202 12171
rect 8241 12141 8275 12171
rect 8314 12141 8348 12171
rect 8387 12141 8421 12171
rect 8460 12141 8494 12171
rect 8533 12141 8567 12171
rect 8606 12141 8640 12171
rect 8680 12141 8714 12171
rect 8754 12141 8788 12171
rect 8828 12141 8862 12171
rect 9422 12141 9456 12171
rect 9501 12141 9535 12171
rect 9580 12141 9614 12171
rect 9659 12141 9693 12171
rect 9739 12141 9773 12171
rect 9819 12141 9853 12171
rect 10007 12141 10041 12171
rect 10082 12141 10116 12171
rect 10157 12141 10191 12171
rect 10233 12141 10267 12171
rect 10483 12141 10517 12171
rect 10558 12141 10592 12171
rect 10633 12141 10667 12171
rect 10709 12141 10743 12171
rect 10785 12141 10819 12171
rect 10861 12141 10895 12171
rect 10937 12141 10971 12171
rect 11013 12141 11047 12171
rect 11089 12141 11094 12171
rect 11094 12141 11123 12171
rect 11165 12141 11199 12175
rect 1651 12069 1676 12103
rect 1676 12069 1685 12103
rect 1743 12069 1745 12103
rect 1745 12069 1777 12103
rect 1836 12069 1849 12103
rect 1849 12069 1870 12103
rect 1929 12069 1952 12103
rect 1952 12069 1963 12103
rect 2287 12069 2297 12103
rect 2297 12069 2321 12103
rect 2363 12069 2366 12103
rect 2366 12069 2397 12103
rect 2439 12069 2470 12103
rect 2470 12069 2473 12103
rect 2515 12069 2539 12103
rect 2539 12069 2549 12103
rect 2592 12069 2608 12103
rect 2608 12069 2626 12103
rect 2669 12069 2677 12103
rect 2677 12069 2703 12103
rect 2746 12069 2780 12103
rect 2823 12069 2849 12103
rect 2849 12069 2857 12103
rect 2900 12069 2918 12103
rect 2918 12069 2934 12103
rect 2977 12069 2987 12103
rect 2987 12069 3011 12103
rect 3054 12069 3056 12103
rect 3056 12069 3088 12103
rect 3131 12069 3160 12103
rect 3160 12069 3165 12103
rect 3208 12069 3229 12103
rect 3229 12069 3242 12103
rect 3285 12069 3298 12103
rect 3298 12069 3319 12103
rect 5077 12069 5111 12103
rect 5154 12069 5188 12103
rect 5231 12069 5265 12103
rect 5308 12069 5342 12103
rect 5385 12069 5419 12103
rect 5463 12069 5497 12103
rect 5541 12069 5575 12103
rect 5619 12069 5653 12103
rect 5697 12069 5731 12103
rect 5775 12069 5809 12103
rect 5853 12069 5887 12103
rect 5931 12069 5965 12103
rect 6889 12069 6923 12103
rect 6971 12069 7005 12103
rect 7053 12069 7087 12103
rect 7135 12069 7169 12103
rect 7218 12069 7252 12103
rect 7301 12069 7335 12103
rect 7384 12069 7418 12103
rect 7803 12069 7837 12103
rect 7876 12069 7910 12103
rect 7949 12069 7983 12103
rect 8022 12069 8056 12103
rect 8095 12069 8129 12103
rect 8168 12069 8202 12103
rect 8241 12069 8275 12103
rect 8314 12069 8348 12103
rect 8387 12069 8421 12103
rect 8460 12069 8494 12103
rect 8533 12069 8567 12103
rect 8606 12069 8640 12103
rect 8680 12069 8714 12103
rect 8754 12069 8788 12103
rect 8828 12069 8862 12103
rect 9422 12069 9456 12103
rect 9501 12069 9535 12103
rect 9580 12069 9614 12103
rect 9659 12069 9693 12103
rect 9739 12069 9773 12103
rect 9819 12069 9853 12103
rect 10007 12069 10041 12103
rect 10082 12069 10116 12103
rect 10157 12069 10191 12103
rect 10233 12069 10267 12103
rect 10483 12069 10517 12103
rect 10558 12069 10592 12103
rect 10633 12069 10667 12103
rect 10709 12069 10743 12103
rect 10785 12069 10819 12103
rect 10861 12069 10895 12103
rect 10937 12069 10971 12103
rect 11013 12069 11047 12103
rect 11089 12069 11094 12103
rect 11094 12069 11123 12103
rect 11165 12069 11199 12103
rect 1651 12001 1676 12031
rect 1676 12001 1685 12031
rect 1743 12001 1745 12031
rect 1745 12001 1777 12031
rect 1836 12001 1849 12031
rect 1849 12001 1870 12031
rect 1929 12001 1952 12031
rect 1952 12001 1963 12031
rect 2287 12001 2297 12031
rect 2297 12001 2321 12031
rect 2363 12001 2366 12031
rect 2366 12001 2397 12031
rect 2439 12001 2470 12031
rect 2470 12001 2473 12031
rect 2515 12001 2539 12031
rect 2539 12001 2549 12031
rect 2592 12001 2608 12031
rect 2608 12001 2626 12031
rect 2669 12001 2677 12031
rect 2677 12001 2703 12031
rect 2746 12001 2780 12031
rect 2823 12001 2849 12031
rect 2849 12001 2857 12031
rect 2900 12001 2918 12031
rect 2918 12001 2934 12031
rect 2977 12001 2987 12031
rect 2987 12001 3011 12031
rect 3054 12001 3056 12031
rect 3056 12001 3088 12031
rect 3131 12001 3160 12031
rect 3160 12001 3165 12031
rect 3208 12001 3229 12031
rect 3229 12001 3242 12031
rect 3285 12001 3298 12031
rect 3298 12001 3319 12031
rect 5077 12001 5111 12031
rect 5154 12001 5188 12031
rect 5231 12001 5265 12031
rect 5308 12001 5342 12031
rect 5385 12001 5419 12031
rect 5463 12001 5497 12031
rect 5541 12001 5575 12031
rect 5619 12001 5653 12031
rect 5697 12001 5731 12031
rect 5775 12001 5809 12031
rect 5853 12001 5887 12031
rect 5931 12001 5965 12031
rect 6889 12001 6923 12031
rect 6971 12001 7005 12031
rect 7053 12001 7087 12031
rect 7135 12001 7169 12031
rect 7218 12001 7252 12031
rect 7301 12001 7335 12031
rect 7384 12001 7418 12031
rect 7803 12001 7837 12031
rect 7876 12001 7910 12031
rect 7949 12001 7983 12031
rect 8022 12001 8056 12031
rect 8095 12001 8129 12031
rect 8168 12001 8202 12031
rect 8241 12001 8275 12031
rect 8314 12001 8348 12031
rect 8387 12001 8421 12031
rect 8460 12001 8494 12031
rect 8533 12001 8567 12031
rect 8606 12001 8640 12031
rect 8680 12001 8714 12031
rect 8754 12001 8788 12031
rect 8828 12001 8862 12031
rect 9422 12001 9456 12031
rect 9501 12001 9535 12031
rect 9580 12001 9614 12031
rect 9659 12001 9693 12031
rect 9739 12001 9773 12031
rect 9819 12001 9853 12031
rect 10007 12001 10041 12031
rect 10082 12001 10116 12031
rect 10157 12001 10191 12031
rect 10233 12001 10267 12031
rect 10483 12001 10517 12031
rect 10558 12001 10592 12031
rect 10633 12001 10667 12031
rect 10709 12001 10743 12031
rect 10785 12001 10819 12031
rect 10861 12001 10895 12031
rect 10937 12001 10971 12031
rect 11013 12001 11047 12031
rect 11089 12001 11094 12031
rect 11094 12001 11123 12031
rect 1651 11997 1685 12001
rect 1743 11997 1777 12001
rect 1836 11997 1870 12001
rect 1929 11997 1963 12001
rect 2287 11997 2321 12001
rect 2363 11997 2397 12001
rect 2439 11997 2473 12001
rect 2515 11997 2549 12001
rect 2592 11997 2626 12001
rect 2669 11997 2703 12001
rect 2746 11997 2780 12001
rect 2823 11997 2857 12001
rect 2900 11997 2934 12001
rect 2977 11997 3011 12001
rect 3054 11997 3088 12001
rect 3131 11997 3165 12001
rect 3208 11997 3242 12001
rect 3285 11997 3319 12001
rect 5077 11997 5111 12001
rect 5154 11997 5188 12001
rect 5231 11997 5265 12001
rect 5308 11997 5342 12001
rect 5385 11997 5419 12001
rect 5463 11997 5497 12001
rect 5541 11997 5575 12001
rect 5619 11997 5653 12001
rect 5697 11997 5731 12001
rect 5775 11997 5809 12001
rect 5853 11997 5887 12001
rect 5931 11997 5965 12001
rect 6889 11997 6923 12001
rect 6971 11997 7005 12001
rect 7053 11997 7087 12001
rect 7135 11997 7169 12001
rect 7218 11997 7252 12001
rect 7301 11997 7335 12001
rect 7384 11997 7418 12001
rect 7803 11997 7837 12001
rect 7876 11997 7910 12001
rect 7949 11997 7983 12001
rect 8022 11997 8056 12001
rect 8095 11997 8129 12001
rect 8168 11997 8202 12001
rect 8241 11997 8275 12001
rect 8314 11997 8348 12001
rect 8387 11997 8421 12001
rect 8460 11997 8494 12001
rect 8533 11997 8567 12001
rect 8606 11997 8640 12001
rect 8680 11997 8714 12001
rect 8754 11997 8788 12001
rect 8828 11997 8862 12001
rect 9422 11997 9456 12001
rect 9501 11997 9535 12001
rect 9580 11997 9614 12001
rect 9659 11997 9693 12001
rect 9739 11997 9773 12001
rect 9819 11997 9853 12001
rect 10007 11997 10041 12001
rect 10082 11997 10116 12001
rect 10157 11997 10191 12001
rect 10233 11997 10267 12001
rect 10483 11997 10517 12001
rect 10558 11997 10592 12001
rect 10633 11997 10667 12001
rect 10709 11997 10743 12001
rect 10785 11997 10819 12001
rect 10861 11997 10895 12001
rect 10937 11997 10971 12001
rect 11013 11997 11047 12001
rect 11089 11997 11123 12001
rect 11165 11997 11199 12031
rect 1185 11689 1219 11723
rect 1268 11689 1302 11723
rect 1630 11689 1661 11723
rect 1661 11689 1664 11723
rect 1713 11689 1729 11723
rect 1729 11689 1747 11723
rect 1796 11689 1797 11723
rect 1797 11689 1830 11723
rect 1879 11689 1899 11723
rect 1899 11689 1913 11723
rect 1962 11689 1967 11723
rect 1967 11689 1996 11723
rect 2230 11689 2239 11723
rect 2239 11689 2264 11723
rect 2302 11689 2307 11723
rect 2307 11689 2336 11723
rect 2374 11689 2375 11723
rect 2375 11689 2408 11723
rect 2446 11689 2477 11723
rect 2477 11689 2480 11723
rect 2518 11689 2545 11723
rect 2545 11689 2552 11723
rect 2591 11689 2613 11723
rect 2613 11689 2625 11723
rect 2664 11689 2681 11723
rect 2681 11689 2698 11723
rect 2737 11689 2749 11723
rect 2749 11689 2771 11723
rect 2810 11689 2841 11723
rect 2841 11689 2844 11723
rect 2883 11689 2909 11723
rect 2909 11689 2917 11723
rect 2956 11689 2977 11723
rect 2977 11689 2990 11723
rect 3029 11689 3045 11723
rect 3045 11689 3063 11723
rect 3102 11689 3113 11723
rect 3113 11689 3136 11723
rect 3175 11689 3181 11723
rect 3181 11689 3209 11723
rect 3248 11689 3249 11723
rect 3249 11689 3282 11723
rect 3321 11689 3351 11723
rect 3351 11689 3355 11723
rect 3577 11689 3589 11723
rect 3589 11689 3611 11723
rect 3693 11689 3725 11723
rect 3725 11689 3727 11723
rect 3765 11689 3793 11723
rect 3793 11689 3799 11723
rect 3843 11689 3861 11723
rect 3861 11689 3877 11723
rect 3921 11689 3929 11723
rect 3929 11689 3955 11723
rect 4000 11689 4031 11723
rect 4031 11689 4034 11723
rect 4079 11689 4099 11723
rect 4099 11689 4113 11723
rect 4158 11689 4167 11723
rect 4167 11689 4192 11723
rect 4499 11689 4507 11723
rect 4507 11689 4533 11723
rect 4573 11689 4575 11723
rect 4575 11689 4607 11723
rect 4647 11689 4677 11723
rect 4677 11689 4681 11723
rect 4721 11689 4745 11723
rect 4745 11689 4755 11723
rect 5061 11689 5085 11723
rect 5085 11689 5095 11723
rect 5145 11689 5153 11723
rect 5153 11689 5179 11723
rect 5230 11689 5255 11723
rect 5255 11689 5264 11723
rect 5315 11689 5323 11723
rect 5323 11689 5349 11723
rect 5400 11689 5425 11723
rect 5425 11689 5434 11723
rect 5485 11689 5519 11723
rect 5557 11689 5591 11723
rect 5629 11689 5663 11723
rect 5703 11689 5722 11723
rect 5722 11689 5737 11723
rect 5777 11689 5790 11723
rect 5790 11689 5811 11723
rect 5851 11689 5858 11723
rect 5858 11689 5885 11723
rect 5925 11689 5926 11723
rect 5926 11689 5959 11723
rect 5999 11689 6028 11723
rect 6028 11689 6033 11723
rect 6339 11689 6368 11723
rect 6368 11689 6373 11723
rect 6413 11689 6436 11723
rect 6436 11689 6447 11723
rect 6487 11689 6504 11723
rect 6504 11689 6521 11723
rect 6561 11689 6572 11723
rect 6572 11689 6595 11723
rect 6901 11689 6912 11723
rect 6912 11689 6935 11723
rect 6976 11689 6980 11723
rect 6980 11689 7010 11723
rect 7051 11689 7082 11723
rect 7082 11689 7085 11723
rect 7126 11689 7150 11723
rect 7150 11689 7160 11723
rect 7201 11689 7218 11723
rect 7218 11689 7235 11723
rect 7276 11689 7286 11723
rect 7286 11689 7310 11723
rect 7351 11689 7354 11723
rect 7354 11689 7385 11723
rect 7423 11689 7456 11723
rect 7456 11689 7457 11723
rect 7826 11689 7830 11723
rect 7830 11689 7860 11723
rect 7901 11689 7923 11723
rect 7923 11689 7935 11723
rect 7976 11689 7991 11723
rect 7991 11689 8010 11723
rect 8051 11689 8059 11723
rect 8059 11689 8085 11723
rect 8126 11689 8127 11723
rect 8127 11689 8160 11723
rect 8201 11689 8229 11723
rect 8229 11689 8235 11723
rect 8276 11689 8297 11723
rect 8297 11689 8310 11723
rect 8352 11689 8365 11723
rect 8365 11689 8386 11723
rect 8428 11689 8433 11723
rect 8433 11689 8462 11723
rect 8504 11689 8535 11723
rect 8535 11689 8538 11723
rect 8580 11689 8603 11723
rect 8603 11689 8614 11723
rect 8656 11689 8671 11723
rect 8671 11689 8690 11723
rect 8732 11689 8739 11723
rect 8739 11689 8766 11723
rect 8808 11689 8841 11723
rect 8841 11689 8842 11723
rect 8884 11689 8909 11723
rect 8909 11689 8918 11723
rect 9347 11689 9351 11723
rect 9351 11689 9381 11723
rect 9427 11689 9453 11723
rect 9453 11689 9461 11723
rect 9507 11689 9521 11723
rect 9521 11689 9541 11723
rect 9587 11689 9589 11723
rect 9589 11689 9621 11723
rect 9667 11689 9691 11723
rect 9691 11689 9701 11723
rect 9747 11689 9759 11723
rect 9759 11689 9781 11723
rect 9827 11689 9861 11723
rect 9899 11689 9929 11723
rect 9929 11689 9933 11723
rect 1185 11616 1219 11650
rect 1185 11543 1219 11577
rect 1185 11470 1219 11504
rect 1185 11397 1219 11431
rect 3693 11621 3717 11650
rect 3717 11621 3727 11650
rect 3693 11616 3727 11621
rect 3693 11553 3717 11577
rect 3717 11553 3727 11577
rect 3693 11543 3727 11553
rect 3693 11485 3717 11504
rect 3717 11485 3727 11504
rect 3693 11470 3727 11485
rect 1185 11324 1219 11358
rect 2246 11395 2280 11429
rect 2319 11395 2353 11429
rect 2392 11395 2426 11429
rect 2465 11395 2499 11429
rect 2538 11395 2572 11429
rect 2246 11323 2280 11357
rect 2319 11323 2353 11357
rect 2392 11323 2426 11357
rect 2465 11323 2499 11357
rect 2538 11323 2572 11357
rect 1185 11251 1219 11285
rect 2246 11251 2280 11285
rect 2319 11251 2353 11285
rect 2392 11251 2426 11285
rect 2465 11251 2499 11285
rect 2538 11251 2572 11285
rect 2611 11251 3221 11429
rect 3693 11417 3717 11431
rect 3717 11417 3727 11431
rect 3693 11397 3727 11417
rect 5557 11621 5591 11651
rect 5557 11617 5591 11621
rect 5557 11553 5591 11579
rect 5557 11545 5591 11553
rect 5557 11485 5591 11507
rect 5557 11473 5591 11485
rect 5557 11417 5591 11435
rect 5557 11401 5591 11417
rect 3693 11349 3717 11359
rect 3717 11349 3727 11359
rect 3693 11325 3727 11349
rect 3693 11281 3717 11287
rect 3717 11281 3727 11287
rect 3693 11253 3727 11281
rect 1185 11179 1219 11213
rect 1185 11107 1219 11141
rect 1185 11035 1219 11069
rect 1185 10963 1219 10997
rect 1185 10891 1219 10925
rect 1185 10819 1219 10853
rect 1185 10747 1219 10781
rect 1185 10675 1219 10709
rect 1185 10603 1219 10637
rect 1185 10531 1219 10565
rect 1185 10459 1219 10493
rect 1185 10387 1219 10421
rect 1396 11224 1430 11228
rect 1396 11194 1430 11224
rect 3506 11224 3540 11228
rect 3506 11194 3540 11224
rect 1396 11151 1430 11154
rect 1396 11120 1430 11151
rect 3506 11151 3540 11154
rect 3506 11120 3540 11151
rect 1396 11078 1430 11080
rect 1396 11046 1430 11078
rect 3506 11078 3540 11080
rect 3506 11046 3540 11078
rect 1396 11005 1430 11006
rect 1396 10972 1430 11005
rect 3506 11005 3540 11006
rect 3506 10972 3540 11005
rect 1396 10898 1430 10932
rect 3506 10898 3540 10932
rect 1396 10825 1430 10858
rect 1396 10824 1430 10825
rect 3506 10825 3540 10858
rect 3506 10824 3540 10825
rect 1396 10752 1430 10784
rect 1396 10750 1430 10752
rect 3506 10752 3540 10784
rect 3506 10750 3540 10752
rect 1396 10678 1430 10710
rect 1396 10676 1430 10678
rect 3506 10678 3540 10710
rect 3506 10676 3540 10678
rect 1396 10604 1430 10636
rect 1396 10602 1430 10604
rect 3506 10604 3540 10636
rect 3506 10602 3540 10604
rect 1396 10530 1430 10561
rect 1396 10527 1430 10530
rect 3506 10530 3540 10561
rect 3506 10527 3540 10530
rect 1396 10456 1430 10486
rect 1396 10452 1430 10456
rect 3506 10456 3540 10486
rect 3506 10452 3540 10456
rect 3693 11213 3717 11215
rect 3717 11213 3727 11215
rect 3693 11181 3727 11213
rect 3693 11111 3727 11143
rect 3693 11109 3717 11111
rect 3717 11109 3727 11111
rect 3693 11043 3727 11071
rect 3693 11037 3717 11043
rect 3717 11037 3727 11043
rect 3693 10975 3727 10999
rect 3693 10965 3717 10975
rect 3717 10965 3727 10975
rect 3693 10907 3727 10927
rect 3693 10893 3717 10907
rect 3717 10893 3727 10907
rect 3693 10839 3727 10855
rect 3693 10821 3717 10839
rect 3717 10821 3727 10839
rect 3693 10771 3727 10783
rect 3693 10749 3717 10771
rect 3717 10749 3727 10771
rect 3693 10703 3727 10711
rect 3693 10677 3717 10703
rect 3717 10677 3727 10703
rect 3693 10635 3727 10639
rect 3693 10605 3717 10635
rect 3717 10605 3727 10635
rect 3693 10533 3717 10567
rect 3717 10533 3727 10567
rect 3693 10465 3717 10495
rect 3717 10465 3727 10495
rect 3693 10461 3727 10465
rect 3693 10397 3717 10423
rect 3717 10397 3727 10423
rect 2246 10362 2280 10396
rect 2319 10362 2353 10396
rect 2392 10362 2426 10396
rect 2465 10362 2499 10396
rect 2538 10362 2572 10396
rect 1185 10315 1219 10349
rect 1185 10243 1219 10277
rect 1185 10171 1219 10205
rect 2246 10290 2280 10324
rect 2319 10290 2353 10324
rect 2392 10290 2426 10324
rect 2465 10290 2499 10324
rect 2538 10290 2572 10324
rect 2246 10218 2280 10252
rect 2319 10218 2353 10252
rect 2392 10218 2426 10252
rect 2465 10218 2499 10252
rect 2538 10218 2572 10252
rect 2611 10218 3221 10396
rect 3693 10389 3727 10397
rect 3693 10329 3717 10351
rect 3717 10329 3727 10351
rect 3693 10317 3727 10329
rect 3693 10261 3717 10279
rect 3717 10261 3727 10279
rect 3693 10245 3727 10261
rect 3693 10193 3717 10207
rect 3717 10193 3727 10207
rect 3693 10173 3727 10193
rect 1185 10099 1219 10133
rect 1185 10027 1219 10061
rect 1185 9955 1219 9989
rect 1185 9883 1219 9917
rect 1185 9811 1219 9845
rect 1185 9739 1219 9773
rect 1185 9667 1219 9701
rect 1185 9595 1219 9629
rect 1185 9523 1219 9557
rect 1185 9451 1219 9485
rect 1185 9379 1219 9413
rect 1396 10138 1430 10142
rect 1396 10108 1430 10138
rect 3506 10138 3540 10142
rect 3506 10108 3540 10138
rect 1396 10065 1430 10068
rect 1396 10034 1430 10065
rect 3506 10065 3540 10068
rect 3506 10034 3540 10065
rect 1396 9992 1430 9994
rect 1396 9960 1430 9992
rect 3506 9992 3540 9994
rect 3506 9960 3540 9992
rect 1396 9919 1430 9920
rect 1396 9886 1430 9919
rect 3506 9919 3540 9920
rect 3506 9886 3540 9919
rect 1396 9812 1430 9846
rect 3506 9812 3540 9846
rect 1396 9739 1430 9772
rect 1396 9738 1430 9739
rect 3506 9739 3540 9772
rect 3506 9738 3540 9739
rect 1396 9666 1430 9698
rect 1396 9664 1430 9666
rect 3506 9666 3540 9698
rect 3506 9664 3540 9666
rect 1396 9592 1430 9624
rect 1396 9590 1430 9592
rect 3506 9592 3540 9624
rect 3506 9590 3540 9592
rect 1396 9518 1430 9550
rect 1396 9516 1430 9518
rect 3506 9518 3540 9550
rect 3506 9516 3540 9518
rect 1396 9444 1430 9475
rect 1396 9441 1430 9444
rect 3506 9444 3540 9475
rect 3506 9441 3540 9444
rect 1396 9370 1430 9400
rect 1396 9366 1430 9370
rect 3506 9370 3540 9400
rect 3506 9366 3540 9370
rect 3693 10125 3717 10135
rect 3717 10125 3727 10135
rect 3693 10101 3727 10125
rect 3693 10057 3717 10063
rect 3717 10057 3727 10063
rect 3693 10029 3727 10057
rect 3693 9989 3717 9991
rect 3717 9989 3727 9991
rect 3693 9957 3727 9989
rect 3693 9887 3727 9919
rect 3693 9885 3717 9887
rect 3717 9885 3727 9887
rect 3693 9819 3727 9847
rect 3693 9813 3717 9819
rect 3717 9813 3727 9819
rect 3693 9751 3727 9775
rect 3693 9741 3717 9751
rect 3717 9741 3727 9751
rect 3693 9683 3727 9703
rect 3693 9669 3717 9683
rect 3717 9669 3727 9683
rect 3693 9615 3727 9631
rect 3693 9597 3717 9615
rect 3717 9597 3727 9615
rect 3693 9547 3727 9559
rect 3693 9525 3717 9547
rect 3717 9525 3727 9547
rect 3693 9479 3727 9487
rect 3693 9453 3717 9479
rect 3717 9453 3727 9479
rect 3693 9411 3727 9415
rect 3693 9381 3717 9411
rect 3717 9381 3727 9411
rect 1185 9307 1219 9341
rect 2246 9309 2280 9343
rect 2319 9309 2353 9343
rect 2392 9309 2426 9343
rect 2465 9309 2499 9343
rect 2538 9309 2572 9343
rect 2611 9309 2645 9343
rect 2683 9309 2717 9343
rect 2755 9309 2789 9343
rect 2827 9309 2861 9343
rect 2899 9309 2933 9343
rect 2971 9309 3005 9343
rect 3043 9309 3077 9343
rect 3115 9309 3149 9343
rect 3187 9309 3221 9343
rect 3693 9309 3717 9343
rect 3717 9309 3727 9343
rect 1185 9235 1219 9269
rect 1185 9163 1219 9197
rect 1185 9091 1219 9125
rect 1185 9019 1219 9053
rect 1185 8947 1219 8981
rect 1185 8875 1219 8909
rect 1185 8803 1219 8837
rect 1185 8731 1219 8765
rect 1185 8659 1219 8693
rect 1185 8587 1219 8621
rect 1185 8515 1219 8549
rect 1396 9282 1430 9286
rect 1396 9252 1430 9282
rect 3506 9282 3540 9286
rect 3506 9252 3540 9282
rect 1396 9209 1430 9212
rect 1396 9178 1430 9209
rect 3506 9209 3540 9212
rect 3506 9178 3540 9209
rect 1396 9136 1430 9138
rect 1396 9104 1430 9136
rect 3506 9136 3540 9138
rect 3506 9104 3540 9136
rect 1396 9063 1430 9064
rect 1396 9030 1430 9063
rect 3506 9063 3540 9064
rect 3506 9030 3540 9063
rect 1396 8956 1430 8990
rect 3506 8956 3540 8990
rect 1396 8883 1430 8916
rect 1396 8882 1430 8883
rect 3506 8883 3540 8916
rect 3506 8882 3540 8883
rect 1396 8810 1430 8842
rect 1396 8808 1430 8810
rect 3506 8810 3540 8842
rect 3506 8808 3540 8810
rect 1396 8736 1430 8768
rect 1396 8734 1430 8736
rect 3506 8736 3540 8768
rect 3506 8734 3540 8736
rect 1396 8662 1430 8694
rect 1396 8660 1430 8662
rect 3506 8662 3540 8694
rect 3506 8660 3540 8662
rect 1396 8588 1430 8619
rect 1396 8585 1430 8588
rect 3506 8588 3540 8619
rect 3506 8585 3540 8588
rect 1396 8514 1430 8544
rect 1396 8510 1430 8514
rect 3506 8514 3540 8544
rect 3506 8510 3540 8514
rect 3693 9241 3717 9271
rect 3717 9241 3727 9271
rect 3693 9237 3727 9241
rect 3693 9173 3717 9199
rect 3717 9173 3727 9199
rect 3693 9165 3727 9173
rect 3693 9105 3717 9127
rect 3717 9105 3727 9127
rect 3693 9093 3727 9105
rect 3693 9037 3717 9055
rect 3717 9037 3727 9055
rect 3693 9021 3727 9037
rect 3693 8969 3717 8983
rect 3717 8969 3727 8983
rect 3693 8949 3727 8969
rect 3693 8901 3717 8911
rect 3717 8901 3727 8911
rect 3693 8877 3727 8901
rect 3693 8833 3717 8839
rect 3717 8833 3727 8839
rect 3693 8805 3727 8833
rect 3693 8765 3717 8767
rect 3717 8765 3727 8767
rect 3693 8733 3727 8765
rect 3693 8663 3727 8695
rect 3693 8661 3717 8663
rect 3717 8661 3727 8663
rect 3693 8595 3727 8623
rect 3693 8589 3717 8595
rect 3717 8589 3727 8595
rect 3693 8527 3727 8551
rect 3693 8517 3717 8527
rect 3717 8517 3727 8527
rect 1185 8443 1219 8477
rect 3693 8459 3727 8479
rect 2246 8423 2280 8457
rect 2319 8423 2353 8457
rect 2392 8423 2426 8457
rect 2465 8423 2499 8457
rect 2538 8423 2572 8457
rect 1185 8371 1219 8405
rect 1185 8299 1219 8333
rect 2246 8351 2280 8385
rect 2319 8351 2353 8385
rect 2392 8351 2426 8385
rect 2465 8351 2499 8385
rect 2538 8351 2572 8385
rect 2246 8279 2280 8313
rect 2319 8279 2353 8313
rect 2392 8279 2426 8313
rect 2465 8279 2499 8313
rect 2538 8279 2572 8313
rect 2611 8279 3221 8457
rect 3693 8445 3717 8459
rect 3717 8445 3727 8459
rect 3693 8391 3727 8407
rect 3693 8373 3717 8391
rect 3717 8373 3727 8391
rect 3693 8323 3727 8335
rect 3693 8301 3717 8323
rect 3717 8301 3727 8323
rect 1185 8227 1219 8261
rect 3693 8255 3727 8263
rect 1185 8155 1219 8189
rect 1185 8083 1219 8117
rect 1185 8011 1219 8045
rect 1185 7939 1219 7973
rect 1185 7867 1219 7901
rect 1185 7795 1219 7829
rect 1185 7723 1219 7757
rect 1185 7651 1219 7685
rect 1185 7579 1219 7613
rect 1185 7507 1219 7541
rect 1185 7435 1219 7469
rect 1185 7363 1219 7397
rect 1396 8222 1430 8252
rect 1396 8218 1430 8222
rect 3506 8222 3540 8252
rect 3506 8218 3540 8222
rect 1396 8153 1430 8180
rect 1396 8146 1430 8153
rect 3506 8153 3540 8180
rect 3506 8146 3540 8153
rect 1396 8084 1430 8108
rect 1396 8074 1430 8084
rect 3506 8084 3540 8108
rect 3506 8074 3540 8084
rect 1396 8015 1430 8036
rect 1396 8002 1430 8015
rect 3506 8015 3540 8036
rect 3506 8002 3540 8015
rect 1396 7946 1430 7964
rect 1396 7930 1430 7946
rect 3506 7946 3540 7964
rect 3506 7930 3540 7946
rect 1396 7877 1430 7892
rect 1396 7858 1430 7877
rect 3506 7877 3540 7892
rect 3506 7858 3540 7877
rect 1396 7808 1430 7820
rect 1396 7786 1430 7808
rect 3506 7808 3540 7820
rect 3506 7786 3540 7808
rect 1396 7739 1430 7748
rect 1396 7714 1430 7739
rect 3506 7739 3540 7748
rect 3506 7714 3540 7739
rect 1396 7670 1430 7676
rect 1396 7642 1430 7670
rect 3506 7670 3540 7676
rect 3506 7642 3540 7670
rect 1396 7601 1430 7604
rect 1396 7570 1430 7601
rect 3506 7601 3540 7604
rect 3506 7570 3540 7601
rect 1396 7498 1430 7531
rect 1396 7497 1430 7498
rect 3506 7498 3540 7531
rect 3506 7497 3540 7498
rect 1396 7428 1430 7458
rect 1396 7424 1430 7428
rect 3506 7428 3540 7458
rect 3506 7424 3540 7428
rect 3693 8229 3717 8255
rect 3717 8229 3727 8255
rect 3693 8187 3727 8191
rect 3693 8157 3717 8187
rect 3717 8157 3727 8187
rect 3693 8085 3717 8119
rect 3717 8085 3727 8119
rect 3693 8017 3717 8047
rect 3717 8017 3727 8047
rect 3693 8013 3727 8017
rect 3693 7949 3717 7975
rect 3717 7949 3727 7975
rect 3693 7941 3727 7949
rect 3693 7881 3717 7903
rect 3717 7881 3727 7903
rect 3693 7869 3727 7881
rect 3693 7813 3717 7831
rect 3717 7813 3727 7831
rect 3693 7797 3727 7813
rect 3693 7745 3717 7759
rect 3717 7745 3727 7759
rect 3693 7725 3727 7745
rect 3693 7677 3717 7687
rect 3717 7677 3727 7687
rect 3693 7653 3727 7677
rect 3693 7609 3717 7615
rect 3717 7609 3727 7615
rect 3693 7581 3727 7609
rect 3693 7541 3717 7543
rect 3717 7541 3727 7543
rect 3693 7509 3727 7541
rect 3693 7439 3727 7471
rect 3693 7437 3717 7439
rect 3717 7437 3727 7439
rect 2246 7367 2280 7401
rect 2319 7367 2353 7401
rect 2392 7367 2426 7401
rect 2465 7367 2499 7401
rect 2538 7367 2572 7401
rect 1185 7291 1219 7325
rect 1185 7219 1219 7253
rect 2246 7295 2280 7329
rect 2319 7295 2353 7329
rect 2392 7295 2426 7329
rect 2465 7295 2499 7329
rect 2538 7295 2572 7329
rect 2246 7223 2280 7257
rect 2319 7223 2353 7257
rect 2392 7223 2426 7257
rect 2465 7223 2499 7257
rect 2538 7223 2572 7257
rect 2611 7223 3221 7401
rect 3693 7371 3727 7399
rect 3693 7365 3717 7371
rect 3717 7365 3727 7371
rect 3693 7303 3727 7327
rect 3693 7293 3717 7303
rect 3717 7293 3727 7303
rect 3693 7235 3727 7255
rect 1185 7147 1219 7181
rect 1185 7075 1219 7109
rect 1185 7003 1219 7037
rect 1185 6931 1219 6965
rect 3693 7221 3717 7235
rect 3717 7221 3727 7235
rect 3693 7167 3727 7183
rect 3693 7149 3717 7167
rect 3717 7149 3727 7167
rect 3693 7099 3727 7111
rect 3693 7077 3717 7099
rect 3717 7077 3727 7099
rect 3693 7031 3727 7039
rect 3693 7005 3717 7031
rect 3717 7005 3727 7031
rect 3693 6963 3727 6967
rect 3693 6933 3717 6963
rect 3717 6933 3727 6963
rect 1185 6859 1219 6893
rect 1185 6787 1219 6821
rect 1185 6715 1219 6749
rect 1185 6643 1219 6677
rect 3693 6861 3717 6895
rect 3717 6861 3727 6895
rect 3693 6793 3717 6823
rect 3717 6793 3727 6823
rect 3693 6789 3727 6793
rect 3693 6725 3717 6751
rect 3717 6725 3727 6751
rect 3693 6717 3727 6725
rect 1185 6571 1219 6605
rect 2022 6635 2056 6669
rect 2095 6635 2129 6669
rect 2168 6635 2202 6669
rect 2241 6635 2275 6669
rect 2314 6635 2348 6669
rect 2022 6563 2056 6597
rect 2095 6563 2129 6597
rect 2168 6563 2202 6597
rect 2241 6563 2275 6597
rect 2314 6563 2348 6597
rect 1185 6499 1219 6533
rect 2022 6491 2056 6525
rect 2095 6491 2129 6525
rect 2168 6491 2202 6525
rect 2241 6491 2275 6525
rect 2314 6491 2348 6525
rect 2387 6491 2997 6669
rect 3693 6657 3717 6679
rect 3717 6657 3727 6679
rect 3693 6645 3727 6657
rect 3693 6589 3717 6607
rect 3717 6589 3727 6607
rect 3693 6573 3727 6589
rect 3693 6521 3717 6535
rect 3717 6521 3727 6535
rect 3693 6501 3727 6521
rect 1185 6427 1219 6461
rect 1185 6355 1219 6389
rect 1185 6283 1219 6317
rect 1185 6211 1219 6245
rect 1185 6139 1219 6173
rect 1185 6067 1219 6101
rect 1185 5995 1219 6029
rect 1185 5923 1219 5957
rect 1185 5851 1219 5885
rect 1185 5779 1219 5813
rect 1185 5707 1219 5741
rect 1396 6464 1430 6468
rect 1396 6434 1430 6464
rect 3506 6464 3540 6468
rect 3506 6434 3540 6464
rect 1396 6391 1430 6394
rect 1396 6360 1430 6391
rect 3506 6391 3540 6394
rect 3506 6360 3540 6391
rect 1396 6318 1430 6320
rect 1396 6286 1430 6318
rect 3506 6318 3540 6320
rect 3506 6286 3540 6318
rect 1396 6245 1430 6246
rect 1396 6212 1430 6245
rect 3506 6245 3540 6246
rect 3506 6212 3540 6245
rect 1396 6138 1430 6172
rect 3506 6138 3540 6172
rect 1396 6065 1430 6098
rect 1396 6064 1430 6065
rect 3506 6065 3540 6098
rect 3506 6064 3540 6065
rect 1396 5992 1430 6024
rect 1396 5990 1430 5992
rect 3506 5992 3540 6024
rect 3506 5990 3540 5992
rect 1396 5918 1430 5950
rect 1396 5916 1430 5918
rect 3506 5918 3540 5950
rect 3506 5916 3540 5918
rect 1396 5844 1430 5876
rect 1396 5842 1430 5844
rect 3506 5844 3540 5876
rect 3506 5842 3540 5844
rect 1396 5770 1430 5801
rect 1396 5767 1430 5770
rect 3506 5770 3540 5801
rect 3506 5767 3540 5770
rect 1396 5696 1430 5726
rect 1396 5692 1430 5696
rect 3506 5696 3540 5726
rect 3506 5692 3540 5696
rect 3693 6453 3717 6463
rect 3717 6453 3727 6463
rect 3693 6429 3727 6453
rect 3693 6385 3717 6391
rect 3717 6385 3727 6391
rect 3693 6357 3727 6385
rect 3693 6317 3717 6319
rect 3717 6317 3727 6319
rect 3693 6285 3727 6317
rect 3693 6215 3727 6247
rect 3693 6213 3717 6215
rect 3717 6213 3727 6215
rect 3693 6147 3727 6175
rect 3693 6141 3717 6147
rect 3717 6141 3727 6147
rect 3693 6079 3727 6103
rect 3693 6069 3717 6079
rect 3717 6069 3727 6079
rect 3693 6011 3727 6031
rect 3693 5997 3717 6011
rect 3717 5997 3727 6011
rect 3693 5943 3727 5959
rect 3693 5925 3717 5943
rect 3717 5925 3727 5943
rect 3693 5875 3727 5887
rect 3693 5853 3717 5875
rect 3717 5853 3727 5875
rect 3693 5807 3727 5815
rect 3693 5781 3717 5807
rect 3717 5781 3727 5807
rect 3693 5739 3727 5743
rect 3693 5709 3717 5739
rect 3717 5709 3727 5739
rect 1185 5635 1219 5669
rect 3693 5637 3717 5671
rect 3717 5637 3727 5671
rect 1185 5563 1219 5597
rect 1185 5491 1219 5525
rect 2022 5576 2056 5610
rect 2095 5576 2129 5610
rect 2168 5576 2202 5610
rect 2241 5576 2275 5610
rect 2314 5576 2348 5610
rect 2022 5504 2056 5538
rect 2095 5504 2129 5538
rect 2168 5504 2202 5538
rect 2241 5504 2275 5538
rect 2314 5504 2348 5538
rect 1185 5419 1219 5453
rect 2022 5432 2056 5466
rect 2095 5432 2129 5466
rect 2168 5432 2202 5466
rect 2241 5432 2275 5466
rect 2314 5432 2348 5466
rect 2387 5432 2997 5610
rect 3693 5569 3717 5599
rect 3717 5569 3727 5599
rect 3693 5565 3727 5569
rect 3693 5501 3717 5527
rect 3717 5501 3727 5527
rect 3693 5493 3727 5501
rect 3693 5433 3717 5455
rect 3717 5433 3727 5455
rect 3693 5421 3727 5433
rect 1185 5347 1219 5381
rect 1185 5275 1219 5309
rect 1185 5203 1219 5237
rect 1185 5131 1219 5165
rect 1185 5059 1219 5093
rect 1185 4987 1219 5021
rect 1185 4915 1219 4949
rect 1185 4843 1219 4877
rect 1185 4771 1219 4805
rect 1185 4699 1219 4733
rect 1185 4627 1219 4661
rect 1396 5378 1430 5382
rect 1396 5348 1430 5378
rect 3506 5378 3540 5382
rect 3506 5348 3540 5378
rect 1396 5305 1430 5308
rect 1396 5274 1430 5305
rect 3506 5305 3540 5308
rect 3506 5274 3540 5305
rect 1396 5232 1430 5234
rect 1396 5200 1430 5232
rect 3506 5232 3540 5234
rect 3506 5200 3540 5232
rect 1396 5159 1430 5160
rect 1396 5126 1430 5159
rect 3506 5159 3540 5160
rect 3506 5126 3540 5159
rect 1396 5052 1430 5086
rect 3506 5052 3540 5086
rect 1396 4979 1430 5012
rect 1396 4978 1430 4979
rect 3506 4979 3540 5012
rect 3506 4978 3540 4979
rect 1396 4906 1430 4938
rect 1396 4904 1430 4906
rect 3506 4906 3540 4938
rect 3506 4904 3540 4906
rect 1396 4832 1430 4864
rect 1396 4830 1430 4832
rect 3506 4832 3540 4864
rect 3506 4830 3540 4832
rect 1396 4758 1430 4790
rect 1396 4756 1430 4758
rect 3506 4758 3540 4790
rect 3506 4756 3540 4758
rect 1396 4684 1430 4715
rect 1396 4681 1430 4684
rect 3506 4684 3540 4715
rect 3506 4681 3540 4684
rect 1396 4610 1430 4640
rect 1396 4606 1430 4610
rect 3506 4610 3540 4640
rect 3506 4606 3540 4610
rect 3693 5365 3717 5383
rect 3717 5365 3727 5383
rect 3693 5349 3727 5365
rect 3693 5297 3717 5311
rect 3717 5297 3727 5311
rect 3693 5277 3727 5297
rect 3693 5229 3717 5239
rect 3717 5229 3727 5239
rect 3693 5205 3727 5229
rect 3693 5161 3717 5167
rect 3717 5161 3727 5167
rect 3693 5133 3727 5161
rect 3693 5093 3717 5095
rect 3717 5093 3727 5095
rect 3693 5061 3727 5093
rect 3693 4991 3727 5023
rect 3693 4989 3717 4991
rect 3717 4989 3727 4991
rect 3693 4923 3727 4951
rect 3693 4917 3717 4923
rect 3717 4917 3727 4923
rect 3693 4855 3727 4879
rect 3693 4845 3717 4855
rect 3717 4845 3727 4855
rect 3693 4787 3727 4807
rect 3693 4773 3717 4787
rect 3717 4773 3727 4787
rect 3693 4719 3727 4735
rect 3693 4701 3717 4719
rect 3717 4701 3727 4719
rect 3693 4651 3727 4663
rect 3693 4629 3717 4651
rect 3717 4629 3727 4651
rect 1185 4555 1219 4589
rect 3693 4583 3727 4591
rect 2022 4549 2056 4583
rect 2095 4549 2129 4583
rect 2168 4549 2202 4583
rect 2241 4549 2275 4583
rect 2314 4549 2348 4583
rect 2387 4549 2421 4583
rect 2459 4549 2493 4583
rect 2531 4549 2565 4583
rect 2603 4549 2637 4583
rect 2675 4549 2709 4583
rect 2747 4549 2781 4583
rect 2819 4549 2853 4583
rect 2891 4549 2925 4583
rect 2963 4549 2997 4583
rect 3693 4557 3717 4583
rect 3717 4557 3727 4583
rect 1185 4483 1219 4517
rect 1185 4411 1219 4445
rect 1185 4339 1219 4373
rect 1185 4267 1219 4301
rect 1185 4195 1219 4229
rect 1185 4123 1219 4157
rect 1185 4051 1219 4085
rect 1185 3979 1219 4013
rect 1185 3907 1219 3941
rect 1185 3835 1219 3869
rect 1185 3763 1219 3797
rect 1396 4522 1430 4526
rect 1396 4492 1430 4522
rect 3506 4522 3540 4526
rect 3506 4492 3540 4522
rect 1396 4449 1430 4452
rect 1396 4418 1430 4449
rect 3506 4449 3540 4452
rect 3506 4418 3540 4449
rect 1396 4376 1430 4378
rect 1396 4344 1430 4376
rect 3506 4376 3540 4378
rect 3506 4344 3540 4376
rect 1396 4303 1430 4304
rect 1396 4270 1430 4303
rect 3506 4303 3540 4304
rect 3506 4270 3540 4303
rect 1396 4196 1430 4230
rect 3506 4196 3540 4230
rect 1396 4123 1430 4156
rect 1396 4122 1430 4123
rect 3506 4123 3540 4156
rect 3506 4122 3540 4123
rect 1396 4050 1430 4082
rect 1396 4048 1430 4050
rect 3506 4050 3540 4082
rect 3506 4048 3540 4050
rect 1396 3976 1430 4008
rect 1396 3974 1430 3976
rect 3506 3976 3540 4008
rect 3506 3974 3540 3976
rect 1396 3902 1430 3934
rect 1396 3900 1430 3902
rect 3506 3902 3540 3934
rect 3506 3900 3540 3902
rect 1396 3828 1430 3859
rect 1396 3825 1430 3828
rect 3506 3828 3540 3859
rect 3506 3825 3540 3828
rect 1396 3754 1430 3784
rect 1396 3750 1430 3754
rect 3506 3754 3540 3784
rect 3506 3750 3540 3754
rect 3693 4515 3727 4519
rect 3693 4485 3717 4515
rect 3717 4485 3727 4515
rect 3693 4413 3717 4447
rect 3717 4413 3727 4447
rect 3693 4345 3717 4375
rect 3717 4345 3727 4375
rect 3693 4341 3727 4345
rect 3693 4277 3717 4303
rect 3717 4277 3727 4303
rect 3693 4269 3727 4277
rect 3693 4209 3717 4231
rect 3717 4209 3727 4231
rect 3693 4197 3727 4209
rect 3693 4141 3717 4159
rect 3717 4141 3727 4159
rect 3693 4125 3727 4141
rect 3693 4073 3717 4087
rect 3717 4073 3727 4087
rect 3693 4053 3727 4073
rect 3693 4005 3717 4015
rect 3717 4005 3727 4015
rect 3693 3981 3727 4005
rect 3693 3937 3717 3943
rect 3717 3937 3727 3943
rect 3693 3909 3727 3937
rect 4038 11328 4068 11362
rect 4068 11328 4072 11362
rect 4150 11328 4170 11362
rect 4170 11328 4184 11362
rect 5070 11328 5088 11362
rect 5088 11328 5104 11362
rect 5150 11328 5156 11362
rect 5156 11328 5184 11362
rect 4000 11239 4034 11252
rect 5274 11290 5308 11324
rect 4000 11218 4034 11239
rect 4000 11170 4034 11180
rect 4000 11146 4034 11170
rect 4538 11214 4572 11248
rect 4610 11214 4644 11248
rect 4682 11214 4716 11248
rect 5274 11239 5308 11251
rect 5274 11217 5308 11239
rect 5274 11170 5308 11178
rect 5274 11144 5308 11170
rect 4000 11101 4034 11108
rect 4000 11074 4034 11101
rect 5274 11101 5308 11105
rect 4538 11056 4572 11090
rect 4610 11056 4644 11090
rect 4682 11056 4716 11090
rect 5274 11071 5308 11101
rect 4000 11032 4034 11036
rect 4000 11002 4034 11032
rect 4000 10963 4034 10964
rect 4000 10930 4034 10963
rect 4000 10860 4034 10892
rect 4000 10858 4034 10860
rect 4000 10791 4034 10820
rect 4000 10786 4034 10791
rect 4000 10722 4034 10748
rect 4000 10714 4034 10722
rect 4000 10653 4034 10676
rect 4000 10642 4034 10653
rect 4000 10584 4034 10604
rect 4000 10570 4034 10584
rect 4000 10515 4034 10532
rect 4000 10498 4034 10515
rect 4000 10446 4034 10460
rect 4000 10426 4034 10446
rect 4000 10377 4034 10388
rect 4000 10354 4034 10377
rect 4000 10308 4034 10316
rect 4000 10282 4034 10308
rect 5192 11029 5226 11033
rect 5192 10999 5226 11029
rect 5192 10956 5226 10959
rect 5192 10925 5226 10956
rect 5192 10883 5226 10885
rect 5192 10851 5226 10883
rect 5192 10810 5226 10811
rect 5192 10777 5226 10810
rect 5192 10703 5226 10737
rect 5192 10630 5226 10663
rect 5192 10629 5226 10630
rect 5192 10557 5226 10589
rect 5192 10555 5226 10557
rect 5192 10483 5226 10515
rect 5192 10481 5226 10483
rect 5192 10409 5226 10441
rect 5192 10407 5226 10409
rect 5192 10335 5226 10366
rect 5192 10332 5226 10335
rect 5192 10261 5226 10291
rect 5192 10257 5226 10261
rect 5274 10998 5308 11032
rect 5274 10929 5308 10959
rect 5274 10925 5308 10929
rect 5274 10860 5308 10886
rect 5274 10852 5308 10860
rect 5274 10791 5308 10813
rect 5274 10779 5308 10791
rect 5274 10722 5308 10740
rect 5274 10706 5308 10722
rect 5274 10653 5308 10667
rect 5274 10633 5308 10653
rect 5274 10584 5308 10594
rect 5274 10560 5308 10584
rect 5274 10515 5308 10521
rect 5274 10487 5308 10515
rect 5274 10446 5308 10448
rect 5274 10414 5308 10446
rect 5274 10342 5308 10375
rect 5274 10341 5308 10342
rect 5274 10273 5308 10302
rect 5274 10268 5308 10273
rect 4000 10239 4034 10244
rect 4000 10210 4034 10239
rect 4840 10200 4874 10234
rect 4912 10200 4946 10234
rect 4984 10200 5018 10234
rect 5274 10204 5308 10229
rect 5274 10195 5308 10204
rect 4000 10170 4034 10172
rect 4000 10138 4034 10170
rect 4000 10066 4034 10100
rect 4000 9997 4034 10028
rect 4000 9994 4034 9997
rect 4000 9928 4034 9956
rect 4000 9922 4034 9928
rect 4000 9859 4034 9884
rect 4000 9850 4034 9859
rect 4000 9790 4034 9812
rect 4000 9778 4034 9790
rect 4000 9721 4034 9740
rect 4000 9706 4034 9721
rect 4000 9652 4034 9668
rect 4000 9634 4034 9652
rect 4000 9583 4034 9596
rect 4000 9562 4034 9583
rect 4000 9514 4034 9524
rect 4000 9490 4034 9514
rect 4000 9445 4034 9452
rect 4000 9418 4034 9445
rect 5192 10173 5226 10177
rect 5192 10143 5226 10173
rect 5192 10100 5226 10103
rect 5192 10069 5226 10100
rect 5192 10027 5226 10029
rect 5192 9995 5226 10027
rect 5192 9954 5226 9955
rect 5192 9921 5226 9954
rect 5192 9847 5226 9881
rect 5192 9774 5226 9807
rect 5192 9773 5226 9774
rect 5192 9701 5226 9733
rect 5192 9699 5226 9701
rect 5192 9627 5226 9659
rect 5192 9625 5226 9627
rect 5192 9553 5226 9585
rect 5192 9551 5226 9553
rect 5192 9479 5226 9510
rect 5192 9476 5226 9479
rect 5192 9405 5226 9435
rect 5192 9401 5226 9405
rect 5274 10135 5308 10156
rect 5274 10122 5308 10135
rect 5274 10066 5308 10083
rect 5274 10049 5308 10066
rect 5274 9997 5308 10010
rect 5274 9976 5308 9997
rect 5274 9928 5308 9937
rect 5274 9903 5308 9928
rect 5274 9859 5308 9864
rect 5274 9830 5308 9859
rect 5274 9790 5308 9791
rect 5274 9757 5308 9790
rect 5274 9687 5308 9718
rect 5274 9684 5308 9687
rect 5274 9618 5308 9645
rect 5274 9611 5308 9618
rect 5274 9549 5308 9572
rect 5274 9538 5308 9549
rect 5274 9480 5308 9499
rect 5274 9465 5308 9480
rect 5274 9411 5308 9426
rect 5274 9392 5308 9411
rect 4000 9376 4034 9380
rect 4000 9346 4034 9376
rect 4538 9344 4572 9378
rect 4610 9344 4644 9378
rect 4682 9344 4716 9378
rect 5274 9342 5308 9353
rect 4000 9307 4034 9308
rect 4000 9274 4034 9307
rect 4000 9204 4034 9236
rect 4000 9202 4034 9204
rect 4000 9135 4034 9164
rect 4000 9130 4034 9135
rect 4000 9066 4034 9092
rect 4000 9058 4034 9066
rect 4000 8997 4034 9020
rect 4000 8986 4034 8997
rect 4000 8928 4034 8948
rect 4000 8914 4034 8928
rect 4000 8859 4034 8876
rect 4000 8842 4034 8859
rect 4000 8790 4034 8804
rect 4000 8770 4034 8790
rect 4000 8721 4034 8732
rect 4000 8698 4034 8721
rect 4000 8652 4034 8660
rect 4000 8626 4034 8652
rect 4000 8583 4034 8588
rect 4000 8554 4034 8583
rect 4082 9317 4116 9321
rect 4082 9287 4116 9317
rect 4082 9244 4116 9247
rect 4082 9213 4116 9244
rect 4082 9171 4116 9173
rect 4082 9139 4116 9171
rect 4082 9098 4116 9099
rect 4082 9065 4116 9098
rect 4082 8991 4116 9025
rect 4082 8918 4116 8951
rect 4082 8917 4116 8918
rect 4082 8845 4116 8877
rect 4082 8843 4116 8845
rect 4082 8771 4116 8803
rect 4082 8769 4116 8771
rect 4082 8697 4116 8729
rect 4082 8695 4116 8697
rect 4082 8623 4116 8654
rect 4082 8620 4116 8623
rect 4082 8549 4116 8579
rect 4082 8545 4116 8549
rect 5274 9319 5308 9342
rect 5274 9273 5308 9280
rect 5274 9246 5308 9273
rect 5274 9204 5308 9207
rect 5274 9173 5308 9204
rect 5274 9100 5308 9134
rect 5274 9031 5308 9061
rect 5274 9027 5308 9031
rect 5274 8962 5308 8988
rect 5274 8954 5308 8962
rect 5274 8893 5308 8915
rect 5274 8881 5308 8893
rect 5274 8824 5308 8842
rect 5274 8808 5308 8824
rect 5274 8755 5308 8769
rect 5274 8735 5308 8755
rect 5274 8686 5308 8696
rect 5274 8662 5308 8686
rect 5274 8617 5308 8623
rect 5274 8589 5308 8617
rect 5274 8548 5308 8550
rect 4000 8514 4034 8516
rect 4000 8482 4034 8514
rect 4236 8488 4270 8522
rect 4308 8488 4342 8522
rect 4380 8488 4414 8522
rect 5274 8516 5308 8548
rect 4000 8410 4034 8444
rect 4000 8341 4034 8372
rect 4000 8338 4034 8341
rect 4000 8272 4034 8300
rect 4000 8266 4034 8272
rect 4000 8203 4034 8228
rect 4000 8194 4034 8203
rect 4000 8134 4034 8156
rect 4000 8122 4034 8134
rect 4000 8065 4034 8084
rect 4000 8050 4034 8065
rect 4000 7996 4034 8012
rect 4000 7978 4034 7996
rect 4000 7927 4034 7940
rect 4000 7906 4034 7927
rect 4000 7858 4034 7868
rect 4000 7834 4034 7858
rect 4000 7789 4034 7796
rect 4000 7762 4034 7789
rect 4000 7720 4034 7724
rect 4000 7690 4034 7720
rect 4082 8461 4116 8465
rect 4082 8431 4116 8461
rect 4082 8388 4116 8391
rect 4082 8357 4116 8388
rect 4082 8315 4116 8317
rect 4082 8283 4116 8315
rect 4082 8242 4116 8243
rect 4082 8209 4116 8242
rect 4082 8135 4116 8169
rect 4082 8062 4116 8095
rect 4082 8061 4116 8062
rect 4082 7989 4116 8021
rect 4082 7987 4116 7989
rect 4082 7915 4116 7947
rect 4082 7913 4116 7915
rect 4082 7841 4116 7873
rect 4082 7839 4116 7841
rect 4082 7767 4116 7798
rect 4082 7764 4116 7767
rect 4082 7693 4116 7723
rect 4082 7689 4116 7693
rect 5274 8445 5308 8477
rect 5274 8443 5308 8445
rect 5274 8376 5308 8404
rect 5274 8370 5308 8376
rect 5274 8307 5308 8331
rect 5274 8297 5308 8307
rect 5274 8238 5308 8258
rect 5274 8224 5308 8238
rect 5274 8169 5308 8185
rect 5274 8151 5308 8169
rect 5274 8100 5308 8112
rect 5274 8078 5308 8100
rect 5274 8031 5308 8040
rect 5274 8006 5308 8031
rect 5274 7962 5308 7968
rect 5274 7934 5308 7962
rect 5274 7893 5308 7896
rect 5274 7862 5308 7893
rect 5274 7790 5308 7824
rect 5274 7720 5308 7752
rect 5274 7718 5308 7720
rect 4000 7651 4034 7652
rect 4000 7618 4034 7651
rect 4538 7632 4572 7666
rect 4610 7632 4644 7666
rect 4682 7632 4716 7666
rect 5274 7651 5308 7680
rect 5274 7646 5308 7651
rect 4000 7549 4034 7580
rect 4000 7546 4034 7549
rect 4000 7481 4034 7508
rect 4000 7474 4034 7481
rect 4000 7413 4034 7436
rect 4000 7402 4034 7413
rect 4000 7345 4034 7364
rect 4000 7330 4034 7345
rect 4000 7277 4034 7292
rect 4000 7258 4034 7277
rect 4000 7209 4034 7220
rect 4000 7186 4034 7209
rect 4000 7141 4034 7147
rect 4000 7113 4034 7141
rect 4000 7073 4034 7074
rect 4000 7040 4034 7073
rect 4000 6971 4034 7001
rect 4000 6967 4034 6971
rect 4000 6903 4034 6928
rect 4000 6894 4034 6903
rect 4000 6835 4034 6855
rect 4000 6821 4034 6835
rect 5192 7605 5226 7609
rect 5192 7575 5226 7605
rect 5192 7532 5226 7535
rect 5192 7501 5226 7532
rect 5192 7459 5226 7461
rect 5192 7427 5226 7459
rect 5192 7386 5226 7387
rect 5192 7353 5226 7386
rect 5192 7279 5226 7313
rect 5192 7206 5226 7239
rect 5192 7205 5226 7206
rect 5192 7133 5226 7165
rect 5192 7131 5226 7133
rect 5192 7059 5226 7091
rect 5192 7057 5226 7059
rect 5192 6985 5226 7017
rect 5192 6983 5226 6985
rect 5192 6911 5226 6942
rect 5192 6908 5226 6911
rect 5192 6837 5226 6867
rect 5192 6833 5226 6837
rect 5274 7583 5308 7608
rect 5274 7574 5308 7583
rect 5274 7515 5308 7536
rect 5274 7502 5308 7515
rect 5274 7447 5308 7464
rect 5274 7430 5308 7447
rect 5274 7379 5308 7392
rect 5274 7358 5308 7379
rect 5274 7311 5308 7320
rect 5274 7286 5308 7311
rect 5274 7243 5308 7248
rect 5274 7214 5308 7243
rect 5274 7175 5308 7176
rect 5274 7142 5308 7175
rect 5274 7073 5308 7104
rect 5274 7070 5308 7073
rect 5274 7005 5308 7032
rect 5274 6998 5308 7005
rect 5274 6937 5308 6960
rect 5274 6926 5308 6937
rect 5274 6869 5308 6888
rect 5274 6854 5308 6869
rect 4000 6767 4034 6782
rect 4840 6776 4874 6810
rect 4912 6776 4946 6810
rect 4984 6776 5018 6810
rect 5274 6801 5308 6816
rect 5274 6782 5308 6801
rect 4000 6748 4034 6767
rect 4000 6699 4034 6709
rect 4000 6675 4034 6699
rect 4000 6631 4034 6636
rect 4000 6602 4034 6631
rect 4000 6529 4034 6563
rect 4000 6461 4034 6490
rect 4000 6456 4034 6461
rect 4000 6393 4034 6417
rect 4000 6383 4034 6393
rect 4000 6325 4034 6344
rect 4000 6310 4034 6325
rect 4000 6257 4034 6271
rect 4000 6237 4034 6257
rect 4000 6189 4034 6198
rect 4000 6164 4034 6189
rect 4000 6121 4034 6125
rect 4000 6091 4034 6121
rect 4000 6019 4034 6052
rect 4000 6018 4034 6019
rect 4000 5951 4034 5979
rect 5192 6749 5226 6753
rect 5192 6719 5226 6749
rect 5192 6676 5226 6679
rect 5192 6645 5226 6676
rect 5192 6603 5226 6605
rect 5192 6571 5226 6603
rect 5192 6530 5226 6531
rect 5192 6497 5226 6530
rect 5192 6423 5226 6457
rect 5192 6350 5226 6383
rect 5192 6349 5226 6350
rect 5192 6277 5226 6309
rect 5192 6275 5226 6277
rect 5192 6203 5226 6235
rect 5192 6201 5226 6203
rect 5192 6129 5226 6161
rect 5192 6127 5226 6129
rect 5192 6055 5226 6086
rect 5192 6052 5226 6055
rect 5192 5981 5226 6011
rect 5192 5977 5226 5981
rect 5274 6733 5308 6744
rect 5274 6710 5308 6733
rect 5274 6665 5308 6672
rect 5274 6638 5308 6665
rect 5274 6597 5308 6600
rect 5274 6566 5308 6597
rect 5274 6495 5308 6528
rect 5274 6494 5308 6495
rect 5274 6427 5308 6456
rect 5274 6422 5308 6427
rect 5274 6359 5308 6384
rect 5274 6350 5308 6359
rect 5274 6291 5308 6312
rect 5274 6278 5308 6291
rect 5274 6223 5308 6240
rect 5274 6206 5308 6223
rect 5274 6155 5308 6168
rect 5274 6134 5308 6155
rect 5274 6087 5308 6096
rect 5274 6062 5308 6087
rect 5274 6019 5308 6024
rect 5274 5990 5308 6019
rect 4000 5945 4034 5951
rect 4538 5920 4572 5954
rect 4610 5920 4644 5954
rect 4682 5920 4716 5954
rect 5274 5951 5308 5952
rect 5274 5918 5308 5951
rect 4000 5883 4034 5906
rect 4000 5872 4034 5883
rect 4000 5815 4034 5833
rect 4000 5799 4034 5815
rect 4000 5747 4034 5760
rect 4000 5726 4034 5747
rect 4000 5679 4034 5687
rect 4000 5653 4034 5679
rect 4000 5611 4034 5614
rect 4000 5580 4034 5611
rect 4000 5509 4034 5541
rect 4000 5507 4034 5509
rect 4000 5441 4034 5468
rect 4000 5434 4034 5441
rect 4000 5373 4034 5395
rect 4000 5361 4034 5373
rect 4000 5305 4034 5322
rect 4000 5288 4034 5305
rect 4000 5237 4034 5249
rect 4000 5215 4034 5237
rect 4000 5169 4034 5176
rect 4000 5142 4034 5169
rect 4082 5893 4116 5897
rect 4082 5863 4116 5893
rect 4082 5820 4116 5823
rect 4082 5789 4116 5820
rect 4082 5747 4116 5749
rect 4082 5715 4116 5747
rect 4082 5674 4116 5675
rect 4082 5641 4116 5674
rect 4082 5567 4116 5601
rect 4082 5494 4116 5527
rect 4082 5493 4116 5494
rect 4082 5421 4116 5453
rect 4082 5419 4116 5421
rect 4082 5347 4116 5379
rect 4082 5345 4116 5347
rect 4082 5273 4116 5305
rect 4082 5271 4116 5273
rect 4082 5199 4116 5230
rect 4082 5196 4116 5199
rect 4082 5125 4116 5155
rect 4082 5121 4116 5125
rect 5274 5849 5308 5880
rect 5274 5846 5308 5849
rect 5274 5781 5308 5808
rect 5274 5774 5308 5781
rect 5274 5713 5308 5736
rect 5274 5702 5308 5713
rect 5274 5645 5308 5664
rect 5274 5630 5308 5645
rect 5274 5577 5308 5592
rect 5274 5558 5308 5577
rect 5274 5509 5308 5520
rect 5274 5486 5308 5509
rect 5274 5441 5308 5448
rect 5274 5414 5308 5441
rect 5274 5373 5308 5376
rect 5274 5342 5308 5373
rect 5274 5271 5308 5304
rect 5274 5270 5308 5271
rect 5274 5203 5308 5232
rect 5274 5198 5308 5203
rect 5274 5135 5308 5160
rect 5274 5126 5308 5135
rect 4000 5101 4034 5103
rect 4000 5069 4034 5101
rect 4236 5064 4270 5098
rect 4308 5064 4342 5098
rect 4380 5064 4414 5098
rect 5274 5067 5308 5088
rect 5274 5054 5308 5067
rect 4000 4999 4034 5030
rect 4000 4996 4034 4999
rect 4000 4931 4034 4957
rect 4000 4923 4034 4931
rect 4000 4863 4034 4884
rect 4000 4850 4034 4863
rect 4000 4795 4034 4811
rect 4000 4777 4034 4795
rect 4000 4727 4034 4738
rect 4000 4704 4034 4727
rect 4000 4659 4034 4665
rect 4000 4631 4034 4659
rect 4000 4591 4034 4592
rect 4000 4558 4034 4591
rect 4000 4489 4034 4519
rect 4000 4485 4034 4489
rect 4000 4421 4034 4446
rect 4000 4412 4034 4421
rect 4000 4353 4034 4373
rect 4000 4339 4034 4353
rect 4000 4285 4034 4300
rect 4000 4266 4034 4285
rect 4082 5037 4116 5041
rect 4082 5007 4116 5037
rect 4082 4964 4116 4967
rect 4082 4933 4116 4964
rect 4082 4891 4116 4893
rect 4082 4859 4116 4891
rect 4082 4818 4116 4819
rect 4082 4785 4116 4818
rect 4082 4711 4116 4745
rect 4082 4638 4116 4671
rect 4082 4637 4116 4638
rect 4082 4565 4116 4597
rect 4082 4563 4116 4565
rect 4082 4491 4116 4523
rect 4082 4489 4116 4491
rect 4082 4417 4116 4449
rect 4082 4415 4116 4417
rect 4082 4343 4116 4374
rect 4082 4340 4116 4343
rect 4082 4269 4116 4299
rect 4082 4265 4116 4269
rect 5274 4999 5308 5016
rect 5274 4982 5308 4999
rect 5274 4931 5308 4944
rect 5274 4910 5308 4931
rect 5274 4863 5308 4872
rect 5274 4838 5308 4863
rect 5274 4795 5308 4800
rect 5274 4766 5308 4795
rect 5274 4727 5308 4728
rect 5274 4694 5308 4727
rect 5274 4625 5308 4656
rect 5274 4622 5308 4625
rect 5274 4557 5308 4584
rect 5274 4550 5308 4557
rect 5274 4489 5308 4512
rect 5274 4478 5308 4489
rect 5274 4421 5308 4440
rect 5274 4406 5308 4421
rect 5274 4353 5308 4368
rect 5274 4334 5308 4353
rect 5274 4285 5308 4296
rect 5274 4262 5308 4285
rect 4000 4217 4034 4227
rect 4000 4193 4034 4217
rect 4538 4208 4572 4242
rect 4610 4208 4644 4242
rect 4682 4208 4716 4242
rect 5274 4217 5308 4224
rect 5274 4190 5308 4217
rect 4000 4149 4034 4154
rect 4000 4120 4034 4149
rect 4000 4047 4034 4081
rect 4538 4050 4572 4084
rect 4610 4050 4644 4084
rect 4682 4050 4716 4084
rect 5274 4149 5308 4152
rect 5274 4118 5308 4149
rect 4000 3974 4034 4008
rect 5274 4046 5308 4080
rect 4138 3936 4170 3970
rect 4170 3936 4172 3970
rect 4224 3936 4238 3970
rect 4238 3936 4258 3970
rect 4310 3936 4340 3970
rect 4340 3936 4344 3970
rect 4397 3936 4408 3970
rect 4408 3936 4431 3970
rect 4843 3936 4850 3970
rect 4850 3936 4877 3970
rect 4921 3936 4952 3970
rect 4952 3936 4955 3970
rect 4999 3936 5020 3970
rect 5020 3936 5033 3970
rect 5078 3936 5088 3970
rect 5088 3936 5112 3970
rect 5157 3936 5190 3970
rect 5190 3936 5191 3970
rect 5236 3936 5270 3970
rect 5557 11349 5591 11363
rect 5557 11329 5591 11349
rect 7423 11621 7431 11650
rect 7431 11621 7457 11650
rect 7423 11616 7457 11621
rect 7423 11553 7431 11577
rect 7431 11553 7457 11577
rect 7423 11543 7457 11553
rect 7423 11485 7431 11504
rect 7431 11485 7457 11504
rect 7423 11470 7457 11485
rect 7423 11417 7431 11431
rect 7431 11417 7457 11431
rect 9899 11621 9929 11650
rect 9929 11621 9933 11650
rect 9899 11616 9933 11621
rect 9899 11553 9929 11577
rect 9929 11553 9933 11577
rect 9899 11543 9933 11553
rect 9899 11485 9929 11504
rect 9929 11485 9933 11504
rect 9899 11470 9933 11485
rect 7423 11397 7457 11417
rect 5557 11281 5591 11291
rect 5557 11257 5591 11281
rect 5557 11213 5591 11219
rect 5557 11185 5591 11213
rect 5557 11145 5591 11147
rect 5557 11113 5591 11145
rect 5557 11043 5591 11075
rect 5557 11041 5591 11043
rect 5557 10975 5591 11003
rect 5557 10969 5591 10975
rect 5557 10907 5591 10931
rect 5557 10897 5591 10907
rect 5557 10839 5591 10859
rect 5557 10825 5591 10839
rect 5557 10771 5591 10787
rect 5557 10753 5591 10771
rect 5557 10703 5591 10715
rect 5557 10681 5591 10703
rect 5557 10635 5591 10643
rect 5557 10609 5591 10635
rect 5557 10567 5591 10571
rect 5557 10537 5591 10567
rect 5557 10465 5591 10499
rect 5557 10397 5591 10427
rect 5557 10393 5591 10397
rect 5557 10329 5591 10355
rect 5557 10321 5591 10329
rect 5557 10261 5591 10283
rect 5557 10249 5591 10261
rect 5557 10193 5591 10211
rect 5557 10177 5591 10193
rect 5557 10125 5591 10139
rect 5557 10105 5591 10125
rect 5557 10057 5591 10067
rect 5557 10033 5591 10057
rect 5557 9989 5591 9995
rect 5557 9961 5591 9989
rect 5557 9921 5591 9923
rect 5557 9889 5591 9921
rect 5557 9819 5591 9851
rect 5557 9817 5591 9819
rect 5557 9751 5591 9779
rect 5557 9745 5591 9751
rect 5557 9683 5591 9707
rect 5557 9673 5591 9683
rect 5557 9615 5591 9635
rect 5557 9601 5591 9615
rect 5557 9547 5591 9563
rect 5557 9529 5591 9547
rect 5557 9479 5591 9491
rect 5557 9457 5591 9479
rect 5557 9411 5591 9419
rect 5557 9385 5591 9411
rect 5557 9343 5591 9347
rect 5557 9313 5591 9343
rect 5557 9241 5591 9275
rect 5557 9173 5591 9203
rect 5557 9169 5591 9173
rect 5557 9105 5591 9131
rect 5557 9097 5591 9105
rect 5557 9037 5591 9059
rect 5557 9025 5591 9037
rect 5557 8969 5591 8987
rect 5557 8953 5591 8969
rect 5557 8901 5591 8915
rect 5557 8881 5591 8901
rect 5557 8833 5591 8843
rect 5557 8809 5591 8833
rect 5557 8765 5591 8771
rect 5557 8737 5591 8765
rect 5557 8697 5591 8699
rect 5557 8665 5591 8697
rect 5557 8595 5591 8627
rect 5557 8593 5591 8595
rect 5557 8527 5591 8555
rect 5557 8521 5591 8527
rect 5557 8459 5591 8483
rect 5557 8449 5591 8459
rect 5557 8391 5591 8411
rect 5557 8377 5591 8391
rect 5557 8323 5591 8339
rect 5557 8305 5591 8323
rect 5557 8255 5591 8267
rect 5557 8233 5591 8255
rect 5557 8187 5591 8195
rect 5557 8161 5591 8187
rect 5557 8119 5591 8123
rect 5557 8089 5591 8119
rect 5557 8017 5591 8051
rect 5557 7949 5591 7979
rect 5557 7945 5591 7949
rect 5557 7881 5591 7907
rect 5557 7873 5591 7881
rect 5557 7813 5591 7835
rect 5557 7801 5591 7813
rect 5557 7745 5591 7763
rect 5557 7729 5591 7745
rect 5557 7677 5591 7691
rect 5557 7657 5591 7677
rect 5557 7609 5591 7619
rect 5557 7585 5591 7609
rect 5557 7541 5591 7547
rect 5557 7513 5591 7541
rect 5557 7473 5591 7475
rect 5557 7441 5591 7473
rect 5557 7371 5591 7403
rect 5557 7369 5591 7371
rect 5557 7303 5591 7331
rect 5557 7297 5591 7303
rect 5557 7235 5591 7259
rect 5557 7225 5591 7235
rect 5557 7167 5591 7187
rect 5557 7153 5591 7167
rect 5557 7099 5591 7115
rect 5557 7081 5591 7099
rect 5557 7031 5591 7043
rect 5557 7009 5591 7031
rect 5557 6963 5591 6971
rect 5557 6937 5591 6963
rect 5557 6895 5591 6899
rect 5557 6865 5591 6895
rect 5557 6793 5591 6826
rect 5557 6792 5591 6793
rect 5557 6725 5591 6753
rect 5557 6719 5591 6725
rect 5557 6657 5591 6680
rect 5557 6646 5591 6657
rect 5557 6589 5591 6607
rect 5557 6573 5591 6589
rect 5557 6521 5591 6534
rect 5557 6500 5591 6521
rect 5557 6453 5591 6461
rect 5557 6427 5591 6453
rect 5557 6385 5591 6388
rect 5557 6354 5591 6385
rect 5557 6283 5591 6315
rect 5557 6281 5591 6283
rect 5557 6215 5591 6242
rect 5557 6208 5591 6215
rect 5557 6147 5591 6169
rect 5557 6135 5591 6147
rect 5557 6079 5591 6096
rect 5557 6062 5591 6079
rect 5557 6011 5591 6023
rect 5557 5989 5591 6011
rect 5557 5943 5591 5950
rect 5557 5916 5591 5943
rect 5557 5875 5591 5877
rect 5557 5843 5591 5875
rect 5557 5773 5591 5804
rect 5557 5770 5591 5773
rect 5557 5705 5591 5731
rect 5557 5697 5591 5705
rect 5557 5637 5591 5658
rect 5557 5624 5591 5637
rect 5557 5569 5591 5585
rect 5557 5551 5591 5569
rect 5557 5501 5591 5512
rect 5557 5478 5591 5501
rect 5557 5433 5591 5439
rect 5557 5405 5591 5433
rect 5557 5365 5591 5366
rect 5557 5332 5591 5365
rect 5557 5263 5591 5293
rect 5557 5259 5591 5263
rect 5557 5195 5591 5220
rect 5557 5186 5591 5195
rect 5557 5127 5591 5147
rect 5557 5113 5591 5127
rect 5557 5059 5591 5074
rect 5557 5040 5591 5059
rect 5557 4991 5591 5001
rect 5557 4967 5591 4991
rect 5557 4923 5591 4928
rect 5557 4894 5591 4923
rect 5557 4821 5591 4855
rect 5557 4753 5591 4782
rect 5557 4748 5591 4753
rect 5557 4685 5591 4709
rect 5557 4675 5591 4685
rect 5557 4617 5591 4636
rect 5557 4602 5591 4617
rect 5557 4549 5591 4563
rect 5557 4529 5591 4549
rect 5557 4481 5591 4490
rect 5557 4456 5591 4481
rect 5557 4413 5591 4417
rect 5557 4383 5591 4413
rect 5557 4311 5591 4344
rect 5557 4310 5591 4311
rect 5557 4243 5591 4271
rect 5557 4237 5591 4243
rect 5557 4175 5591 4198
rect 5557 4164 5591 4175
rect 5557 4107 5591 4125
rect 5557 4091 5591 4107
rect 5557 4039 5591 4052
rect 5557 4018 5591 4039
rect 5557 3971 5591 3979
rect 5557 3945 5591 3971
rect 3693 3869 3717 3871
rect 3717 3869 3727 3871
rect 3693 3837 3727 3869
rect 3693 3767 3727 3799
rect 3693 3765 3717 3767
rect 3717 3765 3727 3767
rect 1185 3691 1219 3725
rect 3693 3699 3727 3727
rect 2022 3663 2056 3697
rect 2095 3663 2129 3697
rect 2168 3663 2202 3697
rect 2241 3663 2275 3697
rect 2314 3663 2348 3697
rect 1185 3619 1219 3653
rect 1185 3547 1219 3581
rect 2022 3591 2056 3625
rect 2095 3591 2129 3625
rect 2168 3591 2202 3625
rect 2241 3591 2275 3625
rect 2314 3591 2348 3625
rect 2387 3591 2997 3697
rect 3693 3693 3717 3699
rect 3717 3693 3727 3699
rect 5557 3903 5591 3906
rect 5557 3872 5591 3903
rect 5878 11328 5908 11362
rect 5908 11328 5912 11362
rect 5990 11328 6010 11362
rect 6010 11328 6024 11362
rect 6910 11328 6928 11362
rect 6928 11328 6944 11362
rect 6990 11328 6996 11362
rect 6996 11328 7024 11362
rect 5840 11239 5874 11252
rect 7114 11290 7148 11324
rect 5840 11218 5874 11239
rect 5840 11170 5874 11180
rect 5840 11146 5874 11170
rect 6378 11214 6412 11248
rect 6450 11214 6484 11248
rect 6522 11214 6556 11248
rect 7114 11239 7148 11251
rect 7114 11217 7148 11239
rect 7114 11170 7148 11178
rect 7114 11144 7148 11170
rect 5840 11101 5874 11108
rect 5840 11074 5874 11101
rect 7114 11101 7148 11105
rect 6378 11056 6412 11090
rect 6450 11056 6484 11090
rect 6522 11056 6556 11090
rect 7114 11071 7148 11101
rect 5840 11032 5874 11036
rect 5840 11002 5874 11032
rect 5840 10963 5874 10964
rect 5840 10930 5874 10963
rect 5840 10860 5874 10892
rect 5840 10858 5874 10860
rect 5840 10791 5874 10820
rect 5840 10786 5874 10791
rect 5840 10722 5874 10748
rect 5840 10714 5874 10722
rect 5840 10653 5874 10676
rect 5840 10642 5874 10653
rect 5840 10584 5874 10604
rect 5840 10570 5874 10584
rect 5840 10515 5874 10532
rect 5840 10498 5874 10515
rect 5840 10446 5874 10460
rect 5840 10426 5874 10446
rect 5840 10377 5874 10388
rect 5840 10354 5874 10377
rect 5840 10308 5874 10316
rect 5840 10282 5874 10308
rect 7032 11029 7066 11033
rect 7032 10999 7066 11029
rect 7032 10956 7066 10959
rect 7032 10925 7066 10956
rect 7032 10883 7066 10885
rect 7032 10851 7066 10883
rect 7032 10810 7066 10811
rect 7032 10777 7066 10810
rect 7032 10703 7066 10737
rect 7032 10630 7066 10663
rect 7032 10629 7066 10630
rect 7032 10557 7066 10589
rect 7032 10555 7066 10557
rect 7032 10483 7066 10515
rect 7032 10481 7066 10483
rect 7032 10409 7066 10441
rect 7032 10407 7066 10409
rect 7032 10335 7066 10366
rect 7032 10332 7066 10335
rect 7032 10261 7066 10291
rect 7032 10257 7066 10261
rect 7114 10998 7148 11032
rect 7114 10929 7148 10959
rect 7114 10925 7148 10929
rect 7114 10860 7148 10886
rect 7114 10852 7148 10860
rect 7114 10791 7148 10813
rect 7114 10779 7148 10791
rect 7114 10722 7148 10740
rect 7114 10706 7148 10722
rect 7114 10653 7148 10667
rect 7114 10633 7148 10653
rect 7114 10584 7148 10594
rect 7114 10560 7148 10584
rect 7114 10515 7148 10521
rect 7114 10487 7148 10515
rect 7114 10446 7148 10448
rect 7114 10414 7148 10446
rect 7114 10342 7148 10375
rect 7114 10341 7148 10342
rect 7114 10273 7148 10302
rect 7114 10268 7148 10273
rect 5840 10239 5874 10244
rect 5840 10210 5874 10239
rect 6680 10200 6714 10234
rect 6752 10200 6786 10234
rect 6824 10200 6858 10234
rect 7114 10204 7148 10229
rect 7114 10195 7148 10204
rect 5840 10170 5874 10172
rect 5840 10138 5874 10170
rect 5840 10066 5874 10100
rect 5840 9997 5874 10028
rect 5840 9994 5874 9997
rect 5840 9928 5874 9956
rect 5840 9922 5874 9928
rect 5840 9859 5874 9884
rect 5840 9850 5874 9859
rect 5840 9790 5874 9812
rect 5840 9778 5874 9790
rect 5840 9721 5874 9740
rect 5840 9706 5874 9721
rect 5840 9652 5874 9668
rect 5840 9634 5874 9652
rect 5840 9583 5874 9596
rect 5840 9562 5874 9583
rect 5840 9514 5874 9524
rect 5840 9490 5874 9514
rect 5840 9445 5874 9452
rect 5840 9418 5874 9445
rect 7032 10173 7066 10177
rect 7032 10143 7066 10173
rect 7032 10100 7066 10103
rect 7032 10069 7066 10100
rect 7032 10027 7066 10029
rect 7032 9995 7066 10027
rect 7032 9954 7066 9955
rect 7032 9921 7066 9954
rect 7032 9847 7066 9881
rect 7032 9774 7066 9807
rect 7032 9773 7066 9774
rect 7032 9701 7066 9733
rect 7032 9699 7066 9701
rect 7032 9627 7066 9659
rect 7032 9625 7066 9627
rect 7032 9553 7066 9585
rect 7032 9551 7066 9553
rect 7032 9479 7066 9510
rect 7032 9476 7066 9479
rect 7032 9405 7066 9435
rect 7032 9401 7066 9405
rect 7114 10135 7148 10156
rect 7114 10122 7148 10135
rect 7114 10066 7148 10083
rect 7114 10049 7148 10066
rect 7114 9997 7148 10010
rect 7114 9976 7148 9997
rect 7114 9928 7148 9937
rect 7114 9903 7148 9928
rect 7114 9859 7148 9864
rect 7114 9830 7148 9859
rect 7114 9790 7148 9791
rect 7114 9757 7148 9790
rect 7114 9687 7148 9718
rect 7114 9684 7148 9687
rect 7114 9618 7148 9645
rect 7114 9611 7148 9618
rect 7114 9549 7148 9572
rect 7114 9538 7148 9549
rect 7114 9480 7148 9499
rect 7114 9465 7148 9480
rect 7114 9411 7148 9426
rect 7114 9392 7148 9411
rect 5840 9376 5874 9380
rect 5840 9346 5874 9376
rect 6378 9344 6412 9378
rect 6450 9344 6484 9378
rect 6522 9344 6556 9378
rect 7114 9342 7148 9353
rect 5840 9307 5874 9308
rect 5840 9274 5874 9307
rect 5840 9204 5874 9236
rect 5840 9202 5874 9204
rect 5840 9135 5874 9164
rect 5840 9130 5874 9135
rect 5840 9066 5874 9092
rect 5840 9058 5874 9066
rect 5840 8997 5874 9020
rect 5840 8986 5874 8997
rect 5840 8928 5874 8948
rect 5840 8914 5874 8928
rect 5840 8859 5874 8876
rect 5840 8842 5874 8859
rect 5840 8790 5874 8804
rect 5840 8770 5874 8790
rect 5840 8721 5874 8732
rect 5840 8698 5874 8721
rect 5840 8652 5874 8660
rect 5840 8626 5874 8652
rect 5840 8583 5874 8588
rect 5840 8554 5874 8583
rect 5922 9317 5956 9321
rect 5922 9287 5956 9317
rect 5922 9244 5956 9247
rect 5922 9213 5956 9244
rect 5922 9171 5956 9173
rect 5922 9139 5956 9171
rect 5922 9098 5956 9099
rect 5922 9065 5956 9098
rect 5922 8991 5956 9025
rect 5922 8918 5956 8951
rect 5922 8917 5956 8918
rect 5922 8845 5956 8877
rect 5922 8843 5956 8845
rect 5922 8771 5956 8803
rect 5922 8769 5956 8771
rect 5922 8697 5956 8729
rect 5922 8695 5956 8697
rect 5922 8623 5956 8654
rect 5922 8620 5956 8623
rect 5922 8549 5956 8579
rect 5922 8545 5956 8549
rect 7114 9319 7148 9342
rect 7114 9273 7148 9280
rect 7114 9246 7148 9273
rect 7114 9204 7148 9207
rect 7114 9173 7148 9204
rect 7114 9100 7148 9134
rect 7114 9031 7148 9061
rect 7114 9027 7148 9031
rect 7114 8962 7148 8988
rect 7114 8954 7148 8962
rect 7114 8893 7148 8915
rect 7114 8881 7148 8893
rect 7114 8824 7148 8842
rect 7114 8808 7148 8824
rect 7114 8755 7148 8769
rect 7114 8735 7148 8755
rect 7114 8686 7148 8696
rect 7114 8662 7148 8686
rect 7114 8617 7148 8623
rect 7114 8589 7148 8617
rect 7114 8548 7148 8550
rect 5840 8514 5874 8516
rect 5840 8482 5874 8514
rect 6076 8488 6110 8522
rect 6148 8488 6182 8522
rect 6220 8488 6254 8522
rect 7114 8516 7148 8548
rect 5840 8410 5874 8444
rect 5840 8341 5874 8372
rect 5840 8338 5874 8341
rect 5840 8272 5874 8300
rect 5840 8266 5874 8272
rect 5840 8203 5874 8228
rect 5840 8194 5874 8203
rect 5840 8134 5874 8156
rect 5840 8122 5874 8134
rect 5840 8065 5874 8084
rect 5840 8050 5874 8065
rect 5840 7996 5874 8012
rect 5840 7978 5874 7996
rect 5840 7927 5874 7940
rect 5840 7906 5874 7927
rect 5840 7858 5874 7868
rect 5840 7834 5874 7858
rect 5840 7789 5874 7796
rect 5840 7762 5874 7789
rect 5840 7720 5874 7724
rect 5840 7690 5874 7720
rect 5922 8461 5956 8465
rect 5922 8431 5956 8461
rect 5922 8388 5956 8391
rect 5922 8357 5956 8388
rect 5922 8315 5956 8317
rect 5922 8283 5956 8315
rect 5922 8242 5956 8243
rect 5922 8209 5956 8242
rect 5922 8135 5956 8169
rect 5922 8062 5956 8095
rect 5922 8061 5956 8062
rect 5922 7989 5956 8021
rect 5922 7987 5956 7989
rect 5922 7915 5956 7947
rect 5922 7913 5956 7915
rect 5922 7841 5956 7873
rect 5922 7839 5956 7841
rect 5922 7767 5956 7798
rect 5922 7764 5956 7767
rect 5922 7693 5956 7723
rect 5922 7689 5956 7693
rect 7114 8445 7148 8477
rect 7114 8443 7148 8445
rect 7114 8376 7148 8404
rect 7114 8370 7148 8376
rect 7114 8307 7148 8331
rect 7114 8297 7148 8307
rect 7114 8238 7148 8258
rect 7114 8224 7148 8238
rect 7114 8169 7148 8185
rect 7114 8151 7148 8169
rect 7114 8100 7148 8112
rect 7114 8078 7148 8100
rect 7114 8031 7148 8040
rect 7114 8006 7148 8031
rect 7114 7962 7148 7968
rect 7114 7934 7148 7962
rect 7114 7893 7148 7896
rect 7114 7862 7148 7893
rect 7114 7790 7148 7824
rect 7114 7720 7148 7752
rect 7114 7718 7148 7720
rect 5840 7651 5874 7652
rect 5840 7618 5874 7651
rect 6378 7632 6412 7666
rect 6450 7632 6484 7666
rect 6522 7632 6556 7666
rect 7114 7651 7148 7680
rect 7114 7646 7148 7651
rect 5840 7549 5874 7580
rect 5840 7546 5874 7549
rect 5840 7481 5874 7508
rect 5840 7474 5874 7481
rect 5840 7413 5874 7436
rect 5840 7402 5874 7413
rect 5840 7345 5874 7364
rect 5840 7330 5874 7345
rect 5840 7277 5874 7292
rect 5840 7258 5874 7277
rect 5840 7209 5874 7220
rect 5840 7186 5874 7209
rect 5840 7141 5874 7147
rect 5840 7113 5874 7141
rect 5840 7073 5874 7074
rect 5840 7040 5874 7073
rect 5840 6971 5874 7001
rect 5840 6967 5874 6971
rect 5840 6903 5874 6928
rect 5840 6894 5874 6903
rect 5840 6835 5874 6855
rect 5840 6821 5874 6835
rect 7032 7605 7066 7609
rect 7032 7575 7066 7605
rect 7032 7532 7066 7535
rect 7032 7501 7066 7532
rect 7032 7459 7066 7461
rect 7032 7427 7066 7459
rect 7032 7386 7066 7387
rect 7032 7353 7066 7386
rect 7032 7279 7066 7313
rect 7032 7206 7066 7239
rect 7032 7205 7066 7206
rect 7032 7133 7066 7165
rect 7032 7131 7066 7133
rect 7032 7059 7066 7091
rect 7032 7057 7066 7059
rect 7032 6985 7066 7017
rect 7032 6983 7066 6985
rect 7032 6911 7066 6942
rect 7032 6908 7066 6911
rect 7032 6837 7066 6867
rect 7032 6833 7066 6837
rect 7114 7583 7148 7608
rect 7114 7574 7148 7583
rect 7114 7515 7148 7536
rect 7114 7502 7148 7515
rect 7114 7447 7148 7464
rect 7114 7430 7148 7447
rect 7114 7379 7148 7392
rect 7114 7358 7148 7379
rect 7114 7311 7148 7320
rect 7114 7286 7148 7311
rect 7114 7243 7148 7248
rect 7114 7214 7148 7243
rect 7114 7175 7148 7176
rect 7114 7142 7148 7175
rect 7114 7073 7148 7104
rect 7114 7070 7148 7073
rect 7114 7005 7148 7032
rect 7114 6998 7148 7005
rect 7114 6937 7148 6960
rect 7114 6926 7148 6937
rect 7114 6869 7148 6888
rect 7114 6854 7148 6869
rect 5840 6767 5874 6782
rect 6680 6776 6714 6810
rect 6752 6776 6786 6810
rect 6824 6776 6858 6810
rect 7114 6801 7148 6816
rect 7114 6782 7148 6801
rect 5840 6748 5874 6767
rect 5840 6699 5874 6709
rect 5840 6675 5874 6699
rect 5840 6631 5874 6636
rect 5840 6602 5874 6631
rect 5840 6529 5874 6563
rect 5840 6461 5874 6490
rect 5840 6456 5874 6461
rect 5840 6393 5874 6417
rect 5840 6383 5874 6393
rect 5840 6325 5874 6344
rect 5840 6310 5874 6325
rect 5840 6257 5874 6271
rect 5840 6237 5874 6257
rect 5840 6189 5874 6198
rect 5840 6164 5874 6189
rect 5840 6121 5874 6125
rect 5840 6091 5874 6121
rect 5840 6019 5874 6052
rect 5840 6018 5874 6019
rect 5840 5951 5874 5979
rect 7032 6749 7066 6753
rect 7032 6719 7066 6749
rect 7032 6676 7066 6679
rect 7032 6645 7066 6676
rect 7032 6603 7066 6605
rect 7032 6571 7066 6603
rect 7032 6530 7066 6531
rect 7032 6497 7066 6530
rect 7032 6423 7066 6457
rect 7032 6350 7066 6383
rect 7032 6349 7066 6350
rect 7032 6277 7066 6309
rect 7032 6275 7066 6277
rect 7032 6203 7066 6235
rect 7032 6201 7066 6203
rect 7032 6129 7066 6161
rect 7032 6127 7066 6129
rect 7032 6055 7066 6086
rect 7032 6052 7066 6055
rect 7032 5981 7066 6011
rect 7032 5977 7066 5981
rect 7114 6733 7148 6744
rect 7114 6710 7148 6733
rect 7114 6665 7148 6672
rect 7114 6638 7148 6665
rect 7114 6597 7148 6600
rect 7114 6566 7148 6597
rect 7114 6495 7148 6528
rect 7114 6494 7148 6495
rect 7114 6427 7148 6456
rect 7114 6422 7148 6427
rect 7114 6359 7148 6384
rect 7114 6350 7148 6359
rect 7114 6291 7148 6312
rect 7114 6278 7148 6291
rect 7114 6223 7148 6240
rect 7114 6206 7148 6223
rect 7114 6155 7148 6168
rect 7114 6134 7148 6155
rect 7114 6087 7148 6096
rect 7114 6062 7148 6087
rect 7114 6019 7148 6024
rect 7114 5990 7148 6019
rect 5840 5945 5874 5951
rect 6378 5920 6412 5954
rect 6450 5920 6484 5954
rect 6522 5920 6556 5954
rect 7114 5951 7148 5952
rect 7114 5918 7148 5951
rect 5840 5883 5874 5906
rect 5840 5872 5874 5883
rect 5840 5815 5874 5833
rect 5840 5799 5874 5815
rect 5840 5747 5874 5760
rect 5840 5726 5874 5747
rect 5840 5679 5874 5687
rect 5840 5653 5874 5679
rect 5840 5611 5874 5614
rect 5840 5580 5874 5611
rect 5840 5509 5874 5541
rect 5840 5507 5874 5509
rect 5840 5441 5874 5468
rect 5840 5434 5874 5441
rect 5840 5373 5874 5395
rect 5840 5361 5874 5373
rect 5840 5305 5874 5322
rect 5840 5288 5874 5305
rect 5840 5237 5874 5249
rect 5840 5215 5874 5237
rect 5840 5169 5874 5176
rect 5840 5142 5874 5169
rect 5922 5893 5956 5897
rect 5922 5863 5956 5893
rect 5922 5820 5956 5823
rect 5922 5789 5956 5820
rect 5922 5747 5956 5749
rect 5922 5715 5956 5747
rect 5922 5674 5956 5675
rect 5922 5641 5956 5674
rect 5922 5567 5956 5601
rect 5922 5494 5956 5527
rect 5922 5493 5956 5494
rect 5922 5421 5956 5453
rect 5922 5419 5956 5421
rect 5922 5347 5956 5379
rect 5922 5345 5956 5347
rect 5922 5273 5956 5305
rect 5922 5271 5956 5273
rect 5922 5199 5956 5230
rect 5922 5196 5956 5199
rect 5922 5125 5956 5155
rect 5922 5121 5956 5125
rect 7114 5849 7148 5880
rect 7114 5846 7148 5849
rect 7114 5781 7148 5808
rect 7114 5774 7148 5781
rect 7114 5713 7148 5736
rect 7114 5702 7148 5713
rect 7114 5645 7148 5664
rect 7114 5630 7148 5645
rect 7114 5577 7148 5592
rect 7114 5558 7148 5577
rect 7114 5509 7148 5520
rect 7114 5486 7148 5509
rect 7114 5441 7148 5448
rect 7114 5414 7148 5441
rect 7114 5373 7148 5376
rect 7114 5342 7148 5373
rect 7114 5271 7148 5304
rect 7114 5270 7148 5271
rect 7114 5203 7148 5232
rect 7114 5198 7148 5203
rect 7114 5135 7148 5160
rect 7114 5126 7148 5135
rect 5840 5101 5874 5103
rect 5840 5069 5874 5101
rect 6076 5064 6110 5098
rect 6148 5064 6182 5098
rect 6220 5064 6254 5098
rect 7114 5067 7148 5088
rect 7114 5054 7148 5067
rect 5840 4999 5874 5030
rect 5840 4996 5874 4999
rect 5840 4931 5874 4957
rect 5840 4923 5874 4931
rect 5840 4863 5874 4884
rect 5840 4850 5874 4863
rect 5840 4795 5874 4811
rect 5840 4777 5874 4795
rect 5840 4727 5874 4738
rect 5840 4704 5874 4727
rect 5840 4659 5874 4665
rect 5840 4631 5874 4659
rect 5840 4591 5874 4592
rect 5840 4558 5874 4591
rect 5840 4489 5874 4519
rect 5840 4485 5874 4489
rect 5840 4421 5874 4446
rect 5840 4412 5874 4421
rect 5840 4353 5874 4373
rect 5840 4339 5874 4353
rect 5840 4285 5874 4300
rect 5840 4266 5874 4285
rect 5922 5037 5956 5041
rect 5922 5007 5956 5037
rect 5922 4964 5956 4967
rect 5922 4933 5956 4964
rect 5922 4891 5956 4893
rect 5922 4859 5956 4891
rect 5922 4818 5956 4819
rect 5922 4785 5956 4818
rect 5922 4711 5956 4745
rect 5922 4638 5956 4671
rect 5922 4637 5956 4638
rect 5922 4565 5956 4597
rect 5922 4563 5956 4565
rect 5922 4491 5956 4523
rect 5922 4489 5956 4491
rect 5922 4417 5956 4449
rect 5922 4415 5956 4417
rect 5922 4343 5956 4374
rect 5922 4340 5956 4343
rect 5922 4269 5956 4299
rect 5922 4265 5956 4269
rect 7114 4999 7148 5016
rect 7114 4982 7148 4999
rect 7114 4931 7148 4944
rect 7114 4910 7148 4931
rect 7114 4863 7148 4872
rect 7114 4838 7148 4863
rect 7114 4795 7148 4800
rect 7114 4766 7148 4795
rect 7114 4727 7148 4728
rect 7114 4694 7148 4727
rect 7114 4625 7148 4656
rect 7114 4622 7148 4625
rect 7114 4557 7148 4584
rect 7114 4550 7148 4557
rect 7114 4489 7148 4512
rect 7114 4478 7148 4489
rect 7114 4421 7148 4440
rect 7114 4406 7148 4421
rect 7114 4353 7148 4368
rect 7114 4334 7148 4353
rect 7114 4285 7148 4296
rect 7114 4262 7148 4285
rect 5840 4217 5874 4227
rect 5840 4193 5874 4217
rect 6378 4208 6412 4242
rect 6450 4208 6484 4242
rect 6522 4208 6556 4242
rect 7114 4217 7148 4224
rect 7114 4190 7148 4217
rect 5840 4149 5874 4154
rect 5840 4120 5874 4149
rect 5840 4047 5874 4081
rect 6378 4050 6412 4084
rect 6450 4050 6484 4084
rect 6522 4050 6556 4084
rect 7114 4149 7148 4152
rect 7114 4118 7148 4149
rect 5840 3974 5874 4008
rect 7114 4046 7148 4080
rect 5978 3936 6010 3970
rect 6010 3936 6012 3970
rect 6064 3936 6078 3970
rect 6078 3936 6098 3970
rect 6150 3936 6180 3970
rect 6180 3936 6184 3970
rect 6237 3936 6248 3970
rect 6248 3936 6271 3970
rect 6671 3936 6690 3970
rect 6690 3936 6705 3970
rect 6752 3936 6758 3970
rect 6758 3936 6786 3970
rect 6833 3936 6860 3970
rect 6860 3936 6867 3970
rect 6914 3936 6928 3970
rect 6928 3936 6948 3970
rect 6995 3936 6996 3970
rect 6996 3936 7029 3970
rect 7076 3936 7110 3970
rect 7423 11349 7431 11359
rect 7431 11349 7457 11359
rect 7423 11325 7457 11349
rect 7423 11281 7431 11287
rect 7431 11281 7457 11287
rect 7423 11253 7457 11281
rect 7927 11251 8537 11429
rect 8576 11395 8610 11429
rect 8649 11395 8683 11429
rect 8722 11395 8756 11429
rect 8795 11395 8829 11429
rect 8868 11395 8902 11429
rect 8576 11323 8610 11357
rect 8649 11323 8683 11357
rect 8722 11323 8756 11357
rect 8795 11323 8829 11357
rect 8868 11323 8902 11357
rect 9899 11417 9929 11431
rect 9929 11417 9933 11431
rect 9899 11397 9933 11417
rect 9899 11349 9929 11358
rect 9929 11349 9933 11358
rect 9899 11324 9933 11349
rect 8576 11251 8610 11285
rect 8649 11251 8683 11285
rect 8722 11251 8756 11285
rect 8795 11251 8829 11285
rect 8868 11251 8902 11285
rect 9899 11281 9929 11285
rect 9929 11281 9933 11285
rect 9899 11251 9933 11281
rect 7423 11213 7431 11215
rect 7431 11213 7457 11215
rect 7423 11181 7457 11213
rect 7423 11111 7457 11143
rect 7423 11109 7431 11111
rect 7431 11109 7457 11111
rect 7423 11043 7457 11071
rect 7423 11037 7431 11043
rect 7431 11037 7457 11043
rect 7423 10975 7457 10999
rect 7423 10965 7431 10975
rect 7431 10965 7457 10975
rect 7423 10907 7457 10927
rect 7423 10893 7431 10907
rect 7431 10893 7457 10907
rect 7423 10839 7457 10855
rect 7423 10821 7431 10839
rect 7431 10821 7457 10839
rect 7423 10771 7457 10783
rect 7423 10749 7431 10771
rect 7431 10749 7457 10771
rect 7423 10703 7457 10711
rect 7423 10677 7431 10703
rect 7431 10677 7457 10703
rect 7423 10635 7457 10639
rect 7423 10605 7431 10635
rect 7431 10605 7457 10635
rect 7423 10533 7431 10567
rect 7431 10533 7457 10567
rect 7423 10465 7431 10495
rect 7431 10465 7457 10495
rect 7423 10461 7457 10465
rect 7608 11224 7642 11228
rect 7608 11194 7642 11224
rect 9718 11224 9752 11228
rect 9718 11194 9752 11224
rect 7608 11151 7642 11154
rect 7608 11120 7642 11151
rect 9718 11151 9752 11154
rect 9718 11120 9752 11151
rect 7608 11078 7642 11080
rect 7608 11046 7642 11078
rect 9718 11078 9752 11080
rect 9718 11046 9752 11078
rect 7608 11005 7642 11006
rect 7608 10972 7642 11005
rect 9718 11005 9752 11006
rect 9718 10972 9752 11005
rect 7608 10898 7642 10932
rect 9718 10898 9752 10932
rect 7608 10825 7642 10858
rect 7608 10824 7642 10825
rect 9718 10825 9752 10858
rect 9718 10824 9752 10825
rect 7608 10752 7642 10784
rect 7608 10750 7642 10752
rect 9718 10752 9752 10784
rect 9718 10750 9752 10752
rect 7608 10678 7642 10710
rect 7608 10676 7642 10678
rect 9718 10678 9752 10710
rect 9718 10676 9752 10678
rect 7608 10604 7642 10636
rect 7608 10602 7642 10604
rect 9718 10604 9752 10636
rect 9718 10602 9752 10604
rect 7608 10530 7642 10561
rect 7608 10527 7642 10530
rect 9718 10530 9752 10561
rect 9718 10527 9752 10530
rect 7608 10456 7642 10486
rect 7608 10452 7642 10456
rect 9718 10456 9752 10486
rect 9718 10452 9752 10456
rect 9899 11179 9933 11212
rect 9899 11178 9929 11179
rect 9929 11178 9933 11179
rect 9899 11111 9933 11139
rect 9899 11105 9929 11111
rect 9929 11105 9933 11111
rect 9899 11043 9933 11066
rect 9899 11032 9929 11043
rect 9929 11032 9933 11043
rect 9899 10975 9933 10993
rect 9899 10959 9929 10975
rect 9929 10959 9933 10975
rect 9899 10907 9933 10920
rect 9899 10886 9929 10907
rect 9929 10886 9933 10907
rect 9899 10839 9933 10847
rect 9899 10813 9929 10839
rect 9929 10813 9933 10839
rect 9899 10771 9933 10774
rect 9899 10740 9929 10771
rect 9929 10740 9933 10771
rect 9899 10669 9929 10701
rect 9929 10669 9933 10701
rect 9899 10667 9933 10669
rect 9899 10601 9929 10628
rect 9929 10601 9933 10628
rect 9899 10594 9933 10601
rect 9899 10533 9929 10555
rect 9929 10533 9933 10555
rect 9899 10521 9933 10533
rect 9899 10465 9929 10482
rect 9929 10465 9933 10482
rect 9899 10448 9933 10465
rect 7423 10397 7431 10423
rect 7431 10397 7457 10423
rect 7423 10389 7457 10397
rect 9899 10397 9929 10409
rect 9929 10397 9933 10409
rect 7423 10329 7431 10351
rect 7431 10329 7457 10351
rect 7423 10317 7457 10329
rect 7423 10261 7431 10279
rect 7431 10261 7457 10279
rect 7423 10245 7457 10261
rect 7927 10218 8537 10396
rect 8576 10362 8610 10396
rect 8649 10362 8683 10396
rect 8722 10362 8756 10396
rect 8795 10362 8829 10396
rect 8868 10362 8902 10396
rect 9899 10375 9933 10397
rect 8576 10290 8610 10324
rect 8649 10290 8683 10324
rect 8722 10290 8756 10324
rect 8795 10290 8829 10324
rect 8868 10290 8902 10324
rect 8576 10218 8610 10252
rect 8649 10218 8683 10252
rect 8722 10218 8756 10252
rect 8795 10218 8829 10252
rect 8868 10218 8902 10252
rect 9899 10329 9929 10336
rect 9929 10329 9933 10336
rect 9899 10302 9933 10329
rect 9899 10261 9929 10263
rect 9929 10261 9933 10263
rect 9899 10229 9933 10261
rect 7423 10193 7431 10207
rect 7431 10193 7457 10207
rect 7423 10173 7457 10193
rect 9899 10159 9933 10190
rect 9899 10156 9929 10159
rect 9929 10156 9933 10159
rect 7423 10125 7431 10135
rect 7431 10125 7457 10135
rect 7423 10101 7457 10125
rect 7423 10057 7431 10063
rect 7431 10057 7457 10063
rect 7423 10029 7457 10057
rect 7423 9989 7431 9991
rect 7431 9989 7457 9991
rect 7423 9957 7457 9989
rect 7423 9887 7457 9919
rect 7423 9885 7431 9887
rect 7431 9885 7457 9887
rect 7423 9819 7457 9847
rect 7423 9813 7431 9819
rect 7431 9813 7457 9819
rect 7423 9751 7457 9775
rect 7423 9741 7431 9751
rect 7431 9741 7457 9751
rect 7423 9683 7457 9703
rect 7423 9669 7431 9683
rect 7431 9669 7457 9683
rect 7423 9615 7457 9631
rect 7423 9597 7431 9615
rect 7431 9597 7457 9615
rect 7423 9547 7457 9559
rect 7423 9525 7431 9547
rect 7431 9525 7457 9547
rect 7423 9479 7457 9487
rect 7423 9453 7431 9479
rect 7431 9453 7457 9479
rect 7423 9411 7457 9415
rect 7423 9381 7431 9411
rect 7431 9381 7457 9411
rect 7608 10138 7642 10142
rect 7608 10108 7642 10138
rect 9718 10138 9752 10142
rect 9718 10108 9752 10138
rect 7608 10065 7642 10068
rect 7608 10034 7642 10065
rect 9718 10065 9752 10068
rect 9718 10034 9752 10065
rect 7608 9992 7642 9994
rect 7608 9960 7642 9992
rect 9718 9992 9752 9994
rect 9718 9960 9752 9992
rect 7608 9919 7642 9920
rect 7608 9886 7642 9919
rect 9718 9919 9752 9920
rect 9718 9886 9752 9919
rect 7608 9812 7642 9846
rect 9718 9812 9752 9846
rect 7608 9739 7642 9772
rect 7608 9738 7642 9739
rect 9718 9739 9752 9772
rect 9718 9738 9752 9739
rect 7608 9666 7642 9698
rect 7608 9664 7642 9666
rect 9718 9666 9752 9698
rect 9718 9664 9752 9666
rect 7608 9592 7642 9624
rect 7608 9590 7642 9592
rect 9718 9592 9752 9624
rect 9718 9590 9752 9592
rect 7608 9518 7642 9550
rect 7608 9516 7642 9518
rect 9718 9518 9752 9550
rect 9718 9516 9752 9518
rect 7608 9444 7642 9475
rect 7608 9441 7642 9444
rect 9718 9444 9752 9475
rect 9718 9441 9752 9444
rect 7608 9370 7642 9400
rect 7608 9366 7642 9370
rect 9718 9370 9752 9400
rect 9718 9366 9752 9370
rect 9899 10091 9933 10117
rect 9899 10083 9929 10091
rect 9929 10083 9933 10091
rect 9899 10023 9933 10044
rect 9899 10010 9929 10023
rect 9929 10010 9933 10023
rect 9899 9955 9933 9971
rect 9899 9937 9929 9955
rect 9929 9937 9933 9955
rect 9899 9887 9933 9898
rect 9899 9864 9929 9887
rect 9929 9864 9933 9887
rect 9899 9819 9933 9825
rect 9899 9791 9929 9819
rect 9929 9791 9933 9819
rect 9899 9751 9933 9752
rect 9899 9718 9929 9751
rect 9929 9718 9933 9751
rect 9899 9649 9929 9679
rect 9929 9649 9933 9679
rect 9899 9645 9933 9649
rect 9899 9581 9929 9606
rect 9929 9581 9933 9606
rect 9899 9572 9933 9581
rect 9899 9513 9929 9533
rect 9929 9513 9933 9533
rect 9899 9499 9933 9513
rect 9899 9445 9929 9460
rect 9929 9445 9933 9460
rect 9899 9426 9933 9445
rect 9899 9377 9929 9387
rect 9929 9377 9933 9387
rect 9899 9353 9933 9377
rect 7423 9309 7431 9343
rect 7431 9309 7457 9343
rect 7927 9309 7961 9343
rect 7999 9309 8033 9343
rect 8071 9309 8105 9343
rect 8143 9309 8177 9343
rect 8215 9309 8249 9343
rect 8287 9309 8321 9343
rect 8359 9309 8393 9343
rect 8431 9309 8465 9343
rect 8503 9309 8537 9343
rect 8576 9309 8610 9343
rect 8649 9309 8683 9343
rect 8722 9309 8756 9343
rect 8795 9309 8829 9343
rect 8868 9309 8902 9343
rect 9899 9309 9929 9314
rect 9929 9309 9933 9314
rect 7423 9241 7431 9271
rect 7431 9241 7457 9271
rect 7423 9237 7457 9241
rect 7423 9173 7431 9199
rect 7431 9173 7457 9199
rect 7423 9165 7457 9173
rect 7423 9105 7431 9127
rect 7431 9105 7457 9127
rect 7423 9093 7457 9105
rect 7423 9037 7431 9055
rect 7431 9037 7457 9055
rect 7423 9021 7457 9037
rect 7423 8969 7431 8983
rect 7431 8969 7457 8983
rect 7423 8949 7457 8969
rect 7423 8901 7431 8911
rect 7431 8901 7457 8911
rect 7423 8877 7457 8901
rect 7423 8833 7431 8839
rect 7431 8833 7457 8839
rect 7423 8805 7457 8833
rect 7423 8765 7431 8767
rect 7431 8765 7457 8767
rect 7423 8733 7457 8765
rect 7423 8663 7457 8695
rect 7423 8661 7431 8663
rect 7431 8661 7457 8663
rect 7423 8595 7457 8623
rect 7423 8589 7431 8595
rect 7431 8589 7457 8595
rect 7423 8527 7457 8551
rect 7423 8517 7431 8527
rect 7431 8517 7457 8527
rect 7608 9282 7642 9286
rect 7608 9252 7642 9282
rect 9718 9282 9752 9286
rect 9718 9252 9752 9282
rect 7608 9209 7642 9212
rect 7608 9178 7642 9209
rect 9718 9209 9752 9212
rect 9718 9178 9752 9209
rect 7608 9136 7642 9138
rect 7608 9104 7642 9136
rect 9718 9136 9752 9138
rect 9718 9104 9752 9136
rect 7608 9063 7642 9064
rect 7608 9030 7642 9063
rect 9718 9063 9752 9064
rect 9718 9030 9752 9063
rect 7608 8956 7642 8990
rect 9718 8956 9752 8990
rect 7608 8883 7642 8916
rect 7608 8882 7642 8883
rect 9718 8883 9752 8916
rect 9718 8882 9752 8883
rect 7608 8810 7642 8842
rect 7608 8808 7642 8810
rect 9718 8810 9752 8842
rect 9718 8808 9752 8810
rect 7608 8736 7642 8768
rect 7608 8734 7642 8736
rect 9718 8736 9752 8768
rect 9718 8734 9752 8736
rect 7608 8662 7642 8694
rect 7608 8660 7642 8662
rect 9718 8662 9752 8694
rect 9718 8660 9752 8662
rect 7608 8588 7642 8619
rect 7608 8585 7642 8588
rect 9718 8588 9752 8619
rect 9718 8585 9752 8588
rect 7608 8514 7642 8544
rect 7608 8510 7642 8514
rect 9718 8514 9752 8544
rect 9718 8510 9752 8514
rect 9899 9280 9933 9309
rect 9899 9207 9933 9241
rect 9899 9139 9933 9168
rect 9899 9134 9929 9139
rect 9929 9134 9933 9139
rect 9899 9071 9933 9095
rect 9899 9061 9929 9071
rect 9929 9061 9933 9071
rect 9899 9003 9933 9022
rect 9899 8988 9929 9003
rect 9929 8988 9933 9003
rect 9899 8935 9933 8949
rect 9899 8915 9929 8935
rect 9929 8915 9933 8935
rect 9899 8867 9933 8876
rect 9899 8842 9929 8867
rect 9929 8842 9933 8867
rect 9899 8799 9933 8803
rect 9899 8769 9929 8799
rect 9929 8769 9933 8799
rect 9899 8697 9929 8730
rect 9929 8697 9933 8730
rect 9899 8696 9933 8697
rect 9899 8629 9929 8657
rect 9929 8629 9933 8657
rect 9899 8623 9933 8629
rect 9899 8561 9929 8584
rect 9929 8561 9933 8584
rect 9899 8550 9933 8561
rect 9899 8493 9929 8511
rect 9929 8493 9933 8511
rect 7423 8459 7457 8479
rect 7423 8445 7431 8459
rect 7431 8445 7457 8459
rect 7927 8449 7961 8483
rect 7999 8449 8033 8483
rect 8071 8449 8105 8483
rect 8143 8449 8177 8483
rect 8215 8449 8249 8483
rect 8287 8449 8321 8483
rect 8359 8449 8393 8483
rect 8431 8449 8465 8483
rect 8503 8449 8537 8483
rect 8576 8449 8610 8483
rect 8649 8449 8683 8483
rect 8722 8449 8756 8483
rect 8795 8449 8829 8483
rect 8868 8449 8902 8483
rect 9899 8477 9933 8493
rect 9899 8425 9929 8438
rect 9929 8425 9933 8438
rect 7423 8391 7457 8407
rect 7423 8373 7431 8391
rect 7431 8373 7457 8391
rect 7423 8323 7457 8335
rect 7423 8301 7431 8323
rect 7431 8301 7457 8323
rect 7423 8255 7457 8263
rect 7423 8229 7431 8255
rect 7431 8229 7457 8255
rect 7927 8253 8537 8359
rect 8576 8325 8610 8359
rect 8649 8325 8683 8359
rect 8722 8325 8756 8359
rect 8795 8325 8829 8359
rect 8868 8325 8902 8359
rect 9899 8404 9933 8425
rect 9899 8357 9929 8365
rect 9929 8357 9933 8365
rect 9899 8331 9933 8357
rect 9899 8289 9929 8292
rect 9929 8289 9933 8292
rect 8576 8253 8610 8287
rect 8649 8253 8683 8287
rect 8722 8253 8756 8287
rect 8795 8253 8829 8287
rect 8868 8253 8902 8287
rect 9899 8258 9933 8289
rect 7423 8187 7457 8191
rect 7423 8157 7431 8187
rect 7431 8157 7457 8187
rect 7423 8085 7431 8119
rect 7431 8085 7457 8119
rect 7423 8017 7431 8047
rect 7431 8017 7457 8047
rect 7423 8013 7457 8017
rect 7423 7949 7431 7975
rect 7431 7949 7457 7975
rect 7423 7941 7457 7949
rect 7423 7881 7431 7903
rect 7431 7881 7457 7903
rect 7423 7869 7457 7881
rect 7423 7813 7431 7831
rect 7431 7813 7457 7831
rect 7423 7797 7457 7813
rect 7423 7745 7431 7759
rect 7431 7745 7457 7759
rect 7423 7725 7457 7745
rect 7423 7677 7431 7687
rect 7431 7677 7457 7687
rect 7423 7653 7457 7677
rect 7423 7609 7431 7615
rect 7431 7609 7457 7615
rect 7423 7581 7457 7609
rect 7423 7541 7431 7543
rect 7431 7541 7457 7543
rect 7423 7509 7457 7541
rect 7423 7439 7457 7471
rect 7423 7437 7431 7439
rect 7431 7437 7457 7439
rect 7608 8196 7642 8200
rect 7608 8166 7642 8196
rect 9718 8196 9752 8200
rect 9718 8166 9752 8196
rect 7608 8123 7642 8126
rect 7608 8092 7642 8123
rect 9718 8123 9752 8126
rect 9718 8092 9752 8123
rect 7608 8050 7642 8052
rect 7608 8018 7642 8050
rect 9718 8050 9752 8052
rect 9718 8018 9752 8050
rect 7608 7977 7642 7978
rect 7608 7944 7642 7977
rect 9718 7977 9752 7978
rect 9718 7944 9752 7977
rect 7608 7870 7642 7904
rect 9718 7870 9752 7904
rect 7608 7797 7642 7830
rect 7608 7796 7642 7797
rect 9718 7797 9752 7830
rect 9718 7796 9752 7797
rect 7608 7724 7642 7756
rect 7608 7722 7642 7724
rect 9718 7724 9752 7756
rect 9718 7722 9752 7724
rect 7608 7650 7642 7682
rect 7608 7648 7642 7650
rect 9718 7650 9752 7682
rect 9718 7648 9752 7650
rect 7608 7576 7642 7608
rect 7608 7574 7642 7576
rect 9718 7576 9752 7608
rect 9718 7574 9752 7576
rect 7608 7502 7642 7533
rect 7608 7499 7642 7502
rect 9718 7502 9752 7533
rect 9718 7499 9752 7502
rect 7608 7428 7642 7458
rect 7608 7424 7642 7428
rect 9718 7428 9752 7458
rect 9718 7424 9752 7428
rect 9899 8187 9933 8219
rect 9899 8185 9929 8187
rect 9929 8185 9933 8187
rect 9899 8119 9933 8146
rect 9899 8112 9929 8119
rect 9929 8112 9933 8119
rect 9899 8051 9933 8073
rect 9899 8039 9929 8051
rect 9929 8039 9933 8051
rect 10317 8006 10337 8040
rect 10337 8006 10351 8040
rect 10389 8006 10405 8040
rect 10405 8006 10423 8040
rect 10461 8006 10473 8040
rect 10473 8006 10495 8040
rect 10533 8006 10541 8040
rect 10541 8006 10567 8040
rect 10605 8006 10609 8040
rect 10609 8006 10639 8040
rect 10677 8006 10711 8040
rect 10749 8006 10779 8040
rect 10779 8006 10783 8040
rect 10821 8006 10847 8040
rect 10847 8006 10855 8040
rect 10893 8006 10915 8040
rect 10915 8006 10927 8040
rect 10965 8006 10983 8040
rect 10983 8006 10999 8040
rect 11037 8006 11051 8040
rect 11051 8006 11071 8040
rect 11109 8006 11119 8040
rect 11119 8006 11143 8040
rect 11181 8006 11187 8040
rect 11187 8006 11215 8040
rect 11253 8006 11255 8040
rect 11255 8006 11287 8040
rect 11325 8006 11357 8040
rect 11357 8006 11359 8040
rect 11397 8006 11425 8040
rect 11425 8006 11431 8040
rect 11469 8006 11493 8040
rect 11493 8006 11503 8040
rect 11541 8006 11561 8040
rect 11561 8006 11575 8040
rect 11613 8006 11629 8040
rect 11629 8006 11647 8040
rect 11685 8006 11697 8040
rect 11697 8006 11719 8040
rect 11757 8006 11765 8040
rect 11765 8006 11791 8040
rect 11829 8006 11833 8040
rect 11833 8006 11863 8040
rect 11901 8006 11935 8040
rect 11973 8006 12003 8040
rect 12003 8006 12007 8040
rect 12045 8006 12071 8040
rect 12071 8006 12079 8040
rect 12117 8006 12139 8040
rect 12139 8006 12151 8040
rect 12189 8006 12207 8040
rect 12207 8006 12223 8040
rect 12261 8006 12275 8040
rect 12275 8006 12295 8040
rect 12333 8006 12343 8040
rect 12343 8006 12367 8040
rect 12405 8006 12411 8040
rect 12411 8006 12439 8040
rect 12478 8006 12479 8040
rect 12479 8006 12512 8040
rect 12551 8006 12581 8040
rect 12581 8006 12585 8040
rect 12624 8006 12649 8040
rect 12649 8006 12658 8040
rect 12697 8006 12717 8040
rect 12717 8006 12731 8040
rect 12770 8006 12785 8040
rect 12785 8006 12804 8040
rect 9899 7983 9933 8000
rect 9899 7966 9929 7983
rect 9929 7966 9933 7983
rect 9899 7915 9933 7927
rect 9899 7893 9929 7915
rect 9929 7893 9933 7915
rect 9899 7847 9933 7854
rect 9899 7820 9929 7847
rect 9929 7820 9933 7847
rect 9899 7779 9933 7782
rect 9899 7748 9929 7779
rect 9929 7748 9933 7779
rect 9899 7677 9929 7710
rect 9929 7677 9933 7710
rect 9899 7676 9933 7677
rect 9899 7609 9929 7638
rect 9929 7609 9933 7638
rect 9899 7604 9933 7609
rect 9899 7541 9929 7566
rect 9929 7541 9933 7566
rect 9899 7532 9933 7541
rect 9899 7473 9929 7494
rect 9929 7473 9933 7494
rect 9899 7460 9933 7473
rect 9899 7405 9929 7422
rect 9929 7405 9933 7422
rect 7423 7371 7457 7399
rect 7423 7365 7431 7371
rect 7431 7365 7457 7371
rect 7423 7303 7457 7327
rect 7423 7293 7431 7303
rect 7431 7293 7457 7303
rect 7423 7235 7457 7255
rect 7423 7221 7431 7235
rect 7431 7221 7457 7235
rect 7927 7223 8537 7401
rect 8576 7367 8610 7401
rect 8649 7367 8683 7401
rect 8722 7367 8756 7401
rect 8795 7367 8829 7401
rect 8868 7367 8902 7401
rect 9899 7388 9933 7405
rect 9899 7337 9929 7350
rect 9929 7337 9933 7350
rect 8576 7295 8610 7329
rect 8649 7295 8683 7329
rect 8722 7295 8756 7329
rect 8795 7295 8829 7329
rect 8868 7295 8902 7329
rect 9899 7316 9933 7337
rect 8576 7223 8610 7257
rect 8649 7223 8683 7257
rect 8722 7223 8756 7257
rect 8795 7223 8829 7257
rect 8868 7223 8902 7257
rect 9899 7269 9929 7278
rect 9929 7269 9933 7278
rect 9899 7244 9933 7269
rect 7423 7167 7457 7183
rect 7423 7149 7431 7167
rect 7431 7149 7457 7167
rect 7423 7099 7457 7111
rect 7423 7077 7431 7099
rect 7431 7077 7457 7099
rect 7423 7031 7457 7039
rect 7423 7005 7431 7031
rect 7431 7005 7457 7031
rect 7423 6963 7457 6967
rect 9899 7201 9929 7206
rect 9929 7201 9933 7206
rect 9899 7172 9933 7201
rect 9899 7133 9929 7134
rect 9929 7133 9933 7134
rect 9899 7100 9933 7133
rect 9899 7031 9933 7062
rect 9899 7028 9929 7031
rect 9929 7028 9933 7031
rect 9899 6963 9933 6990
rect 7423 6933 7431 6963
rect 7431 6933 7457 6963
rect 9899 6956 9929 6963
rect 9929 6956 9933 6963
rect 7423 6861 7431 6895
rect 7431 6861 7457 6895
rect 7423 6793 7431 6823
rect 7431 6793 7457 6823
rect 7423 6789 7457 6793
rect 7423 6725 7431 6751
rect 7431 6725 7457 6751
rect 7423 6717 7457 6725
rect 7423 6657 7431 6679
rect 7431 6657 7457 6679
rect 9899 6895 9933 6918
rect 9899 6884 9929 6895
rect 9929 6884 9933 6895
rect 9899 6827 9933 6846
rect 9899 6812 9929 6827
rect 9929 6812 9933 6827
rect 9899 6759 9933 6774
rect 9899 6740 9929 6759
rect 9929 6740 9933 6759
rect 9899 6691 9933 6702
rect 7423 6645 7457 6657
rect 7423 6589 7431 6607
rect 7431 6589 7457 6607
rect 7423 6573 7457 6589
rect 7423 6521 7431 6535
rect 7431 6521 7457 6535
rect 7423 6501 7457 6521
rect 8151 6491 8761 6669
rect 8800 6635 8834 6669
rect 8873 6635 8907 6669
rect 8946 6635 8980 6669
rect 9019 6635 9053 6669
rect 9092 6635 9126 6669
rect 9899 6668 9929 6691
rect 9929 6668 9933 6691
rect 8800 6563 8834 6597
rect 8873 6563 8907 6597
rect 8946 6563 8980 6597
rect 9019 6563 9053 6597
rect 9092 6563 9126 6597
rect 9899 6623 9933 6630
rect 9899 6596 9929 6623
rect 9929 6596 9933 6623
rect 9899 6555 9933 6558
rect 8800 6491 8834 6525
rect 8873 6491 8907 6525
rect 8946 6491 8980 6525
rect 9019 6491 9053 6525
rect 9092 6491 9126 6525
rect 9899 6524 9929 6555
rect 9929 6524 9933 6555
rect 7423 6453 7431 6463
rect 7431 6453 7457 6463
rect 7423 6429 7457 6453
rect 7423 6385 7431 6391
rect 7431 6385 7457 6391
rect 7423 6357 7457 6385
rect 7423 6317 7431 6319
rect 7431 6317 7457 6319
rect 7423 6285 7457 6317
rect 7423 6215 7457 6247
rect 7423 6213 7431 6215
rect 7431 6213 7457 6215
rect 7423 6147 7457 6175
rect 7423 6141 7431 6147
rect 7431 6141 7457 6147
rect 7423 6079 7457 6103
rect 7423 6069 7431 6079
rect 7431 6069 7457 6079
rect 7423 6011 7457 6031
rect 7423 5997 7431 6011
rect 7431 5997 7457 6011
rect 7423 5943 7457 5959
rect 7423 5925 7431 5943
rect 7431 5925 7457 5943
rect 7423 5875 7457 5887
rect 7423 5853 7431 5875
rect 7431 5853 7457 5875
rect 7423 5807 7457 5815
rect 7423 5781 7431 5807
rect 7431 5781 7457 5807
rect 7423 5739 7457 5743
rect 7423 5709 7431 5739
rect 7431 5709 7457 5739
rect 7423 5637 7431 5671
rect 7431 5637 7457 5671
rect 7608 6464 7642 6468
rect 7608 6434 7642 6464
rect 9718 6464 9752 6468
rect 9718 6434 9752 6464
rect 7608 6361 7642 6392
rect 7608 6358 7642 6361
rect 9718 6361 9752 6392
rect 9718 6358 9752 6361
rect 7608 6292 7642 6316
rect 7608 6282 7642 6292
rect 9718 6292 9752 6316
rect 9718 6282 9752 6292
rect 7608 6223 7642 6239
rect 7608 6205 7642 6223
rect 9718 6223 9752 6239
rect 9718 6205 9752 6223
rect 7608 6154 7642 6162
rect 7608 6128 7642 6154
rect 9718 6154 9752 6162
rect 9718 6128 9752 6154
rect 7608 6051 7642 6085
rect 9718 6051 9752 6085
rect 7608 5981 7642 6008
rect 7608 5974 7642 5981
rect 9718 5981 9752 6008
rect 9718 5974 9752 5981
rect 7608 5912 7642 5931
rect 7608 5897 7642 5912
rect 9718 5912 9752 5931
rect 9718 5897 9752 5912
rect 7608 5843 7642 5854
rect 7608 5820 7642 5843
rect 9718 5843 9752 5854
rect 9718 5820 9752 5843
rect 7608 5774 7642 5777
rect 7608 5743 7642 5774
rect 9718 5774 9752 5777
rect 9718 5743 9752 5774
rect 7608 5670 7642 5700
rect 7608 5666 7642 5670
rect 9718 5670 9752 5700
rect 9718 5666 9752 5670
rect 9899 6453 9929 6486
rect 9929 6453 9933 6486
rect 9899 6452 9933 6453
rect 9899 6385 9929 6414
rect 9929 6385 9933 6414
rect 9899 6380 9933 6385
rect 9899 6317 9929 6342
rect 9929 6317 9933 6342
rect 9899 6308 9933 6317
rect 9899 6249 9929 6270
rect 9929 6249 9933 6270
rect 9899 6236 9933 6249
rect 9899 6181 9929 6198
rect 9929 6181 9933 6198
rect 9899 6164 9933 6181
rect 9899 6113 9929 6126
rect 9929 6113 9933 6126
rect 9899 6092 9933 6113
rect 9899 6045 9929 6054
rect 9929 6045 9933 6054
rect 9899 6020 9933 6045
rect 9899 5977 9929 5982
rect 9929 5977 9933 5982
rect 9899 5948 9933 5977
rect 9899 5909 9929 5910
rect 9929 5909 9933 5910
rect 9899 5876 9933 5909
rect 9899 5807 9933 5838
rect 9899 5804 9929 5807
rect 9929 5804 9933 5807
rect 9899 5739 9933 5766
rect 9899 5732 9929 5739
rect 9929 5732 9933 5739
rect 9899 5671 9933 5694
rect 9899 5660 9929 5671
rect 9929 5660 9933 5671
rect 7423 5569 7431 5599
rect 7431 5569 7457 5599
rect 7423 5565 7457 5569
rect 7423 5501 7431 5527
rect 7431 5501 7457 5527
rect 7423 5493 7457 5501
rect 7423 5433 7431 5455
rect 7431 5433 7457 5455
rect 7423 5421 7457 5433
rect 8151 5432 8761 5610
rect 8800 5576 8834 5610
rect 8873 5576 8907 5610
rect 8946 5576 8980 5610
rect 9019 5576 9053 5610
rect 9092 5576 9126 5610
rect 9899 5603 9933 5622
rect 9899 5588 9929 5603
rect 9929 5588 9933 5603
rect 8800 5504 8834 5538
rect 8873 5504 8907 5538
rect 8946 5504 8980 5538
rect 9019 5504 9053 5538
rect 9092 5504 9126 5538
rect 8800 5432 8834 5466
rect 8873 5432 8907 5466
rect 8946 5432 8980 5466
rect 9019 5432 9053 5466
rect 9092 5432 9126 5466
rect 9899 5535 9933 5550
rect 9899 5516 9929 5535
rect 9929 5516 9933 5535
rect 9899 5467 9933 5478
rect 9899 5444 9929 5467
rect 9929 5444 9933 5467
rect 9899 5399 9933 5406
rect 7423 5365 7431 5383
rect 7431 5365 7457 5383
rect 7423 5349 7457 5365
rect 7423 5297 7431 5311
rect 7431 5297 7457 5311
rect 7423 5277 7457 5297
rect 7423 5229 7431 5239
rect 7431 5229 7457 5239
rect 7423 5205 7457 5229
rect 7423 5161 7431 5167
rect 7431 5161 7457 5167
rect 7423 5133 7457 5161
rect 7423 5093 7431 5095
rect 7431 5093 7457 5095
rect 7423 5061 7457 5093
rect 7423 4991 7457 5023
rect 7423 4989 7431 4991
rect 7431 4989 7457 4991
rect 7423 4923 7457 4951
rect 7423 4917 7431 4923
rect 7431 4917 7457 4923
rect 7423 4855 7457 4879
rect 7423 4845 7431 4855
rect 7431 4845 7457 4855
rect 7423 4787 7457 4807
rect 7423 4773 7431 4787
rect 7431 4773 7457 4787
rect 7423 4719 7457 4735
rect 7423 4701 7431 4719
rect 7431 4701 7457 4719
rect 7423 4651 7457 4663
rect 7423 4629 7431 4651
rect 7431 4629 7457 4651
rect 7608 5378 7642 5382
rect 7608 5348 7642 5378
rect 9718 5378 9752 5382
rect 9718 5348 9752 5378
rect 7608 5305 7642 5308
rect 7608 5274 7642 5305
rect 9718 5305 9752 5308
rect 9718 5274 9752 5305
rect 7608 5232 7642 5234
rect 7608 5200 7642 5232
rect 9718 5232 9752 5234
rect 9718 5200 9752 5232
rect 7608 5159 7642 5160
rect 7608 5126 7642 5159
rect 9718 5159 9752 5160
rect 9718 5126 9752 5159
rect 7608 5052 7642 5086
rect 9718 5052 9752 5086
rect 7608 4979 7642 5012
rect 7608 4978 7642 4979
rect 9718 4979 9752 5012
rect 9718 4978 9752 4979
rect 7608 4906 7642 4938
rect 7608 4904 7642 4906
rect 9718 4906 9752 4938
rect 9718 4904 9752 4906
rect 7608 4832 7642 4864
rect 7608 4830 7642 4832
rect 9718 4832 9752 4864
rect 9718 4830 9752 4832
rect 7608 4758 7642 4790
rect 7608 4756 7642 4758
rect 9718 4758 9752 4790
rect 9718 4756 9752 4758
rect 7608 4684 7642 4715
rect 7608 4681 7642 4684
rect 9718 4684 9752 4715
rect 9718 4681 9752 4684
rect 7608 4610 7642 4640
rect 7608 4606 7642 4610
rect 9718 4610 9752 4640
rect 9718 4606 9752 4610
rect 9899 5372 9929 5399
rect 9929 5372 9933 5399
rect 9899 5331 9933 5334
rect 9899 5300 9929 5331
rect 9929 5300 9933 5331
rect 9899 5229 9929 5262
rect 9929 5229 9933 5262
rect 9899 5228 9933 5229
rect 9899 5161 9929 5190
rect 9929 5161 9933 5190
rect 9899 5156 9933 5161
rect 9899 5093 9929 5118
rect 9929 5093 9933 5118
rect 9899 5084 9933 5093
rect 9899 5025 9929 5046
rect 9929 5025 9933 5046
rect 9899 5012 9933 5025
rect 9899 4957 9929 4974
rect 9929 4957 9933 4974
rect 9899 4940 9933 4957
rect 9899 4889 9929 4902
rect 9929 4889 9933 4902
rect 9899 4868 9933 4889
rect 9899 4821 9929 4830
rect 9929 4821 9933 4830
rect 9899 4796 9933 4821
rect 9899 4753 9929 4758
rect 9929 4753 9933 4758
rect 9899 4724 9933 4753
rect 9899 4685 9929 4686
rect 9929 4685 9933 4686
rect 9899 4652 9933 4685
rect 7423 4583 7457 4591
rect 9899 4583 9933 4614
rect 7423 4557 7431 4583
rect 7431 4557 7457 4583
rect 8151 4549 8185 4583
rect 8223 4549 8257 4583
rect 8295 4549 8329 4583
rect 8367 4549 8401 4583
rect 8439 4549 8473 4583
rect 8511 4549 8545 4583
rect 8583 4549 8617 4583
rect 8655 4549 8689 4583
rect 8727 4549 8761 4583
rect 8800 4549 8834 4583
rect 8873 4549 8907 4583
rect 8946 4549 8980 4583
rect 9019 4549 9053 4583
rect 9092 4549 9126 4583
rect 9899 4580 9929 4583
rect 9929 4580 9933 4583
rect 7423 4515 7457 4519
rect 7423 4485 7431 4515
rect 7431 4485 7457 4515
rect 7423 4413 7431 4447
rect 7431 4413 7457 4447
rect 7423 4345 7431 4375
rect 7431 4345 7457 4375
rect 7423 4341 7457 4345
rect 7423 4277 7431 4303
rect 7431 4277 7457 4303
rect 7423 4269 7457 4277
rect 7423 4209 7431 4231
rect 7431 4209 7457 4231
rect 7423 4197 7457 4209
rect 7423 4141 7431 4159
rect 7431 4141 7457 4159
rect 7423 4125 7457 4141
rect 7423 4073 7431 4087
rect 7431 4073 7457 4087
rect 7423 4053 7457 4073
rect 7423 4005 7431 4015
rect 7431 4005 7457 4015
rect 7423 3981 7457 4005
rect 7423 3937 7431 3943
rect 7431 3937 7457 3943
rect 5557 3801 5591 3833
rect 5557 3799 5591 3801
rect 5557 3726 5591 3760
rect 7423 3909 7457 3937
rect 7423 3869 7431 3871
rect 7431 3869 7457 3871
rect 7423 3837 7457 3869
rect 7423 3767 7457 3799
rect 7423 3765 7431 3767
rect 7431 3765 7457 3767
rect 7608 4522 7642 4526
rect 7608 4492 7642 4522
rect 9718 4522 9752 4526
rect 9718 4492 9752 4522
rect 7608 4449 7642 4452
rect 7608 4418 7642 4449
rect 9718 4449 9752 4452
rect 9718 4418 9752 4449
rect 7608 4376 7642 4378
rect 7608 4344 7642 4376
rect 9718 4376 9752 4378
rect 9718 4344 9752 4376
rect 7608 4303 7642 4304
rect 7608 4270 7642 4303
rect 9718 4303 9752 4304
rect 9718 4270 9752 4303
rect 7608 4196 7642 4230
rect 9718 4196 9752 4230
rect 7608 4123 7642 4156
rect 7608 4122 7642 4123
rect 9718 4123 9752 4156
rect 9718 4122 9752 4123
rect 7608 4050 7642 4082
rect 7608 4048 7642 4050
rect 9718 4050 9752 4082
rect 9718 4048 9752 4050
rect 7608 3976 7642 4008
rect 7608 3974 7642 3976
rect 9718 3976 9752 4008
rect 9718 3974 9752 3976
rect 7608 3902 7642 3934
rect 7608 3900 7642 3902
rect 9718 3902 9752 3934
rect 9718 3900 9752 3902
rect 7608 3828 7642 3859
rect 7608 3825 7642 3828
rect 9718 3828 9752 3859
rect 9718 3825 9752 3828
rect 7608 3754 7642 3784
rect 7608 3750 7642 3754
rect 9718 3754 9752 3784
rect 9718 3750 9752 3754
rect 9899 4515 9933 4542
rect 9899 4508 9929 4515
rect 9929 4508 9933 4515
rect 9899 4447 9933 4470
rect 9899 4436 9929 4447
rect 9929 4436 9933 4447
rect 9899 4379 9933 4398
rect 9899 4364 9929 4379
rect 9929 4364 9933 4379
rect 9899 4311 9933 4326
rect 9899 4292 9929 4311
rect 9929 4292 9933 4311
rect 9899 4243 9933 4254
rect 9899 4220 9929 4243
rect 9929 4220 9933 4243
rect 9899 4175 9933 4182
rect 9899 4148 9929 4175
rect 9929 4148 9933 4175
rect 9899 4107 9933 4110
rect 9899 4076 9929 4107
rect 9929 4076 9933 4107
rect 9899 4005 9929 4038
rect 9929 4005 9933 4038
rect 9899 4004 9933 4005
rect 9899 3937 9929 3966
rect 9929 3937 9933 3966
rect 9899 3932 9933 3937
rect 9899 3869 9929 3894
rect 9929 3869 9933 3894
rect 9899 3860 9933 3869
rect 9899 3801 9929 3822
rect 9929 3801 9933 3822
rect 9899 3788 9933 3801
rect 7423 3699 7457 3727
rect 7423 3693 7431 3699
rect 7431 3693 7457 3699
rect 9899 3733 9929 3750
rect 9929 3733 9933 3750
rect 9899 3716 9933 3733
rect 3693 3631 3727 3655
rect 5557 3653 5591 3687
rect 3693 3621 3717 3631
rect 3717 3621 3727 3631
rect 3693 3563 3727 3583
rect 3693 3549 3717 3563
rect 3717 3549 3727 3563
rect 1185 3475 1219 3509
rect 2022 3493 2056 3527
rect 2095 3493 2129 3527
rect 2168 3493 2202 3527
rect 2241 3493 2275 3527
rect 2314 3493 2348 3527
rect 2387 3493 2421 3527
rect 2459 3493 2493 3527
rect 2531 3493 2565 3527
rect 2603 3493 2637 3527
rect 2675 3493 2709 3527
rect 2747 3493 2781 3527
rect 2819 3493 2853 3527
rect 2891 3493 2925 3527
rect 2963 3493 2997 3527
rect 3693 3495 3727 3511
rect 3693 3477 3717 3495
rect 3717 3477 3727 3495
rect 1185 3403 1219 3437
rect 1185 3331 1219 3365
rect 1185 3259 1219 3293
rect 1185 3187 1219 3221
rect 1185 3115 1219 3149
rect 1185 3043 1219 3077
rect 1185 2971 1219 3005
rect 1185 2899 1219 2933
rect 1185 2827 1219 2861
rect 1185 2755 1219 2789
rect 1185 2683 1219 2717
rect 1396 3436 1430 3440
rect 1396 3406 1430 3436
rect 3506 3436 3540 3440
rect 3506 3406 3540 3436
rect 1396 3363 1430 3366
rect 1396 3332 1430 3363
rect 3506 3363 3540 3366
rect 3506 3332 3540 3363
rect 1396 3290 1430 3292
rect 1396 3258 1430 3290
rect 3506 3290 3540 3292
rect 3506 3258 3540 3290
rect 1396 3217 1430 3218
rect 1396 3184 1430 3217
rect 3506 3217 3540 3218
rect 3506 3184 3540 3217
rect 1396 3110 1430 3144
rect 3506 3110 3540 3144
rect 1396 3037 1430 3070
rect 1396 3036 1430 3037
rect 3506 3037 3540 3070
rect 3506 3036 3540 3037
rect 1396 2964 1430 2996
rect 1396 2962 1430 2964
rect 3506 2964 3540 2996
rect 3506 2962 3540 2964
rect 1396 2890 1430 2922
rect 1396 2888 1430 2890
rect 3506 2890 3540 2922
rect 3506 2888 3540 2890
rect 1396 2816 1430 2848
rect 1396 2814 1430 2816
rect 3506 2816 3540 2848
rect 3506 2814 3540 2816
rect 1396 2742 1430 2773
rect 1396 2739 1430 2742
rect 3506 2742 3540 2773
rect 3506 2739 3540 2742
rect 1396 2668 1430 2698
rect 1396 2664 1430 2668
rect 3506 2668 3540 2698
rect 3506 2664 3540 2668
rect 3693 3427 3727 3439
rect 3693 3405 3717 3427
rect 3717 3405 3727 3427
rect 7423 3631 7457 3655
rect 7423 3621 7431 3631
rect 7431 3621 7457 3631
rect 7423 3563 7457 3583
rect 8151 3591 8761 3697
rect 8800 3663 8834 3697
rect 8873 3663 8907 3697
rect 8946 3663 8980 3697
rect 9019 3663 9053 3697
rect 9092 3663 9126 3697
rect 9899 3665 9929 3678
rect 9929 3665 9933 3678
rect 9899 3644 9933 3665
rect 8800 3591 8834 3625
rect 8873 3591 8907 3625
rect 8946 3591 8980 3625
rect 9019 3591 9053 3625
rect 9092 3591 9126 3625
rect 9899 3597 9929 3606
rect 9929 3597 9933 3606
rect 9899 3572 9933 3597
rect 7423 3549 7431 3563
rect 7431 3549 7457 3563
rect 9899 3529 9929 3534
rect 9929 3529 9933 3534
rect 7423 3495 7457 3511
rect 7423 3477 7431 3495
rect 7431 3477 7457 3495
rect 8151 3493 8185 3527
rect 8223 3493 8257 3527
rect 8295 3493 8329 3527
rect 8367 3493 8401 3527
rect 8439 3493 8473 3527
rect 8511 3493 8545 3527
rect 8583 3493 8617 3527
rect 8655 3493 8689 3527
rect 8727 3493 8761 3527
rect 8800 3493 8834 3527
rect 8873 3493 8907 3527
rect 8946 3493 8980 3527
rect 9019 3493 9053 3527
rect 9092 3493 9126 3527
rect 9899 3500 9933 3529
rect 9899 3461 9929 3462
rect 9929 3461 9933 3462
rect 7423 3427 7457 3439
rect 7423 3405 7431 3427
rect 7431 3405 7457 3427
rect 3693 3359 3727 3367
rect 3693 3333 3717 3359
rect 3717 3333 3727 3359
rect 3693 3291 3727 3295
rect 3693 3261 3717 3291
rect 3717 3261 3727 3291
rect 3693 3189 3717 3223
rect 3717 3189 3727 3223
rect 3693 3121 3717 3151
rect 3717 3121 3727 3151
rect 3693 3117 3727 3121
rect 3693 3053 3717 3079
rect 3717 3053 3727 3079
rect 3693 3045 3727 3053
rect 3693 2985 3717 3007
rect 3717 2985 3727 3007
rect 3693 2973 3727 2985
rect 3693 2917 3717 2935
rect 3717 2917 3727 2935
rect 3693 2901 3727 2917
rect 3693 2849 3717 2863
rect 3717 2849 3727 2863
rect 3693 2829 3727 2849
rect 3693 2781 3717 2791
rect 3717 2781 3727 2791
rect 3693 2757 3727 2781
rect 3693 2713 3717 2719
rect 3717 2713 3727 2719
rect 3693 2685 3727 2713
rect 1185 2611 1219 2645
rect 3693 2645 3717 2647
rect 3717 2645 3727 2647
rect 2022 2607 2056 2641
rect 2095 2607 2129 2641
rect 2168 2607 2202 2641
rect 2241 2607 2275 2641
rect 2314 2607 2348 2641
rect 1185 2543 1219 2573
rect 1185 2539 1219 2543
rect 1185 2475 1219 2501
rect 1185 2467 1219 2475
rect 2022 2535 2056 2569
rect 2095 2535 2129 2569
rect 2168 2535 2202 2569
rect 2241 2535 2275 2569
rect 2314 2535 2348 2569
rect 2022 2463 2056 2497
rect 2095 2463 2129 2497
rect 2168 2463 2202 2497
rect 2241 2463 2275 2497
rect 2314 2463 2348 2497
rect 2387 2463 2997 2641
rect 3693 2613 3727 2645
rect 3693 2543 3727 2575
rect 3693 2541 3717 2543
rect 3717 2541 3727 2543
rect 3693 2475 3727 2503
rect 3693 2469 3717 2475
rect 3717 2469 3727 2475
rect 1185 2407 1219 2429
rect 1185 2395 1219 2407
rect 1185 2339 1219 2357
rect 1185 2323 1219 2339
rect 1185 2271 1219 2285
rect 1185 2251 1219 2271
rect 1185 2203 1219 2213
rect 3693 2407 3727 2431
rect 3693 2397 3717 2407
rect 3717 2397 3727 2407
rect 3693 2339 3727 2359
rect 3693 2325 3717 2339
rect 3717 2325 3727 2339
rect 3693 2271 3727 2287
rect 3693 2253 3717 2271
rect 3717 2253 3727 2271
rect 3693 2203 3727 2215
rect 1185 2179 1219 2203
rect 3693 2181 3717 2203
rect 3717 2181 3727 2203
rect 5413 3098 5447 3132
rect 5493 3098 5527 3132
rect 5573 3098 5607 3132
rect 1185 2135 1219 2141
rect 1185 2107 1219 2135
rect 1185 2067 1219 2069
rect 1185 2035 1219 2067
rect 1185 1965 1219 1997
rect 1185 1963 1219 1965
rect 1185 1897 1219 1925
rect 1185 1891 1219 1897
rect 3773 2026 3807 2060
rect 3845 2026 3879 2060
rect 3773 1951 3807 1985
rect 3845 1951 3879 1985
rect 3773 1896 3807 1910
rect 3845 1896 3879 1910
rect 1185 1829 1219 1853
rect 1185 1819 1219 1829
rect 1185 1761 1219 1781
rect 1185 1747 1219 1761
rect 3773 1876 3777 1896
rect 3777 1876 3807 1896
rect 3845 1876 3879 1896
rect 3773 1827 3807 1835
rect 3845 1827 3879 1835
rect 3773 1801 3777 1827
rect 3777 1801 3807 1827
rect 3845 1801 3879 1827
rect 1185 1693 1219 1709
rect 1185 1675 1219 1693
rect 1185 1625 1219 1637
rect 1185 1603 1219 1625
rect 1185 1557 1219 1565
rect 1185 1531 1219 1557
rect 1185 1489 1219 1493
rect 1185 1459 1219 1489
rect 1185 1387 1219 1421
rect 1185 1319 1219 1349
rect 1185 1315 1219 1319
rect 1185 1251 1219 1277
rect 1185 1243 1219 1251
rect 1185 1183 1219 1205
rect 1185 1171 1219 1183
rect 1185 1115 1219 1133
rect 1185 1099 1219 1115
rect 1185 1047 1219 1061
rect 1185 1027 1219 1047
rect 1185 979 1219 989
rect 1185 955 1219 979
rect 1396 1743 1430 1747
rect 1396 1713 1430 1743
rect 3506 1743 3540 1747
rect 3506 1713 3540 1743
rect 1396 1670 1430 1673
rect 1396 1639 1430 1670
rect 3506 1670 3540 1673
rect 3506 1639 3540 1670
rect 1396 1597 1430 1599
rect 1396 1565 1430 1597
rect 3506 1597 3540 1599
rect 3506 1565 3540 1597
rect 1396 1524 1430 1525
rect 1396 1491 1430 1524
rect 3506 1524 3540 1525
rect 3506 1491 3540 1524
rect 1396 1417 1430 1451
rect 3506 1417 3540 1451
rect 1396 1344 1430 1377
rect 1396 1343 1430 1344
rect 3506 1344 3540 1377
rect 3506 1343 3540 1344
rect 1396 1271 1430 1303
rect 1396 1269 1430 1271
rect 3506 1271 3540 1303
rect 3506 1269 3540 1271
rect 1396 1197 1430 1229
rect 1396 1195 1430 1197
rect 3506 1197 3540 1229
rect 3506 1195 3540 1197
rect 1396 1123 1430 1155
rect 1396 1121 1430 1123
rect 3506 1123 3540 1155
rect 3506 1121 3540 1123
rect 1396 1049 1430 1080
rect 1396 1046 1430 1049
rect 3506 1049 3540 1080
rect 3506 1046 3540 1049
rect 1396 975 1430 1005
rect 1396 971 1430 975
rect 3506 975 3540 1005
rect 3506 971 3540 975
rect 3773 1758 3807 1760
rect 3845 1758 3879 1760
rect 3773 1726 3777 1758
rect 3777 1726 3807 1758
rect 3845 1726 3879 1758
rect 3773 1655 3777 1685
rect 3777 1655 3807 1685
rect 3845 1655 3879 1685
rect 3773 1651 3807 1655
rect 3845 1651 3879 1655
rect 3773 1586 3777 1610
rect 3777 1586 3807 1610
rect 3845 1586 3879 1610
rect 3773 1576 3807 1586
rect 3845 1576 3879 1586
rect 3773 1517 3777 1535
rect 3777 1517 3807 1535
rect 3845 1517 3879 1535
rect 3773 1501 3807 1517
rect 3845 1501 3879 1517
rect 3773 1448 3777 1460
rect 3777 1448 3807 1460
rect 3845 1448 3879 1460
rect 3773 1426 3807 1448
rect 3845 1426 3879 1448
rect 3773 1379 3777 1385
rect 3777 1379 3807 1385
rect 3845 1379 3879 1385
rect 3773 1351 3807 1379
rect 3845 1351 3879 1379
rect 3773 1276 3807 1310
rect 3845 1276 3879 1310
rect 3773 1204 3807 1235
rect 3845 1204 3879 1235
rect 3773 1201 3777 1204
rect 3777 1201 3807 1204
rect 3845 1201 3879 1204
rect 3773 1134 3807 1160
rect 3845 1134 3879 1160
rect 3773 1126 3777 1134
rect 3777 1126 3807 1134
rect 3845 1126 3879 1134
rect 5194 3020 5228 3036
rect 5194 3002 5228 3020
rect 5194 2952 5228 2964
rect 5194 2930 5228 2952
rect 5194 2858 5228 2892
rect 5194 2786 5228 2820
rect 5194 2730 5228 2748
rect 5194 2714 5228 2730
rect 5194 2662 5228 2676
rect 5194 2642 5228 2662
rect 5194 2570 5228 2604
rect 5194 2508 5228 2532
rect 5194 2498 5228 2508
rect 5194 2440 5228 2459
rect 5194 2425 5228 2440
rect 5194 2352 5228 2386
rect 5194 2279 5228 2313
rect 5194 2218 5228 2240
rect 5194 2206 5228 2218
rect 5194 2150 5228 2167
rect 5194 2133 5228 2150
rect 5194 2060 5228 2094
rect 5194 1996 5228 2021
rect 5194 1987 5228 1996
rect 5194 1928 5228 1948
rect 5194 1914 5228 1928
rect 5194 1841 5228 1875
rect 5194 1768 5228 1802
rect 5194 1706 5228 1729
rect 5194 1695 5228 1706
rect 5194 1638 5228 1656
rect 5194 1622 5228 1638
rect 5194 1549 5228 1583
rect 5194 1484 5228 1510
rect 5194 1476 5228 1484
rect 5194 1416 5228 1437
rect 5194 1403 5228 1416
rect 5194 1330 5228 1364
rect 5194 1257 5228 1291
rect 5194 1194 5228 1218
rect 5194 1184 5228 1194
rect 5194 1126 5228 1145
rect 5194 1111 5228 1126
rect 5712 3014 5746 3048
rect 5712 2946 5746 2976
rect 5712 2942 5746 2946
rect 5553 2862 5587 2896
rect 5627 2862 5661 2896
rect 5701 2862 5735 2896
rect 5413 2627 5447 2661
rect 5493 2627 5527 2661
rect 5573 2627 5607 2661
rect 5563 2520 5597 2544
rect 5563 2510 5597 2520
rect 5563 2451 5597 2471
rect 5563 2437 5597 2451
rect 5563 2382 5597 2398
rect 5563 2364 5597 2382
rect 5563 2313 5597 2325
rect 5563 2291 5597 2313
rect 5563 2244 5597 2252
rect 5563 2218 5597 2244
rect 5563 2175 5597 2179
rect 5563 2145 5597 2175
rect 5563 2072 5597 2106
rect 5563 2003 5597 2033
rect 5563 1999 5597 2003
rect 5563 1934 5597 1960
rect 5563 1926 5597 1934
rect 5563 1865 5597 1887
rect 5563 1853 5597 1865
rect 5563 1796 5597 1814
rect 5563 1780 5597 1796
rect 5563 1727 5597 1740
rect 5563 1706 5597 1727
rect 5563 1658 5597 1666
rect 5563 1632 5597 1658
rect 5563 1589 5597 1592
rect 5563 1558 5597 1589
rect 5563 1485 5597 1518
rect 5563 1484 5597 1485
rect 5563 1416 5597 1444
rect 5563 1410 5597 1416
rect 5563 1346 5597 1370
rect 5563 1336 5597 1346
rect 5563 1276 5597 1296
rect 5563 1262 5597 1276
rect 5563 1206 5597 1222
rect 5563 1188 5597 1206
rect 5563 1136 5597 1148
rect 3773 1064 3807 1085
rect 3845 1064 3879 1085
rect 3773 1051 3777 1064
rect 3777 1051 3807 1064
rect 3845 1051 3879 1064
rect 5563 1114 5597 1136
rect 7032 3020 7066 3036
rect 7032 3002 7066 3020
rect 7032 2952 7066 2964
rect 7032 2930 7066 2952
rect 7032 2858 7066 2892
rect 7032 2786 7066 2820
rect 7032 2730 7066 2748
rect 7032 2714 7066 2730
rect 7032 2662 7066 2676
rect 7032 2642 7066 2662
rect 7032 2570 7066 2604
rect 7032 2508 7066 2532
rect 7032 2498 7066 2508
rect 7032 2440 7066 2459
rect 7032 2425 7066 2440
rect 7032 2352 7066 2386
rect 7032 2279 7066 2313
rect 7032 2218 7066 2240
rect 7032 2206 7066 2218
rect 7032 2150 7066 2167
rect 7032 2133 7066 2150
rect 7032 2060 7066 2094
rect 7032 1996 7066 2021
rect 7032 1987 7066 1996
rect 7032 1928 7066 1948
rect 7032 1914 7066 1928
rect 7032 1841 7066 1875
rect 7032 1768 7066 1802
rect 7032 1706 7066 1729
rect 7032 1695 7066 1706
rect 7032 1638 7066 1656
rect 7032 1622 7066 1638
rect 7032 1549 7066 1583
rect 7032 1484 7066 1510
rect 7032 1476 7066 1484
rect 7032 1416 7066 1437
rect 7032 1403 7066 1416
rect 7032 1330 7066 1364
rect 7032 1257 7066 1291
rect 7032 1194 7066 1218
rect 7032 1184 7066 1194
rect 7032 1126 7066 1145
rect 7032 1111 7066 1126
rect 7423 3359 7457 3367
rect 7423 3333 7431 3359
rect 7431 3333 7457 3359
rect 7423 3291 7457 3295
rect 7423 3261 7431 3291
rect 7431 3261 7457 3291
rect 7423 3189 7431 3223
rect 7431 3189 7457 3223
rect 7423 3121 7431 3151
rect 7431 3121 7457 3151
rect 7423 3117 7457 3121
rect 7423 3053 7431 3079
rect 7431 3053 7457 3079
rect 7423 3045 7457 3053
rect 7423 2985 7431 3007
rect 7431 2985 7457 3007
rect 7423 2973 7457 2985
rect 7423 2917 7431 2935
rect 7431 2917 7457 2935
rect 7423 2901 7457 2917
rect 7423 2849 7431 2863
rect 7431 2849 7457 2863
rect 7423 2829 7457 2849
rect 7423 2781 7431 2791
rect 7431 2781 7457 2791
rect 7423 2757 7457 2781
rect 7423 2713 7431 2719
rect 7431 2713 7457 2719
rect 7423 2685 7457 2713
rect 7608 3436 7642 3440
rect 7608 3406 7642 3436
rect 9718 3436 9752 3440
rect 9718 3406 9752 3436
rect 7608 3363 7642 3366
rect 7608 3332 7642 3363
rect 9718 3363 9752 3366
rect 9718 3332 9752 3363
rect 7608 3290 7642 3292
rect 7608 3258 7642 3290
rect 9718 3290 9752 3292
rect 9718 3258 9752 3290
rect 7608 3217 7642 3218
rect 7608 3184 7642 3217
rect 9718 3217 9752 3218
rect 9718 3184 9752 3217
rect 7608 3110 7642 3144
rect 9718 3110 9752 3144
rect 7608 3037 7642 3070
rect 7608 3036 7642 3037
rect 9718 3037 9752 3070
rect 9718 3036 9752 3037
rect 7608 2964 7642 2996
rect 7608 2962 7642 2964
rect 9718 2964 9752 2996
rect 9718 2962 9752 2964
rect 7608 2890 7642 2922
rect 7608 2888 7642 2890
rect 9718 2890 9752 2922
rect 9718 2888 9752 2890
rect 7608 2816 7642 2848
rect 7608 2814 7642 2816
rect 9718 2816 9752 2848
rect 9718 2814 9752 2816
rect 7608 2742 7642 2773
rect 7608 2739 7642 2742
rect 9718 2742 9752 2773
rect 9718 2739 9752 2742
rect 7608 2668 7642 2698
rect 7608 2664 7642 2668
rect 9718 2668 9752 2698
rect 9718 2664 9752 2668
rect 9899 3428 9933 3461
rect 9899 3359 9933 3390
rect 9899 3356 9929 3359
rect 9929 3356 9933 3359
rect 9899 3291 9933 3318
rect 9899 3284 9929 3291
rect 9929 3284 9933 3291
rect 9899 3223 9933 3246
rect 9899 3212 9929 3223
rect 9929 3212 9933 3223
rect 9899 3155 9933 3174
rect 9899 3140 9929 3155
rect 9929 3140 9933 3155
rect 9899 3087 9933 3102
rect 9899 3068 9929 3087
rect 9929 3068 9933 3087
rect 9899 3019 9933 3030
rect 9899 2996 9929 3019
rect 9929 2996 9933 3019
rect 9899 2951 9933 2958
rect 9899 2924 9929 2951
rect 9929 2924 9933 2951
rect 9899 2883 9933 2886
rect 9899 2852 9929 2883
rect 9929 2852 9933 2883
rect 9899 2781 9929 2814
rect 9929 2781 9933 2814
rect 9899 2780 9933 2781
rect 9899 2713 9929 2742
rect 9929 2713 9933 2742
rect 9899 2708 9933 2713
rect 7423 2645 7431 2647
rect 7431 2645 7457 2647
rect 7423 2613 7457 2645
rect 9899 2645 9929 2670
rect 9929 2645 9933 2670
rect 7423 2543 7457 2575
rect 7423 2541 7431 2543
rect 7431 2541 7457 2543
rect 7423 2475 7457 2503
rect 7423 2469 7431 2475
rect 7431 2469 7457 2475
rect 8151 2463 8761 2641
rect 8800 2607 8834 2641
rect 8873 2607 8907 2641
rect 8946 2607 8980 2641
rect 9019 2607 9053 2641
rect 9092 2607 9126 2641
rect 9899 2636 9933 2645
rect 9899 2577 9929 2598
rect 9929 2577 9933 2598
rect 8800 2535 8834 2569
rect 8873 2535 8907 2569
rect 8946 2535 8980 2569
rect 9019 2535 9053 2569
rect 9092 2535 9126 2569
rect 9899 2564 9933 2577
rect 8800 2463 8834 2497
rect 8873 2463 8907 2497
rect 8946 2463 8980 2497
rect 9019 2463 9053 2497
rect 9092 2463 9126 2497
rect 9899 2509 9929 2526
rect 9929 2509 9933 2526
rect 9899 2492 9933 2509
rect 7423 2407 7457 2431
rect 7423 2397 7431 2407
rect 7431 2397 7457 2407
rect 7423 2339 7457 2359
rect 7423 2325 7431 2339
rect 7431 2325 7457 2339
rect 7423 2271 7457 2287
rect 7423 2253 7431 2271
rect 7431 2253 7457 2271
rect 7423 2203 7457 2215
rect 9899 2441 9929 2454
rect 9929 2441 9933 2454
rect 9899 2420 9933 2441
rect 9899 2373 9929 2382
rect 9929 2373 9933 2382
rect 9899 2348 9933 2373
rect 9899 2305 9929 2310
rect 9929 2305 9933 2310
rect 9899 2276 9933 2305
rect 9899 2237 9929 2238
rect 9929 2237 9933 2238
rect 9899 2204 9933 2237
rect 7423 2181 7431 2203
rect 7431 2181 7457 2203
rect 9899 2135 9933 2166
rect 9899 2132 9929 2135
rect 9929 2132 9933 2135
rect 9899 2067 9933 2094
rect 9899 2060 9929 2067
rect 9929 2060 9933 2067
rect 7271 2026 7305 2060
rect 7343 2026 7377 2060
rect 7271 1951 7305 1985
rect 7343 1951 7377 1985
rect 9899 1999 9933 2022
rect 9899 1988 9929 1999
rect 9929 1988 9933 1999
rect 9899 1931 9933 1950
rect 7271 1896 7305 1910
rect 7343 1896 7377 1910
rect 7271 1876 7275 1896
rect 7275 1876 7305 1896
rect 7343 1876 7377 1896
rect 9899 1916 9929 1931
rect 9929 1916 9933 1931
rect 7271 1827 7305 1835
rect 7343 1827 7377 1835
rect 7271 1801 7275 1827
rect 7275 1801 7305 1827
rect 7343 1801 7377 1827
rect 7271 1758 7305 1760
rect 7343 1758 7377 1760
rect 9899 1863 9933 1878
rect 9899 1844 9929 1863
rect 9929 1844 9933 1863
rect 9899 1795 9933 1806
rect 9899 1772 9929 1795
rect 9929 1772 9933 1795
rect 7271 1726 7275 1758
rect 7275 1726 7305 1758
rect 7343 1726 7377 1758
rect 7271 1655 7275 1685
rect 7275 1655 7305 1685
rect 7343 1655 7377 1685
rect 7271 1651 7305 1655
rect 7343 1651 7377 1655
rect 7271 1586 7275 1610
rect 7275 1586 7305 1610
rect 7343 1586 7377 1610
rect 7271 1576 7305 1586
rect 7343 1576 7377 1586
rect 7271 1517 7275 1535
rect 7275 1517 7305 1535
rect 7343 1517 7377 1535
rect 7271 1501 7305 1517
rect 7343 1501 7377 1517
rect 7271 1448 7275 1460
rect 7275 1448 7305 1460
rect 7343 1448 7377 1460
rect 7271 1426 7305 1448
rect 7343 1426 7377 1448
rect 7271 1379 7275 1385
rect 7275 1379 7305 1385
rect 7343 1379 7377 1385
rect 7271 1351 7305 1379
rect 7343 1351 7377 1379
rect 7271 1276 7305 1310
rect 7343 1276 7377 1310
rect 7271 1204 7305 1235
rect 7343 1204 7377 1235
rect 7271 1201 7275 1204
rect 7275 1201 7305 1204
rect 7343 1201 7377 1204
rect 7271 1134 7305 1160
rect 7343 1134 7377 1160
rect 5563 1066 5597 1074
rect 5563 1040 5597 1066
rect 3773 994 3807 1010
rect 3845 994 3879 1010
rect 1185 911 1219 917
rect 1185 883 1219 911
rect 3773 976 3777 994
rect 3777 976 3807 994
rect 3845 976 3879 994
rect 3773 924 3807 935
rect 3845 924 3879 935
rect 3773 901 3777 924
rect 3777 901 3807 924
rect 3845 901 3879 924
rect 1185 843 1219 845
rect 1185 811 1219 843
rect 3506 829 3540 863
rect 1624 792 1633 826
rect 1633 792 1658 826
rect 1716 792 1733 826
rect 1733 792 1750 826
rect 7271 1126 7275 1134
rect 7275 1126 7305 1134
rect 7343 1126 7377 1134
rect 7271 1064 7305 1085
rect 7343 1064 7377 1085
rect 7271 1051 7275 1064
rect 7275 1051 7305 1064
rect 7343 1051 7377 1064
rect 5563 996 5597 1000
rect 5563 966 5597 996
rect 5563 892 5597 926
rect 3773 854 3807 860
rect 3845 854 3879 860
rect 3773 826 3777 854
rect 3777 826 3807 854
rect 3845 826 3879 854
rect 1185 741 1219 773
rect 2060 766 2094 800
rect 3175 766 3178 800
rect 3178 766 3209 800
rect 3247 766 3280 800
rect 3280 766 3281 800
rect 3506 766 3526 791
rect 3526 766 3540 791
rect 3773 784 3807 785
rect 3845 784 3879 785
rect 1185 739 1219 741
rect 1185 673 1219 701
rect 1185 667 1219 673
rect 1185 605 1219 629
rect 1185 595 1219 605
rect 1185 537 1219 557
rect 1538 692 1572 726
rect 1538 620 1572 654
rect 1538 548 1572 582
rect 1794 674 1828 708
rect 1794 602 1828 636
rect 1185 523 1219 537
rect 1794 530 1828 564
rect 1904 674 1938 708
rect 1904 602 1938 636
rect 3506 757 3540 766
rect 3773 751 3777 784
rect 3777 751 3807 784
rect 3845 751 3879 784
rect 2060 694 2094 728
rect 2060 622 2094 656
rect 2316 674 2350 708
rect 1904 530 1938 564
rect 2316 602 2350 636
rect 2316 530 2350 564
rect 2572 696 2606 730
rect 2572 624 2606 658
rect 2572 552 2606 586
rect 2828 674 2862 708
rect 2828 602 2862 636
rect 2828 530 2862 564
rect 3084 696 3118 730
rect 7271 994 7305 1010
rect 7343 994 7377 1010
rect 7271 976 7275 994
rect 7275 976 7305 994
rect 7343 976 7377 994
rect 7608 1743 7642 1747
rect 7608 1713 7642 1743
rect 9718 1743 9752 1747
rect 9718 1713 9752 1743
rect 7608 1670 7642 1673
rect 7608 1639 7642 1670
rect 9718 1670 9752 1673
rect 9718 1639 9752 1670
rect 7608 1597 7642 1599
rect 7608 1565 7642 1597
rect 9718 1597 9752 1599
rect 9718 1565 9752 1597
rect 7608 1524 7642 1525
rect 7608 1491 7642 1524
rect 9718 1524 9752 1525
rect 9718 1491 9752 1524
rect 7608 1417 7642 1451
rect 9718 1417 9752 1451
rect 7608 1344 7642 1377
rect 7608 1343 7642 1344
rect 9718 1344 9752 1377
rect 9718 1343 9752 1344
rect 7608 1271 7642 1303
rect 7608 1269 7642 1271
rect 9718 1271 9752 1303
rect 9718 1269 9752 1271
rect 7608 1197 7642 1229
rect 7608 1195 7642 1197
rect 9718 1197 9752 1229
rect 9718 1195 9752 1197
rect 7608 1123 7642 1155
rect 7608 1121 7642 1123
rect 9718 1123 9752 1155
rect 9718 1121 9752 1123
rect 7608 1049 7642 1080
rect 7608 1046 7642 1049
rect 9718 1049 9752 1080
rect 9718 1046 9752 1049
rect 7608 975 7642 1005
rect 7608 971 7642 975
rect 9718 975 9752 1005
rect 9718 971 9752 975
rect 9899 1727 9933 1734
rect 9899 1700 9929 1727
rect 9929 1700 9933 1727
rect 9899 1659 9933 1662
rect 9899 1628 9929 1659
rect 9929 1628 9933 1659
rect 9899 1557 9929 1590
rect 9929 1557 9933 1590
rect 9899 1556 9933 1557
rect 9899 1489 9929 1518
rect 9929 1489 9933 1518
rect 9899 1484 9933 1489
rect 9899 1421 9929 1446
rect 9929 1421 9933 1446
rect 9899 1412 9933 1421
rect 9899 1353 9929 1374
rect 9929 1353 9933 1374
rect 9899 1340 9933 1353
rect 9899 1285 9929 1302
rect 9929 1285 9933 1302
rect 9899 1268 9933 1285
rect 9899 1217 9929 1230
rect 9929 1217 9933 1230
rect 9899 1196 9933 1217
rect 9899 1149 9929 1158
rect 9929 1149 9933 1158
rect 9899 1124 9933 1149
rect 9899 1081 9929 1086
rect 9929 1081 9933 1086
rect 9899 1052 9933 1081
rect 9899 1013 9929 1014
rect 9929 1013 9933 1014
rect 9899 980 9933 1013
rect 7271 924 7305 935
rect 7343 924 7377 935
rect 7271 901 7275 924
rect 7275 901 7305 924
rect 7343 901 7377 924
rect 5563 822 5597 852
rect 5563 818 5597 822
rect 5563 752 5597 778
rect 5563 744 5597 752
rect 3084 624 3118 658
rect 3506 671 3540 705
rect 3506 599 3540 633
rect 3773 680 3777 710
rect 3777 680 3807 710
rect 3845 680 3879 710
rect 3773 676 3807 680
rect 3845 676 3879 680
rect 3773 610 3777 634
rect 3777 610 3807 634
rect 3845 610 3879 634
rect 3773 600 3807 610
rect 3845 600 3879 610
rect 3084 552 3118 586
rect 3268 519 3302 553
rect 3340 519 3374 553
rect 3773 540 3777 558
rect 3777 540 3807 558
rect 3845 540 3879 558
rect 3773 524 3807 540
rect 3845 524 3879 540
rect 5192 678 5226 692
rect 5192 658 5226 678
rect 5192 576 5226 600
rect 5192 566 5226 576
rect 9899 911 9933 942
rect 9899 908 9929 911
rect 9929 908 9933 911
rect 7271 854 7305 860
rect 7343 854 7377 860
rect 7271 826 7275 854
rect 7275 826 7305 854
rect 7343 826 7377 854
rect 7271 784 7305 785
rect 7343 784 7377 785
rect 7271 751 7275 784
rect 7275 751 7305 784
rect 7343 751 7377 784
rect 7587 826 7621 860
rect 9899 843 9933 870
rect 9899 836 9929 843
rect 9929 836 9933 843
rect 7587 754 7621 788
rect 9054 766 9088 800
rect 9899 775 9933 798
rect 5563 682 5597 704
rect 5563 670 5597 682
rect 5563 612 5597 630
rect 5563 596 5597 612
rect 5563 542 5597 556
rect 1185 469 1219 485
rect 1185 451 1219 469
rect 3773 470 3777 482
rect 3777 470 3807 482
rect 3845 470 3879 482
rect 3773 448 3807 470
rect 3845 448 3879 470
rect 5563 522 5597 542
rect 7032 678 7066 692
rect 7032 658 7066 678
rect 7032 610 7066 620
rect 7032 586 7066 610
rect 7032 542 7066 547
rect 7032 513 7066 542
rect 7271 680 7275 710
rect 7275 680 7305 710
rect 7343 680 7377 710
rect 7271 676 7305 680
rect 7343 676 7377 680
rect 7271 610 7275 634
rect 7275 610 7305 634
rect 7343 610 7377 634
rect 7271 600 7305 610
rect 7343 600 7377 610
rect 7618 674 7652 708
rect 7618 602 7652 636
rect 8030 696 8064 730
rect 8030 624 8064 658
rect 7271 540 7275 558
rect 7275 540 7305 558
rect 7343 540 7377 558
rect 7774 544 7808 578
rect 7846 544 7880 578
rect 8030 552 8064 586
rect 8286 674 8320 708
rect 8286 602 8320 636
rect 7271 524 7305 540
rect 7343 524 7377 540
rect 8286 530 8320 564
rect 8542 696 8576 730
rect 8542 624 8576 658
rect 8542 552 8576 586
rect 8798 674 8832 708
rect 8798 602 8832 636
rect 9054 694 9088 728
rect 9054 622 9088 656
rect 9210 674 9244 708
rect 8798 530 8832 564
rect 9210 602 9244 636
rect 9210 530 9244 564
rect 9899 764 9929 775
rect 9929 764 9933 775
rect 9899 707 9933 726
rect 9899 692 9929 707
rect 9929 692 9933 707
rect 9899 639 9933 654
rect 9899 620 9929 639
rect 9929 620 9933 639
rect 9899 571 9933 582
rect 9899 548 9929 571
rect 9929 548 9933 571
rect 5563 472 5597 482
rect 5563 448 5597 472
rect 7271 470 7275 482
rect 7275 470 7305 482
rect 7343 470 7377 482
rect 9899 503 9933 510
rect 7271 448 7305 470
rect 7343 448 7377 470
rect 9899 476 9929 503
rect 9929 476 9933 503
rect 1185 401 1219 413
rect 1185 379 1219 401
rect 1185 333 1219 341
rect 1185 307 1219 333
rect 1185 265 1219 269
rect 1185 235 1219 265
rect 10205 7671 10239 7699
rect 10277 7671 10283 7705
rect 10283 7671 10311 7705
rect 10349 7671 10351 7705
rect 10351 7671 10383 7705
rect 10421 7671 10453 7705
rect 10453 7671 10455 7705
rect 10493 7671 10521 7705
rect 10521 7671 10527 7705
rect 10565 7671 10589 7705
rect 10589 7671 10599 7705
rect 10637 7671 10657 7705
rect 10657 7671 10671 7705
rect 10709 7671 10725 7705
rect 10725 7671 10743 7705
rect 10782 7671 10793 7705
rect 10793 7671 10816 7705
rect 10855 7671 10861 7705
rect 10861 7671 10889 7705
rect 10928 7671 10929 7705
rect 10929 7671 10962 7705
rect 11001 7671 11031 7705
rect 11031 7671 11035 7705
rect 11074 7671 11099 7705
rect 11099 7671 11108 7705
rect 11147 7671 11167 7705
rect 11167 7671 11181 7705
rect 11220 7671 11235 7705
rect 11235 7671 11254 7705
rect 11293 7671 11303 7705
rect 11303 7671 11327 7705
rect 11366 7671 11371 7705
rect 11371 7671 11400 7705
rect 11439 7671 11473 7705
rect 11512 7671 11541 7705
rect 11541 7671 11546 7705
rect 11585 7671 11609 7705
rect 11609 7671 11619 7705
rect 11658 7671 11677 7705
rect 11677 7671 11692 7705
rect 11731 7671 11745 7705
rect 11745 7671 11765 7705
rect 11804 7671 11813 7705
rect 11813 7671 11838 7705
rect 11877 7671 11881 7705
rect 11881 7671 11911 7705
rect 11950 7671 11983 7705
rect 11983 7671 11984 7705
rect 12023 7671 12051 7705
rect 12051 7671 12057 7705
rect 12096 7671 12119 7705
rect 12119 7671 12130 7705
rect 12169 7671 12187 7705
rect 12187 7671 12203 7705
rect 12242 7671 12255 7705
rect 12255 7671 12276 7705
rect 12315 7671 12323 7705
rect 12323 7671 12349 7705
rect 12388 7671 12391 7705
rect 12391 7671 12422 7705
rect 12461 7671 12493 7705
rect 12493 7671 12495 7705
rect 12534 7671 12561 7705
rect 12561 7671 12568 7705
rect 12607 7671 12629 7705
rect 12629 7671 12641 7705
rect 12680 7671 12697 7705
rect 12697 7671 12714 7705
rect 12753 7671 12765 7705
rect 12765 7671 12787 7705
rect 10205 7665 10212 7671
rect 10212 7665 10239 7671
rect 10205 7603 10239 7627
rect 10205 7593 10212 7603
rect 10212 7593 10239 7603
rect 10205 7535 10239 7555
rect 10205 7521 10212 7535
rect 10212 7521 10239 7535
rect 10205 7467 10239 7483
rect 10205 7449 10212 7467
rect 10212 7449 10239 7467
rect 10205 7399 10239 7411
rect 10205 7377 10212 7399
rect 10212 7377 10239 7399
rect 10205 7331 10239 7339
rect 10205 7305 10212 7331
rect 10212 7305 10239 7331
rect 10205 7263 10239 7267
rect 10205 7233 10212 7263
rect 10212 7233 10239 7263
rect 10205 7161 10212 7195
rect 10212 7161 10239 7195
rect 10205 7093 10212 7123
rect 10212 7093 10239 7123
rect 10205 7089 10239 7093
rect 10205 7025 10212 7051
rect 10212 7025 10239 7051
rect 10205 7017 10239 7025
rect 10205 6957 10212 6979
rect 10212 6957 10239 6979
rect 10205 6945 10239 6957
rect 10205 6889 10212 6907
rect 10212 6889 10239 6907
rect 10205 6873 10239 6889
rect 10205 6821 10212 6835
rect 10212 6821 10239 6835
rect 10205 6801 10239 6821
rect 10205 6753 10212 6763
rect 10212 6753 10239 6763
rect 10205 6729 10239 6753
rect 10205 6685 10212 6691
rect 10212 6685 10239 6691
rect 10205 6657 10239 6685
rect 10205 6617 10212 6619
rect 10212 6617 10239 6619
rect 10205 6585 10239 6617
rect 10205 6515 10239 6547
rect 10205 6513 10212 6515
rect 10212 6513 10239 6515
rect 10205 6447 10239 6475
rect 10205 6441 10212 6447
rect 10212 6441 10239 6447
rect 10205 6379 10239 6403
rect 10205 6369 10212 6379
rect 10212 6369 10239 6379
rect 10205 6311 10239 6331
rect 10205 6297 10212 6311
rect 10212 6297 10239 6311
rect 10205 6243 10239 6259
rect 10205 6225 10212 6243
rect 10212 6225 10239 6243
rect 10205 6175 10239 6187
rect 10205 6153 10212 6175
rect 10212 6153 10239 6175
rect 10205 6107 10239 6115
rect 10205 6081 10212 6107
rect 10212 6081 10239 6107
rect 10205 6039 10239 6043
rect 10205 6009 10212 6039
rect 10212 6009 10239 6039
rect 10205 5937 10212 5971
rect 10212 5937 10239 5971
rect 10205 5869 10212 5899
rect 10212 5869 10239 5899
rect 10205 5865 10239 5869
rect 10205 5801 10212 5827
rect 10212 5801 10239 5827
rect 10205 5793 10239 5801
rect 10205 5733 10212 5755
rect 10212 5733 10239 5755
rect 10205 5721 10239 5733
rect 10205 5665 10212 5683
rect 10212 5665 10239 5683
rect 10205 5649 10239 5665
rect 10205 5597 10212 5611
rect 10212 5597 10239 5611
rect 10205 5577 10239 5597
rect 10205 5529 10212 5539
rect 10212 5529 10239 5539
rect 10205 5505 10239 5529
rect 10205 5461 10212 5467
rect 10212 5461 10239 5467
rect 10205 5433 10239 5461
rect 10205 5393 10212 5395
rect 10212 5393 10239 5395
rect 10205 5361 10239 5393
rect 10205 5291 10239 5323
rect 10205 5289 10212 5291
rect 10212 5289 10239 5291
rect 10205 5223 10239 5251
rect 10205 5217 10212 5223
rect 10212 5217 10239 5223
rect 10205 5155 10239 5179
rect 10205 5145 10212 5155
rect 10212 5145 10239 5155
rect 10205 5087 10239 5107
rect 10205 5073 10212 5087
rect 10212 5073 10239 5087
rect 10205 5019 10239 5035
rect 10205 5001 10212 5019
rect 10212 5001 10239 5019
rect 10205 4951 10239 4963
rect 10205 4929 10212 4951
rect 10212 4929 10239 4951
rect 10205 4883 10239 4891
rect 10205 4857 10212 4883
rect 10212 4857 10239 4883
rect 10205 4815 10239 4819
rect 10205 4785 10212 4815
rect 10212 4785 10239 4815
rect 10205 4713 10212 4747
rect 10212 4713 10239 4747
rect 10205 4645 10212 4675
rect 10212 4645 10239 4675
rect 10205 4641 10239 4645
rect 10205 4577 10212 4603
rect 10212 4577 10239 4603
rect 10205 4569 10239 4577
rect 10205 4509 10212 4531
rect 10212 4509 10239 4531
rect 10205 4497 10239 4509
rect 10205 4441 10212 4459
rect 10212 4441 10239 4459
rect 10205 4425 10239 4441
rect 10205 4373 10212 4387
rect 10212 4373 10239 4387
rect 10205 4353 10239 4373
rect 10205 4305 10212 4315
rect 10212 4305 10239 4315
rect 10205 4281 10239 4305
rect 10205 4237 10212 4243
rect 10212 4237 10239 4243
rect 10205 4209 10239 4237
rect 10205 4169 10212 4171
rect 10212 4169 10239 4171
rect 10205 4137 10239 4169
rect 10205 4067 10239 4099
rect 10205 4065 10212 4067
rect 10212 4065 10239 4067
rect 10205 3999 10239 4027
rect 10205 3993 10212 3999
rect 10212 3993 10239 3999
rect 10205 3931 10239 3955
rect 10205 3921 10212 3931
rect 10212 3921 10239 3931
rect 10205 3863 10239 3883
rect 10205 3849 10212 3863
rect 10212 3849 10239 3863
rect 10205 3795 10239 3811
rect 10205 3777 10212 3795
rect 10212 3777 10239 3795
rect 10205 3727 10239 3739
rect 10205 3705 10212 3727
rect 10212 3705 10239 3727
rect 10205 3659 10239 3667
rect 10205 3633 10212 3659
rect 10212 3633 10239 3659
rect 10205 3591 10239 3595
rect 10205 3561 10212 3591
rect 10212 3561 10239 3591
rect 10205 3489 10212 3523
rect 10212 3489 10239 3523
rect 10205 3421 10212 3451
rect 10212 3421 10239 3451
rect 10205 3417 10239 3421
rect 10205 3353 10212 3379
rect 10212 3353 10239 3379
rect 10205 3345 10239 3353
rect 10205 3285 10212 3307
rect 10212 3285 10239 3307
rect 10205 3273 10239 3285
rect 10205 3217 10212 3235
rect 10212 3217 10239 3235
rect 10205 3201 10239 3217
rect 10205 3149 10212 3163
rect 10212 3149 10239 3163
rect 10205 3129 10239 3149
rect 10205 3081 10212 3091
rect 10212 3081 10239 3091
rect 10205 3057 10239 3081
rect 10205 3013 10212 3019
rect 10212 3013 10239 3019
rect 10205 2985 10239 3013
rect 10205 2945 10212 2947
rect 10212 2945 10239 2947
rect 10205 2913 10239 2945
rect 10205 2843 10239 2875
rect 10205 2841 10212 2843
rect 10212 2841 10239 2843
rect 10205 2775 10239 2803
rect 10205 2769 10212 2775
rect 10212 2769 10239 2775
rect 10205 2707 10239 2731
rect 10205 2697 10212 2707
rect 10212 2697 10239 2707
rect 10205 2639 10239 2659
rect 10205 2625 10212 2639
rect 10212 2625 10239 2639
rect 10205 2571 10239 2587
rect 10205 2553 10212 2571
rect 10212 2553 10239 2571
rect 10205 2503 10239 2515
rect 10205 2481 10212 2503
rect 10212 2481 10239 2503
rect 10205 2435 10239 2443
rect 10205 2409 10212 2435
rect 10212 2409 10239 2435
rect 10205 2367 10239 2371
rect 10205 2337 10212 2367
rect 10212 2337 10239 2367
rect 10205 2265 10212 2299
rect 10212 2265 10239 2299
rect 10205 2197 10212 2227
rect 10212 2197 10239 2227
rect 10205 2193 10239 2197
rect 10205 2129 10212 2155
rect 10212 2129 10239 2155
rect 10205 2121 10239 2129
rect 10205 2061 10212 2083
rect 10212 2061 10239 2083
rect 10205 2049 10239 2061
rect 10205 1993 10212 2011
rect 10212 1993 10239 2011
rect 10205 1977 10239 1993
rect 10205 1925 10212 1939
rect 10212 1925 10239 1939
rect 10205 1905 10239 1925
rect 10205 1857 10212 1867
rect 10212 1857 10239 1867
rect 10205 1833 10239 1857
rect 10205 1789 10212 1795
rect 10212 1789 10239 1795
rect 10205 1761 10239 1789
rect 10205 1721 10212 1723
rect 10212 1721 10239 1723
rect 10205 1689 10239 1721
rect 10205 1619 10239 1651
rect 10205 1617 10212 1619
rect 10212 1617 10239 1619
rect 10205 1551 10239 1579
rect 10205 1545 10212 1551
rect 10212 1545 10239 1551
rect 10205 1483 10239 1507
rect 10205 1473 10212 1483
rect 10212 1473 10239 1483
rect 10205 1415 10239 1435
rect 10205 1401 10212 1415
rect 10212 1401 10239 1415
rect 10205 1347 10239 1363
rect 10205 1329 10212 1347
rect 10212 1329 10239 1347
rect 10205 1279 10239 1291
rect 10205 1257 10212 1279
rect 10212 1257 10239 1279
rect 10205 1211 10239 1219
rect 10205 1185 10212 1211
rect 10212 1185 10239 1211
rect 10205 1143 10239 1147
rect 10205 1113 10212 1143
rect 10212 1113 10239 1143
rect 10205 1041 10212 1075
rect 10212 1041 10239 1075
rect 10205 973 10212 1003
rect 10212 973 10239 1003
rect 10205 969 10239 973
rect 10205 905 10212 930
rect 10212 905 10239 930
rect 10205 896 10239 905
rect 10205 837 10212 857
rect 10212 837 10239 857
rect 10205 823 10239 837
rect 10205 769 10212 784
rect 10212 769 10239 784
rect 10205 750 10239 769
rect 10205 701 10212 711
rect 10212 701 10239 711
rect 10205 677 10239 701
rect 10205 633 10212 638
rect 10212 633 10239 638
rect 10205 604 10239 633
rect 10205 531 10239 565
rect 10205 458 10239 492
rect 13069 7156 13103 7160
rect 13069 7126 13103 7156
rect 13069 7054 13103 7088
rect 13069 6986 13103 7016
rect 13069 6982 13103 6986
rect 13069 6918 13103 6944
rect 13069 6910 13103 6918
rect 13069 6850 13103 6872
rect 13069 6838 13103 6850
rect 13069 6782 13103 6800
rect 13069 6766 13103 6782
rect 13069 6714 13103 6728
rect 13069 6694 13103 6714
rect 13069 6646 13103 6656
rect 13069 6622 13103 6646
rect 13069 6578 13103 6584
rect 13069 6550 13103 6578
rect 13069 6510 13103 6512
rect 13069 6478 13103 6510
rect 13069 6408 13103 6440
rect 13069 6406 13103 6408
rect 13069 6340 13103 6368
rect 13069 6334 13103 6340
rect 13069 6272 13103 6296
rect 13069 6262 13103 6272
rect 13069 6204 13103 6224
rect 13069 6190 13103 6204
rect 13069 6136 13103 6152
rect 13069 6118 13103 6136
rect 13069 6068 13103 6080
rect 13069 6046 13103 6068
rect 13069 6000 13103 6008
rect 13069 5974 13103 6000
rect 13069 5932 13103 5936
rect 13069 5902 13103 5932
rect 13069 5830 13103 5864
rect 13069 5762 13103 5792
rect 13069 5758 13103 5762
rect 13069 5694 13103 5720
rect 13069 5686 13103 5694
rect 13069 5626 13103 5648
rect 13069 5614 13103 5626
rect 13069 5558 13103 5576
rect 13069 5542 13103 5558
rect 13069 5490 13103 5504
rect 13069 5470 13103 5490
rect 13069 5422 13103 5432
rect 13069 5398 13103 5422
rect 13069 5354 13103 5360
rect 13069 5326 13103 5354
rect 13069 5286 13103 5288
rect 13069 5254 13103 5286
rect 13069 5184 13103 5216
rect 13069 5182 13103 5184
rect 13069 5116 13103 5144
rect 13069 5110 13103 5116
rect 13069 5048 13103 5072
rect 13069 5038 13103 5048
rect 13069 4980 13103 5000
rect 13069 4966 13103 4980
rect 13069 4912 13103 4928
rect 13069 4894 13103 4912
rect 13069 4844 13103 4856
rect 13069 4822 13103 4844
rect 13069 4776 13103 4784
rect 13069 4750 13103 4776
rect 13069 4708 13103 4712
rect 13069 4678 13103 4708
rect 13069 4606 13103 4640
rect 13069 4538 13103 4568
rect 13069 4534 13103 4538
rect 13069 4470 13103 4496
rect 13069 4462 13103 4470
rect 13069 4402 13103 4424
rect 13069 4390 13103 4402
rect 13069 4334 13103 4352
rect 13069 4318 13103 4334
rect 13069 4266 13103 4280
rect 13069 4246 13103 4266
rect 13069 4198 13103 4208
rect 13069 4174 13103 4198
rect 13069 4130 13103 4136
rect 13069 4102 13103 4130
rect 13069 4062 13103 4064
rect 13069 4030 13103 4062
rect 13069 3960 13103 3992
rect 13069 3958 13103 3960
rect 13069 3892 13103 3920
rect 13069 3886 13103 3892
rect 13069 3824 13103 3848
rect 13069 3814 13103 3824
rect 13069 3756 13103 3776
rect 13069 3742 13103 3756
rect 13069 3688 13103 3704
rect 13069 3670 13103 3688
rect 13069 3620 13103 3632
rect 13069 3598 13103 3620
rect 13069 3552 13103 3560
rect 13069 3526 13103 3552
rect 13069 3484 13103 3488
rect 13069 3454 13103 3484
rect 13069 3382 13103 3416
rect 13069 3314 13103 3344
rect 13069 3310 13103 3314
rect 13069 3246 13103 3272
rect 13069 3238 13103 3246
rect 13069 3178 13103 3200
rect 13069 3166 13103 3178
rect 13069 3110 13103 3128
rect 13069 3094 13103 3110
rect 13069 3042 13103 3056
rect 13069 3022 13103 3042
rect 13069 2974 13103 2984
rect 13069 2950 13103 2974
rect 13069 2906 13103 2912
rect 13069 2878 13103 2906
rect 13069 2838 13103 2840
rect 13069 2806 13103 2838
rect 13069 2736 13103 2768
rect 13069 2734 13103 2736
rect 13069 2668 13103 2696
rect 13069 2662 13103 2668
rect 13069 2600 13103 2623
rect 13069 2589 13103 2600
rect 13069 2532 13103 2550
rect 13069 2516 13103 2532
rect 13069 2464 13103 2477
rect 13069 2443 13103 2464
rect 13069 2396 13103 2404
rect 13069 2370 13103 2396
rect 13069 2328 13103 2331
rect 13069 2297 13103 2328
rect 13069 2226 13103 2258
rect 13069 2224 13103 2226
rect 13069 2158 13103 2185
rect 13069 2151 13103 2158
rect 13069 2090 13103 2112
rect 13069 2078 13103 2090
rect 13069 2022 13103 2039
rect 13069 2005 13103 2022
rect 13069 1954 13103 1966
rect 13069 1932 13103 1954
rect 13069 1886 13103 1893
rect 13069 1859 13103 1886
rect 13069 1818 13103 1820
rect 13069 1786 13103 1818
rect 13069 1716 13103 1747
rect 13069 1713 13103 1716
rect 13069 1648 13103 1674
rect 13069 1640 13103 1648
rect 13069 1580 13103 1601
rect 13069 1567 13103 1580
rect 13069 1512 13103 1528
rect 13069 1494 13103 1512
rect 13069 1444 13103 1455
rect 13069 1421 13103 1444
rect 13069 1376 13103 1382
rect 13069 1348 13103 1376
rect 13069 1308 13103 1309
rect 13069 1275 13103 1308
rect 13069 1206 13103 1236
rect 13069 1202 13103 1206
rect 13069 1138 13103 1163
rect 13069 1129 13103 1138
rect 13069 1070 13103 1090
rect 13069 1056 13103 1070
rect 13069 1002 13103 1017
rect 13069 983 13103 1002
rect 13069 934 13103 944
rect 13069 910 13103 934
rect 13069 866 13103 871
rect 13069 837 13103 866
rect 13069 764 13103 798
rect 13069 696 13103 725
rect 13069 691 13103 696
rect 13069 628 13103 652
rect 13069 618 13103 628
rect 13069 560 13103 579
rect 13069 545 13103 560
rect 13069 492 13103 506
rect 10277 446 10280 480
rect 10280 446 10311 480
rect 10350 446 10382 480
rect 10382 446 10384 480
rect 10423 446 10450 480
rect 10450 446 10457 480
rect 10496 446 10518 480
rect 10518 446 10530 480
rect 10569 446 10586 480
rect 10586 446 10603 480
rect 10642 446 10676 480
rect 10715 446 10724 480
rect 10724 446 10749 480
rect 10788 446 10792 480
rect 10792 446 10822 480
rect 10861 446 10894 480
rect 10894 446 10895 480
rect 10934 446 10962 480
rect 10962 446 10968 480
rect 11007 446 11030 480
rect 11030 446 11041 480
rect 11080 446 11098 480
rect 11098 446 11114 480
rect 11153 446 11166 480
rect 11166 446 11187 480
rect 11226 446 11234 480
rect 11234 446 11260 480
rect 11299 446 11302 480
rect 11302 446 11333 480
rect 11372 446 11404 480
rect 11404 446 11406 480
rect 11445 446 11472 480
rect 11472 446 11479 480
rect 11518 446 11540 480
rect 11540 446 11552 480
rect 11591 446 11608 480
rect 11608 446 11625 480
rect 11664 446 11676 480
rect 11676 446 11698 480
rect 11737 446 11744 480
rect 11744 446 11771 480
rect 11810 446 11812 480
rect 11812 446 11844 480
rect 11883 446 11914 480
rect 11914 446 11917 480
rect 11956 446 11982 480
rect 11982 446 11990 480
rect 12029 446 12050 480
rect 12050 446 12063 480
rect 12102 446 12118 480
rect 12118 446 12136 480
rect 12175 446 12186 480
rect 12186 446 12209 480
rect 12248 446 12254 480
rect 12254 446 12282 480
rect 12321 446 12322 480
rect 12322 446 12355 480
rect 12393 446 12424 480
rect 12424 446 12427 480
rect 12465 446 12492 480
rect 12492 446 12499 480
rect 12537 446 12560 480
rect 12560 446 12571 480
rect 12609 446 12628 480
rect 12628 446 12643 480
rect 12681 446 12696 480
rect 12696 446 12715 480
rect 12753 446 12764 480
rect 12764 446 12787 480
rect 13069 472 13103 492
rect 9899 435 9933 438
rect 9899 404 9929 435
rect 9929 404 9933 435
rect 9899 333 9929 366
rect 9929 333 9933 366
rect 9899 332 9933 333
rect 9899 265 9929 294
rect 9929 265 9933 294
rect 9899 260 9933 265
rect 9899 197 9929 222
rect 9929 197 9933 222
rect 13069 424 13103 433
rect 13069 399 13103 424
rect 13069 356 13103 360
rect 13069 326 13103 356
rect 13069 253 13103 287
rect 1185 163 1219 197
rect 1257 163 1282 197
rect 1282 163 1291 197
rect 1329 163 1350 197
rect 1350 163 1363 197
rect 1401 163 1418 197
rect 1418 163 1435 197
rect 1473 163 1486 197
rect 1486 163 1507 197
rect 1545 163 1554 197
rect 1554 163 1579 197
rect 1617 163 1622 197
rect 1622 163 1651 197
rect 1689 163 1690 197
rect 1690 163 1723 197
rect 1761 163 1792 197
rect 1792 163 1795 197
rect 1833 163 1860 197
rect 1860 163 1867 197
rect 1905 163 1928 197
rect 1928 163 1939 197
rect 1977 163 1996 197
rect 1996 163 2011 197
rect 2049 163 2064 197
rect 2064 163 2083 197
rect 2121 163 2132 197
rect 2132 163 2155 197
rect 2193 163 2200 197
rect 2200 163 2227 197
rect 2265 163 2268 197
rect 2268 163 2299 197
rect 2337 163 2370 197
rect 2370 163 2371 197
rect 2409 163 2438 197
rect 2438 163 2443 197
rect 2481 163 2506 197
rect 2506 163 2515 197
rect 2553 163 2574 197
rect 2574 163 2587 197
rect 2625 163 2642 197
rect 2642 163 2659 197
rect 2697 163 2710 197
rect 2710 163 2731 197
rect 2769 163 2778 197
rect 2778 163 2803 197
rect 2841 163 2846 197
rect 2846 163 2875 197
rect 2913 163 2914 197
rect 2914 163 2947 197
rect 2985 163 3016 197
rect 3016 163 3019 197
rect 3057 163 3084 197
rect 3084 163 3091 197
rect 3129 163 3152 197
rect 3152 163 3163 197
rect 3201 163 3220 197
rect 3220 163 3235 197
rect 3273 163 3288 197
rect 3288 163 3307 197
rect 3345 163 3356 197
rect 3356 163 3379 197
rect 3417 163 3424 197
rect 3424 163 3451 197
rect 3489 163 3492 197
rect 3492 163 3523 197
rect 3561 163 3594 197
rect 3594 163 3595 197
rect 3633 163 3662 197
rect 3662 163 3667 197
rect 3705 163 3730 197
rect 3730 163 3739 197
rect 3777 163 3798 197
rect 3798 163 3811 197
rect 3849 163 3866 197
rect 3866 163 3883 197
rect 3921 163 3934 197
rect 3934 163 3955 197
rect 3993 163 4002 197
rect 4002 163 4027 197
rect 4065 163 4070 197
rect 4070 163 4099 197
rect 4137 163 4138 197
rect 4138 163 4171 197
rect 4209 163 4240 197
rect 4240 163 4243 197
rect 4281 163 4308 197
rect 4308 163 4315 197
rect 4353 163 4376 197
rect 4376 163 4387 197
rect 4425 163 4444 197
rect 4444 163 4459 197
rect 4497 163 4512 197
rect 4512 163 4531 197
rect 4569 163 4580 197
rect 4580 163 4603 197
rect 4641 163 4648 197
rect 4648 163 4675 197
rect 4713 163 4716 197
rect 4716 163 4747 197
rect 4785 163 4818 197
rect 4818 163 4819 197
rect 4857 163 4886 197
rect 4886 163 4891 197
rect 4929 163 4954 197
rect 4954 163 4963 197
rect 5001 163 5022 197
rect 5022 163 5035 197
rect 5073 163 5090 197
rect 5090 163 5107 197
rect 5145 163 5158 197
rect 5158 163 5179 197
rect 5217 163 5226 197
rect 5226 163 5251 197
rect 5289 163 5294 197
rect 5294 163 5323 197
rect 5361 163 5362 197
rect 5362 163 5395 197
rect 5433 163 5464 197
rect 5464 163 5467 197
rect 5505 163 5532 197
rect 5532 163 5539 197
rect 5577 163 5600 197
rect 5600 163 5611 197
rect 5649 163 5668 197
rect 5668 163 5683 197
rect 5721 163 5736 197
rect 5736 163 5755 197
rect 5793 163 5804 197
rect 5804 163 5827 197
rect 5865 163 5872 197
rect 5872 163 5899 197
rect 5937 163 5940 197
rect 5940 163 5971 197
rect 6009 163 6042 197
rect 6042 163 6043 197
rect 6081 163 6110 197
rect 6110 163 6115 197
rect 6153 163 6178 197
rect 6178 163 6187 197
rect 6225 163 6246 197
rect 6246 163 6259 197
rect 6297 163 6314 197
rect 6314 163 6331 197
rect 6369 163 6382 197
rect 6382 163 6403 197
rect 6441 163 6450 197
rect 6450 163 6475 197
rect 6513 163 6518 197
rect 6518 163 6547 197
rect 6585 163 6586 197
rect 6586 163 6619 197
rect 6657 163 6688 197
rect 6688 163 6691 197
rect 6729 163 6756 197
rect 6756 163 6763 197
rect 6801 163 6824 197
rect 6824 163 6835 197
rect 6873 163 6892 197
rect 6892 163 6907 197
rect 6945 163 6960 197
rect 6960 163 6979 197
rect 7017 163 7028 197
rect 7028 163 7051 197
rect 7089 163 7096 197
rect 7096 163 7123 197
rect 7161 163 7164 197
rect 7164 163 7195 197
rect 7233 163 7266 197
rect 7266 163 7267 197
rect 7305 163 7334 197
rect 7334 163 7339 197
rect 7377 163 7402 197
rect 7402 163 7411 197
rect 7449 163 7470 197
rect 7470 163 7483 197
rect 7521 163 7538 197
rect 7538 163 7555 197
rect 7593 163 7606 197
rect 7606 163 7627 197
rect 7665 163 7674 197
rect 7674 163 7699 197
rect 7737 163 7742 197
rect 7742 163 7771 197
rect 7809 163 7810 197
rect 7810 163 7843 197
rect 7881 163 7912 197
rect 7912 163 7915 197
rect 7953 163 7980 197
rect 7980 163 7987 197
rect 8025 163 8048 197
rect 8048 163 8059 197
rect 8097 163 8116 197
rect 8116 163 8131 197
rect 8169 163 8184 197
rect 8184 163 8203 197
rect 8241 163 8252 197
rect 8252 163 8275 197
rect 8313 163 8320 197
rect 8320 163 8347 197
rect 8385 163 8388 197
rect 8388 163 8419 197
rect 8457 163 8490 197
rect 8490 163 8491 197
rect 8529 163 8558 197
rect 8558 163 8563 197
rect 8601 163 8626 197
rect 8626 163 8635 197
rect 8673 163 8694 197
rect 8694 163 8707 197
rect 8745 163 8762 197
rect 8762 163 8779 197
rect 8817 163 8830 197
rect 8830 163 8851 197
rect 8889 163 8898 197
rect 8898 163 8923 197
rect 8961 163 8966 197
rect 8966 163 8995 197
rect 9033 163 9034 197
rect 9034 163 9067 197
rect 9105 163 9136 197
rect 9136 163 9139 197
rect 9177 163 9204 197
rect 9204 163 9211 197
rect 9249 163 9272 197
rect 9272 163 9283 197
rect 9321 163 9340 197
rect 9340 163 9355 197
rect 9393 163 9408 197
rect 9408 163 9427 197
rect 9465 163 9476 197
rect 9476 163 9499 197
rect 9537 163 9544 197
rect 9544 163 9571 197
rect 9609 163 9612 197
rect 9612 163 9643 197
rect 9681 163 9714 197
rect 9714 163 9715 197
rect 9754 163 9782 197
rect 9782 163 9788 197
rect 9827 163 9850 197
rect 9850 163 9861 197
rect 9899 188 9933 197
rect 9971 163 10005 197
rect 10044 163 10077 197
rect 10077 163 10078 197
rect 10117 163 10145 197
rect 10145 163 10151 197
rect 10189 163 10213 197
rect 10213 163 10223 197
rect 10261 163 10281 197
rect 10281 163 10295 197
rect 10333 163 10349 197
rect 10349 163 10367 197
rect 10405 163 10417 197
rect 10417 163 10439 197
rect 10477 163 10485 197
rect 10485 163 10511 197
rect 10549 163 10553 197
rect 10553 163 10583 197
rect 10621 163 10655 197
rect 10693 163 10723 197
rect 10723 163 10727 197
rect 10765 163 10791 197
rect 10791 163 10799 197
rect 10837 163 10859 197
rect 10859 163 10871 197
rect 10909 163 10927 197
rect 10927 163 10943 197
rect 10981 163 10995 197
rect 10995 163 11015 197
rect 11053 163 11063 197
rect 11063 163 11087 197
rect 11125 163 11131 197
rect 11131 163 11159 197
rect 11197 163 11199 197
rect 11199 163 11231 197
rect 11269 163 11301 197
rect 11301 163 11303 197
rect 11341 163 11369 197
rect 11369 163 11375 197
rect 11413 163 11437 197
rect 11437 163 11447 197
rect 11485 163 11505 197
rect 11505 163 11519 197
rect 11557 163 11573 197
rect 11573 163 11591 197
rect 11629 163 11641 197
rect 11641 163 11663 197
rect 11701 163 11709 197
rect 11709 163 11735 197
rect 11773 163 11777 197
rect 11777 163 11807 197
rect 11845 163 11879 197
rect 11917 163 11947 197
rect 11947 163 11951 197
rect 11989 163 12015 197
rect 12015 163 12023 197
rect 12061 163 12083 197
rect 12083 163 12095 197
rect 12133 163 12151 197
rect 12151 163 12167 197
rect 12205 163 12219 197
rect 12219 163 12239 197
rect 12277 163 12287 197
rect 12287 163 12311 197
rect 12349 163 12355 197
rect 12355 163 12383 197
rect 12421 163 12423 197
rect 12423 163 12455 197
rect 12493 163 12525 197
rect 12525 163 12527 197
rect 12565 163 12593 197
rect 12593 163 12599 197
rect 12637 163 12661 197
rect 12661 163 12671 197
rect 12709 163 12729 197
rect 12729 163 12743 197
rect 12781 163 12797 197
rect 12797 163 12815 197
rect 12853 163 12865 197
rect 12865 163 12887 197
rect 12925 163 12933 197
rect 12933 163 12959 197
rect 12997 163 13001 197
rect 13001 163 13031 197
rect 13069 180 13103 214
<< metal1 >>
rect 1191 14234 11117 14240
rect 1191 14200 1235 14234
rect 1269 14200 1308 14234
rect 1342 14200 1381 14234
rect 1415 14200 1454 14234
rect 1488 14200 1527 14234
rect 1561 14200 1600 14234
rect 1634 14200 1673 14234
rect 1707 14200 1746 14234
rect 1780 14200 1819 14234
rect 1853 14200 1892 14234
rect 1926 14200 1965 14234
rect 1999 14200 2038 14234
rect 2072 14200 2111 14234
rect 2145 14200 2183 14234
rect 2217 14200 2255 14234
rect 2289 14200 2327 14234
rect 2361 14200 2399 14234
rect 2433 14200 2471 14234
rect 2505 14200 2543 14234
rect 2577 14200 2615 14234
rect 2649 14200 2687 14234
rect 2721 14200 2759 14234
rect 2793 14200 2831 14234
rect 2865 14200 2903 14234
rect 2937 14200 2975 14234
rect 3009 14200 3047 14234
rect 3081 14200 3119 14234
rect 3153 14200 3191 14234
rect 3225 14200 3263 14234
rect 3297 14200 3335 14234
rect 3369 14200 3407 14234
rect 3441 14200 3479 14234
rect 3513 14200 3551 14234
rect 3585 14200 3623 14234
rect 3657 14200 3695 14234
rect 3729 14200 3767 14234
rect 3801 14200 3839 14234
rect 3873 14200 3911 14234
rect 3945 14200 3983 14234
rect 4017 14200 4055 14234
rect 4089 14200 4127 14234
rect 4161 14200 4199 14234
rect 4233 14200 4271 14234
rect 4305 14200 4343 14234
rect 4377 14200 4415 14234
rect 4449 14200 4487 14234
rect 4521 14200 4559 14234
rect 4593 14200 4631 14234
rect 4665 14200 4703 14234
rect 4737 14200 4775 14234
rect 4809 14200 4847 14234
rect 4881 14200 4919 14234
rect 4953 14200 4991 14234
rect 5025 14200 5063 14234
rect 5097 14200 5135 14234
rect 5169 14200 5207 14234
rect 5241 14200 5279 14234
rect 5313 14200 5351 14234
rect 5385 14200 5423 14234
rect 5457 14200 5495 14234
rect 5529 14200 5567 14234
rect 5601 14200 5639 14234
rect 5673 14200 5711 14234
rect 5745 14200 5783 14234
rect 5817 14200 5855 14234
rect 5889 14200 5927 14234
rect 5961 14200 5999 14234
rect 6033 14200 6071 14234
rect 6105 14200 6143 14234
rect 6177 14200 6215 14234
rect 6249 14200 6287 14234
rect 6321 14200 6359 14234
rect 6393 14200 6431 14234
rect 6465 14200 6503 14234
rect 6537 14200 6575 14234
rect 6609 14200 6647 14234
rect 6681 14200 6719 14234
rect 6753 14200 6791 14234
rect 6825 14200 6863 14234
rect 6897 14200 6935 14234
rect 6969 14200 7007 14234
rect 7041 14200 7079 14234
rect 7113 14200 7151 14234
rect 7185 14200 7223 14234
rect 7257 14200 7295 14234
rect 7329 14200 7367 14234
rect 7401 14200 7439 14234
rect 7473 14200 7511 14234
rect 7545 14200 7583 14234
rect 7617 14200 7655 14234
rect 7689 14200 7727 14234
rect 7761 14200 7799 14234
rect 7833 14200 7871 14234
rect 7905 14200 7943 14234
rect 7977 14200 8015 14234
rect 8049 14200 8087 14234
rect 8121 14200 8159 14234
rect 8193 14200 8231 14234
rect 8265 14200 8303 14234
rect 8337 14200 8375 14234
rect 8409 14200 8447 14234
rect 8481 14200 8519 14234
rect 8553 14200 8591 14234
rect 8625 14200 8663 14234
rect 8697 14200 8735 14234
rect 8769 14200 8807 14234
rect 8841 14200 8879 14234
rect 8913 14200 8951 14234
rect 8985 14200 9023 14234
rect 9057 14200 9095 14234
rect 9129 14200 9167 14234
rect 9201 14200 9239 14234
rect 9273 14200 9311 14234
rect 9345 14200 9383 14234
rect 9417 14200 9455 14234
rect 9489 14200 9527 14234
rect 9561 14200 9599 14234
rect 9633 14200 9671 14234
rect 9705 14200 9743 14234
rect 9777 14200 9815 14234
rect 9849 14200 9887 14234
rect 9921 14200 9959 14234
rect 9993 14200 10031 14234
rect 10065 14200 10103 14234
rect 10137 14200 10175 14234
rect 10209 14200 10247 14234
rect 10281 14200 10319 14234
rect 10353 14200 10391 14234
rect 10425 14200 10463 14234
rect 10497 14200 10535 14234
rect 10569 14200 10607 14234
rect 10641 14200 10679 14234
rect 10713 14200 10751 14234
rect 10785 14200 10823 14234
rect 10857 14200 10895 14234
rect 10929 14200 10967 14234
rect 11001 14200 11117 14234
rect 1191 14196 11117 14200
rect 1191 14194 11077 14196
rect 1191 14124 1237 14194
tri 1237 14169 1262 14194 nw
tri 9334 14169 9359 14194 ne
tri 4336 14162 4340 14166 se
rect 4340 14162 7303 14166
tri 7303 14162 7307 14166 sw
tri 4318 14144 4336 14162 se
rect 4336 14144 7307 14162
rect 1191 14090 1197 14124
rect 1231 14090 1237 14124
rect 1972 14132 3079 14138
rect 1191 14052 1237 14090
rect 1191 14018 1197 14052
rect 1231 14018 1237 14052
rect 1191 13980 1237 14018
rect 1191 13946 1197 13980
rect 1231 13946 1237 13980
rect 1191 13908 1237 13946
rect 1751 14093 1797 14105
rect 1751 14059 1757 14093
rect 1791 14059 1797 14093
rect 1751 14018 1797 14059
rect 1751 13984 1757 14018
rect 1791 13984 1797 14018
rect 1751 13943 1797 13984
rect 1191 13874 1197 13908
rect 1231 13874 1237 13908
rect 1191 13836 1237 13874
rect 1191 13802 1197 13836
rect 1231 13802 1237 13836
rect 1191 13764 1237 13802
rect 1191 13730 1197 13764
rect 1231 13730 1237 13764
rect 1191 13692 1237 13730
rect 1191 13658 1197 13692
rect 1231 13658 1237 13692
rect 1191 13620 1237 13658
rect 1191 13586 1197 13620
rect 1231 13586 1237 13620
rect 1191 13548 1237 13586
rect 1191 13514 1197 13548
rect 1231 13514 1237 13548
rect 1191 13476 1237 13514
rect 1191 13442 1197 13476
rect 1231 13442 1237 13476
rect 1191 13404 1237 13442
rect 1191 13370 1197 13404
rect 1231 13370 1237 13404
rect 1191 13332 1237 13370
rect 1191 13298 1197 13332
rect 1231 13298 1237 13332
rect 1191 13260 1237 13298
rect 1191 13226 1197 13260
rect 1231 13226 1237 13260
rect 1191 13188 1237 13226
rect 1191 13154 1197 13188
rect 1231 13154 1237 13188
rect 1191 13116 1237 13154
rect 1191 13082 1197 13116
rect 1231 13082 1237 13116
rect 1191 13043 1237 13082
rect 1191 13009 1197 13043
rect 1231 13009 1237 13043
rect 1191 12970 1237 13009
rect 1191 12936 1197 12970
rect 1231 12936 1237 12970
rect 1191 12897 1237 12936
rect 1191 12863 1197 12897
rect 1231 12863 1237 12897
rect 1191 12824 1237 12863
rect 1191 12790 1197 12824
rect 1231 12790 1237 12824
rect 1191 12751 1237 12790
rect 1191 12717 1197 12751
rect 1231 12717 1237 12751
rect 1191 12678 1237 12717
rect 1191 12644 1197 12678
rect 1231 12644 1237 12678
rect 1191 12605 1237 12644
rect 1191 12571 1197 12605
rect 1231 12571 1237 12605
rect 1191 12532 1237 12571
rect 1191 12498 1197 12532
rect 1231 12498 1237 12532
rect 1191 12459 1237 12498
rect 1191 12425 1197 12459
rect 1231 12425 1237 12459
rect 1191 12386 1237 12425
rect 1191 12352 1197 12386
rect 1231 12352 1237 12386
tri 1179 12233 1191 12245 se
rect 1191 12233 1237 12352
rect 1179 12225 1237 12233
tri 1176 11842 1179 11845 se
rect 1179 11842 1225 12225
tri 1225 12213 1237 12225 nw
rect 1342 13881 1348 13933
rect 1400 13881 1413 13933
rect 1465 13881 1471 13933
rect 1751 13909 1757 13943
rect 1791 13909 1797 13943
rect 1342 13874 1418 13881
tri 1418 13874 1425 13881 nw
rect 1342 13873 1417 13874
tri 1417 13873 1418 13874 nw
rect 1342 13868 1412 13873
tri 1412 13868 1417 13873 nw
rect 1751 13868 1797 13909
rect 1342 13044 1400 13868
tri 1400 13856 1412 13868 nw
rect 1342 13010 1357 13044
rect 1391 13010 1400 13044
rect 1342 12972 1400 13010
rect 1342 12938 1357 12972
rect 1391 12938 1400 12972
rect 1342 12900 1400 12938
rect 1342 12866 1357 12900
rect 1391 12866 1400 12900
rect 1342 12828 1400 12866
rect 1342 12794 1357 12828
rect 1391 12794 1400 12828
rect 1342 12755 1400 12794
rect 1342 12721 1357 12755
rect 1391 12721 1400 12755
rect 1342 12682 1400 12721
rect 1342 12648 1357 12682
rect 1391 12648 1400 12682
rect 1342 12609 1400 12648
rect 1342 12575 1357 12609
rect 1391 12575 1400 12609
rect 1342 12536 1400 12575
rect 1342 12502 1357 12536
rect 1391 12502 1400 12536
tri 1225 11842 1228 11845 sw
rect 1176 11836 1228 11842
rect 1176 11763 1228 11784
tri 1228 11729 1253 11754 sw
rect 1228 11723 1314 11729
rect 1228 11711 1268 11723
rect 1176 11690 1185 11711
rect 1219 11690 1268 11711
rect 1228 11689 1268 11690
rect 1302 11689 1314 11723
rect 1228 11683 1314 11689
tri 1228 11658 1253 11683 nw
rect 1176 11617 1185 11638
rect 1219 11617 1228 11638
tri 1337 11579 1342 11584 se
rect 1342 11579 1400 12502
rect 1604 13835 1656 13841
rect 1604 13767 1656 13783
rect 1604 13699 1656 13715
rect 1604 13631 1656 13647
rect 1604 13563 1656 13579
rect 1604 13044 1656 13511
rect 1604 13010 1613 13044
rect 1647 13010 1656 13044
rect 1604 12972 1656 13010
rect 1604 12938 1613 12972
rect 1647 12938 1656 12972
rect 1604 12900 1656 12938
rect 1604 12866 1613 12900
rect 1647 12866 1656 12900
rect 1604 12828 1656 12866
rect 1604 12794 1613 12828
rect 1647 12794 1656 12828
rect 1604 12755 1656 12794
rect 1604 12721 1613 12755
rect 1647 12721 1656 12755
rect 1604 12682 1656 12721
rect 1604 12648 1613 12682
rect 1647 12648 1656 12682
rect 1604 12609 1656 12648
rect 1604 12575 1613 12609
rect 1647 12575 1656 12609
rect 1604 12536 1656 12575
rect 1604 12502 1613 12536
rect 1647 12502 1656 12536
rect 1604 12490 1656 12502
rect 1751 13834 1757 13868
rect 1791 13834 1797 13868
rect 1751 13793 1797 13834
rect 1751 13759 1757 13793
rect 1791 13759 1797 13793
rect 1751 13718 1797 13759
rect 1751 13684 1757 13718
rect 1791 13684 1797 13718
rect 1751 13643 1797 13684
rect 1751 13609 1757 13643
rect 1791 13609 1797 13643
rect 1751 13568 1797 13609
rect 1751 13534 1757 13568
rect 1791 13534 1797 13568
rect 1751 13493 1797 13534
rect 1751 13459 1757 13493
rect 1791 13459 1797 13493
rect 1751 13418 1797 13459
rect 1751 13384 1757 13418
rect 1791 13384 1797 13418
rect 1751 13343 1797 13384
rect 1751 13309 1757 13343
rect 1791 13309 1797 13343
rect 1751 13268 1797 13309
rect 1751 13234 1757 13268
rect 1791 13234 1797 13268
rect 1751 13193 1797 13234
rect 1751 13159 1757 13193
rect 1791 13159 1797 13193
rect 1751 13119 1797 13159
rect 1751 13085 1757 13119
rect 1791 13085 1797 13119
rect 1751 13045 1797 13085
rect 1751 13011 1757 13045
rect 1791 13011 1797 13045
rect 1751 12971 1797 13011
rect 1751 12937 1757 12971
rect 1791 12937 1797 12971
rect 1751 12897 1797 12937
rect 1751 12863 1757 12897
rect 1791 12863 1797 12897
rect 1751 12823 1797 12863
rect 1751 12789 1757 12823
rect 1791 12789 1797 12823
rect 1751 12749 1797 12789
rect 1751 12715 1757 12749
rect 1791 12715 1797 12749
rect 1751 12675 1797 12715
rect 1751 12641 1757 12675
rect 1791 12641 1797 12675
rect 1751 12601 1797 12641
rect 1751 12567 1757 12601
rect 1791 12567 1797 12601
rect 1751 12527 1797 12567
rect 1751 12493 1757 12527
rect 1791 12493 1797 12527
rect 1751 12481 1797 12493
rect 1972 14098 1984 14132
rect 2018 14098 2059 14132
rect 2093 14098 2134 14132
rect 2168 14098 2209 14132
rect 2243 14098 2284 14132
rect 2318 14098 2359 14132
rect 2393 14098 2434 14132
rect 2468 14098 2509 14132
rect 2543 14098 2584 14132
rect 2618 14098 2659 14132
rect 2693 14098 2734 14132
rect 2768 14098 2809 14132
rect 2843 14098 2884 14132
rect 2918 14098 2959 14132
rect 2993 14098 3033 14132
rect 3067 14098 3079 14132
rect 1972 14018 3079 14098
rect 3281 14093 3327 14105
rect 3281 14059 3287 14093
rect 3321 14059 3327 14093
tri 3079 14018 3100 14039 sw
tri 3260 14018 3281 14039 se
rect 3281 14018 3327 14059
rect 1972 14014 3100 14018
tri 3100 14014 3104 14018 sw
tri 3256 14014 3260 14018 se
rect 3260 14014 3287 14018
rect 1972 13962 3212 14014
rect 3214 14013 3250 14014
rect 3213 13963 3251 14013
rect 3252 13984 3287 14014
rect 3321 13984 3327 14018
rect 3214 13962 3250 13963
rect 3252 13962 3327 13984
rect 1972 13946 3088 13962
tri 3088 13946 3104 13962 nw
tri 3256 13946 3272 13962 ne
rect 3272 13946 3327 13962
rect 1972 13943 3085 13946
tri 3085 13943 3088 13946 nw
tri 3272 13943 3275 13946 ne
rect 3275 13943 3327 13946
rect 1972 13361 3079 13943
tri 3079 13937 3085 13943 nw
tri 3275 13937 3281 13943 ne
rect 1972 13309 1996 13361
rect 2048 13309 2073 13361
rect 2125 13309 2150 13361
rect 2202 13309 2227 13361
rect 2279 13309 2304 13361
rect 2356 13309 2384 13361
rect 2436 13309 2461 13361
rect 2513 13309 2538 13361
rect 2590 13309 2615 13361
rect 2667 13309 2692 13361
rect 2744 13309 2769 13361
rect 2821 13309 2843 13361
rect 2895 13309 2918 13361
rect 2970 13309 2993 13361
rect 3045 13309 3079 13361
rect 1972 13293 3079 13309
rect 1972 13241 1996 13293
rect 2048 13241 2073 13293
rect 2125 13241 2150 13293
rect 2202 13241 2227 13293
rect 2279 13241 2304 13293
rect 2356 13241 2384 13293
rect 2436 13241 2461 13293
rect 2513 13241 2538 13293
rect 2590 13241 2615 13293
rect 2667 13241 2692 13293
rect 2744 13241 2769 13293
rect 2821 13241 2843 13293
rect 2895 13241 2918 13293
rect 2970 13241 2993 13293
rect 3045 13241 3079 13293
rect 1972 13225 3079 13241
rect 1972 13173 1996 13225
rect 2048 13173 2073 13225
rect 2125 13173 2150 13225
rect 2202 13173 2227 13225
rect 2279 13173 2304 13225
rect 2356 13173 2384 13225
rect 2436 13173 2461 13225
rect 2513 13173 2538 13225
rect 2590 13173 2615 13225
rect 2667 13173 2692 13225
rect 2744 13173 2769 13225
rect 2821 13173 2843 13225
rect 2895 13173 2918 13225
rect 2970 13173 2993 13225
rect 3045 13173 3079 13225
rect 1972 13157 3079 13173
rect 1972 13105 1996 13157
rect 2048 13105 2073 13157
rect 2125 13105 2150 13157
rect 2202 13105 2227 13157
rect 2279 13105 2304 13157
rect 2356 13105 2384 13157
rect 2436 13105 2461 13157
rect 2513 13105 2538 13157
rect 2590 13105 2615 13157
rect 2667 13105 2692 13157
rect 2744 13105 2769 13157
rect 2821 13105 2843 13157
rect 2895 13105 2918 13157
rect 2970 13105 2993 13157
rect 3045 13105 3079 13157
rect 1972 13089 3079 13105
rect 1972 13037 1996 13089
rect 2048 13037 2073 13089
rect 2125 13037 2150 13089
rect 2202 13037 2227 13089
rect 2279 13037 2304 13089
rect 2356 13037 2384 13089
rect 2436 13037 2461 13089
rect 2513 13037 2538 13089
rect 2590 13037 2615 13089
rect 2667 13037 2692 13089
rect 2744 13037 2769 13089
rect 2821 13037 2843 13089
rect 2895 13037 2918 13089
rect 2970 13037 2993 13089
rect 3045 13037 3079 13089
rect 1972 12482 3079 13037
rect 3281 13909 3287 13943
rect 3321 13909 3327 13943
rect 3281 13868 3327 13909
rect 3281 13834 3287 13868
rect 3321 13834 3327 13868
rect 3281 13793 3327 13834
rect 3688 13980 3890 14144
rect 3688 13946 3700 13980
rect 3734 13946 3772 13980
rect 3806 13946 3844 13980
rect 3878 13946 3890 13980
rect 3281 13759 3287 13793
rect 3321 13759 3327 13793
rect 3281 13718 3327 13759
rect 3281 13684 3287 13718
rect 3321 13684 3327 13718
rect 3281 13643 3327 13684
rect 3281 13609 3287 13643
rect 3321 13609 3327 13643
rect 3281 13568 3327 13609
rect 3281 13534 3287 13568
rect 3321 13534 3327 13568
rect 3281 13493 3327 13534
rect 3281 13459 3287 13493
rect 3321 13459 3327 13493
rect 3281 13418 3327 13459
rect 3281 13384 3287 13418
rect 3321 13384 3327 13418
rect 3281 13343 3327 13384
rect 3281 13309 3287 13343
rect 3321 13309 3327 13343
rect 3281 13268 3327 13309
rect 3281 13234 3287 13268
rect 3321 13234 3327 13268
rect 3281 13193 3327 13234
rect 3281 13159 3287 13193
rect 3321 13159 3327 13193
rect 3281 13119 3327 13159
rect 3281 13085 3287 13119
rect 3321 13085 3327 13119
rect 3281 13045 3327 13085
tri 3264 13011 3281 13028 se
rect 3281 13011 3287 13045
rect 3321 13011 3327 13045
tri 3256 13003 3264 13011 se
rect 3264 13003 3327 13011
rect 3135 12997 3214 13003
rect 3187 12951 3214 12997
rect 3215 12952 3216 13002
rect 3252 12952 3253 13002
rect 3254 12971 3327 13003
rect 3254 12951 3287 12971
rect 3187 12945 3198 12951
rect 3135 12937 3198 12945
tri 3198 12937 3212 12951 nw
tri 3256 12937 3270 12951 ne
rect 3270 12937 3287 12951
rect 3321 12937 3327 12971
rect 3135 12933 3190 12937
rect 3187 12929 3190 12933
tri 3190 12929 3198 12937 nw
tri 3270 12929 3278 12937 ne
rect 3278 12929 3327 12937
rect 3187 12927 3188 12929
tri 3188 12927 3190 12929 nw
tri 3278 12927 3280 12929 ne
rect 3280 12927 3327 12929
tri 3187 12926 3188 12927 nw
tri 3280 12926 3281 12927 ne
rect 3135 12875 3187 12881
rect 3281 12897 3327 12927
rect 1428 12458 1447 12467
rect 1428 12424 1440 12458
rect 1428 12415 1447 12424
rect 1499 12415 1511 12467
rect 1563 12415 1575 12467
rect 1972 12448 1984 12482
rect 2018 12448 2059 12482
rect 2093 12448 2134 12482
rect 2168 12448 2209 12482
rect 2243 12448 2284 12482
rect 2318 12448 2359 12482
rect 2393 12448 2434 12482
rect 2468 12448 2509 12482
rect 2543 12448 2584 12482
rect 2618 12448 2659 12482
rect 2693 12448 2734 12482
rect 2768 12448 2809 12482
rect 2843 12448 2884 12482
rect 2918 12448 2959 12482
rect 2993 12448 3033 12482
rect 3067 12448 3079 12482
rect 3281 12863 3287 12897
rect 3321 12863 3327 12897
rect 3281 12823 3327 12863
rect 3281 12789 3287 12823
rect 3321 12789 3327 12823
rect 3281 12749 3327 12789
rect 3281 12715 3287 12749
rect 3321 12715 3327 12749
rect 3281 12675 3327 12715
rect 3281 12641 3287 12675
rect 3321 12641 3327 12675
rect 3281 12601 3327 12641
rect 3281 12567 3287 12601
rect 3321 12567 3327 12601
rect 3281 12527 3327 12567
rect 3281 12493 3287 12527
rect 3321 12493 3327 12527
rect 3281 12481 3327 12493
rect 3407 13568 3609 13833
rect 3407 13534 3419 13568
rect 3453 13534 3491 13568
rect 3525 13534 3563 13568
rect 3597 13534 3609 13568
rect 3407 13056 3609 13534
rect 3407 13022 3419 13056
rect 3453 13022 3491 13056
rect 3525 13022 3563 13056
rect 3597 13022 3609 13056
rect 3407 12643 3609 13022
rect 3407 12591 3477 12643
rect 3529 12591 3609 12643
rect 3407 12579 3609 12591
rect 3407 12527 3477 12579
rect 3529 12574 3609 12579
rect 3529 12567 3602 12574
tri 3602 12567 3609 12574 nw
rect 3688 13824 3890 13946
rect 3688 13790 3700 13824
rect 3734 13790 3772 13824
rect 3806 13790 3844 13824
rect 3878 13790 3890 13824
rect 3688 13361 3890 13790
rect 3740 13309 3762 13361
rect 3814 13309 3838 13361
rect 3688 13293 3700 13309
rect 3734 13293 3772 13309
rect 3806 13293 3844 13309
rect 3878 13293 3890 13309
rect 3740 13241 3762 13293
rect 3814 13241 3838 13293
rect 3688 13225 3890 13241
rect 3740 13173 3762 13225
rect 3814 13173 3838 13225
rect 3688 13157 3890 13173
rect 3740 13105 3762 13157
rect 3814 13105 3838 13157
rect 3688 13089 3890 13105
rect 3740 13037 3762 13089
rect 3814 13037 3838 13089
rect 3688 12800 3890 13037
rect 3688 12766 3700 12800
rect 3734 12766 3772 12800
rect 3806 12766 3844 12800
rect 3878 12766 3890 12800
rect 3688 12644 3890 12766
rect 3688 12610 3700 12644
rect 3734 12610 3772 12644
rect 3806 12610 3844 12644
rect 3878 12610 3890 12644
rect 3529 12560 3595 12567
tri 3595 12560 3602 12567 nw
rect 3529 12550 3585 12560
tri 3585 12550 3595 12560 nw
rect 3529 12527 3551 12550
rect 3407 12516 3551 12527
tri 3551 12516 3585 12550 nw
rect 3688 12528 3890 12610
rect 3969 13740 4171 14144
tri 4306 14132 4318 14144 se
rect 4318 14132 7307 14144
tri 7307 14132 7337 14162 sw
tri 4272 14098 4306 14132 se
rect 4306 14120 7337 14132
rect 4306 14098 4450 14120
tri 4450 14098 4472 14120 nw
tri 7179 14098 7201 14120 ne
rect 7201 14098 7337 14120
tri 7337 14098 7371 14132 sw
tri 4267 14093 4272 14098 se
rect 4272 14093 4447 14098
tri 4447 14095 4450 14098 nw
tri 7201 14095 7204 14098 ne
tri 4248 14074 4267 14093 se
rect 4267 14074 4447 14093
rect 7204 14093 7371 14098
tri 7371 14093 7376 14098 sw
rect 3969 13706 4131 13740
rect 4165 13706 4171 13740
rect 3969 13652 4171 13706
rect 3969 13618 4131 13652
rect 4165 13618 4171 13652
rect 3969 13485 4171 13618
rect 3969 13451 4131 13485
rect 4165 13451 4171 13485
rect 3969 13397 4171 13451
rect 3969 13363 4131 13397
rect 4165 13363 4171 13397
rect 3969 13228 4171 13363
rect 3969 13194 4131 13228
rect 4165 13194 4171 13228
rect 3969 13140 4171 13194
rect 3969 13106 4131 13140
rect 4165 13106 4171 13140
rect 3969 13003 4171 13106
rect 3969 12951 3975 13003
rect 4027 12951 4039 13003
rect 4091 12951 4103 13003
rect 4155 12972 4171 13003
rect 3969 12938 4131 12951
rect 4165 12938 4171 12972
rect 3969 12884 4171 12938
rect 3969 12850 4131 12884
rect 4165 12850 4171 12884
rect 3969 12528 4171 12850
tri 4245 14071 4248 14074 se
rect 4248 14071 4447 14074
rect 4245 13834 4447 14071
rect 4245 13800 4251 13834
rect 4285 13800 4447 13834
rect 4245 13746 4447 13800
rect 4245 13712 4251 13746
rect 4285 13712 4447 13746
rect 4245 13662 4447 13712
rect 4245 13628 4257 13662
rect 4291 13628 4329 13662
rect 4363 13628 4401 13662
rect 4435 13628 4447 13662
rect 4245 12810 4447 13628
rect 4245 12776 4251 12810
rect 4285 12776 4447 12810
rect 4245 12722 4447 12776
rect 4245 12688 4251 12722
rect 4285 12688 4447 12722
rect 1972 12442 3079 12448
tri 1500 12386 1529 12415 ne
tri 1335 11577 1337 11579 se
rect 1337 11577 1400 11579
rect 1176 11544 1185 11565
rect 1219 11544 1228 11565
tri 1318 11560 1335 11577 se
rect 1335 11560 1400 11577
tri 1301 11543 1318 11560 se
rect 1318 11543 1383 11560
tri 1383 11543 1400 11560 nw
rect 1176 11470 1185 11492
rect 1219 11470 1228 11492
rect 1176 11412 1185 11418
tri 1176 11409 1179 11412 ne
rect 1179 11397 1185 11412
rect 1219 11412 1228 11418
rect 1219 11397 1225 11412
tri 1225 11409 1228 11412 nw
tri 1278 11520 1301 11543 se
rect 1301 11520 1347 11543
rect 1278 11507 1347 11520
tri 1347 11507 1383 11543 nw
rect 1278 11504 1344 11507
tri 1344 11504 1347 11507 nw
rect 1179 11358 1225 11397
rect 1179 11324 1185 11358
rect 1219 11324 1225 11358
rect 1179 11285 1225 11324
rect 1179 11251 1185 11285
rect 1219 11251 1225 11285
rect 1179 11213 1225 11251
rect 1179 11179 1185 11213
rect 1219 11179 1225 11213
rect 1179 11141 1225 11179
rect 1179 11107 1185 11141
rect 1219 11107 1225 11141
rect 1179 11069 1225 11107
rect 1179 11035 1185 11069
rect 1219 11035 1225 11069
rect 1179 10997 1225 11035
rect 1179 10963 1185 10997
rect 1219 10963 1225 10997
rect 1179 10925 1225 10963
rect 1179 10891 1185 10925
rect 1219 10891 1225 10925
rect 1179 10853 1225 10891
rect 1179 10819 1185 10853
rect 1219 10819 1225 10853
rect 1179 10781 1225 10819
rect 1179 10747 1185 10781
rect 1219 10747 1225 10781
rect 1179 10709 1225 10747
rect 1179 10675 1185 10709
rect 1219 10675 1225 10709
rect 1179 10637 1225 10675
rect 1179 10603 1185 10637
rect 1219 10603 1225 10637
rect 1179 10565 1225 10603
rect 1179 10531 1185 10565
rect 1219 10531 1225 10565
rect 1179 10493 1225 10531
rect 1179 10459 1185 10493
rect 1219 10459 1225 10493
rect 1179 10421 1225 10459
rect 1179 10387 1185 10421
rect 1219 10387 1225 10421
rect 1179 10349 1225 10387
rect 1179 10315 1185 10349
rect 1219 10315 1225 10349
tri 1160 10290 1179 10309 se
rect 1179 10290 1225 10315
tri 1147 10277 1160 10290 se
rect 1160 10277 1225 10290
tri 1117 10247 1147 10277 se
rect 1147 10247 1185 10277
rect 1117 10243 1185 10247
rect 1219 10252 1225 10277
tri 1225 10252 1228 10255 sw
rect 1219 10247 1228 10252
tri 1228 10247 1233 10252 sw
rect 1219 10243 1233 10247
rect 1117 10241 1233 10243
rect 1169 10189 1181 10241
rect 1117 10171 1185 10189
rect 1219 10171 1233 10189
rect 1117 10133 1233 10171
rect 1117 10114 1185 10133
rect 1219 10114 1233 10133
rect 1169 10062 1181 10114
rect 1117 10061 1233 10062
rect 1117 10027 1185 10061
rect 1219 10056 1233 10061
rect 1219 10027 1225 10056
tri 1225 10048 1233 10056 nw
rect 1117 9989 1225 10027
rect 1117 9955 1185 9989
rect 1219 9955 1225 9989
rect 1117 9917 1225 9955
rect 1117 9883 1185 9917
rect 1219 9883 1225 9917
rect 1117 9845 1225 9883
rect 1117 9811 1185 9845
rect 1219 9811 1225 9845
rect 1117 9773 1225 9811
rect 1117 9739 1185 9773
rect 1219 9739 1225 9773
rect 1117 9701 1225 9739
rect 1117 9667 1185 9701
rect 1219 9667 1225 9701
rect 1117 9629 1225 9667
rect 1117 9595 1185 9629
rect 1219 9595 1225 9629
rect 1117 9557 1225 9595
rect 1117 9523 1185 9557
rect 1219 9523 1225 9557
rect 1117 9485 1225 9523
rect 1117 9451 1185 9485
rect 1219 9451 1225 9485
rect 1117 9413 1225 9451
rect 1117 9379 1185 9413
rect 1219 9379 1225 9413
rect 1117 9341 1225 9379
rect 1117 9307 1185 9341
rect 1219 9307 1225 9341
rect 1117 9269 1225 9307
rect 1117 9235 1185 9269
rect 1219 9235 1225 9269
rect 1117 9197 1225 9235
rect 1117 9163 1185 9197
rect 1219 9163 1225 9197
rect 1117 9125 1225 9163
rect 1117 9091 1185 9125
rect 1219 9091 1225 9125
rect 1117 9053 1225 9091
rect 1117 9019 1185 9053
rect 1219 9019 1225 9053
rect 1117 8981 1225 9019
rect 1117 8947 1185 8981
rect 1219 8947 1225 8981
rect 1117 8909 1225 8947
rect 1117 8875 1185 8909
rect 1219 8875 1225 8909
rect 1117 8837 1225 8875
rect 1117 8803 1185 8837
rect 1219 8803 1225 8837
rect 1117 8765 1225 8803
rect 1117 8731 1185 8765
rect 1219 8731 1225 8765
rect 1117 8693 1225 8731
rect 1117 8659 1185 8693
rect 1219 8659 1225 8693
rect 1117 8621 1225 8659
rect 1117 8587 1185 8621
rect 1219 8587 1225 8621
rect 1117 8549 1225 8587
rect 1117 8515 1185 8549
rect 1219 8515 1225 8549
rect 1117 8477 1225 8515
rect 1117 8443 1185 8477
rect 1219 8443 1225 8477
rect 1117 8405 1225 8443
rect 1117 8371 1185 8405
rect 1219 8371 1225 8405
rect 1117 8333 1225 8371
rect 1117 8299 1185 8333
rect 1219 8299 1225 8333
rect 1117 8261 1225 8299
rect 1117 8227 1185 8261
rect 1219 8227 1225 8261
rect 1117 8189 1225 8227
rect 1117 8155 1185 8189
rect 1219 8155 1225 8189
rect 1117 8152 1225 8155
tri 1225 8152 1233 8160 sw
rect 1117 8146 1233 8152
rect 1117 8017 1185 8030
rect 1219 8017 1233 8030
rect 1169 7965 1181 8017
rect 1117 7939 1185 7965
rect 1219 7959 1233 7965
rect 1219 7939 1225 7959
tri 1225 7951 1233 7959 nw
rect 1117 7901 1225 7939
rect 1117 7867 1185 7901
rect 1219 7867 1225 7901
rect 1117 7829 1225 7867
rect 1117 7795 1185 7829
rect 1219 7795 1225 7829
rect 1117 7757 1225 7795
rect 1117 7723 1185 7757
rect 1219 7723 1225 7757
rect 1117 7685 1225 7723
rect 1117 7651 1185 7685
rect 1219 7651 1225 7685
rect 1117 7613 1225 7651
rect 1117 7579 1185 7613
rect 1219 7579 1225 7613
rect 1117 7541 1225 7579
rect 1117 7507 1185 7541
rect 1219 7507 1225 7541
rect 1117 7469 1225 7507
rect 1117 7435 1185 7469
rect 1219 7435 1225 7469
rect 1117 7397 1225 7435
rect 1117 7363 1185 7397
rect 1219 7363 1225 7397
rect 1117 7325 1225 7363
rect 1117 7291 1185 7325
rect 1219 7291 1225 7325
rect 1117 7253 1225 7291
rect 1117 7219 1185 7253
rect 1219 7219 1225 7253
rect 1117 7181 1225 7219
rect 1117 7147 1185 7181
rect 1219 7147 1225 7181
rect 1117 7109 1225 7147
rect 1117 7075 1185 7109
rect 1219 7075 1225 7109
rect 1117 7037 1225 7075
rect 1117 7003 1185 7037
rect 1219 7003 1225 7037
rect 1117 6965 1225 7003
rect 1117 6931 1185 6965
rect 1219 6931 1225 6965
rect 1117 6893 1225 6931
rect 1117 6859 1185 6893
rect 1219 6859 1225 6893
rect 1117 6821 1225 6859
rect 1117 6787 1185 6821
rect 1219 6787 1225 6821
rect 1117 6749 1225 6787
rect 1117 6715 1185 6749
rect 1219 6715 1225 6749
rect 1117 6677 1225 6715
rect 1117 6643 1185 6677
rect 1219 6643 1225 6677
rect 1117 6605 1225 6643
rect 1117 6571 1185 6605
rect 1219 6571 1225 6605
rect 1117 6533 1225 6571
rect 1117 6499 1185 6533
rect 1219 6499 1225 6533
rect 1117 6461 1225 6499
rect 1117 6427 1185 6461
rect 1219 6427 1225 6461
rect 1117 6389 1225 6427
rect 1117 6355 1185 6389
rect 1219 6355 1225 6389
rect 1117 6317 1225 6355
rect 1117 6283 1185 6317
rect 1219 6283 1225 6317
rect 1117 6245 1225 6283
rect 1117 6211 1185 6245
rect 1219 6211 1225 6245
rect 1117 6173 1225 6211
rect 1117 6139 1185 6173
rect 1219 6139 1225 6173
rect 1117 6101 1225 6139
rect 1117 6067 1185 6101
rect 1219 6067 1225 6101
rect 1117 6029 1225 6067
rect 1117 5995 1185 6029
rect 1219 5995 1225 6029
rect 1117 5957 1225 5995
rect 1117 5923 1185 5957
rect 1219 5923 1225 5957
rect 1117 5885 1225 5923
rect 1117 5851 1185 5885
rect 1219 5851 1225 5885
rect 1117 5813 1225 5851
rect 1117 5779 1185 5813
rect 1219 5779 1225 5813
rect 1117 5741 1225 5779
rect 1117 5707 1185 5741
rect 1219 5707 1225 5741
rect 1117 5669 1225 5707
rect 1117 5635 1185 5669
rect 1219 5635 1225 5669
rect 1117 5597 1225 5635
rect 1117 5563 1185 5597
rect 1219 5563 1225 5597
rect 1117 5525 1225 5563
rect 1117 5491 1185 5525
rect 1219 5491 1225 5525
rect 1117 5453 1225 5491
rect 1117 5419 1185 5453
rect 1219 5419 1225 5453
rect 1117 5381 1225 5419
rect 1117 5347 1185 5381
rect 1219 5347 1225 5381
rect 1117 5309 1225 5347
rect 1117 5275 1185 5309
rect 1219 5275 1225 5309
rect 1117 5237 1225 5275
rect 1117 5203 1185 5237
rect 1219 5203 1225 5237
rect 1117 5165 1225 5203
rect 1117 5131 1185 5165
rect 1219 5131 1225 5165
rect 1117 5093 1225 5131
rect 1117 5059 1185 5093
rect 1219 5059 1225 5093
rect 1117 5021 1225 5059
rect 1117 4987 1185 5021
rect 1219 4987 1225 5021
rect 1117 4949 1225 4987
rect 1117 4915 1185 4949
rect 1219 4915 1225 4949
rect 1117 4893 1225 4915
tri 1225 4893 1226 4894 sw
rect 1117 4886 1226 4893
tri 1226 4886 1233 4893 sw
rect 1117 4880 1233 4886
rect 1169 4828 1181 4880
rect 1117 4814 1233 4828
rect 1169 4762 1181 4814
rect 1117 4756 1233 4762
rect 1117 4733 1225 4756
tri 1225 4748 1233 4756 nw
rect 1117 4699 1185 4733
rect 1219 4699 1225 4733
rect 1117 4661 1225 4699
rect 1117 4627 1185 4661
rect 1219 4627 1225 4661
rect 1117 4589 1225 4627
rect 1117 4555 1185 4589
rect 1219 4555 1225 4589
rect 1117 4517 1225 4555
rect 1117 4483 1185 4517
rect 1219 4483 1225 4517
rect 1117 4445 1225 4483
rect 1117 4411 1185 4445
rect 1219 4411 1225 4445
rect 1117 4373 1225 4411
rect 1117 4339 1185 4373
rect 1219 4339 1225 4373
rect 1117 4301 1225 4339
rect 1117 4267 1185 4301
rect 1219 4267 1225 4301
rect 1117 4229 1225 4267
rect 1117 4195 1185 4229
rect 1219 4195 1225 4229
rect 1117 4157 1225 4195
rect 1117 4123 1185 4157
rect 1219 4123 1225 4157
rect 1117 4085 1225 4123
rect 1117 4051 1185 4085
rect 1219 4051 1225 4085
rect 1117 4013 1225 4051
rect 1117 3979 1185 4013
rect 1219 3979 1225 4013
rect 1117 3941 1225 3979
rect 1117 3907 1185 3941
rect 1219 3907 1225 3941
rect 1117 3869 1225 3907
rect 1117 3835 1185 3869
rect 1219 3835 1225 3869
rect 1117 3797 1225 3835
rect 1117 3763 1185 3797
rect 1219 3763 1225 3797
rect 1117 3725 1225 3763
rect 1117 3691 1185 3725
rect 1219 3691 1225 3725
rect 1117 3653 1225 3691
rect 1117 3619 1185 3653
rect 1219 3619 1225 3653
rect 1117 3581 1225 3619
rect 1117 3547 1185 3581
rect 1219 3547 1225 3581
rect 1117 3509 1225 3547
rect 1117 3475 1185 3509
rect 1219 3475 1225 3509
rect 1117 3437 1225 3475
rect 1117 3403 1185 3437
rect 1219 3403 1225 3437
rect 1117 3365 1225 3403
rect 1117 3331 1185 3365
rect 1219 3331 1225 3365
rect 1117 3293 1225 3331
rect 1117 3259 1185 3293
rect 1219 3259 1225 3293
rect 1117 3221 1225 3259
rect 1117 3187 1185 3221
rect 1219 3187 1225 3221
rect 1117 3149 1225 3187
rect 1117 3115 1185 3149
rect 1219 3115 1225 3149
rect 1117 3077 1225 3115
rect 1117 3043 1185 3077
rect 1219 3043 1225 3077
rect 1117 3005 1225 3043
rect 1117 2971 1185 3005
rect 1219 2971 1225 3005
rect 1117 2933 1225 2971
rect 1117 2899 1185 2933
rect 1219 2899 1225 2933
rect 1117 2861 1225 2899
rect 1117 2827 1185 2861
rect 1219 2827 1225 2861
rect 1117 2789 1225 2827
rect 1117 2755 1185 2789
rect 1219 2755 1225 2789
rect 1117 2717 1225 2755
rect 1117 2683 1185 2717
rect 1219 2683 1225 2717
rect 1117 2645 1225 2683
rect 1117 2611 1185 2645
rect 1219 2611 1225 2645
rect 1117 2573 1225 2611
rect 1117 2539 1185 2573
rect 1219 2539 1225 2573
rect 1117 2501 1225 2539
rect 1117 2467 1185 2501
rect 1219 2467 1225 2501
rect 1117 2429 1225 2467
rect 1117 2395 1185 2429
rect 1219 2395 1225 2429
rect 1117 2357 1225 2395
rect 1117 2323 1185 2357
rect 1219 2323 1225 2357
rect 1117 2285 1225 2323
rect 1117 2251 1185 2285
rect 1219 2251 1225 2285
rect 1117 2213 1225 2251
rect 1117 2179 1185 2213
rect 1219 2179 1225 2213
rect 1117 2141 1225 2179
rect 1117 2107 1185 2141
rect 1219 2107 1225 2141
rect 1117 2069 1225 2107
rect 1117 2035 1185 2069
rect 1219 2035 1225 2069
rect 1117 1997 1225 2035
rect 1117 1963 1185 1997
rect 1219 1963 1225 1997
rect 1278 2036 1336 11504
tri 1336 11496 1344 11504 nw
rect 1529 11486 1575 12415
rect 2048 12270 2178 12276
rect 1639 12175 1975 12181
rect 1639 12141 1651 12175
rect 1685 12141 1743 12175
rect 1777 12141 1836 12175
rect 1870 12141 1929 12175
rect 1963 12141 1975 12175
rect 1639 12120 1975 12141
rect 1639 12103 1758 12120
rect 1874 12103 1975 12120
rect 1639 12069 1651 12103
rect 1685 12069 1743 12103
rect 1874 12069 1929 12103
rect 1963 12069 1975 12103
rect 1639 12031 1758 12069
rect 1874 12031 1975 12069
rect 1639 11997 1651 12031
rect 1685 11997 1743 12031
rect 1874 12004 1929 12031
rect 1777 11997 1836 12004
rect 1870 11997 1929 12004
rect 1963 11997 1975 12031
rect 1639 11991 1975 11997
rect 2164 12154 2178 12270
rect 1618 11680 1624 11732
rect 1676 11680 1689 11732
rect 1741 11723 1754 11732
rect 1806 11723 1819 11732
rect 1871 11723 1884 11732
rect 1747 11689 1754 11723
rect 1871 11689 1879 11723
rect 1741 11680 1754 11689
rect 1806 11680 1819 11689
rect 1871 11680 1884 11689
rect 1936 11680 1950 11732
rect 2002 11680 2008 11732
tri 1575 11486 1592 11503 sw
rect 1529 11483 1592 11486
tri 1529 11470 1542 11483 ne
rect 1542 11470 1592 11483
tri 1592 11470 1608 11486 sw
tri 1542 11435 1577 11470 ne
rect 1577 11435 1608 11470
tri 1608 11435 1643 11470 sw
tri 1577 11431 1581 11435 ne
rect 1581 11431 1643 11435
tri 1643 11431 1647 11435 sw
tri 1581 11429 1583 11431 ne
rect 1583 11429 1647 11431
tri 1647 11429 1649 11431 sw
tri 1583 11420 1592 11429 ne
rect 1592 11420 1649 11429
tri 1649 11420 1658 11429 sw
tri 1592 11400 1612 11420 ne
rect 1384 11228 1436 11240
rect 1384 11194 1396 11228
rect 1430 11194 1436 11228
rect 1384 11154 1436 11194
rect 1384 11120 1396 11154
rect 1430 11120 1436 11154
rect 1384 11080 1436 11120
rect 1384 11046 1396 11080
rect 1430 11046 1436 11080
rect 1384 11006 1436 11046
rect 1384 10972 1396 11006
rect 1430 10972 1436 11006
rect 1384 10932 1436 10972
rect 1384 10898 1396 10932
rect 1430 10898 1436 10932
rect 1384 10858 1436 10898
rect 1384 10824 1396 10858
rect 1430 10824 1436 10858
rect 1384 10784 1436 10824
rect 1384 10750 1396 10784
rect 1430 10750 1436 10784
rect 1384 10710 1436 10750
rect 1384 10676 1396 10710
rect 1430 10676 1436 10710
rect 1384 10636 1436 10676
rect 1384 10602 1396 10636
rect 1430 10602 1436 10636
rect 1384 10561 1436 10602
rect 1384 10527 1396 10561
rect 1430 10527 1436 10561
rect 1384 10486 1436 10527
rect 1384 10452 1396 10486
rect 1430 10452 1436 10486
rect 1384 10142 1436 10452
rect 1384 10108 1396 10142
rect 1430 10108 1436 10142
rect 1384 10068 1436 10108
rect 1384 10034 1396 10068
rect 1430 10034 1436 10068
rect 1384 9994 1436 10034
rect 1384 9960 1396 9994
rect 1430 9960 1436 9994
rect 1384 9920 1436 9960
rect 1384 9886 1396 9920
rect 1430 9886 1436 9920
rect 1384 9849 1436 9886
rect 1384 9783 1436 9797
rect 1384 9698 1436 9731
rect 1384 9664 1396 9698
rect 1430 9664 1436 9698
rect 1384 9624 1436 9664
rect 1384 9590 1396 9624
rect 1430 9590 1436 9624
rect 1384 9550 1436 9590
rect 1384 9516 1396 9550
rect 1430 9516 1436 9550
rect 1384 9475 1436 9516
rect 1384 9441 1396 9475
rect 1430 9441 1436 9475
rect 1384 9400 1436 9441
rect 1384 9366 1396 9400
rect 1430 9366 1436 9400
rect 1384 9286 1436 9366
rect 1384 9252 1396 9286
rect 1430 9252 1436 9286
rect 1384 9212 1436 9252
rect 1384 9178 1396 9212
rect 1430 9178 1436 9212
rect 1384 9138 1436 9178
rect 1384 9104 1396 9138
rect 1430 9104 1436 9138
rect 1384 9064 1436 9104
rect 1384 9030 1396 9064
rect 1430 9030 1436 9064
rect 1384 8990 1436 9030
rect 1384 8956 1396 8990
rect 1430 8956 1436 8990
rect 1384 8916 1436 8956
rect 1384 8882 1396 8916
rect 1430 8882 1436 8916
rect 1384 8842 1436 8882
rect 1384 8808 1396 8842
rect 1430 8808 1436 8842
rect 1384 8768 1436 8808
rect 1384 8734 1396 8768
rect 1430 8734 1436 8768
rect 1384 8694 1436 8734
rect 1384 8660 1396 8694
rect 1430 8660 1436 8694
rect 1384 8619 1436 8660
rect 1384 8585 1396 8619
rect 1430 8585 1436 8619
rect 1384 8544 1436 8585
rect 1384 8510 1396 8544
rect 1430 8510 1436 8544
rect 1384 8252 1436 8510
rect 1384 8218 1396 8252
rect 1430 8218 1436 8252
rect 1384 8180 1436 8218
rect 1384 8146 1396 8180
rect 1430 8146 1436 8180
rect 1384 8108 1436 8146
rect 1384 8074 1396 8108
rect 1430 8074 1436 8108
rect 1384 8036 1436 8074
rect 1384 8002 1396 8036
rect 1430 8002 1436 8036
rect 1384 7964 1436 8002
rect 1384 7930 1396 7964
rect 1430 7930 1436 7964
rect 1384 7892 1436 7930
rect 1384 7858 1396 7892
rect 1430 7858 1436 7892
rect 1384 7820 1436 7858
rect 1384 7786 1396 7820
rect 1430 7786 1436 7820
rect 1384 7748 1436 7786
rect 1384 7714 1396 7748
rect 1430 7714 1436 7748
rect 1384 7676 1436 7714
rect 1384 7642 1396 7676
rect 1430 7642 1436 7676
rect 1384 7604 1436 7642
rect 1384 7570 1396 7604
rect 1430 7570 1436 7604
rect 1384 7531 1436 7570
rect 1384 7497 1396 7531
rect 1430 7497 1436 7531
rect 1384 7458 1436 7497
rect 1384 7424 1396 7458
rect 1430 7424 1436 7458
rect 1384 7412 1436 7424
rect 1384 6474 1436 6480
rect 1384 6408 1436 6422
rect 1384 6320 1436 6356
rect 1384 6286 1396 6320
rect 1430 6286 1436 6320
rect 1384 6246 1436 6286
rect 1384 6212 1396 6246
rect 1430 6212 1436 6246
rect 1384 6172 1436 6212
rect 1384 6138 1396 6172
rect 1430 6138 1436 6172
rect 1384 6098 1436 6138
rect 1384 6064 1396 6098
rect 1430 6064 1436 6098
rect 1384 6024 1436 6064
rect 1384 5990 1396 6024
rect 1430 5990 1436 6024
rect 1384 5950 1436 5990
rect 1384 5916 1396 5950
rect 1430 5916 1436 5950
rect 1384 5876 1436 5916
rect 1384 5842 1396 5876
rect 1430 5842 1436 5876
rect 1384 5801 1436 5842
rect 1384 5767 1396 5801
rect 1430 5767 1436 5801
rect 1384 5726 1436 5767
rect 1384 5692 1396 5726
rect 1430 5692 1436 5726
rect 1384 5382 1436 5692
rect 1384 5348 1396 5382
rect 1430 5348 1436 5382
rect 1384 5308 1436 5348
rect 1384 5274 1396 5308
rect 1430 5274 1436 5308
rect 1384 5234 1436 5274
rect 1384 5200 1396 5234
rect 1430 5200 1436 5234
rect 1384 5160 1436 5200
rect 1384 5126 1396 5160
rect 1430 5126 1436 5160
rect 1384 5086 1436 5126
rect 1384 5052 1396 5086
rect 1430 5052 1436 5086
rect 1384 5012 1436 5052
rect 1384 4978 1396 5012
rect 1430 4978 1436 5012
rect 1384 4938 1436 4978
rect 1384 4904 1396 4938
rect 1430 4904 1436 4938
rect 1384 4864 1436 4904
rect 1384 4830 1396 4864
rect 1430 4830 1436 4864
rect 1384 4790 1436 4830
rect 1384 4756 1396 4790
rect 1430 4756 1436 4790
rect 1384 4715 1436 4756
rect 1384 4681 1396 4715
rect 1430 4681 1436 4715
rect 1384 4640 1436 4681
rect 1384 4606 1396 4640
rect 1430 4606 1436 4640
rect 1384 4526 1436 4606
rect 1384 4492 1396 4526
rect 1430 4492 1436 4526
rect 1384 4452 1436 4492
rect 1384 4418 1396 4452
rect 1430 4418 1436 4452
rect 1384 4378 1436 4418
rect 1384 4344 1396 4378
rect 1430 4344 1436 4378
rect 1384 4304 1436 4344
rect 1384 4270 1396 4304
rect 1430 4270 1436 4304
rect 1384 4230 1436 4270
rect 1384 4196 1396 4230
rect 1430 4196 1436 4230
rect 1384 4156 1436 4196
rect 1384 4122 1396 4156
rect 1430 4122 1436 4156
rect 1384 4082 1436 4122
rect 1384 4048 1396 4082
rect 1430 4048 1436 4082
rect 1384 4008 1436 4048
rect 1384 3974 1396 4008
rect 1430 3974 1436 4008
rect 1384 3934 1436 3974
rect 1384 3900 1396 3934
rect 1430 3900 1436 3934
rect 1384 3859 1436 3900
rect 1384 3825 1396 3859
rect 1430 3825 1436 3859
rect 1384 3784 1436 3825
rect 1384 3750 1396 3784
rect 1430 3750 1436 3784
rect 1384 3440 1436 3750
rect 1384 3406 1396 3440
rect 1430 3406 1436 3440
rect 1384 3366 1436 3406
rect 1384 3332 1396 3366
rect 1430 3332 1436 3366
rect 1384 3292 1436 3332
rect 1384 3258 1396 3292
rect 1430 3258 1436 3292
rect 1384 3218 1436 3258
rect 1384 3184 1396 3218
rect 1430 3184 1436 3218
rect 1384 3144 1436 3184
rect 1384 3110 1396 3144
rect 1430 3110 1436 3144
rect 1384 3070 1436 3110
rect 1384 3036 1396 3070
rect 1430 3036 1436 3070
rect 1384 2996 1436 3036
rect 1384 2962 1396 2996
rect 1430 2962 1436 2996
rect 1384 2922 1436 2962
rect 1384 2888 1396 2922
rect 1430 2888 1436 2922
rect 1384 2848 1436 2888
rect 1384 2814 1396 2848
rect 1430 2814 1436 2848
rect 1384 2773 1436 2814
rect 1384 2739 1396 2773
rect 1430 2739 1436 2773
rect 1384 2698 1436 2739
rect 1384 2664 1396 2698
rect 1430 2664 1436 2698
rect 1384 2652 1436 2664
tri 1336 2036 1338 2038 sw
rect 1278 2026 1338 2036
tri 1338 2026 1348 2036 sw
rect 1278 2021 1348 2026
tri 1348 2021 1353 2026 sw
rect 1278 2014 1353 2021
tri 1278 1987 1305 2014 ne
rect 1305 1987 1353 2014
tri 1353 1987 1387 2021 sw
tri 1305 1985 1307 1987 ne
rect 1307 1985 1387 1987
tri 1387 1985 1389 1987 sw
rect 1117 1925 1225 1963
tri 1307 1954 1338 1985 ne
rect 1338 1954 1389 1985
tri 1389 1954 1420 1985 sw
tri 1338 1951 1341 1954 ne
rect 1341 1951 1420 1954
tri 1420 1951 1423 1954 sw
tri 1341 1948 1344 1951 ne
rect 1344 1948 1423 1951
tri 1423 1948 1426 1951 sw
rect 1117 1891 1185 1925
rect 1219 1891 1225 1925
tri 1344 1914 1378 1948 ne
rect 1378 1914 1426 1948
tri 1426 1914 1460 1948 sw
tri 1378 1910 1382 1914 ne
rect 1382 1910 1460 1914
tri 1460 1910 1464 1914 sw
rect 1117 1853 1225 1891
tri 1382 1876 1416 1910 ne
rect 1416 1876 1464 1910
tri 1464 1876 1498 1910 sw
tri 1416 1875 1417 1876 ne
rect 1417 1875 1498 1876
tri 1498 1875 1499 1876 sw
tri 1417 1872 1420 1875 ne
rect 1420 1872 1499 1875
tri 1499 1872 1502 1875 sw
rect 1117 1819 1185 1853
rect 1219 1819 1225 1853
tri 1420 1841 1451 1872 ne
rect 1451 1841 1502 1872
tri 1502 1841 1533 1872 sw
tri 1451 1835 1457 1841 ne
rect 1457 1835 1533 1841
tri 1533 1835 1539 1841 sw
rect 1117 1781 1225 1819
tri 1457 1801 1491 1835 ne
rect 1491 1801 1539 1835
tri 1539 1801 1573 1835 sw
tri 1491 1790 1502 1801 ne
rect 1502 1790 1573 1801
tri 1573 1790 1584 1801 sw
rect 1117 1747 1185 1781
rect 1219 1747 1225 1781
tri 1502 1768 1524 1790 ne
rect 1524 1768 1584 1790
tri 1524 1766 1526 1768 ne
rect 1117 1709 1225 1747
rect 1117 1675 1185 1709
rect 1219 1675 1225 1709
rect 1117 1637 1225 1675
rect 1117 1603 1185 1637
rect 1219 1603 1225 1637
rect 1117 1565 1225 1603
rect 1117 1531 1185 1565
rect 1219 1531 1225 1565
rect 1117 1493 1225 1531
rect 1117 1459 1185 1493
rect 1219 1459 1225 1493
rect 1117 1421 1225 1459
rect 1117 1387 1185 1421
rect 1219 1387 1225 1421
rect 1117 1349 1225 1387
rect 1117 1315 1185 1349
rect 1219 1315 1225 1349
rect 1117 1277 1225 1315
rect 1117 1243 1185 1277
rect 1219 1243 1225 1277
rect 1117 1205 1225 1243
rect 1117 1171 1185 1205
rect 1219 1171 1225 1205
rect 1117 1133 1225 1171
rect 1117 1099 1185 1133
rect 1219 1099 1225 1133
rect 1117 1061 1225 1099
rect 1117 1027 1185 1061
rect 1219 1027 1225 1061
rect 1117 989 1225 1027
rect 1117 955 1185 989
rect 1219 955 1225 989
rect 1384 1747 1436 1759
rect 1384 1713 1396 1747
rect 1430 1713 1436 1747
rect 1384 1673 1436 1713
rect 1384 1639 1396 1673
rect 1430 1639 1436 1673
rect 1384 1599 1436 1639
rect 1384 1565 1396 1599
rect 1430 1565 1436 1599
rect 1384 1525 1436 1565
rect 1384 1491 1396 1525
rect 1430 1491 1436 1525
rect 1384 1451 1436 1491
rect 1384 1417 1396 1451
rect 1430 1417 1436 1451
rect 1384 1377 1436 1417
rect 1384 1343 1396 1377
rect 1430 1343 1436 1377
rect 1384 1303 1436 1343
rect 1384 1269 1396 1303
rect 1430 1269 1436 1303
rect 1384 1229 1436 1269
rect 1384 1195 1396 1229
rect 1430 1195 1436 1229
rect 1384 1185 1436 1195
rect 1384 1121 1396 1133
rect 1430 1121 1436 1133
rect 1384 1046 1396 1069
rect 1430 1046 1436 1069
rect 1384 1005 1436 1046
rect 1384 971 1396 1005
rect 1430 971 1436 1005
rect 1384 959 1436 971
rect 1117 917 1225 955
rect 1117 883 1185 917
rect 1219 883 1225 917
rect 1117 845 1225 883
rect 1117 811 1185 845
rect 1219 811 1225 845
rect 1117 773 1225 811
rect 1117 739 1185 773
rect 1219 739 1225 773
rect 1117 701 1225 739
rect 1117 667 1185 701
rect 1219 667 1225 701
rect 1117 629 1225 667
rect 1117 595 1185 629
rect 1219 595 1225 629
rect 1117 557 1225 595
rect 1117 523 1185 557
rect 1219 523 1225 557
rect 1526 918 1584 1768
rect 1526 866 1532 918
rect 1526 854 1584 866
rect 1526 802 1532 854
rect 1526 726 1584 802
rect 1526 692 1538 726
rect 1572 692 1584 726
rect 1526 654 1584 692
rect 1526 620 1538 654
rect 1572 620 1584 654
rect 1526 582 1584 620
rect 1526 548 1538 582
rect 1572 548 1584 582
rect 1526 542 1584 548
rect 1612 832 1658 11420
rect 2048 6789 2178 12154
rect 2275 12175 3331 12181
rect 2275 12141 2287 12175
rect 2321 12141 2363 12175
rect 2397 12141 2439 12175
rect 2473 12141 2515 12175
rect 2549 12141 2592 12175
rect 2626 12141 2669 12175
rect 2703 12141 2746 12175
rect 2780 12141 2823 12175
rect 2857 12141 2900 12175
rect 2934 12141 2977 12175
rect 3011 12141 3054 12175
rect 3088 12141 3131 12175
rect 3165 12141 3208 12175
rect 3242 12141 3285 12175
rect 3319 12141 3331 12175
rect 2275 12120 3331 12141
rect 2275 12103 2720 12120
rect 2836 12103 3331 12120
rect 2275 12069 2287 12103
rect 2321 12069 2363 12103
rect 2397 12069 2439 12103
rect 2473 12069 2515 12103
rect 2549 12069 2592 12103
rect 2626 12069 2669 12103
rect 2703 12069 2720 12103
rect 2857 12069 2900 12103
rect 2934 12069 2977 12103
rect 3011 12069 3054 12103
rect 3088 12069 3131 12103
rect 3165 12069 3208 12103
rect 3242 12069 3285 12103
rect 3319 12069 3331 12103
rect 2275 12031 2720 12069
rect 2836 12031 3331 12069
rect 2275 11997 2287 12031
rect 2321 11997 2363 12031
rect 2397 11997 2439 12031
rect 2473 11997 2515 12031
rect 2549 11997 2592 12031
rect 2626 11997 2669 12031
rect 2703 12004 2720 12031
rect 2703 11997 2746 12004
rect 2780 11997 2823 12004
rect 2857 11997 2900 12031
rect 2934 11997 2977 12031
rect 3011 11997 3054 12031
rect 3088 11997 3131 12031
rect 3165 11997 3208 12031
rect 3242 11997 3285 12031
rect 3319 11997 3331 12031
rect 2275 11991 3331 11997
rect 2218 11680 2224 11732
rect 2276 11680 2292 11732
rect 2344 11680 2360 11732
rect 2412 11680 2428 11732
rect 2480 11680 2496 11732
rect 2548 11723 2564 11732
rect 2616 11723 2632 11732
rect 2684 11723 2700 11732
rect 2752 11723 2768 11732
rect 2820 11723 2836 11732
rect 2888 11723 2904 11732
rect 2956 11723 2972 11732
rect 3024 11723 3040 11732
rect 3092 11723 3108 11732
rect 2552 11689 2564 11723
rect 2625 11689 2632 11723
rect 2698 11689 2700 11723
rect 3024 11689 3029 11723
rect 3092 11689 3102 11723
rect 2548 11680 2564 11689
rect 2616 11680 2632 11689
rect 2684 11680 2700 11689
rect 2752 11680 2768 11689
rect 2820 11680 2836 11689
rect 2888 11680 2904 11689
rect 2956 11680 2972 11689
rect 3024 11680 3040 11689
rect 3092 11680 3108 11689
rect 3160 11680 3175 11732
rect 3227 11680 3242 11732
rect 3294 11680 3309 11732
rect 3361 11680 3367 11732
tri 3401 11651 3407 11657 se
rect 3407 11651 3537 12516
tri 3537 12502 3551 12516 nw
rect 3600 12386 4143 12392
rect 3600 12352 3612 12386
rect 3646 12352 3693 12386
rect 3727 12352 3774 12386
rect 3808 12352 3855 12386
rect 3889 12352 3936 12386
rect 3970 12352 4017 12386
rect 4051 12352 4097 12386
rect 4131 12352 4143 12386
rect 3600 12346 4143 12352
tri 3604 12321 3629 12346 ne
rect 3629 11887 3675 12346
tri 3675 12321 3700 12346 nw
rect 3761 12004 3767 12120
rect 3883 12004 3889 12120
tri 3629 11856 3660 11887 ne
rect 3660 11849 3675 11887
tri 3675 11849 3733 11907 sw
rect 3660 11836 3733 11849
rect 3660 11784 3681 11836
rect 3660 11762 3733 11784
tri 3635 11729 3660 11754 se
rect 3660 11729 3681 11762
rect 3565 11723 3681 11729
tri 3733 11729 3758 11754 sw
rect 3733 11723 4204 11729
rect 3565 11689 3577 11723
rect 3611 11710 3681 11723
rect 3733 11710 3765 11723
rect 3611 11689 3693 11710
rect 3727 11689 3765 11710
rect 3799 11689 3843 11723
rect 3877 11689 3921 11723
rect 3955 11689 4000 11723
rect 4034 11689 4079 11723
rect 4113 11689 4158 11723
rect 4192 11689 4204 11723
rect 3565 11688 4204 11689
rect 3565 11683 3681 11688
tri 3635 11658 3660 11683 ne
tri 3400 11650 3401 11651 se
rect 3401 11650 3537 11651
tri 3366 11616 3400 11650 se
rect 3400 11616 3537 11650
tri 3334 11584 3366 11616 se
rect 3366 11603 3537 11616
rect 3366 11584 3513 11603
rect 3334 11579 3513 11584
tri 3513 11579 3537 11603 nw
rect 3660 11636 3681 11683
rect 3733 11683 4204 11688
tri 3733 11658 3758 11683 nw
rect 3660 11616 3693 11636
rect 3727 11616 3733 11636
rect 3660 11614 3733 11616
rect 3334 11577 3511 11579
tri 3511 11577 3513 11579 nw
rect 3334 11543 3477 11577
tri 3477 11543 3511 11577 nw
rect 3660 11562 3681 11614
rect 3660 11543 3693 11562
rect 3727 11543 3733 11562
rect 2234 11429 3233 11435
rect 2234 11395 2246 11429
rect 2280 11395 2319 11429
rect 2353 11395 2392 11429
rect 2426 11395 2465 11429
rect 2499 11395 2538 11429
rect 2572 11395 2611 11429
rect 2234 11357 2611 11395
rect 2234 11323 2246 11357
rect 2280 11323 2319 11357
rect 2353 11323 2392 11357
rect 2426 11323 2465 11357
rect 2499 11323 2538 11357
rect 2572 11323 2611 11357
rect 2234 11285 2611 11323
rect 2234 11251 2246 11285
rect 2280 11251 2319 11285
rect 2353 11251 2392 11285
rect 2426 11251 2465 11285
rect 2499 11251 2538 11285
rect 2572 11251 2611 11285
rect 3221 11251 3233 11429
rect 2234 10396 3233 11251
rect 2234 10362 2246 10396
rect 2280 10362 2319 10396
rect 2353 10362 2392 10396
rect 2426 10362 2465 10396
rect 2499 10362 2538 10396
rect 2572 10362 2611 10396
rect 2234 10324 2611 10362
rect 2234 10290 2246 10324
rect 2280 10290 2319 10324
rect 2353 10290 2392 10324
rect 2426 10290 2465 10324
rect 2499 10290 2538 10324
rect 2572 10290 2611 10324
rect 2234 10252 2611 10290
rect 2234 10218 2246 10252
rect 2280 10218 2319 10252
rect 2353 10218 2392 10252
rect 2426 10218 2465 10252
rect 2499 10218 2538 10252
rect 2572 10218 2611 10252
rect 3221 10218 3233 10396
rect 2234 9343 3233 10218
rect 2234 9309 2246 9343
rect 2280 9309 2319 9343
rect 2353 9309 2392 9343
rect 2426 9309 2465 9343
rect 2499 9309 2538 9343
rect 2572 9309 2611 9343
rect 2645 9309 2683 9343
rect 2717 9309 2755 9343
rect 2789 9309 2827 9343
rect 2861 9309 2899 9343
rect 2933 9309 2971 9343
rect 3005 9309 3043 9343
rect 3077 9309 3115 9343
rect 3149 9309 3187 9343
rect 3221 9309 3233 9343
rect 2234 8457 3233 9309
rect 2234 8423 2246 8457
rect 2280 8423 2319 8457
rect 2353 8423 2392 8457
rect 2426 8423 2465 8457
rect 2499 8423 2538 8457
rect 2572 8423 2611 8457
rect 2234 8385 2611 8423
rect 2234 8351 2246 8385
rect 2280 8351 2319 8385
rect 2353 8351 2392 8385
rect 2426 8351 2465 8385
rect 2499 8351 2538 8385
rect 2572 8351 2611 8385
rect 2234 8313 2611 8351
rect 2234 8279 2246 8313
rect 2280 8279 2319 8313
rect 2353 8279 2392 8313
rect 2426 8279 2465 8313
rect 2499 8279 2538 8313
rect 2572 8279 2611 8313
rect 3221 8279 3233 8457
rect 2234 7584 3233 8279
rect 2234 7532 2983 7584
rect 3035 7532 3047 7584
rect 3099 7532 3111 7584
rect 3163 7532 3175 7584
rect 3227 7532 3233 7584
rect 2234 7401 3233 7532
rect 2234 7367 2246 7401
rect 2280 7367 2319 7401
rect 2353 7367 2392 7401
rect 2426 7367 2465 7401
rect 2499 7367 2538 7401
rect 2572 7367 2611 7401
rect 2234 7329 2611 7367
rect 2234 7295 2246 7329
rect 2280 7295 2319 7329
rect 2353 7295 2392 7329
rect 2426 7295 2465 7329
rect 2499 7295 2538 7329
rect 2572 7295 2611 7329
rect 2234 7257 2611 7295
rect 2234 7223 2246 7257
rect 2280 7223 2319 7257
rect 2353 7223 2392 7257
rect 2426 7223 2465 7257
rect 2499 7223 2538 7257
rect 2572 7223 2611 7257
rect 3221 7223 3233 7401
rect 2234 7207 3233 7223
tri 2178 6789 2206 6817 sw
rect 2048 6782 2206 6789
tri 2206 6782 2213 6789 sw
rect 2048 6751 2213 6782
tri 2213 6751 2244 6782 sw
rect 2048 6717 2244 6751
tri 2244 6717 2278 6751 sw
tri 2045 6710 2048 6713 se
rect 2048 6710 2278 6717
tri 2278 6710 2285 6717 sw
tri 2044 6709 2045 6710 se
rect 2045 6709 2285 6710
tri 2285 6709 2286 6710 sw
tri 2014 6679 2044 6709 se
rect 2044 6679 2286 6709
tri 2286 6679 2316 6709 sw
tri 2010 6675 2014 6679 se
rect 2014 6675 2316 6679
tri 2316 6675 2320 6679 sw
rect 2010 6669 3009 6675
rect 2010 6635 2022 6669
rect 2056 6635 2095 6669
rect 2129 6635 2168 6669
rect 2202 6635 2241 6669
rect 2275 6635 2314 6669
rect 2348 6635 2387 6669
rect 2010 6597 2387 6635
rect 2010 6563 2022 6597
rect 2056 6563 2095 6597
rect 2129 6563 2168 6597
rect 2202 6563 2241 6597
rect 2275 6563 2314 6597
rect 2348 6563 2387 6597
rect 2010 6525 2387 6563
rect 2010 6491 2022 6525
rect 2056 6491 2095 6525
rect 2129 6491 2168 6525
rect 2202 6491 2241 6525
rect 2275 6491 2314 6525
rect 2348 6491 2387 6525
rect 2997 6491 3009 6669
rect 2010 5610 3009 6491
rect 2010 5576 2022 5610
rect 2056 5576 2095 5610
rect 2129 5576 2168 5610
rect 2202 5576 2241 5610
rect 2275 5576 2314 5610
rect 2348 5576 2387 5610
rect 2010 5538 2387 5576
rect 2010 5504 2022 5538
rect 2056 5504 2095 5538
rect 2129 5504 2168 5538
rect 2202 5504 2241 5538
rect 2275 5504 2314 5538
rect 2348 5504 2387 5538
rect 2010 5466 2387 5504
rect 2010 5432 2022 5466
rect 2056 5432 2095 5466
rect 2129 5432 2168 5466
rect 2202 5432 2241 5466
rect 2275 5432 2314 5466
rect 2348 5432 2387 5466
rect 2997 5432 3009 5610
rect 2010 4583 3009 5432
rect 2010 4549 2022 4583
rect 2056 4549 2095 4583
rect 2129 4549 2168 4583
rect 2202 4549 2241 4583
rect 2275 4549 2314 4583
rect 2348 4549 2387 4583
rect 2421 4549 2459 4583
rect 2493 4549 2531 4583
rect 2565 4549 2603 4583
rect 2637 4549 2675 4583
rect 2709 4549 2747 4583
rect 2781 4549 2819 4583
rect 2853 4549 2891 4583
rect 2925 4549 2963 4583
rect 2997 4549 3009 4583
rect 2010 3697 3009 4549
rect 2010 3663 2022 3697
rect 2056 3663 2095 3697
rect 2129 3663 2168 3697
rect 2202 3663 2241 3697
rect 2275 3663 2314 3697
rect 2348 3663 2387 3697
rect 2010 3625 2387 3663
rect 2010 3591 2022 3625
rect 2056 3591 2095 3625
rect 2129 3591 2168 3625
rect 2202 3591 2241 3625
rect 2275 3591 2314 3625
rect 2348 3591 2387 3625
rect 2997 3591 3009 3697
rect 2010 3527 3009 3591
rect 2010 3493 2022 3527
rect 2056 3493 2095 3527
rect 2129 3493 2168 3527
rect 2202 3493 2241 3527
rect 2275 3493 2314 3527
rect 2348 3493 2387 3527
rect 2421 3493 2459 3527
rect 2493 3493 2531 3527
rect 2565 3493 2603 3527
rect 2637 3493 2675 3527
rect 2709 3493 2747 3527
rect 2781 3493 2819 3527
rect 2853 3493 2891 3527
rect 2925 3493 2963 3527
rect 2997 3493 3009 3527
rect 2010 2641 3009 3493
rect 2010 2607 2022 2641
rect 2056 2607 2095 2641
rect 2129 2607 2168 2641
rect 2202 2607 2241 2641
rect 2275 2607 2314 2641
rect 2348 2607 2387 2641
rect 2010 2569 2387 2607
rect 2010 2535 2022 2569
rect 2056 2535 2095 2569
rect 2129 2535 2168 2569
rect 2202 2535 2241 2569
rect 2275 2535 2314 2569
rect 2348 2535 2387 2569
rect 2010 2497 2387 2535
rect 2010 2463 2022 2497
rect 2056 2463 2095 2497
rect 2129 2463 2168 2497
rect 2202 2463 2241 2497
rect 2275 2463 2314 2497
rect 2348 2463 2387 2497
rect 2997 2463 3009 2641
rect 2010 2447 3009 2463
rect 3334 3961 3464 11543
tri 3464 11530 3477 11543 nw
rect 3660 11540 3733 11543
rect 3660 11488 3681 11540
rect 3660 11470 3693 11488
rect 3727 11470 3733 11488
rect 3660 11467 3733 11470
rect 3660 11430 3681 11467
tri 4234 11435 4245 11446 se
rect 4245 11435 4447 12688
rect 4526 14074 4728 14080
rect 4526 14040 4538 14074
rect 4572 14040 4610 14074
rect 4644 14040 4682 14074
rect 4716 14040 4728 14074
rect 4526 13918 4728 14040
rect 4526 13884 4538 13918
rect 4572 13884 4610 13918
rect 4644 13884 4682 13918
rect 4716 13884 4728 13918
rect 4526 13406 4728 13884
rect 4526 13372 4538 13406
rect 4572 13372 4610 13406
rect 4644 13372 4682 13406
rect 4716 13372 4728 13406
rect 4526 13361 4728 13372
rect 4578 13309 4601 13361
rect 4653 13309 4676 13361
rect 4526 13293 4728 13309
rect 4578 13241 4601 13293
rect 4653 13241 4676 13293
rect 4526 13225 4728 13241
rect 4578 13173 4601 13225
rect 4653 13173 4676 13225
rect 4526 13157 4728 13173
rect 4578 13105 4601 13157
rect 4653 13105 4676 13157
rect 4526 13089 4728 13105
rect 4578 13037 4601 13089
rect 4653 13037 4676 13089
rect 4526 12894 4728 13037
rect 4526 12860 4538 12894
rect 4572 12860 4610 12894
rect 4644 12860 4682 12894
rect 4716 12860 4728 12894
rect 4526 12685 4728 12860
tri 4526 12675 4536 12685 ne
rect 4536 12675 4728 12685
tri 4536 12660 4551 12675 ne
rect 4551 12660 4728 12675
tri 4551 12650 4561 12660 ne
rect 4561 12650 4728 12660
rect 4475 12638 4521 12650
rect 4475 12604 4481 12638
rect 4515 12604 4521 12638
tri 4561 12626 4585 12650 ne
rect 4585 12626 4728 12650
tri 4585 12615 4596 12626 ne
rect 4475 12550 4521 12604
rect 4475 12516 4481 12550
rect 4515 12516 4521 12550
rect 4475 12504 4521 12516
tri 4521 12504 4527 12510 sw
rect 4475 12270 4527 12504
rect 4596 12482 4728 12626
rect 4596 12448 4608 12482
rect 4642 12448 4682 12482
rect 4716 12448 4728 12482
rect 4596 12442 4728 12448
rect 4807 14074 6338 14080
rect 4807 14040 6218 14074
rect 6252 14040 6292 14074
rect 6326 14040 6338 14074
rect 4807 14034 6338 14040
rect 4807 14018 5018 14034
tri 5018 14018 5034 14034 nw
rect 4807 13149 5009 14018
tri 5009 14009 5018 14018 nw
tri 6009 14000 6015 14006 se
rect 6015 14000 6149 14006
tri 5975 13966 6009 14000 se
rect 6009 13966 6029 14000
rect 6063 13966 6103 14000
rect 6137 13966 6149 14000
tri 5962 13953 5975 13966 se
rect 5975 13960 6149 13966
rect 5975 13953 6036 13960
tri 6036 13953 6043 13960 nw
rect 5962 13946 6029 13953
tri 6029 13946 6036 13953 nw
rect 5962 13943 6026 13946
tri 6026 13943 6029 13946 nw
rect 5256 13881 5262 13933
rect 5314 13881 5326 13933
rect 5378 13881 5390 13933
rect 5442 13921 5454 13933
rect 5506 13921 5518 13933
rect 5570 13921 5582 13933
rect 5634 13921 5646 13933
rect 5450 13887 5454 13921
rect 5634 13887 5638 13921
rect 5442 13881 5454 13887
rect 5506 13881 5518 13887
rect 5570 13881 5582 13887
rect 5634 13881 5646 13887
rect 5698 13881 5710 13933
rect 5762 13881 5774 13933
rect 5826 13881 5832 13933
rect 4807 13115 4819 13149
rect 4853 13115 4891 13149
rect 4925 13115 4963 13149
rect 4997 13115 5009 13149
rect 4807 13003 5009 13115
rect 4807 12951 4813 13003
rect 4865 12951 4877 13003
rect 4929 12951 4941 13003
rect 4993 12951 5009 13003
rect 4475 12206 4527 12218
rect 4475 12148 4527 12154
rect 4487 11680 4493 11732
rect 4545 11680 4565 11732
rect 4617 11680 4637 11732
rect 4689 11680 4709 11732
rect 4761 11680 4767 11732
tri 3660 11415 3675 11430 ne
rect 3675 11415 3681 11430
tri 3675 11403 3687 11415 ne
rect 3687 11397 3693 11415
rect 3727 11397 3733 11415
rect 3687 11359 3733 11397
tri 4224 11425 4234 11435 se
rect 4234 11425 4447 11435
rect 3687 11325 3693 11359
rect 3727 11325 3733 11359
rect 3687 11287 3733 11325
rect 3687 11253 3693 11287
rect 3727 11253 3733 11287
rect 3500 11228 3552 11240
rect 3500 11194 3506 11228
rect 3540 11194 3552 11228
rect 3500 11154 3552 11194
rect 3500 11120 3506 11154
rect 3540 11120 3552 11154
rect 3500 11080 3552 11120
rect 3500 11046 3506 11080
rect 3540 11046 3552 11080
rect 3500 11006 3552 11046
rect 3500 10972 3506 11006
rect 3540 10972 3552 11006
rect 3500 10932 3552 10972
rect 3500 10898 3506 10932
rect 3540 10898 3552 10932
rect 3500 10858 3552 10898
rect 3500 10824 3506 10858
rect 3540 10824 3552 10858
rect 3500 10784 3552 10824
rect 3500 10750 3506 10784
rect 3540 10750 3552 10784
rect 3500 10710 3552 10750
rect 3500 10676 3506 10710
rect 3540 10676 3552 10710
rect 3500 10636 3552 10676
rect 3500 10602 3506 10636
rect 3540 10602 3552 10636
rect 3500 10561 3552 10602
rect 3500 10527 3506 10561
rect 3540 10527 3552 10561
rect 3500 10486 3552 10527
rect 3500 10452 3506 10486
rect 3540 10452 3552 10486
rect 3500 10142 3552 10452
rect 3687 11215 3733 11253
rect 3687 11181 3693 11215
rect 3727 11181 3733 11215
rect 3687 11143 3733 11181
rect 3687 11109 3693 11143
rect 3727 11109 3733 11143
rect 3687 11071 3733 11109
rect 3687 11037 3693 11071
rect 3727 11037 3733 11071
rect 3687 10999 3733 11037
rect 3687 10965 3693 10999
rect 3727 10965 3733 10999
rect 3687 10927 3733 10965
rect 3687 10893 3693 10927
rect 3727 10893 3733 10927
rect 3687 10855 3733 10893
rect 3687 10821 3693 10855
rect 3727 10821 3733 10855
rect 3687 10783 3733 10821
rect 3687 10749 3693 10783
rect 3727 10749 3733 10783
rect 3687 10711 3733 10749
rect 3687 10677 3693 10711
rect 3727 10677 3733 10711
rect 3687 10639 3733 10677
rect 3687 10605 3693 10639
rect 3727 10605 3733 10639
rect 3687 10567 3733 10605
rect 3687 10533 3693 10567
rect 3727 10533 3733 10567
rect 3687 10495 3733 10533
rect 3687 10461 3693 10495
rect 3727 10461 3733 10495
rect 3687 10423 3733 10461
rect 3687 10389 3693 10423
rect 3727 10389 3733 10423
rect 3687 10351 3733 10389
rect 3687 10317 3693 10351
rect 3727 10317 3733 10351
rect 3687 10279 3733 10317
rect 3500 10108 3506 10142
rect 3540 10108 3552 10142
rect 3500 10068 3552 10108
rect 3500 10034 3506 10068
rect 3540 10034 3552 10068
tri 3681 10249 3687 10255 se
rect 3687 10249 3693 10279
rect 3681 10245 3693 10249
rect 3727 10245 3733 10279
rect 3681 10243 3733 10245
rect 3681 10179 3693 10191
rect 3727 10179 3733 10191
rect 3681 10114 3693 10127
rect 3727 10114 3733 10127
rect 3681 10056 3693 10062
tri 3681 10050 3687 10056 ne
rect 3500 9994 3552 10034
rect 3500 9960 3506 9994
rect 3540 9960 3552 9994
rect 3500 9920 3552 9960
rect 3500 9886 3506 9920
rect 3540 9886 3552 9920
rect 3500 9849 3552 9886
rect 3500 9783 3552 9797
rect 3500 9698 3552 9731
rect 3500 9664 3506 9698
rect 3540 9664 3552 9698
rect 3500 9624 3552 9664
rect 3500 9590 3506 9624
rect 3540 9590 3552 9624
rect 3500 9550 3552 9590
rect 3500 9516 3506 9550
rect 3540 9516 3552 9550
rect 3500 9475 3552 9516
rect 3500 9441 3506 9475
rect 3540 9441 3552 9475
rect 3500 9400 3552 9441
rect 3500 9366 3506 9400
rect 3540 9366 3552 9400
rect 3500 9286 3552 9366
rect 3500 9252 3506 9286
rect 3540 9252 3552 9286
rect 3500 9212 3552 9252
rect 3500 9178 3506 9212
rect 3540 9178 3552 9212
rect 3500 9138 3552 9178
rect 3500 9104 3506 9138
rect 3540 9104 3552 9138
rect 3500 9064 3552 9104
rect 3500 9030 3506 9064
rect 3540 9030 3552 9064
rect 3500 8990 3552 9030
rect 3500 8956 3506 8990
rect 3540 8956 3552 8990
rect 3500 8916 3552 8956
rect 3500 8882 3506 8916
rect 3540 8882 3552 8916
rect 3500 8842 3552 8882
rect 3500 8808 3506 8842
rect 3540 8808 3552 8842
rect 3500 8768 3552 8808
rect 3500 8734 3506 8768
rect 3540 8734 3552 8768
rect 3500 8694 3552 8734
rect 3500 8660 3506 8694
rect 3540 8660 3552 8694
rect 3500 8619 3552 8660
rect 3500 8585 3506 8619
rect 3540 8585 3552 8619
rect 3500 8544 3552 8585
rect 3500 8510 3506 8544
rect 3540 8510 3552 8544
rect 3500 8252 3552 8510
rect 3500 8218 3506 8252
rect 3540 8218 3552 8252
rect 3500 8180 3552 8218
rect 3500 8146 3506 8180
rect 3540 8146 3552 8180
rect 3687 10029 3693 10056
rect 3727 10029 3733 10062
rect 3687 9991 3733 10029
rect 3687 9957 3693 9991
rect 3727 9957 3733 9991
rect 3687 9919 3733 9957
rect 3687 9885 3693 9919
rect 3727 9885 3733 9919
rect 3687 9847 3733 9885
rect 3687 9813 3693 9847
rect 3727 9813 3733 9847
rect 3687 9775 3733 9813
rect 3687 9741 3693 9775
rect 3727 9741 3733 9775
rect 3687 9703 3733 9741
rect 3687 9669 3693 9703
rect 3727 9669 3733 9703
rect 3687 9631 3733 9669
rect 3687 9597 3693 9631
rect 3727 9597 3733 9631
rect 3687 9559 3733 9597
rect 3687 9525 3693 9559
rect 3727 9525 3733 9559
rect 3687 9487 3733 9525
rect 3687 9453 3693 9487
rect 3727 9453 3733 9487
rect 3687 9415 3733 9453
rect 3687 9381 3693 9415
rect 3727 9381 3733 9415
rect 3687 9343 3733 9381
rect 3687 9309 3693 9343
rect 3727 9309 3733 9343
rect 3687 9271 3733 9309
rect 3687 9237 3693 9271
rect 3727 9237 3733 9271
rect 3687 9199 3733 9237
rect 3687 9165 3693 9199
rect 3727 9165 3733 9199
rect 3687 9127 3733 9165
rect 3687 9093 3693 9127
rect 3727 9093 3733 9127
rect 3687 9055 3733 9093
rect 3687 9021 3693 9055
rect 3727 9021 3733 9055
rect 3687 8983 3733 9021
rect 3687 8949 3693 8983
rect 3727 8949 3733 8983
rect 3687 8911 3733 8949
rect 3687 8877 3693 8911
rect 3727 8877 3733 8911
rect 3687 8839 3733 8877
rect 3687 8805 3693 8839
rect 3727 8805 3733 8839
rect 3687 8767 3733 8805
rect 3687 8733 3693 8767
rect 3727 8733 3733 8767
rect 3687 8695 3733 8733
rect 3687 8661 3693 8695
rect 3727 8661 3733 8695
rect 3687 8623 3733 8661
rect 3687 8589 3693 8623
rect 3727 8589 3733 8623
rect 3687 8551 3733 8589
rect 3687 8517 3693 8551
rect 3727 8517 3733 8551
rect 3687 8479 3733 8517
rect 3687 8445 3693 8479
rect 3727 8445 3733 8479
rect 3687 8407 3733 8445
rect 3687 8373 3693 8407
rect 3727 8373 3733 8407
rect 3687 8335 3733 8373
rect 3687 8301 3693 8335
rect 3727 8301 3733 8335
rect 3687 8263 3733 8301
rect 3687 8229 3693 8263
rect 3727 8229 3733 8263
rect 3687 8191 3733 8229
tri 3686 8157 3687 8158 se
rect 3687 8157 3693 8191
rect 3727 8157 3733 8191
tri 3685 8156 3686 8157 se
rect 3686 8156 3733 8157
rect 3500 8108 3552 8146
rect 3500 8074 3506 8108
rect 3540 8074 3552 8108
rect 3500 8036 3552 8074
rect 3500 8002 3506 8036
rect 3540 8002 3552 8036
rect 3500 7964 3552 8002
rect 3500 7930 3506 7964
rect 3540 7930 3552 7964
tri 3681 8152 3685 8156 se
rect 3685 8152 3733 8156
rect 3681 8146 3733 8152
rect 3681 8085 3693 8094
rect 3727 8085 3733 8094
rect 3681 8082 3733 8085
rect 3681 8017 3693 8030
rect 3727 8017 3733 8030
rect 3681 7959 3693 7965
tri 3681 7953 3687 7959 ne
rect 3500 7892 3552 7930
rect 3500 7858 3506 7892
rect 3540 7858 3552 7892
rect 3500 7820 3552 7858
rect 3500 7786 3506 7820
rect 3540 7786 3552 7820
rect 3500 7748 3552 7786
rect 3500 7714 3506 7748
rect 3540 7714 3552 7748
rect 3500 7676 3552 7714
rect 3500 7642 3506 7676
rect 3540 7642 3552 7676
rect 3500 7604 3552 7642
rect 3500 7570 3506 7604
rect 3540 7570 3552 7604
rect 3500 7531 3552 7570
rect 3500 7497 3506 7531
rect 3540 7497 3552 7531
rect 3500 7458 3552 7497
rect 3500 7424 3506 7458
rect 3540 7424 3552 7458
rect 3500 7412 3552 7424
rect 3687 7941 3693 7959
rect 3727 7941 3733 7965
rect 3687 7903 3733 7941
rect 3687 7869 3693 7903
rect 3727 7869 3733 7903
rect 3687 7831 3733 7869
rect 3687 7797 3693 7831
rect 3727 7797 3733 7831
rect 3687 7759 3733 7797
rect 3687 7725 3693 7759
rect 3727 7725 3733 7759
rect 3687 7687 3733 7725
rect 3687 7653 3693 7687
rect 3727 7653 3733 7687
rect 3687 7615 3733 7653
rect 3687 7581 3693 7615
rect 3727 7581 3733 7615
rect 3687 7543 3733 7581
rect 3687 7509 3693 7543
rect 3727 7509 3733 7543
rect 3687 7471 3733 7509
rect 3687 7437 3693 7471
rect 3727 7437 3733 7471
rect 3687 7399 3733 7437
rect 3687 7365 3693 7399
rect 3727 7365 3733 7399
rect 3687 7327 3733 7365
rect 3687 7293 3693 7327
rect 3727 7293 3733 7327
rect 3687 7255 3733 7293
rect 3687 7221 3693 7255
rect 3727 7221 3733 7255
rect 3687 7183 3733 7221
rect 3687 7149 3693 7183
rect 3727 7149 3733 7183
rect 3687 7111 3733 7149
rect 3687 7077 3693 7111
rect 3727 7077 3733 7111
rect 3687 7039 3733 7077
rect 3687 7005 3693 7039
rect 3727 7005 3733 7039
rect 3687 6967 3733 7005
rect 3687 6933 3693 6967
rect 3727 6933 3733 6967
rect 3687 6895 3733 6933
rect 3687 6861 3693 6895
rect 3727 6861 3733 6895
rect 3687 6823 3733 6861
rect 3687 6789 3693 6823
rect 3727 6789 3733 6823
rect 3687 6751 3733 6789
rect 3687 6717 3693 6751
rect 3727 6717 3733 6751
rect 3687 6679 3733 6717
rect 3687 6645 3693 6679
rect 3727 6645 3733 6679
rect 3687 6607 3733 6645
rect 3687 6573 3693 6607
rect 3727 6573 3733 6607
rect 3687 6535 3733 6573
rect 3687 6501 3693 6535
rect 3727 6501 3733 6535
rect 3334 3909 3340 3961
rect 3392 3909 3404 3961
rect 3456 3909 3464 3961
tri 2023 2431 2039 2447 ne
rect 2039 2431 2304 2447
tri 2304 2431 2320 2447 nw
tri 2039 2422 2048 2431 ne
rect 2048 2397 2270 2431
tri 2270 2397 2304 2431 nw
rect 2048 2386 2259 2397
tri 2259 2386 2270 2397 nw
rect 2048 2359 2232 2386
tri 2232 2359 2259 2386 nw
rect 2048 2325 2198 2359
tri 2198 2325 2232 2359 nw
rect 2048 2313 2186 2325
tri 2186 2313 2198 2325 nw
tri 2027 1195 2048 1216 se
rect 2048 1195 2178 2313
tri 2178 2305 2186 2313 nw
tri 2023 1191 2027 1195 se
rect 2027 1191 2178 1195
rect 1933 1185 1984 1191
rect 1933 1121 1984 1133
rect 1933 1063 1984 1069
rect 1985 1064 1986 1190
rect 2022 1064 2023 1190
rect 2024 1063 2178 1191
tri 2023 1046 2040 1063 ne
rect 2040 1046 2178 1063
tri 2040 1040 2046 1046 ne
rect 2046 1040 2178 1046
tri 2046 1038 2048 1040 ne
tri 1658 832 1683 857 sw
rect 1612 826 1762 832
rect 1612 792 1624 826
rect 1658 792 1716 826
rect 1750 792 1762 826
rect 1612 786 1762 792
rect 2048 800 2178 1040
rect 1612 766 1689 786
tri 1689 766 1709 786 nw
rect 2048 766 2060 800
rect 2094 766 2178 800
rect 1612 757 1680 766
tri 1680 757 1689 766 nw
rect 1612 751 1674 757
tri 1674 751 1680 757 nw
rect 1612 744 1667 751
tri 1667 744 1674 751 nw
rect 1117 485 1225 523
rect 1117 451 1185 485
rect 1219 451 1225 485
rect 1117 413 1225 451
rect 1612 482 1658 744
tri 1658 735 1667 744 nw
rect 1782 708 1955 736
rect 1782 674 1794 708
rect 1828 674 1904 708
rect 1938 674 1955 708
rect 1782 636 1955 674
rect 1782 602 1794 636
rect 1828 624 1904 636
rect 1938 624 1955 636
rect 1828 602 1833 624
rect 1782 564 1833 602
rect 1782 530 1794 564
rect 1828 530 1833 564
rect 1782 508 1833 530
rect 1949 508 1955 624
rect 2048 728 2178 766
rect 2048 694 2060 728
rect 2094 694 2178 728
rect 2048 682 2178 694
rect 2048 674 2170 682
tri 2170 674 2178 682 nw
rect 2303 1588 3009 1838
rect 2303 1536 2354 1588
rect 2406 1536 2420 1588
rect 2472 1536 2486 1588
rect 2538 1536 2552 1588
rect 2604 1536 2618 1588
rect 2670 1536 2684 1588
rect 2736 1536 2749 1588
rect 2801 1536 2814 1588
rect 2866 1536 2879 1588
rect 2931 1536 2944 1588
rect 2996 1536 3009 1588
rect 2303 1524 3009 1536
rect 2303 1472 2354 1524
rect 2406 1472 2420 1524
rect 2472 1472 2486 1524
rect 2538 1472 2552 1524
rect 2604 1472 2618 1524
rect 2670 1472 2684 1524
rect 2736 1472 2749 1524
rect 2801 1472 2814 1524
rect 2866 1472 2879 1524
rect 2931 1472 2944 1524
rect 2996 1472 3009 1524
rect 2303 1460 3009 1472
rect 2303 1408 2354 1460
rect 2406 1408 2420 1460
rect 2472 1408 2486 1460
rect 2538 1408 2552 1460
rect 2604 1408 2618 1460
rect 2670 1408 2684 1460
rect 2736 1408 2749 1460
rect 2801 1408 2814 1460
rect 2866 1408 2879 1460
rect 2931 1408 2944 1460
rect 2996 1408 3009 1460
rect 2303 1396 3009 1408
rect 2303 1344 2354 1396
rect 2406 1344 2420 1396
rect 2472 1344 2486 1396
rect 2538 1344 2552 1396
rect 2604 1344 2618 1396
rect 2670 1344 2684 1396
rect 2736 1344 2749 1396
rect 2801 1344 2814 1396
rect 2866 1344 2879 1396
rect 2931 1344 2944 1396
rect 2996 1344 3009 1396
rect 2303 1332 3009 1344
rect 2303 1280 2354 1332
rect 2406 1280 2420 1332
rect 2472 1280 2486 1332
rect 2538 1280 2552 1332
rect 2604 1280 2618 1332
rect 2670 1280 2684 1332
rect 2736 1280 2749 1332
rect 2801 1280 2814 1332
rect 2866 1280 2879 1332
rect 2931 1280 2944 1332
rect 2996 1280 3009 1332
rect 2303 1195 3009 1280
tri 3009 1195 3030 1216 sw
rect 2303 1191 3030 1195
tri 3030 1191 3034 1195 sw
rect 2303 1063 3033 1191
rect 3035 1190 3071 1191
rect 3034 1064 3072 1190
rect 3073 1185 3125 1191
rect 3073 1121 3125 1133
rect 3035 1063 3071 1064
rect 3073 1063 3125 1069
rect 2303 1046 3017 1063
tri 3017 1046 3034 1063 nw
rect 2303 1040 3011 1046
tri 3011 1040 3017 1046 nw
rect 2303 899 3009 1040
tri 3009 1038 3011 1040 nw
rect 3334 1007 3464 3909
rect 3500 6474 3552 6480
rect 3500 6408 3552 6422
rect 3500 6320 3552 6356
rect 3500 6286 3506 6320
rect 3540 6286 3552 6320
rect 3500 6246 3552 6286
rect 3500 6212 3506 6246
rect 3540 6212 3552 6246
rect 3500 6172 3552 6212
rect 3500 6138 3506 6172
rect 3540 6138 3552 6172
rect 3500 6098 3552 6138
rect 3500 6064 3506 6098
rect 3540 6064 3552 6098
rect 3500 6024 3552 6064
rect 3500 5990 3506 6024
rect 3540 5990 3552 6024
rect 3500 5950 3552 5990
rect 3500 5916 3506 5950
rect 3540 5916 3552 5950
rect 3500 5876 3552 5916
rect 3500 5842 3506 5876
rect 3540 5842 3552 5876
rect 3500 5801 3552 5842
rect 3500 5767 3506 5801
rect 3540 5767 3552 5801
rect 3500 5726 3552 5767
rect 3500 5692 3506 5726
rect 3540 5692 3552 5726
rect 3500 5382 3552 5692
rect 3500 5348 3506 5382
rect 3540 5348 3552 5382
rect 3500 5308 3552 5348
rect 3500 5274 3506 5308
rect 3540 5274 3552 5308
rect 3500 5234 3552 5274
rect 3500 5200 3506 5234
rect 3540 5200 3552 5234
rect 3500 5160 3552 5200
rect 3500 5126 3506 5160
rect 3540 5126 3552 5160
rect 3500 5086 3552 5126
rect 3500 5052 3506 5086
rect 3540 5052 3552 5086
rect 3500 5012 3552 5052
rect 3500 4978 3506 5012
rect 3540 4978 3552 5012
rect 3500 4938 3552 4978
rect 3500 4904 3506 4938
rect 3540 4904 3552 4938
rect 3500 4864 3552 4904
rect 3687 6463 3733 6501
rect 3687 6429 3693 6463
rect 3727 6429 3733 6463
rect 3687 6391 3733 6429
rect 3687 6357 3693 6391
rect 3727 6357 3733 6391
rect 3687 6319 3733 6357
rect 3687 6285 3693 6319
rect 3727 6285 3733 6319
rect 3687 6247 3733 6285
rect 3687 6213 3693 6247
rect 3727 6213 3733 6247
rect 3687 6175 3733 6213
rect 3687 6141 3693 6175
rect 3727 6141 3733 6175
rect 3687 6103 3733 6141
rect 3687 6069 3693 6103
rect 3727 6069 3733 6103
rect 3687 6031 3733 6069
rect 3687 5997 3693 6031
rect 3727 5997 3733 6031
rect 3687 5959 3733 5997
rect 3687 5925 3693 5959
rect 3727 5925 3733 5959
rect 3687 5887 3733 5925
rect 3687 5853 3693 5887
rect 3727 5853 3733 5887
rect 3687 5815 3733 5853
rect 3687 5781 3693 5815
rect 3727 5781 3733 5815
rect 3687 5743 3733 5781
rect 3687 5709 3693 5743
rect 3727 5709 3733 5743
rect 3687 5671 3733 5709
rect 3687 5637 3693 5671
rect 3727 5637 3733 5671
rect 3687 5599 3733 5637
rect 3687 5565 3693 5599
rect 3727 5565 3733 5599
rect 3687 5527 3733 5565
rect 3687 5493 3693 5527
rect 3727 5493 3733 5527
rect 3687 5455 3733 5493
rect 3687 5421 3693 5455
rect 3727 5421 3733 5455
rect 3687 5383 3733 5421
rect 3687 5349 3693 5383
rect 3727 5349 3733 5383
rect 3687 5311 3733 5349
rect 3687 5277 3693 5311
rect 3727 5277 3733 5311
rect 3687 5239 3733 5277
rect 3687 5205 3693 5239
rect 3727 5205 3733 5239
rect 3687 5167 3733 5205
rect 3687 5133 3693 5167
rect 3727 5133 3733 5167
rect 3687 5095 3733 5133
rect 3687 5061 3693 5095
rect 3727 5061 3733 5095
rect 3687 5023 3733 5061
rect 3687 4989 3693 5023
rect 3727 4989 3733 5023
rect 3687 4951 3733 4989
rect 3687 4917 3693 4951
rect 3727 4917 3733 4951
rect 3500 4830 3506 4864
rect 3540 4830 3552 4864
rect 3500 4790 3552 4830
rect 3500 4756 3506 4790
rect 3540 4756 3552 4790
rect 3500 4715 3552 4756
tri 3681 4886 3687 4892 se
rect 3687 4886 3733 4917
rect 3681 4880 3733 4886
rect 3681 4814 3733 4828
rect 3681 4756 3733 4762
tri 3681 4750 3687 4756 ne
rect 3500 4681 3506 4715
rect 3540 4681 3552 4715
rect 3500 4640 3552 4681
rect 3500 4606 3506 4640
rect 3540 4606 3552 4640
rect 3500 4526 3552 4606
rect 3500 4492 3506 4526
rect 3540 4492 3552 4526
rect 3500 4452 3552 4492
rect 3500 4418 3506 4452
rect 3540 4418 3552 4452
rect 3500 4378 3552 4418
rect 3500 4344 3506 4378
rect 3540 4344 3552 4378
rect 3500 4304 3552 4344
rect 3500 4270 3506 4304
rect 3540 4270 3552 4304
rect 3500 4230 3552 4270
rect 3500 4196 3506 4230
rect 3540 4196 3552 4230
rect 3500 4156 3552 4196
rect 3500 4122 3506 4156
rect 3540 4122 3552 4156
rect 3500 4082 3552 4122
rect 3500 4048 3506 4082
rect 3540 4048 3552 4082
rect 3500 4008 3552 4048
rect 3500 3974 3506 4008
rect 3540 3974 3552 4008
rect 3500 3934 3552 3974
rect 3500 3900 3506 3934
rect 3540 3900 3552 3934
rect 3500 3859 3552 3900
rect 3500 3825 3506 3859
rect 3540 3825 3552 3859
rect 3500 3784 3552 3825
rect 3500 3750 3506 3784
rect 3540 3750 3552 3784
rect 3500 3440 3552 3750
rect 3500 3406 3506 3440
rect 3540 3406 3552 3440
rect 3500 3366 3552 3406
rect 3500 3332 3506 3366
rect 3540 3332 3552 3366
rect 3500 3292 3552 3332
rect 3500 3258 3506 3292
rect 3540 3258 3552 3292
rect 3500 3218 3552 3258
rect 3500 3184 3506 3218
rect 3540 3184 3552 3218
rect 3500 3144 3552 3184
rect 3500 3110 3506 3144
rect 3540 3110 3552 3144
rect 3500 3070 3552 3110
rect 3500 3036 3506 3070
rect 3540 3036 3552 3070
rect 3500 2996 3552 3036
rect 3500 2962 3506 2996
rect 3540 2962 3552 2996
rect 3500 2922 3552 2962
rect 3500 2888 3506 2922
rect 3540 2888 3552 2922
rect 3500 2848 3552 2888
rect 3500 2814 3506 2848
rect 3540 2814 3552 2848
rect 3500 2773 3552 2814
rect 3500 2739 3506 2773
rect 3540 2739 3552 2773
rect 3500 2698 3552 2739
rect 3500 2664 3506 2698
rect 3540 2664 3552 2698
rect 3500 2652 3552 2664
rect 3687 4735 3733 4756
rect 3687 4701 3693 4735
rect 3727 4701 3733 4735
rect 3687 4663 3733 4701
rect 3687 4629 3693 4663
rect 3727 4629 3733 4663
rect 3687 4591 3733 4629
rect 3687 4557 3693 4591
rect 3727 4557 3733 4591
rect 3687 4519 3733 4557
rect 3687 4485 3693 4519
rect 3727 4485 3733 4519
rect 3687 4447 3733 4485
rect 3687 4413 3693 4447
rect 3727 4413 3733 4447
rect 3687 4375 3733 4413
rect 3687 4341 3693 4375
rect 3727 4341 3733 4375
rect 3687 4303 3733 4341
rect 3687 4269 3693 4303
rect 3727 4269 3733 4303
rect 3687 4231 3733 4269
rect 3687 4197 3693 4231
rect 3727 4197 3733 4231
rect 3687 4159 3733 4197
rect 3687 4125 3693 4159
rect 3727 4125 3733 4159
rect 3687 4087 3733 4125
rect 3687 4053 3693 4087
rect 3727 4053 3733 4087
rect 3687 4015 3733 4053
rect 3687 3981 3693 4015
rect 3727 3981 3733 4015
rect 3687 3943 3733 3981
rect 3687 3909 3693 3943
rect 3727 3909 3733 3943
rect 3687 3871 3733 3909
rect 3687 3837 3693 3871
rect 3727 3837 3733 3871
rect 3687 3799 3733 3837
rect 3687 3765 3693 3799
rect 3727 3765 3733 3799
rect 3687 3727 3733 3765
rect 3687 3693 3693 3727
rect 3727 3693 3733 3727
rect 3687 3655 3733 3693
rect 3687 3621 3693 3655
rect 3727 3621 3733 3655
rect 3687 3583 3733 3621
rect 3687 3549 3693 3583
rect 3727 3549 3733 3583
rect 3687 3511 3733 3549
rect 3687 3477 3693 3511
rect 3727 3477 3733 3511
rect 3687 3439 3733 3477
rect 3687 3405 3693 3439
rect 3727 3405 3733 3439
rect 3687 3367 3733 3405
rect 3687 3333 3693 3367
rect 3727 3333 3733 3367
rect 3687 3295 3733 3333
rect 3687 3261 3693 3295
rect 3727 3261 3733 3295
rect 3687 3223 3733 3261
rect 3687 3189 3693 3223
rect 3727 3189 3733 3223
rect 3687 3151 3733 3189
rect 3687 3117 3693 3151
rect 3727 3117 3733 3151
rect 3687 3079 3733 3117
rect 3687 3045 3693 3079
rect 3727 3045 3733 3079
rect 3687 3007 3733 3045
rect 3687 2973 3693 3007
rect 3727 2973 3733 3007
rect 3687 2935 3733 2973
rect 3687 2901 3693 2935
rect 3727 2901 3733 2935
rect 3687 2863 3733 2901
rect 3687 2829 3693 2863
rect 3727 2829 3733 2863
rect 3687 2791 3733 2829
rect 3687 2757 3693 2791
rect 3727 2757 3733 2791
rect 3687 2719 3733 2757
rect 3687 2685 3693 2719
rect 3727 2685 3733 2719
rect 3687 2647 3733 2685
rect 3687 2613 3693 2647
rect 3727 2613 3733 2647
rect 3687 2575 3733 2613
rect 3687 2541 3693 2575
rect 3727 2541 3733 2575
rect 3687 2503 3733 2541
rect 3687 2469 3693 2503
rect 3727 2469 3733 2503
rect 3687 2431 3733 2469
rect 3687 2397 3693 2431
rect 3727 2397 3733 2431
rect 3687 2359 3733 2397
rect 3687 2325 3693 2359
rect 3727 2325 3733 2359
rect 3687 2287 3733 2325
rect 3687 2253 3693 2287
rect 3727 2253 3733 2287
rect 3687 2215 3733 2253
rect 3687 2181 3693 2215
rect 3727 2181 3733 2215
rect 3687 2169 3733 2181
rect 3761 7341 3928 11368
rect 3930 11367 3966 11368
rect 3761 7161 3768 7341
rect 3884 7161 3928 7341
rect 3761 6819 3928 7161
rect 3761 6639 3768 6819
rect 3884 6639 3928 6819
rect 3761 5638 3928 6639
rect 3761 5458 3768 5638
rect 3884 5458 3928 5638
rect 3761 4203 3928 5458
rect 3761 4023 3768 4203
rect 3884 4023 3928 4203
rect 3761 3930 3928 4023
rect 3929 3931 3967 11367
rect 3968 11362 4196 11368
rect 3968 11328 4038 11362
rect 4072 11328 4150 11362
rect 4184 11328 4196 11362
rect 3968 11322 4196 11328
rect 4224 11362 4447 11425
rect 3968 11252 4040 11322
tri 4040 11297 4065 11322 nw
rect 3968 11218 4000 11252
rect 4034 11218 4040 11252
rect 3968 11180 4040 11218
rect 3968 11146 4000 11180
rect 4034 11146 4040 11180
rect 3968 11108 4040 11146
rect 3968 11074 4000 11108
rect 4034 11074 4040 11108
rect 3968 11036 4040 11074
rect 3968 11002 4000 11036
rect 4034 11002 4040 11036
rect 3968 10964 4040 11002
rect 3968 10930 4000 10964
rect 4034 10930 4040 10964
rect 3968 10892 4040 10930
rect 3968 10858 4000 10892
rect 4034 10858 4040 10892
rect 3968 10820 4040 10858
rect 3968 10786 4000 10820
rect 4034 10786 4040 10820
rect 3968 10748 4040 10786
rect 3968 10714 4000 10748
rect 4034 10714 4040 10748
rect 3968 10676 4040 10714
rect 3968 10642 4000 10676
rect 4034 10642 4040 10676
rect 3968 10604 4040 10642
rect 3968 10570 4000 10604
rect 4034 10570 4040 10604
rect 3968 10532 4040 10570
rect 3968 10498 4000 10532
rect 4034 10498 4040 10532
rect 3968 10460 4040 10498
rect 3968 10426 4000 10460
rect 4034 10426 4040 10460
rect 3968 10388 4040 10426
rect 3968 10354 4000 10388
rect 4034 10354 4040 10388
rect 3968 10316 4040 10354
rect 3968 10282 4000 10316
rect 4034 10282 4040 10316
rect 3968 10244 4040 10282
rect 3968 10210 4000 10244
rect 4034 10210 4040 10244
rect 3968 10172 4040 10210
rect 3968 10138 4000 10172
rect 4034 10138 4040 10172
rect 3968 10100 4040 10138
rect 3968 10066 4000 10100
rect 4034 10066 4040 10100
rect 3968 10028 4040 10066
rect 3968 9994 4000 10028
rect 4034 9994 4040 10028
rect 3968 9956 4040 9994
rect 3968 9922 4000 9956
rect 4034 9922 4040 9956
rect 3968 9884 4040 9922
rect 3968 9850 4000 9884
rect 4034 9850 4040 9884
rect 3968 9812 4040 9850
rect 3968 9778 4000 9812
rect 4034 9778 4040 9812
rect 3968 9740 4040 9778
rect 3968 9706 4000 9740
rect 4034 9706 4040 9740
rect 3968 9668 4040 9706
rect 3968 9634 4000 9668
rect 4034 9634 4040 9668
rect 3968 9596 4040 9634
rect 3968 9562 4000 9596
rect 4034 9562 4040 9596
rect 3968 9524 4040 9562
rect 3968 9490 4000 9524
rect 4034 9490 4040 9524
rect 3968 9452 4040 9490
rect 3968 9418 4000 9452
rect 4034 9418 4040 9452
rect 3968 9380 4040 9418
rect 3968 9346 4000 9380
rect 4034 9346 4040 9380
rect 3968 9308 4040 9346
rect 3968 9274 4000 9308
rect 4034 9274 4040 9308
rect 3968 9236 4040 9274
rect 3968 9202 4000 9236
rect 4034 9202 4040 9236
rect 3968 9164 4040 9202
rect 3968 9130 4000 9164
rect 4034 9130 4040 9164
rect 3968 9092 4040 9130
rect 3968 9058 4000 9092
rect 4034 9058 4040 9092
rect 3968 9020 4040 9058
rect 3968 8986 4000 9020
rect 4034 8986 4040 9020
rect 3968 8948 4040 8986
rect 3968 8914 4000 8948
rect 4034 8914 4040 8948
rect 3968 8876 4040 8914
rect 3968 8842 4000 8876
rect 4034 8842 4040 8876
rect 3968 8804 4040 8842
rect 3968 8770 4000 8804
rect 4034 8770 4040 8804
rect 3968 8732 4040 8770
rect 3968 8698 4000 8732
rect 4034 8698 4040 8732
rect 3968 8660 4040 8698
rect 3968 8626 4000 8660
rect 4034 8626 4040 8660
rect 3968 8588 4040 8626
rect 3968 8554 4000 8588
rect 4034 8554 4040 8588
rect 3968 8516 4040 8554
rect 3968 8482 4000 8516
rect 4034 8482 4040 8516
rect 3968 8444 4040 8482
rect 3968 8410 4000 8444
rect 4034 8410 4040 8444
rect 3968 8372 4040 8410
rect 3968 8338 4000 8372
rect 4034 8338 4040 8372
rect 3968 8300 4040 8338
rect 3968 8266 4000 8300
rect 4034 8266 4040 8300
rect 3968 8228 4040 8266
rect 3968 8194 4000 8228
rect 4034 8194 4040 8228
rect 3968 8156 4040 8194
rect 3968 8122 4000 8156
rect 4034 8122 4040 8156
rect 3968 8084 4040 8122
rect 3968 8050 4000 8084
rect 4034 8050 4040 8084
rect 3968 8012 4040 8050
rect 3968 7978 4000 8012
rect 4034 7978 4040 8012
rect 3968 7940 4040 7978
rect 3968 7906 4000 7940
rect 4034 7906 4040 7940
rect 3968 7868 4040 7906
rect 3968 7834 4000 7868
rect 4034 7834 4040 7868
rect 3968 7796 4040 7834
rect 3968 7762 4000 7796
rect 4034 7762 4040 7796
rect 3968 7724 4040 7762
rect 3968 7690 4000 7724
rect 4034 7690 4040 7724
rect 3968 7652 4040 7690
rect 3968 7618 4000 7652
rect 4034 7618 4040 7652
rect 3968 7580 4040 7618
rect 3968 7546 4000 7580
rect 4034 7546 4040 7580
rect 3968 7508 4040 7546
rect 3968 7474 4000 7508
rect 4034 7474 4040 7508
rect 3968 7436 4040 7474
rect 3968 7402 4000 7436
rect 4034 7402 4040 7436
rect 3968 7364 4040 7402
rect 3968 7330 4000 7364
rect 4034 7330 4040 7364
rect 3968 7292 4040 7330
rect 3968 7258 4000 7292
rect 4034 7258 4040 7292
rect 3968 7220 4040 7258
rect 3968 7186 4000 7220
rect 4034 7186 4040 7220
rect 3968 7147 4040 7186
rect 3968 7113 4000 7147
rect 4034 7113 4040 7147
rect 3968 7074 4040 7113
rect 3968 7040 4000 7074
rect 4034 7040 4040 7074
rect 3968 7001 4040 7040
rect 3968 6967 4000 7001
rect 4034 6967 4040 7001
rect 3968 6928 4040 6967
rect 3968 6894 4000 6928
rect 4034 6894 4040 6928
rect 3968 6855 4040 6894
rect 3968 6821 4000 6855
rect 4034 6821 4040 6855
rect 3968 6782 4040 6821
rect 3968 6748 4000 6782
rect 4034 6748 4040 6782
rect 3968 6709 4040 6748
rect 3968 6675 4000 6709
rect 4034 6675 4040 6709
rect 3968 6636 4040 6675
rect 3968 6602 4000 6636
rect 4034 6602 4040 6636
rect 3968 6563 4040 6602
rect 3968 6529 4000 6563
rect 4034 6529 4040 6563
rect 3968 6490 4040 6529
rect 3968 6456 4000 6490
rect 4034 6456 4040 6490
rect 3968 6417 4040 6456
rect 3968 6383 4000 6417
rect 4034 6383 4040 6417
rect 3968 6344 4040 6383
rect 3968 6310 4000 6344
rect 4034 6310 4040 6344
rect 3968 6271 4040 6310
rect 3968 6237 4000 6271
rect 4034 6237 4040 6271
rect 3968 6198 4040 6237
rect 3968 6164 4000 6198
rect 4034 6164 4040 6198
rect 3968 6125 4040 6164
rect 3968 6091 4000 6125
rect 4034 6091 4040 6125
rect 3968 6052 4040 6091
rect 3968 6018 4000 6052
rect 4034 6018 4040 6052
rect 3968 5979 4040 6018
rect 3968 5945 4000 5979
rect 4034 5945 4040 5979
rect 3968 5906 4040 5945
rect 3968 5872 4000 5906
rect 4034 5872 4040 5906
rect 3968 5833 4040 5872
rect 3968 5799 4000 5833
rect 4034 5799 4040 5833
rect 3968 5760 4040 5799
rect 3968 5726 4000 5760
rect 4034 5726 4040 5760
rect 3968 5687 4040 5726
rect 3968 5653 4000 5687
rect 4034 5653 4040 5687
rect 3968 5614 4040 5653
rect 3968 5580 4000 5614
rect 4034 5580 4040 5614
rect 3968 5541 4040 5580
rect 3968 5507 4000 5541
rect 4034 5507 4040 5541
rect 3968 5468 4040 5507
rect 3968 5434 4000 5468
rect 4034 5434 4040 5468
rect 3968 5395 4040 5434
rect 3968 5361 4000 5395
rect 4034 5361 4040 5395
rect 3968 5322 4040 5361
rect 3968 5288 4000 5322
rect 4034 5288 4040 5322
rect 3968 5249 4040 5288
rect 3968 5215 4000 5249
rect 4034 5215 4040 5249
rect 3968 5176 4040 5215
rect 3968 5142 4000 5176
rect 4034 5142 4040 5176
rect 3968 5103 4040 5142
rect 3968 5069 4000 5103
rect 4034 5069 4040 5103
rect 3968 5030 4040 5069
rect 3968 4996 4000 5030
rect 4034 4996 4040 5030
rect 3968 4957 4040 4996
rect 3968 4923 4000 4957
rect 4034 4923 4040 4957
rect 3968 4884 4040 4923
rect 3968 4850 4000 4884
rect 4034 4850 4040 4884
rect 3968 4811 4040 4850
rect 3968 4777 4000 4811
rect 4034 4777 4040 4811
rect 3968 4738 4040 4777
rect 3968 4704 4000 4738
rect 4034 4704 4040 4738
rect 3968 4665 4040 4704
rect 3968 4631 4000 4665
rect 4034 4631 4040 4665
rect 3968 4592 4040 4631
rect 3968 4558 4000 4592
rect 4034 4558 4040 4592
rect 3968 4519 4040 4558
rect 3968 4485 4000 4519
rect 4034 4485 4040 4519
rect 3968 4446 4040 4485
rect 3968 4412 4000 4446
rect 4034 4412 4040 4446
rect 3968 4373 4040 4412
rect 3968 4339 4000 4373
rect 4034 4339 4040 4373
rect 3968 4300 4040 4339
rect 3968 4266 4000 4300
rect 4034 4266 4040 4300
rect 3968 4227 4040 4266
rect 4070 9321 4122 11045
rect 4070 9287 4082 9321
rect 4116 9287 4122 9321
rect 4070 9247 4122 9287
rect 4070 9213 4082 9247
rect 4116 9213 4122 9247
rect 4070 9173 4122 9213
rect 4070 9139 4082 9173
rect 4116 9139 4122 9173
rect 4070 9099 4122 9139
rect 4070 9065 4082 9099
rect 4116 9065 4122 9099
rect 4070 9025 4122 9065
rect 4070 8991 4082 9025
rect 4116 8991 4122 9025
rect 4070 8983 4122 8991
rect 4070 8917 4082 8931
rect 4116 8917 4122 8931
rect 4070 8843 4082 8865
rect 4116 8843 4122 8865
rect 4070 8803 4122 8843
rect 4070 8769 4082 8803
rect 4116 8769 4122 8803
rect 4070 8729 4122 8769
rect 4070 8695 4082 8729
rect 4116 8695 4122 8729
rect 4070 8654 4122 8695
rect 4070 8620 4082 8654
rect 4116 8620 4122 8654
rect 4070 8579 4122 8620
rect 4070 8545 4082 8579
rect 4116 8545 4122 8579
rect 4070 8465 4122 8545
rect 4070 8431 4082 8465
rect 4116 8431 4122 8465
rect 4070 8391 4122 8431
rect 4070 8357 4082 8391
rect 4116 8357 4122 8391
rect 4070 8317 4122 8357
rect 4070 8283 4082 8317
rect 4116 8283 4122 8317
rect 4070 8243 4122 8283
rect 4070 8209 4082 8243
rect 4116 8209 4122 8243
rect 4070 8169 4122 8209
rect 4070 8135 4082 8169
rect 4116 8135 4122 8169
rect 4070 8095 4122 8135
rect 4070 8061 4082 8095
rect 4116 8061 4122 8095
rect 4070 8021 4122 8061
rect 4070 7987 4082 8021
rect 4116 7987 4122 8021
rect 4070 7947 4122 7987
rect 4070 7913 4082 7947
rect 4116 7913 4122 7947
rect 4070 7873 4122 7913
rect 4070 7839 4082 7873
rect 4116 7839 4122 7873
rect 4070 7798 4122 7839
rect 4070 7764 4082 7798
rect 4116 7764 4122 7798
rect 4070 7723 4122 7764
rect 4070 7689 4082 7723
rect 4116 7689 4122 7723
rect 4070 5897 4122 7689
rect 4070 5863 4082 5897
rect 4116 5863 4122 5897
rect 4070 5823 4122 5863
rect 4070 5789 4082 5823
rect 4116 5789 4122 5823
rect 4070 5749 4122 5789
rect 4070 5715 4082 5749
rect 4116 5715 4122 5749
rect 4070 5675 4122 5715
rect 4070 5641 4082 5675
rect 4116 5641 4122 5675
rect 4070 5601 4122 5641
rect 4070 5567 4082 5601
rect 4116 5567 4122 5601
rect 4070 5527 4122 5567
rect 4070 5493 4082 5527
rect 4116 5493 4122 5527
rect 4070 5453 4122 5493
rect 4070 5419 4082 5453
rect 4116 5419 4122 5453
rect 4070 5379 4122 5419
rect 4070 5345 4082 5379
rect 4116 5345 4122 5379
rect 4070 5305 4122 5345
rect 4070 5282 4082 5305
rect 4116 5282 4122 5305
rect 4070 5216 4082 5230
rect 4116 5216 4122 5230
rect 4070 5155 4122 5164
rect 4070 5121 4082 5155
rect 4116 5121 4122 5155
rect 4070 5041 4122 5121
rect 4070 5007 4082 5041
rect 4116 5007 4122 5041
rect 4070 4967 4122 5007
rect 4070 4933 4082 4967
rect 4116 4933 4122 4967
rect 4070 4893 4122 4933
rect 4070 4859 4082 4893
rect 4116 4859 4122 4893
rect 4070 4819 4122 4859
rect 4070 4785 4082 4819
rect 4116 4785 4122 4819
rect 4070 4745 4122 4785
rect 4070 4711 4082 4745
rect 4116 4711 4122 4745
rect 4070 4671 4122 4711
rect 4070 4637 4082 4671
rect 4116 4637 4122 4671
rect 4070 4597 4122 4637
rect 4070 4563 4082 4597
rect 4116 4563 4122 4597
rect 4070 4523 4122 4563
rect 4070 4489 4082 4523
rect 4116 4489 4122 4523
rect 4070 4449 4122 4489
rect 4070 4415 4082 4449
rect 4116 4415 4122 4449
rect 4070 4374 4122 4415
rect 4070 4340 4082 4374
rect 4116 4340 4122 4374
rect 4070 4299 4122 4340
rect 4070 4265 4082 4299
rect 4116 4265 4122 4299
rect 4070 4249 4122 4265
rect 4224 8522 4426 11362
tri 4426 11341 4447 11362 nw
rect 4807 11435 5009 12951
rect 5215 13835 5267 13841
rect 5215 13767 5267 13783
rect 5215 13699 5267 13715
rect 5215 13643 5224 13647
rect 5258 13643 5267 13647
rect 5215 13631 5267 13643
rect 5215 13568 5224 13579
rect 5258 13568 5267 13579
rect 5215 13563 5267 13568
rect 5215 13493 5224 13511
rect 5258 13493 5267 13511
rect 5215 13452 5267 13493
rect 5215 13418 5224 13452
rect 5258 13418 5267 13452
rect 5215 13377 5267 13418
rect 5215 13343 5224 13377
rect 5258 13343 5267 13377
rect 5215 13302 5267 13343
rect 5215 13268 5224 13302
rect 5258 13268 5267 13302
rect 5215 13227 5267 13268
rect 5215 13193 5224 13227
rect 5258 13193 5267 13227
rect 5215 13152 5267 13193
rect 5215 13118 5224 13152
rect 5258 13118 5267 13152
rect 5215 13077 5267 13118
rect 5215 13043 5224 13077
rect 5258 13043 5267 13077
rect 5215 13002 5267 13043
rect 5215 12968 5224 13002
rect 5258 12968 5267 13002
rect 5215 12927 5267 12968
rect 5215 12893 5224 12927
rect 5258 12893 5267 12927
rect 5215 12881 5267 12893
rect 5371 13827 5423 13839
rect 5371 13793 5380 13827
rect 5414 13793 5423 13827
rect 5371 13752 5423 13793
rect 5371 13718 5380 13752
rect 5414 13718 5423 13752
rect 5371 13677 5423 13718
rect 5371 13643 5380 13677
rect 5414 13643 5423 13677
rect 5371 13602 5423 13643
rect 5371 13568 5380 13602
rect 5414 13568 5423 13602
rect 5371 13527 5423 13568
rect 5371 13493 5380 13527
rect 5414 13493 5423 13527
rect 5371 13452 5423 13493
rect 5371 13418 5380 13452
rect 5414 13418 5423 13452
rect 5371 13377 5423 13418
rect 5371 13361 5380 13377
rect 5414 13361 5423 13377
rect 5371 13302 5423 13309
rect 5371 13293 5380 13302
rect 5414 13293 5423 13302
rect 5371 13227 5423 13241
rect 5371 13225 5380 13227
rect 5414 13225 5423 13227
rect 5371 13157 5423 13173
rect 5371 13089 5423 13105
rect 5371 13002 5423 13037
rect 5371 12968 5380 13002
rect 5414 12968 5423 13002
rect 5371 12927 5423 12968
rect 5371 12893 5380 12927
rect 5414 12893 5423 12927
rect 5371 12881 5423 12893
rect 5527 13835 5579 13841
rect 5527 13767 5579 13783
rect 5527 13699 5579 13715
rect 5527 13643 5536 13647
rect 5570 13643 5579 13647
rect 5527 13631 5579 13643
rect 5527 13568 5536 13579
rect 5570 13568 5579 13579
rect 5527 13563 5579 13568
rect 5527 13493 5536 13511
rect 5570 13493 5579 13511
rect 5527 13452 5579 13493
rect 5527 13418 5536 13452
rect 5570 13418 5579 13452
rect 5527 13377 5579 13418
rect 5527 13343 5536 13377
rect 5570 13343 5579 13377
rect 5527 13302 5579 13343
rect 5527 13268 5536 13302
rect 5570 13268 5579 13302
rect 5527 13227 5579 13268
rect 5527 13193 5536 13227
rect 5570 13193 5579 13227
rect 5527 13152 5579 13193
rect 5527 13118 5536 13152
rect 5570 13118 5579 13152
rect 5527 13077 5579 13118
rect 5527 13043 5536 13077
rect 5570 13043 5579 13077
rect 5527 13002 5579 13043
rect 5527 12968 5536 13002
rect 5570 12968 5579 13002
rect 5527 12927 5579 12968
rect 5527 12893 5536 12927
rect 5570 12893 5579 12927
rect 5527 12881 5579 12893
rect 5683 13827 5735 13839
rect 5683 13793 5692 13827
rect 5726 13793 5735 13827
rect 5683 13752 5735 13793
rect 5683 13718 5692 13752
rect 5726 13718 5735 13752
rect 5683 13677 5735 13718
rect 5683 13643 5692 13677
rect 5726 13643 5735 13677
rect 5683 13602 5735 13643
rect 5683 13568 5692 13602
rect 5726 13568 5735 13602
rect 5683 13527 5735 13568
rect 5683 13493 5692 13527
rect 5726 13493 5735 13527
rect 5683 13452 5735 13493
rect 5683 13418 5692 13452
rect 5726 13418 5735 13452
rect 5683 13377 5735 13418
rect 5683 13361 5692 13377
rect 5726 13361 5735 13377
rect 5683 13302 5735 13309
rect 5683 13293 5692 13302
rect 5726 13293 5735 13302
rect 5683 13227 5735 13241
rect 5683 13225 5692 13227
rect 5726 13225 5735 13227
rect 5683 13157 5735 13173
rect 5683 13089 5735 13105
rect 5683 13002 5735 13037
rect 5683 12968 5692 13002
rect 5726 12968 5735 13002
rect 5683 12927 5735 12968
rect 5683 12893 5692 12927
rect 5726 12893 5735 12927
rect 5683 12881 5735 12893
rect 5839 13835 5891 13841
rect 5839 13767 5891 13783
rect 5839 13699 5891 13715
rect 5839 13643 5848 13647
rect 5882 13643 5891 13647
rect 5839 13631 5891 13643
rect 5839 13568 5848 13579
rect 5882 13568 5891 13579
rect 5839 13563 5891 13568
rect 5839 13493 5848 13511
rect 5882 13493 5891 13511
rect 5839 13452 5891 13493
rect 5839 13418 5848 13452
rect 5882 13418 5891 13452
rect 5839 13377 5891 13418
rect 5839 13343 5848 13377
rect 5882 13343 5891 13377
rect 5839 13302 5891 13343
rect 5839 13268 5848 13302
rect 5882 13268 5891 13302
rect 5839 13227 5891 13268
rect 5839 13193 5848 13227
rect 5882 13193 5891 13227
rect 5839 13152 5891 13193
rect 5839 13118 5848 13152
rect 5882 13118 5891 13152
rect 5839 13077 5891 13118
rect 5839 13043 5848 13077
rect 5882 13043 5891 13077
rect 5839 13002 5891 13043
rect 5839 12968 5848 13002
rect 5882 12968 5891 13002
rect 5839 12927 5891 12968
rect 5839 12893 5848 12927
rect 5882 12893 5891 12927
tri 5830 12688 5839 12697 se
rect 5839 12688 5891 12893
tri 5817 12675 5830 12688 se
rect 5830 12675 5891 12688
tri 5814 12672 5817 12675 se
rect 5817 12672 5891 12675
rect 5435 12660 5499 12672
rect 5435 12643 5457 12660
rect 5491 12643 5499 12660
rect 5435 12591 5447 12643
rect 5435 12579 5499 12591
rect 5435 12527 5447 12579
rect 5435 12526 5457 12527
rect 5491 12526 5499 12527
rect 5435 12514 5499 12526
rect 5604 12660 5891 12672
rect 5604 12626 5614 12660
rect 5648 12643 5891 12660
rect 5648 12638 5886 12643
tri 5886 12638 5891 12643 nw
rect 5648 12626 5854 12638
rect 5604 12606 5854 12626
tri 5854 12606 5886 12638 nw
rect 5604 12604 5852 12606
tri 5852 12604 5854 12606 nw
tri 5960 12604 5962 12606 se
rect 5962 12604 6014 13943
tri 6014 13931 6026 13943 nw
rect 5604 12601 5849 12604
tri 5849 12601 5852 12604 nw
tri 5957 12601 5960 12604 se
rect 5960 12601 6014 12604
rect 5604 12567 5815 12601
tri 5815 12567 5849 12601 nw
tri 5923 12567 5957 12601 se
rect 5957 12584 6014 12601
rect 5957 12567 5997 12584
tri 5997 12567 6014 12584 nw
rect 6085 13834 6287 13926
rect 6085 13800 6091 13834
rect 6125 13800 6287 13834
rect 6085 13746 6287 13800
rect 6085 13712 6091 13746
rect 6125 13712 6287 13746
rect 6085 13662 6287 13712
rect 6085 13628 6097 13662
rect 6131 13628 6169 13662
rect 6203 13628 6241 13662
rect 6275 13628 6287 13662
rect 6085 12810 6287 13628
rect 6085 12776 6091 12810
rect 6125 12776 6287 12810
rect 6085 12722 6287 12776
rect 6085 12688 6091 12722
rect 6125 12688 6287 12722
rect 5604 12560 5801 12567
rect 5604 12526 5614 12560
rect 5648 12553 5801 12560
tri 5801 12553 5815 12567 nw
tri 5909 12553 5923 12567 se
rect 5923 12553 5983 12567
tri 5983 12553 5997 12567 nw
rect 5648 12550 5798 12553
tri 5798 12550 5801 12553 nw
tri 5906 12550 5909 12553 se
rect 5909 12550 5980 12553
tri 5980 12550 5983 12553 nw
rect 5648 12526 5764 12550
rect 5604 12516 5764 12526
tri 5764 12516 5798 12550 nw
tri 5888 12532 5906 12550 se
rect 5906 12532 5962 12550
tri 5962 12532 5980 12550 nw
tri 5872 12516 5888 12532 se
rect 5888 12516 5946 12532
tri 5946 12516 5962 12532 nw
rect 5604 12514 5762 12516
tri 5762 12514 5764 12516 nw
tri 5870 12514 5872 12516 se
rect 5872 12514 5923 12516
tri 5860 12504 5870 12514 se
rect 5870 12504 5923 12514
tri 5849 12493 5860 12504 se
rect 5860 12493 5923 12504
tri 5923 12493 5946 12516 nw
tri 5838 12482 5849 12493 se
rect 5849 12482 5912 12493
tri 5912 12482 5923 12493 nw
tri 5823 12467 5838 12482 se
rect 5838 12467 5897 12482
tri 5897 12467 5912 12482 nw
rect 5488 12415 5495 12467
rect 5547 12415 5559 12467
rect 5611 12448 5878 12467
tri 5878 12448 5897 12467 nw
rect 5611 12441 5871 12448
tri 5871 12441 5878 12448 nw
rect 5611 12420 5850 12441
tri 5850 12420 5871 12441 nw
rect 5611 12415 5845 12420
tri 5845 12415 5850 12420 nw
rect 5075 12381 6057 12387
rect 5075 12347 5087 12381
rect 5121 12347 5162 12381
rect 5196 12347 5237 12381
rect 5271 12347 5312 12381
rect 5346 12347 5386 12381
rect 5420 12347 5460 12381
rect 5494 12347 5534 12381
rect 5568 12347 5608 12381
rect 5642 12347 5682 12381
rect 5716 12347 5756 12381
rect 5790 12347 5830 12381
rect 5864 12347 5904 12381
rect 5938 12347 5978 12381
rect 6012 12347 6057 12381
rect 5075 12341 6057 12347
tri 5980 12316 6005 12341 ne
rect 5065 12175 5977 12181
rect 5065 12141 5077 12175
rect 5111 12141 5154 12175
rect 5188 12141 5231 12175
rect 5265 12141 5308 12175
rect 5342 12141 5385 12175
rect 5419 12141 5463 12175
rect 5497 12141 5541 12175
rect 5575 12141 5619 12175
rect 5653 12141 5697 12175
rect 5731 12141 5775 12175
rect 5809 12141 5853 12175
rect 5887 12141 5931 12175
rect 5965 12141 5977 12175
rect 5065 12120 5977 12141
rect 5065 12103 5478 12120
rect 5594 12103 5977 12120
rect 5065 12069 5077 12103
rect 5111 12069 5154 12103
rect 5188 12069 5231 12103
rect 5265 12069 5308 12103
rect 5342 12069 5385 12103
rect 5419 12069 5463 12103
rect 5594 12069 5619 12103
rect 5653 12069 5697 12103
rect 5731 12069 5775 12103
rect 5809 12069 5853 12103
rect 5887 12069 5931 12103
rect 5965 12069 5977 12103
rect 5065 12031 5478 12069
rect 5594 12031 5977 12069
rect 5065 11997 5077 12031
rect 5111 11997 5154 12031
rect 5188 11997 5231 12031
rect 5265 11997 5308 12031
rect 5342 11997 5385 12031
rect 5419 11997 5463 12031
rect 5594 12004 5619 12031
rect 5497 11997 5541 12004
rect 5575 11997 5619 12004
rect 5653 11997 5697 12031
rect 5731 11997 5775 12031
rect 5809 11997 5853 12031
rect 5887 11997 5931 12031
rect 5965 11997 5977 12031
rect 5065 11991 5977 11997
tri 5980 11735 6005 11760 se
rect 6005 11735 6057 12341
tri 5545 11732 5548 11735 se
rect 5548 11732 6057 11735
rect 5049 11680 5055 11732
rect 5107 11680 5122 11732
rect 5174 11723 5189 11732
rect 5241 11723 5256 11732
rect 5308 11723 5323 11732
rect 5179 11689 5189 11723
rect 5308 11689 5315 11723
rect 5174 11680 5189 11689
rect 5241 11680 5256 11689
rect 5308 11680 5323 11689
rect 5375 11680 5390 11732
rect 5442 11680 5457 11732
rect 5509 11723 5524 11732
rect 5576 11723 5591 11732
rect 5643 11723 5657 11732
rect 5709 11723 5723 11732
rect 5775 11723 5789 11732
rect 5841 11723 5855 11732
rect 5519 11689 5524 11723
rect 5775 11689 5777 11723
rect 5841 11689 5851 11723
rect 5509 11680 5524 11689
rect 5576 11680 5591 11689
rect 5643 11680 5657 11689
rect 5709 11680 5723 11689
rect 5775 11680 5789 11689
rect 5841 11680 5855 11689
rect 5907 11680 5921 11732
rect 5973 11680 5987 11732
rect 6039 11680 6057 11732
tri 5523 11655 5548 11680 ne
rect 5548 11651 5600 11680
tri 5600 11655 5625 11680 nw
rect 5548 11617 5557 11651
rect 5591 11617 5600 11651
rect 5548 11579 5600 11617
rect 5548 11545 5557 11579
rect 5591 11545 5600 11579
rect 5548 11507 5600 11545
rect 5548 11473 5557 11507
rect 5591 11473 5600 11507
tri 5009 11435 5020 11446 sw
rect 5548 11435 5600 11473
rect 4807 11425 5020 11435
tri 5020 11425 5030 11435 sw
rect 4807 11362 5030 11425
rect 5548 11401 5557 11435
rect 5591 11401 5600 11435
tri 6070 11431 6085 11446 se
rect 6085 11431 6287 12688
rect 6366 13918 6568 14080
rect 6366 13884 6378 13918
rect 6412 13884 6450 13918
rect 6484 13884 6522 13918
rect 6556 13884 6568 13918
rect 6366 13835 6568 13884
rect 6418 13783 6442 13835
rect 6494 13783 6516 13835
rect 6366 13767 6568 13783
rect 6418 13715 6442 13767
rect 6494 13715 6516 13767
rect 6366 13699 6568 13715
rect 6418 13647 6442 13699
rect 6494 13647 6516 13699
rect 6366 13631 6568 13647
rect 6418 13579 6442 13631
rect 6494 13579 6516 13631
rect 6366 13563 6568 13579
rect 6418 13511 6442 13563
rect 6494 13511 6516 13563
rect 6366 13406 6568 13511
rect 6366 13372 6378 13406
rect 6412 13372 6450 13406
rect 6484 13372 6522 13406
rect 6556 13372 6568 13406
rect 6366 12894 6568 13372
rect 6366 12860 6378 12894
rect 6412 12860 6450 12894
rect 6484 12860 6522 12894
rect 6556 12860 6568 12894
rect 6366 12685 6568 12860
tri 6366 12675 6376 12685 ne
rect 6376 12675 6568 12685
tri 6376 12650 6401 12675 ne
rect 6401 12650 6568 12675
rect 6315 12638 6361 12650
tri 6401 12644 6407 12650 ne
rect 6407 12644 6568 12650
rect 6315 12604 6321 12638
rect 6355 12604 6361 12638
tri 6407 12615 6436 12644 ne
rect 6315 12550 6361 12604
rect 6315 12516 6321 12550
rect 6355 12516 6361 12550
rect 6315 12504 6361 12516
tri 6361 12504 6367 12510 sw
rect 6315 12270 6367 12504
rect 6436 12482 6568 12644
rect 6436 12448 6448 12482
rect 6482 12448 6522 12482
rect 6556 12448 6568 12482
rect 6436 12442 6568 12448
rect 6647 13149 6849 14080
rect 6647 13115 6659 13149
rect 6693 13115 6731 13149
rect 6765 13115 6803 13149
rect 6837 13115 6849 13149
rect 6647 13003 6849 13115
rect 6647 12951 6653 13003
rect 6705 12951 6717 13003
rect 6769 12951 6781 13003
rect 6833 12951 6849 13003
rect 6315 12206 6367 12218
rect 6315 12148 6367 12154
rect 6327 11680 6333 11732
rect 6385 11680 6405 11732
rect 6457 11680 6477 11732
rect 6529 11680 6549 11732
rect 6601 11680 6607 11732
tri 4807 11341 4828 11362 ne
rect 4224 8488 4236 8522
rect 4270 8488 4308 8522
rect 4342 8488 4380 8522
rect 4414 8488 4426 8522
rect 4224 5098 4426 8488
rect 4224 5064 4236 5098
rect 4270 5064 4308 5098
rect 4342 5064 4380 5098
rect 4414 5064 4426 5098
rect 3968 4193 4000 4227
rect 4034 4193 4040 4227
rect 3968 4154 4040 4193
rect 3968 4120 4000 4154
rect 4034 4120 4040 4154
rect 3968 4081 4040 4120
rect 3968 4047 4000 4081
rect 4034 4047 4040 4081
rect 4224 4052 4426 5064
rect 4526 11248 4728 11254
rect 4526 11214 4538 11248
rect 4572 11214 4610 11248
rect 4644 11214 4682 11248
rect 4716 11214 4728 11248
rect 4526 11090 4728 11214
rect 4526 11056 4538 11090
rect 4572 11056 4610 11090
rect 4644 11056 4682 11090
rect 4716 11056 4728 11090
rect 4526 9378 4728 11056
rect 4526 9344 4538 9378
rect 4572 9344 4610 9378
rect 4644 9344 4682 9378
rect 4716 9344 4728 9378
rect 4526 7666 4728 9344
rect 4526 7632 4538 7666
rect 4572 7632 4610 7666
rect 4644 7632 4682 7666
rect 4716 7632 4728 7666
rect 4526 5954 4728 7632
rect 4526 5920 4538 5954
rect 4572 5920 4610 5954
rect 4644 5920 4682 5954
rect 4716 5920 4728 5954
rect 4526 4242 4728 5920
rect 4526 4208 4538 4242
rect 4572 4208 4610 4242
rect 4644 4208 4682 4242
rect 4716 4208 4728 4242
rect 4526 4084 4728 4208
rect 3968 4008 4040 4047
rect 3968 3974 4000 4008
rect 4034 3979 4040 4008
rect 4526 4050 4538 4084
rect 4572 4050 4610 4084
rect 4644 4050 4682 4084
rect 4716 4050 4728 4084
rect 4828 10234 5030 11362
rect 5058 11362 5320 11368
rect 5322 11367 5358 11368
rect 5058 11328 5070 11362
rect 5104 11328 5150 11362
rect 5184 11328 5320 11362
rect 5058 11324 5320 11328
rect 5058 11322 5274 11324
tri 5243 11297 5268 11322 ne
rect 5268 11290 5274 11322
rect 5308 11290 5320 11324
rect 5268 11251 5320 11290
rect 5268 11217 5274 11251
rect 5308 11217 5320 11251
rect 5268 11178 5320 11217
rect 5268 11144 5274 11178
rect 5308 11144 5320 11178
rect 5268 11105 5320 11144
rect 5268 11071 5274 11105
rect 5308 11071 5320 11105
rect 4828 10200 4840 10234
rect 4874 10200 4912 10234
rect 4946 10200 4984 10234
rect 5018 10200 5030 10234
rect 4828 9849 5030 10200
rect 4828 9797 4850 9849
rect 4902 9797 4930 9849
rect 4982 9797 5030 9849
rect 4828 9783 5030 9797
rect 4828 9731 4850 9783
rect 4902 9731 4930 9783
rect 4982 9731 5030 9783
rect 4828 6810 5030 9731
rect 4828 6776 4840 6810
rect 4874 6776 4912 6810
rect 4946 6776 4984 6810
rect 5018 6776 5030 6810
rect 4828 4052 5030 6776
rect 5186 11033 5238 11045
rect 5186 10999 5192 11033
rect 5226 10999 5238 11033
rect 5186 10967 5238 10999
rect 5186 10901 5238 10915
rect 5186 10811 5238 10849
rect 5186 10777 5192 10811
rect 5226 10777 5238 10811
rect 5186 10737 5238 10777
rect 5186 10703 5192 10737
rect 5226 10703 5238 10737
rect 5186 10663 5238 10703
rect 5186 10629 5192 10663
rect 5226 10629 5238 10663
rect 5186 10589 5238 10629
rect 5186 10555 5192 10589
rect 5226 10555 5238 10589
rect 5186 10515 5238 10555
rect 5186 10481 5192 10515
rect 5226 10481 5238 10515
rect 5186 10441 5238 10481
rect 5186 10407 5192 10441
rect 5226 10407 5238 10441
rect 5186 10366 5238 10407
rect 5186 10332 5192 10366
rect 5226 10332 5238 10366
rect 5186 10291 5238 10332
rect 5186 10257 5192 10291
rect 5226 10257 5238 10291
rect 5186 10177 5238 10257
rect 5186 10143 5192 10177
rect 5226 10143 5238 10177
rect 5186 10103 5238 10143
rect 5186 10069 5192 10103
rect 5226 10069 5238 10103
rect 5186 10029 5238 10069
rect 5186 9995 5192 10029
rect 5226 9995 5238 10029
rect 5186 9955 5238 9995
rect 5186 9921 5192 9955
rect 5226 9921 5238 9955
rect 5186 9881 5238 9921
rect 5186 9847 5192 9881
rect 5226 9847 5238 9881
rect 5186 9807 5238 9847
rect 5186 9773 5192 9807
rect 5226 9773 5238 9807
rect 5186 9733 5238 9773
rect 5186 9699 5192 9733
rect 5226 9699 5238 9733
rect 5186 9659 5238 9699
rect 5186 9625 5192 9659
rect 5226 9625 5238 9659
rect 5186 9585 5238 9625
rect 5186 9551 5192 9585
rect 5226 9551 5238 9585
rect 5186 9510 5238 9551
rect 5186 9476 5192 9510
rect 5226 9476 5238 9510
rect 5186 9435 5238 9476
rect 5186 9401 5192 9435
rect 5226 9401 5238 9435
rect 5186 7609 5238 9401
rect 5186 7575 5192 7609
rect 5226 7575 5238 7609
rect 5186 7535 5238 7575
rect 5186 7501 5192 7535
rect 5226 7501 5238 7535
rect 5186 7461 5238 7501
rect 5186 7427 5192 7461
rect 5226 7427 5238 7461
rect 5186 7387 5238 7427
rect 5186 7353 5192 7387
rect 5226 7353 5238 7387
rect 5186 7313 5238 7353
rect 5186 7279 5192 7313
rect 5226 7279 5238 7313
rect 5186 7239 5238 7279
rect 5186 7205 5192 7239
rect 5226 7205 5238 7239
rect 5186 7165 5238 7205
rect 5186 7131 5192 7165
rect 5226 7131 5238 7165
rect 5186 7091 5238 7131
rect 5186 7057 5192 7091
rect 5226 7057 5238 7091
rect 5186 7043 5238 7057
rect 5186 6983 5192 6991
rect 5226 6983 5238 6991
rect 5186 6977 5238 6983
rect 5186 6908 5192 6925
rect 5226 6908 5238 6925
rect 5186 6867 5238 6908
rect 5186 6833 5192 6867
rect 5226 6833 5238 6867
rect 5186 6753 5238 6833
rect 5186 6719 5192 6753
rect 5226 6719 5238 6753
rect 5186 6679 5238 6719
rect 5186 6645 5192 6679
rect 5226 6645 5238 6679
rect 5186 6605 5238 6645
rect 5186 6571 5192 6605
rect 5226 6571 5238 6605
rect 5186 6531 5238 6571
rect 5186 6497 5192 6531
rect 5226 6497 5238 6531
rect 5186 6457 5238 6497
rect 5186 6423 5192 6457
rect 5226 6423 5238 6457
rect 5186 6383 5238 6423
rect 5186 6349 5192 6383
rect 5226 6349 5238 6383
rect 5186 6309 5238 6349
rect 5186 6275 5192 6309
rect 5226 6275 5238 6309
rect 5186 6235 5238 6275
rect 5186 6201 5192 6235
rect 5226 6201 5238 6235
rect 5186 6161 5238 6201
rect 5186 6127 5192 6161
rect 5226 6127 5238 6161
rect 5186 6086 5238 6127
rect 5186 6052 5192 6086
rect 5226 6052 5238 6086
rect 5186 6011 5238 6052
rect 5186 5977 5192 6011
rect 5226 5977 5238 6011
rect 5186 4249 5238 5977
rect 5268 11032 5320 11071
rect 5268 10998 5274 11032
rect 5308 10998 5320 11032
rect 5268 10959 5320 10998
rect 5268 10925 5274 10959
rect 5308 10925 5320 10959
rect 5268 10886 5320 10925
rect 5268 10852 5274 10886
rect 5308 10852 5320 10886
rect 5268 10813 5320 10852
rect 5268 10779 5274 10813
rect 5308 10779 5320 10813
rect 5268 10740 5320 10779
rect 5268 10706 5274 10740
rect 5308 10706 5320 10740
rect 5268 10667 5320 10706
rect 5268 10633 5274 10667
rect 5308 10633 5320 10667
rect 5268 10594 5320 10633
rect 5268 10560 5274 10594
rect 5308 10560 5320 10594
rect 5268 10521 5320 10560
rect 5268 10487 5274 10521
rect 5308 10487 5320 10521
rect 5268 10448 5320 10487
rect 5268 10414 5274 10448
rect 5308 10414 5320 10448
rect 5268 10375 5320 10414
rect 5268 10341 5274 10375
rect 5308 10341 5320 10375
rect 5268 10302 5320 10341
rect 5268 10268 5274 10302
rect 5308 10268 5320 10302
rect 5268 10229 5320 10268
rect 5268 10195 5274 10229
rect 5308 10195 5320 10229
rect 5268 10156 5320 10195
rect 5268 10122 5274 10156
rect 5308 10122 5320 10156
rect 5268 10083 5320 10122
rect 5268 10049 5274 10083
rect 5308 10049 5320 10083
rect 5268 10010 5320 10049
rect 5268 9976 5274 10010
rect 5308 9976 5320 10010
rect 5268 9937 5320 9976
rect 5268 9903 5274 9937
rect 5308 9903 5320 9937
rect 5268 9864 5320 9903
rect 5268 9830 5274 9864
rect 5308 9830 5320 9864
rect 5268 9791 5320 9830
rect 5268 9757 5274 9791
rect 5308 9757 5320 9791
rect 5268 9718 5320 9757
rect 5268 9684 5274 9718
rect 5308 9684 5320 9718
rect 5268 9645 5320 9684
rect 5268 9611 5274 9645
rect 5308 9611 5320 9645
rect 5268 9572 5320 9611
rect 5268 9538 5274 9572
rect 5308 9538 5320 9572
rect 5268 9499 5320 9538
rect 5268 9465 5274 9499
rect 5308 9465 5320 9499
rect 5268 9426 5320 9465
rect 5268 9392 5274 9426
rect 5308 9392 5320 9426
rect 5268 9353 5320 9392
rect 5268 9319 5274 9353
rect 5308 9319 5320 9353
rect 5268 9280 5320 9319
rect 5268 9246 5274 9280
rect 5308 9246 5320 9280
rect 5268 9207 5320 9246
rect 5268 9173 5274 9207
rect 5308 9173 5320 9207
rect 5268 9134 5320 9173
rect 5268 9100 5274 9134
rect 5308 9100 5320 9134
rect 5268 9061 5320 9100
rect 5268 9027 5274 9061
rect 5308 9027 5320 9061
rect 5268 8988 5320 9027
rect 5268 8954 5274 8988
rect 5308 8954 5320 8988
rect 5268 8915 5320 8954
rect 5268 8881 5274 8915
rect 5308 8881 5320 8915
rect 5268 8842 5320 8881
rect 5268 8808 5274 8842
rect 5308 8808 5320 8842
rect 5268 8769 5320 8808
rect 5268 8735 5274 8769
rect 5308 8735 5320 8769
rect 5268 8696 5320 8735
rect 5268 8662 5274 8696
rect 5308 8662 5320 8696
rect 5268 8623 5320 8662
rect 5268 8589 5274 8623
rect 5308 8589 5320 8623
rect 5268 8550 5320 8589
rect 5268 8516 5274 8550
rect 5308 8516 5320 8550
rect 5268 8477 5320 8516
rect 5268 8443 5274 8477
rect 5308 8443 5320 8477
rect 5268 8404 5320 8443
rect 5268 8370 5274 8404
rect 5308 8370 5320 8404
rect 5268 8331 5320 8370
rect 5268 8297 5274 8331
rect 5308 8297 5320 8331
rect 5268 8258 5320 8297
rect 5268 8224 5274 8258
rect 5308 8224 5320 8258
rect 5268 8185 5320 8224
rect 5268 8151 5274 8185
rect 5308 8151 5320 8185
rect 5268 8112 5320 8151
rect 5268 8078 5274 8112
rect 5308 8078 5320 8112
rect 5268 8040 5320 8078
rect 5268 8006 5274 8040
rect 5308 8006 5320 8040
rect 5268 7968 5320 8006
rect 5268 7934 5274 7968
rect 5308 7934 5320 7968
rect 5268 7896 5320 7934
rect 5268 7862 5274 7896
rect 5308 7862 5320 7896
rect 5268 7824 5320 7862
rect 5268 7790 5274 7824
rect 5308 7790 5320 7824
rect 5268 7752 5320 7790
rect 5268 7718 5274 7752
rect 5308 7718 5320 7752
rect 5268 7680 5320 7718
rect 5268 7646 5274 7680
rect 5308 7646 5320 7680
rect 5268 7608 5320 7646
rect 5268 7574 5274 7608
rect 5308 7574 5320 7608
rect 5268 7536 5320 7574
rect 5268 7502 5274 7536
rect 5308 7502 5320 7536
rect 5268 7464 5320 7502
rect 5268 7430 5274 7464
rect 5308 7430 5320 7464
rect 5268 7392 5320 7430
rect 5268 7358 5274 7392
rect 5308 7358 5320 7392
rect 5268 7320 5320 7358
rect 5268 7286 5274 7320
rect 5308 7286 5320 7320
rect 5268 7248 5320 7286
rect 5268 7214 5274 7248
rect 5308 7214 5320 7248
rect 5268 7176 5320 7214
rect 5268 7142 5274 7176
rect 5308 7142 5320 7176
rect 5268 7104 5320 7142
rect 5268 7070 5274 7104
rect 5308 7070 5320 7104
rect 5268 7032 5320 7070
rect 5268 6998 5274 7032
rect 5308 6998 5320 7032
rect 5268 6960 5320 6998
rect 5268 6926 5274 6960
rect 5308 6926 5320 6960
rect 5268 6888 5320 6926
rect 5268 6854 5274 6888
rect 5308 6854 5320 6888
rect 5268 6816 5320 6854
rect 5268 6782 5274 6816
rect 5308 6782 5320 6816
rect 5268 6744 5320 6782
rect 5268 6710 5274 6744
rect 5308 6710 5320 6744
rect 5268 6672 5320 6710
rect 5268 6638 5274 6672
rect 5308 6638 5320 6672
rect 5268 6600 5320 6638
rect 5268 6566 5274 6600
rect 5308 6566 5320 6600
rect 5268 6528 5320 6566
rect 5268 6494 5274 6528
rect 5308 6494 5320 6528
rect 5268 6456 5320 6494
rect 5268 6422 5274 6456
rect 5308 6422 5320 6456
rect 5268 6384 5320 6422
rect 5268 6350 5274 6384
rect 5308 6350 5320 6384
rect 5268 6312 5320 6350
rect 5268 6278 5274 6312
rect 5308 6278 5320 6312
rect 5268 6240 5320 6278
rect 5268 6206 5274 6240
rect 5308 6206 5320 6240
rect 5268 6168 5320 6206
rect 5268 6134 5274 6168
rect 5308 6134 5320 6168
rect 5268 6096 5320 6134
rect 5268 6062 5274 6096
rect 5308 6062 5320 6096
rect 5268 6024 5320 6062
rect 5268 5990 5274 6024
rect 5308 5990 5320 6024
rect 5268 5952 5320 5990
rect 5268 5918 5274 5952
rect 5308 5918 5320 5952
rect 5268 5880 5320 5918
rect 5268 5846 5274 5880
rect 5308 5846 5320 5880
rect 5268 5808 5320 5846
rect 5268 5774 5274 5808
rect 5308 5774 5320 5808
rect 5268 5736 5320 5774
rect 5268 5702 5274 5736
rect 5308 5702 5320 5736
rect 5268 5664 5320 5702
rect 5268 5630 5274 5664
rect 5308 5630 5320 5664
rect 5268 5592 5320 5630
rect 5268 5558 5274 5592
rect 5308 5558 5320 5592
rect 5268 5520 5320 5558
rect 5268 5486 5274 5520
rect 5308 5486 5320 5520
rect 5268 5448 5320 5486
rect 5268 5414 5274 5448
rect 5308 5414 5320 5448
rect 5268 5376 5320 5414
rect 5268 5342 5274 5376
rect 5308 5342 5320 5376
rect 5268 5304 5320 5342
rect 5268 5270 5274 5304
rect 5308 5270 5320 5304
rect 5268 5232 5320 5270
rect 5268 5198 5274 5232
rect 5308 5198 5320 5232
rect 5268 5160 5320 5198
rect 5268 5126 5274 5160
rect 5308 5126 5320 5160
rect 5268 5088 5320 5126
rect 5268 5054 5274 5088
rect 5308 5054 5320 5088
rect 5268 5016 5320 5054
rect 5268 4982 5274 5016
rect 5308 4982 5320 5016
rect 5268 4944 5320 4982
rect 5268 4910 5274 4944
rect 5308 4910 5320 4944
rect 5268 4872 5320 4910
rect 5268 4838 5274 4872
rect 5308 4838 5320 4872
rect 5268 4800 5320 4838
rect 5268 4766 5274 4800
rect 5308 4766 5320 4800
rect 5268 4728 5320 4766
rect 5268 4694 5274 4728
rect 5308 4694 5320 4728
rect 5268 4656 5320 4694
rect 5268 4622 5274 4656
rect 5308 4622 5320 4656
rect 5268 4584 5320 4622
rect 5268 4550 5274 4584
rect 5308 4550 5320 4584
rect 5268 4512 5320 4550
rect 5268 4478 5274 4512
rect 5308 4478 5320 4512
rect 5268 4440 5320 4478
rect 5268 4406 5274 4440
rect 5308 4406 5320 4440
rect 5268 4368 5320 4406
rect 5268 4334 5274 4368
rect 5308 4334 5320 4368
rect 5268 4296 5320 4334
rect 5268 4262 5274 4296
rect 5308 4262 5320 4296
rect 5268 4224 5320 4262
rect 5268 4190 5274 4224
rect 5308 4190 5320 4224
rect 5268 4152 5320 4190
rect 5268 4118 5274 4152
rect 5308 4118 5320 4152
rect 5268 4080 5320 4118
tri 4040 3979 4062 4001 sw
tri 4504 3979 4526 4001 se
rect 4526 3979 4728 4050
rect 5268 4046 5274 4080
rect 5308 4046 5320 4080
tri 4728 3979 4750 4001 sw
tri 5246 3979 5268 4001 se
rect 5268 3979 5320 4046
rect 4034 3976 4062 3979
tri 4062 3976 4065 3979 sw
tri 4501 3976 4504 3979 se
rect 4504 3976 4750 3979
tri 4750 3976 4753 3979 sw
tri 5243 3976 5246 3979 se
rect 5246 3976 5320 3979
rect 4034 3974 4453 3976
rect 3968 3970 4453 3974
rect 3968 3936 4138 3970
rect 4172 3936 4224 3970
rect 4258 3936 4310 3970
rect 4344 3936 4397 3970
rect 4431 3936 4453 3970
rect 3930 3930 3966 3931
rect 3968 3930 4453 3936
rect 4454 3931 4455 3975
rect 4491 3931 4492 3975
rect 4493 3930 4769 3976
rect 4770 3931 4771 3975
rect 4807 3931 4808 3975
rect 4809 3970 5320 3976
rect 4809 3936 4843 3970
rect 4877 3936 4921 3970
rect 4955 3936 4999 3970
rect 5033 3936 5078 3970
rect 5112 3936 5157 3970
rect 5191 3936 5236 3970
rect 5270 3936 5320 3970
rect 4809 3930 5320 3936
rect 5321 3931 5359 11367
rect 5360 4203 5483 11368
rect 5360 4023 5367 4203
rect 5322 3930 5358 3931
rect 5360 3930 5483 4023
rect 5548 11363 5600 11401
tri 6064 11425 6070 11431 se
rect 6070 11425 6287 11431
rect 5548 11329 5557 11363
rect 5591 11329 5600 11363
rect 5548 11291 5600 11329
rect 5548 11257 5557 11291
rect 5591 11257 5600 11291
rect 5548 11219 5600 11257
rect 5548 11185 5557 11219
rect 5591 11185 5600 11219
rect 5548 11147 5600 11185
rect 5548 11113 5557 11147
rect 5591 11113 5600 11147
rect 5548 11075 5600 11113
rect 5548 11041 5557 11075
rect 5591 11041 5600 11075
rect 5548 11003 5600 11041
rect 5548 10969 5557 11003
rect 5591 10969 5600 11003
rect 5548 10931 5600 10969
rect 5548 10897 5557 10931
rect 5591 10897 5600 10931
rect 5548 10859 5600 10897
rect 5548 10825 5557 10859
rect 5591 10825 5600 10859
rect 5548 10787 5600 10825
rect 5548 10753 5557 10787
rect 5591 10753 5600 10787
rect 5548 10715 5600 10753
rect 5548 10681 5557 10715
rect 5591 10681 5600 10715
rect 5548 10643 5600 10681
rect 5548 10609 5557 10643
rect 5591 10609 5600 10643
rect 5548 10571 5600 10609
rect 5548 10537 5557 10571
rect 5591 10537 5600 10571
rect 5548 10499 5600 10537
rect 5548 10465 5557 10499
rect 5591 10465 5600 10499
rect 5548 10427 5600 10465
rect 5548 10393 5557 10427
rect 5591 10393 5600 10427
rect 5548 10355 5600 10393
rect 5548 10321 5557 10355
rect 5591 10321 5600 10355
rect 5548 10283 5600 10321
rect 5548 10249 5557 10283
rect 5591 10249 5600 10283
rect 5548 10243 5600 10249
rect 5548 10179 5557 10191
rect 5591 10179 5600 10191
rect 5548 10114 5557 10127
rect 5591 10114 5600 10127
rect 5548 10033 5557 10062
rect 5591 10033 5600 10062
rect 5548 9995 5600 10033
rect 5548 9961 5557 9995
rect 5591 9961 5600 9995
rect 5548 9923 5600 9961
rect 5548 9889 5557 9923
rect 5591 9889 5600 9923
rect 5548 9851 5600 9889
rect 5548 9817 5557 9851
rect 5591 9817 5600 9851
rect 5548 9779 5600 9817
rect 5548 9745 5557 9779
rect 5591 9745 5600 9779
rect 5548 9707 5600 9745
rect 5548 9673 5557 9707
rect 5591 9673 5600 9707
rect 5548 9635 5600 9673
rect 5548 9601 5557 9635
rect 5591 9601 5600 9635
rect 5548 9563 5600 9601
rect 5548 9529 5557 9563
rect 5591 9529 5600 9563
rect 5548 9491 5600 9529
rect 5548 9457 5557 9491
rect 5591 9457 5600 9491
rect 5548 9419 5600 9457
rect 5548 9385 5557 9419
rect 5591 9385 5600 9419
rect 5548 9347 5600 9385
rect 5548 9313 5557 9347
rect 5591 9313 5600 9347
rect 5548 9275 5600 9313
rect 5548 9241 5557 9275
rect 5591 9241 5600 9275
rect 5548 9203 5600 9241
rect 5548 9169 5557 9203
rect 5591 9169 5600 9203
rect 5548 9131 5600 9169
rect 5548 9097 5557 9131
rect 5591 9097 5600 9131
rect 5548 9059 5600 9097
rect 5548 9025 5557 9059
rect 5591 9025 5600 9059
rect 5548 8987 5600 9025
rect 5548 8953 5557 8987
rect 5591 8953 5600 8987
rect 5548 8915 5600 8953
rect 5548 8881 5557 8915
rect 5591 8881 5600 8915
rect 5548 8843 5600 8881
rect 5548 8809 5557 8843
rect 5591 8809 5600 8843
rect 5548 8771 5600 8809
rect 5548 8737 5557 8771
rect 5591 8737 5600 8771
rect 5548 8699 5600 8737
rect 5548 8665 5557 8699
rect 5591 8665 5600 8699
rect 5548 8627 5600 8665
rect 5548 8593 5557 8627
rect 5591 8593 5600 8627
rect 5548 8555 5600 8593
rect 5548 8521 5557 8555
rect 5591 8521 5600 8555
rect 5548 8483 5600 8521
rect 5548 8449 5557 8483
rect 5591 8449 5600 8483
rect 5548 8411 5600 8449
rect 5548 8377 5557 8411
rect 5591 8377 5600 8411
rect 5548 8339 5600 8377
rect 5548 8305 5557 8339
rect 5591 8305 5600 8339
rect 5548 8267 5600 8305
rect 5548 8233 5557 8267
rect 5591 8233 5600 8267
rect 5548 8195 5600 8233
rect 5548 8161 5557 8195
rect 5591 8161 5600 8195
rect 5548 8146 5600 8161
rect 5548 8089 5557 8094
rect 5591 8089 5600 8094
rect 5548 8082 5600 8089
rect 5548 8017 5557 8030
rect 5591 8017 5600 8030
rect 5548 7945 5557 7965
rect 5591 7945 5600 7965
rect 5548 7907 5600 7945
rect 5548 7873 5557 7907
rect 5591 7873 5600 7907
rect 5548 7835 5600 7873
rect 5548 7801 5557 7835
rect 5591 7801 5600 7835
rect 5548 7763 5600 7801
rect 5548 7729 5557 7763
rect 5591 7729 5600 7763
rect 5548 7691 5600 7729
rect 5548 7657 5557 7691
rect 5591 7657 5600 7691
rect 5548 7619 5600 7657
rect 5548 7585 5557 7619
rect 5591 7585 5600 7619
rect 5548 7547 5600 7585
rect 5548 7513 5557 7547
rect 5591 7513 5600 7547
rect 5548 7475 5600 7513
rect 5548 7441 5557 7475
rect 5591 7441 5600 7475
rect 5548 7403 5600 7441
rect 5548 7369 5557 7403
rect 5591 7369 5600 7403
rect 5548 7331 5600 7369
rect 5548 7297 5557 7331
rect 5591 7297 5600 7331
rect 5548 7259 5600 7297
rect 5548 7225 5557 7259
rect 5591 7225 5600 7259
rect 5548 7187 5600 7225
rect 5548 7153 5557 7187
rect 5591 7153 5600 7187
rect 5548 7115 5600 7153
rect 5548 7081 5557 7115
rect 5591 7081 5600 7115
rect 5548 7043 5600 7081
rect 5548 7009 5557 7043
rect 5591 7009 5600 7043
rect 5548 6971 5600 7009
rect 5548 6937 5557 6971
rect 5591 6937 5600 6971
rect 5548 6899 5600 6937
rect 5548 6865 5557 6899
rect 5591 6865 5600 6899
rect 5548 6826 5600 6865
rect 5548 6792 5557 6826
rect 5591 6792 5600 6826
rect 5548 6753 5600 6792
rect 5548 6719 5557 6753
rect 5591 6719 5600 6753
rect 5548 6680 5600 6719
rect 5548 6646 5557 6680
rect 5591 6646 5600 6680
rect 5548 6607 5600 6646
rect 5548 6573 5557 6607
rect 5591 6573 5600 6607
rect 5548 6534 5600 6573
rect 5548 6500 5557 6534
rect 5591 6500 5600 6534
rect 5548 6461 5600 6500
rect 5548 6427 5557 6461
rect 5591 6427 5600 6461
rect 5548 6388 5600 6427
rect 5548 6354 5557 6388
rect 5591 6354 5600 6388
rect 5548 6315 5600 6354
rect 5548 6281 5557 6315
rect 5591 6281 5600 6315
rect 5548 6242 5600 6281
rect 5548 6208 5557 6242
rect 5591 6208 5600 6242
rect 5548 6169 5600 6208
rect 5548 6135 5557 6169
rect 5591 6135 5600 6169
rect 5548 6096 5600 6135
rect 5548 6062 5557 6096
rect 5591 6062 5600 6096
rect 5548 6023 5600 6062
rect 5548 5989 5557 6023
rect 5591 5989 5600 6023
rect 5548 5950 5600 5989
rect 5548 5916 5557 5950
rect 5591 5916 5600 5950
rect 5548 5877 5600 5916
rect 5548 5843 5557 5877
rect 5591 5843 5600 5877
rect 5548 5804 5600 5843
rect 5548 5770 5557 5804
rect 5591 5770 5600 5804
rect 5548 5731 5600 5770
rect 5548 5697 5557 5731
rect 5591 5697 5600 5731
rect 5548 5658 5600 5697
rect 5548 5624 5557 5658
rect 5591 5624 5600 5658
rect 5548 5585 5600 5624
rect 5548 5551 5557 5585
rect 5591 5551 5600 5585
rect 5548 5512 5600 5551
rect 5548 5478 5557 5512
rect 5591 5478 5600 5512
rect 5548 5439 5600 5478
rect 5548 5405 5557 5439
rect 5591 5405 5600 5439
rect 5548 5366 5600 5405
rect 5548 5332 5557 5366
rect 5591 5332 5600 5366
rect 5548 5293 5600 5332
rect 5548 5259 5557 5293
rect 5591 5259 5600 5293
rect 5548 5220 5600 5259
rect 5548 5186 5557 5220
rect 5591 5186 5600 5220
rect 5548 5147 5600 5186
rect 5548 5113 5557 5147
rect 5591 5113 5600 5147
rect 5548 5074 5600 5113
rect 5548 5040 5557 5074
rect 5591 5040 5600 5074
rect 5548 5001 5600 5040
rect 5548 4967 5557 5001
rect 5591 4967 5600 5001
rect 5548 4928 5600 4967
rect 5548 4894 5557 4928
rect 5591 4894 5600 4928
rect 5548 4880 5600 4894
rect 5548 4821 5557 4828
rect 5591 4821 5600 4828
rect 5548 4814 5600 4821
rect 5548 4748 5557 4762
rect 5591 4748 5600 4762
rect 5548 4709 5600 4748
rect 5548 4675 5557 4709
rect 5591 4675 5600 4709
rect 5548 4636 5600 4675
rect 5548 4602 5557 4636
rect 5591 4602 5600 4636
rect 5548 4563 5600 4602
rect 5548 4529 5557 4563
rect 5591 4529 5600 4563
rect 5548 4490 5600 4529
rect 5548 4456 5557 4490
rect 5591 4456 5600 4490
rect 5548 4417 5600 4456
rect 5548 4383 5557 4417
rect 5591 4383 5600 4417
rect 5548 4344 5600 4383
rect 5548 4310 5557 4344
rect 5591 4310 5600 4344
rect 5548 4271 5600 4310
rect 5548 4237 5557 4271
rect 5591 4237 5600 4271
rect 5548 4198 5600 4237
rect 5548 4164 5557 4198
rect 5591 4164 5600 4198
rect 5548 4125 5600 4164
rect 5548 4091 5557 4125
rect 5591 4091 5600 4125
rect 5548 4052 5600 4091
rect 5548 4018 5557 4052
rect 5591 4018 5600 4052
rect 5548 3979 5600 4018
rect 5548 3945 5557 3979
rect 5591 3945 5600 3979
rect 3761 3909 3895 3930
tri 3895 3909 3916 3930 nw
tri 4501 3909 4522 3930 ne
rect 4522 3909 4732 3930
tri 4732 3909 4753 3930 nw
rect 3761 3906 3892 3909
tri 3892 3906 3895 3909 nw
tri 4522 3906 4525 3909 ne
rect 4525 3906 4729 3909
tri 4729 3906 4732 3909 nw
rect 5548 3906 5600 3945
rect 5678 7341 5788 11368
rect 5790 11367 5826 11368
rect 5789 7341 5827 11367
rect 5794 7161 5827 7341
rect 5678 6819 5788 7161
rect 5789 6819 5827 7161
rect 5794 6639 5827 6819
rect 5678 5638 5788 6639
rect 5789 5638 5827 6639
rect 5794 5458 5827 5638
rect 5678 4203 5788 5458
rect 5789 4203 5827 5458
rect 5794 4023 5827 4203
rect 5678 3930 5788 4023
rect 5789 3931 5827 4023
rect 5828 11362 6036 11368
rect 5828 11328 5878 11362
rect 5912 11328 5990 11362
rect 6024 11328 6036 11362
rect 5828 11322 6036 11328
rect 6064 11362 6287 11425
rect 5828 11252 5880 11322
tri 5880 11297 5905 11322 nw
rect 5828 11218 5840 11252
rect 5874 11218 5880 11252
rect 5828 11180 5880 11218
rect 5828 11146 5840 11180
rect 5874 11146 5880 11180
rect 5828 11108 5880 11146
rect 5828 11074 5840 11108
rect 5874 11074 5880 11108
rect 5828 11036 5880 11074
rect 5828 11002 5840 11036
rect 5874 11002 5880 11036
rect 5828 10964 5880 11002
rect 5828 10930 5840 10964
rect 5874 10930 5880 10964
rect 5828 10892 5880 10930
rect 5828 10858 5840 10892
rect 5874 10858 5880 10892
rect 5828 10820 5880 10858
rect 5828 10786 5840 10820
rect 5874 10786 5880 10820
rect 5828 10748 5880 10786
rect 5828 10714 5840 10748
rect 5874 10714 5880 10748
rect 5828 10676 5880 10714
rect 5828 10642 5840 10676
rect 5874 10642 5880 10676
rect 5828 10604 5880 10642
rect 5828 10570 5840 10604
rect 5874 10570 5880 10604
rect 5828 10532 5880 10570
rect 5828 10498 5840 10532
rect 5874 10498 5880 10532
rect 5828 10460 5880 10498
rect 5828 10426 5840 10460
rect 5874 10426 5880 10460
rect 5828 10388 5880 10426
rect 5828 10354 5840 10388
rect 5874 10354 5880 10388
rect 5828 10316 5880 10354
rect 5828 10282 5840 10316
rect 5874 10282 5880 10316
rect 5828 10244 5880 10282
rect 5828 10210 5840 10244
rect 5874 10210 5880 10244
rect 5828 10172 5880 10210
rect 5828 10138 5840 10172
rect 5874 10138 5880 10172
rect 5828 10100 5880 10138
rect 5828 10066 5840 10100
rect 5874 10066 5880 10100
rect 5828 10028 5880 10066
rect 5828 9994 5840 10028
rect 5874 9994 5880 10028
rect 5828 9956 5880 9994
rect 5828 9922 5840 9956
rect 5874 9922 5880 9956
rect 5828 9884 5880 9922
rect 5828 9850 5840 9884
rect 5874 9850 5880 9884
rect 5828 9812 5880 9850
rect 5828 9778 5840 9812
rect 5874 9778 5880 9812
rect 5828 9740 5880 9778
rect 5828 9706 5840 9740
rect 5874 9706 5880 9740
rect 5828 9668 5880 9706
rect 5828 9634 5840 9668
rect 5874 9634 5880 9668
rect 5828 9596 5880 9634
rect 5828 9562 5840 9596
rect 5874 9562 5880 9596
rect 5828 9524 5880 9562
rect 5828 9490 5840 9524
rect 5874 9490 5880 9524
rect 5828 9452 5880 9490
rect 5828 9418 5840 9452
rect 5874 9418 5880 9452
rect 5828 9380 5880 9418
rect 5828 9346 5840 9380
rect 5874 9346 5880 9380
rect 5828 9308 5880 9346
rect 5828 9274 5840 9308
rect 5874 9274 5880 9308
rect 5828 9236 5880 9274
rect 5828 9202 5840 9236
rect 5874 9202 5880 9236
rect 5828 9164 5880 9202
rect 5828 9130 5840 9164
rect 5874 9130 5880 9164
rect 5828 9092 5880 9130
rect 5828 9058 5840 9092
rect 5874 9058 5880 9092
rect 5828 9020 5880 9058
rect 5828 8986 5840 9020
rect 5874 8986 5880 9020
rect 5828 8948 5880 8986
rect 5828 8914 5840 8948
rect 5874 8914 5880 8948
rect 5828 8876 5880 8914
rect 5828 8842 5840 8876
rect 5874 8842 5880 8876
rect 5828 8804 5880 8842
rect 5828 8770 5840 8804
rect 5874 8770 5880 8804
rect 5828 8732 5880 8770
rect 5828 8698 5840 8732
rect 5874 8698 5880 8732
rect 5828 8660 5880 8698
rect 5828 8626 5840 8660
rect 5874 8626 5880 8660
rect 5828 8588 5880 8626
rect 5828 8554 5840 8588
rect 5874 8554 5880 8588
rect 5828 8516 5880 8554
rect 5828 8482 5840 8516
rect 5874 8482 5880 8516
rect 5828 8444 5880 8482
rect 5828 8410 5840 8444
rect 5874 8410 5880 8444
rect 5828 8372 5880 8410
rect 5828 8338 5840 8372
rect 5874 8338 5880 8372
rect 5828 8300 5880 8338
rect 5828 8266 5840 8300
rect 5874 8266 5880 8300
rect 5828 8228 5880 8266
rect 5828 8194 5840 8228
rect 5874 8194 5880 8228
rect 5828 8156 5880 8194
rect 5828 8122 5840 8156
rect 5874 8122 5880 8156
rect 5828 8084 5880 8122
rect 5828 8050 5840 8084
rect 5874 8050 5880 8084
rect 5828 8012 5880 8050
rect 5828 7978 5840 8012
rect 5874 7978 5880 8012
rect 5828 7940 5880 7978
rect 5828 7906 5840 7940
rect 5874 7906 5880 7940
rect 5828 7868 5880 7906
rect 5828 7834 5840 7868
rect 5874 7834 5880 7868
rect 5828 7796 5880 7834
rect 5828 7762 5840 7796
rect 5874 7762 5880 7796
rect 5828 7724 5880 7762
rect 5828 7690 5840 7724
rect 5874 7690 5880 7724
rect 5828 7652 5880 7690
rect 5828 7618 5840 7652
rect 5874 7618 5880 7652
rect 5828 7580 5880 7618
rect 5828 7546 5840 7580
rect 5874 7546 5880 7580
rect 5828 7508 5880 7546
rect 5828 7474 5840 7508
rect 5874 7474 5880 7508
rect 5828 7436 5880 7474
rect 5828 7402 5840 7436
rect 5874 7402 5880 7436
rect 5828 7364 5880 7402
rect 5828 7330 5840 7364
rect 5874 7330 5880 7364
rect 5828 7292 5880 7330
rect 5828 7258 5840 7292
rect 5874 7258 5880 7292
rect 5828 7220 5880 7258
rect 5828 7186 5840 7220
rect 5874 7186 5880 7220
rect 5828 7147 5880 7186
rect 5828 7113 5840 7147
rect 5874 7113 5880 7147
rect 5828 7074 5880 7113
rect 5828 7040 5840 7074
rect 5874 7040 5880 7074
rect 5828 7001 5880 7040
rect 5828 6967 5840 7001
rect 5874 6967 5880 7001
rect 5828 6928 5880 6967
rect 5828 6894 5840 6928
rect 5874 6894 5880 6928
rect 5828 6855 5880 6894
rect 5828 6821 5840 6855
rect 5874 6821 5880 6855
rect 5828 6782 5880 6821
rect 5828 6748 5840 6782
rect 5874 6748 5880 6782
rect 5828 6709 5880 6748
rect 5828 6675 5840 6709
rect 5874 6675 5880 6709
rect 5828 6636 5880 6675
rect 5828 6602 5840 6636
rect 5874 6602 5880 6636
rect 5828 6563 5880 6602
rect 5828 6529 5840 6563
rect 5874 6529 5880 6563
rect 5828 6490 5880 6529
rect 5828 6456 5840 6490
rect 5874 6456 5880 6490
rect 5828 6417 5880 6456
rect 5828 6383 5840 6417
rect 5874 6383 5880 6417
rect 5828 6344 5880 6383
rect 5828 6310 5840 6344
rect 5874 6310 5880 6344
rect 5828 6271 5880 6310
rect 5828 6237 5840 6271
rect 5874 6237 5880 6271
rect 5828 6198 5880 6237
rect 5828 6164 5840 6198
rect 5874 6164 5880 6198
rect 5828 6125 5880 6164
rect 5828 6091 5840 6125
rect 5874 6091 5880 6125
rect 5828 6052 5880 6091
rect 5828 6018 5840 6052
rect 5874 6018 5880 6052
rect 5828 5979 5880 6018
rect 5828 5945 5840 5979
rect 5874 5945 5880 5979
rect 5828 5906 5880 5945
rect 5828 5872 5840 5906
rect 5874 5872 5880 5906
rect 5828 5833 5880 5872
rect 5828 5799 5840 5833
rect 5874 5799 5880 5833
rect 5828 5760 5880 5799
rect 5828 5726 5840 5760
rect 5874 5726 5880 5760
rect 5828 5687 5880 5726
rect 5828 5653 5840 5687
rect 5874 5653 5880 5687
rect 5828 5614 5880 5653
rect 5828 5580 5840 5614
rect 5874 5580 5880 5614
rect 5828 5541 5880 5580
rect 5828 5507 5840 5541
rect 5874 5507 5880 5541
rect 5828 5468 5880 5507
rect 5828 5434 5840 5468
rect 5874 5434 5880 5468
rect 5828 5395 5880 5434
rect 5828 5361 5840 5395
rect 5874 5361 5880 5395
rect 5828 5322 5880 5361
rect 5828 5288 5840 5322
rect 5874 5288 5880 5322
rect 5828 5249 5880 5288
rect 5828 5215 5840 5249
rect 5874 5215 5880 5249
rect 5828 5176 5880 5215
rect 5828 5142 5840 5176
rect 5874 5142 5880 5176
rect 5828 5103 5880 5142
rect 5828 5069 5840 5103
rect 5874 5069 5880 5103
rect 5828 5030 5880 5069
rect 5828 4996 5840 5030
rect 5874 4996 5880 5030
rect 5828 4957 5880 4996
rect 5828 4923 5840 4957
rect 5874 4923 5880 4957
rect 5828 4884 5880 4923
rect 5828 4850 5840 4884
rect 5874 4850 5880 4884
rect 5828 4811 5880 4850
rect 5828 4777 5840 4811
rect 5874 4777 5880 4811
rect 5828 4738 5880 4777
rect 5828 4704 5840 4738
rect 5874 4704 5880 4738
rect 5828 4665 5880 4704
rect 5828 4631 5840 4665
rect 5874 4631 5880 4665
rect 5828 4592 5880 4631
rect 5828 4558 5840 4592
rect 5874 4558 5880 4592
rect 5828 4519 5880 4558
rect 5828 4485 5840 4519
rect 5874 4485 5880 4519
rect 5828 4446 5880 4485
rect 5828 4412 5840 4446
rect 5874 4412 5880 4446
rect 5828 4373 5880 4412
rect 5828 4339 5840 4373
rect 5874 4339 5880 4373
rect 5828 4300 5880 4339
rect 5828 4266 5840 4300
rect 5874 4266 5880 4300
rect 5828 4227 5880 4266
rect 5910 9321 5962 11045
rect 5910 9287 5922 9321
rect 5956 9287 5962 9321
rect 5910 9247 5962 9287
rect 5910 9213 5922 9247
rect 5956 9213 5962 9247
rect 5910 9173 5962 9213
rect 5910 9139 5922 9173
rect 5956 9139 5962 9173
rect 5910 9099 5962 9139
rect 5910 9065 5922 9099
rect 5956 9065 5962 9099
rect 5910 9025 5962 9065
rect 5910 8991 5922 9025
rect 5956 8991 5962 9025
rect 5910 8983 5962 8991
rect 5910 8917 5922 8931
rect 5956 8917 5962 8931
rect 5910 8843 5922 8865
rect 5956 8843 5962 8865
rect 5910 8803 5962 8843
rect 5910 8769 5922 8803
rect 5956 8769 5962 8803
rect 5910 8729 5962 8769
rect 5910 8695 5922 8729
rect 5956 8695 5962 8729
rect 5910 8654 5962 8695
rect 5910 8620 5922 8654
rect 5956 8620 5962 8654
rect 5910 8579 5962 8620
rect 5910 8545 5922 8579
rect 5956 8545 5962 8579
rect 5910 8465 5962 8545
rect 5910 8431 5922 8465
rect 5956 8431 5962 8465
rect 5910 8391 5962 8431
rect 5910 8357 5922 8391
rect 5956 8357 5962 8391
rect 5910 8317 5962 8357
rect 5910 8283 5922 8317
rect 5956 8283 5962 8317
rect 5910 8243 5962 8283
rect 5910 8209 5922 8243
rect 5956 8209 5962 8243
rect 5910 8169 5962 8209
rect 5910 8135 5922 8169
rect 5956 8135 5962 8169
rect 5910 8095 5962 8135
rect 5910 8061 5922 8095
rect 5956 8061 5962 8095
rect 5910 8021 5962 8061
rect 5910 7987 5922 8021
rect 5956 7987 5962 8021
rect 5910 7947 5962 7987
rect 5910 7913 5922 7947
rect 5956 7913 5962 7947
rect 5910 7873 5962 7913
rect 5910 7839 5922 7873
rect 5956 7839 5962 7873
rect 5910 7798 5962 7839
rect 5910 7764 5922 7798
rect 5956 7764 5962 7798
rect 5910 7723 5962 7764
rect 5910 7689 5922 7723
rect 5956 7689 5962 7723
rect 5910 5897 5962 7689
rect 5910 5863 5922 5897
rect 5956 5863 5962 5897
rect 5910 5823 5962 5863
rect 5910 5789 5922 5823
rect 5956 5789 5962 5823
rect 5910 5749 5962 5789
rect 5910 5715 5922 5749
rect 5956 5715 5962 5749
rect 5910 5675 5962 5715
rect 5910 5641 5922 5675
rect 5956 5641 5962 5675
rect 5910 5601 5962 5641
rect 5910 5567 5922 5601
rect 5956 5567 5962 5601
rect 5910 5527 5962 5567
rect 5910 5493 5922 5527
rect 5956 5493 5962 5527
rect 5910 5453 5962 5493
rect 5910 5419 5922 5453
rect 5956 5419 5962 5453
rect 5910 5379 5962 5419
rect 5910 5345 5922 5379
rect 5956 5345 5962 5379
rect 5910 5305 5962 5345
rect 5910 5282 5922 5305
rect 5956 5282 5962 5305
rect 5910 5216 5922 5230
rect 5956 5216 5962 5230
rect 5910 5155 5962 5164
rect 5910 5121 5922 5155
rect 5956 5121 5962 5155
rect 5910 5041 5962 5121
rect 5910 5007 5922 5041
rect 5956 5007 5962 5041
rect 5910 4967 5962 5007
rect 5910 4933 5922 4967
rect 5956 4933 5962 4967
rect 5910 4893 5962 4933
rect 5910 4859 5922 4893
rect 5956 4859 5962 4893
rect 5910 4819 5962 4859
rect 5910 4785 5922 4819
rect 5956 4785 5962 4819
rect 5910 4745 5962 4785
rect 5910 4711 5922 4745
rect 5956 4711 5962 4745
rect 5910 4671 5962 4711
rect 5910 4637 5922 4671
rect 5956 4637 5962 4671
rect 5910 4597 5962 4637
rect 5910 4563 5922 4597
rect 5956 4563 5962 4597
rect 5910 4523 5962 4563
rect 5910 4489 5922 4523
rect 5956 4489 5962 4523
rect 5910 4449 5962 4489
rect 5910 4415 5922 4449
rect 5956 4415 5962 4449
rect 5910 4374 5962 4415
rect 5910 4340 5922 4374
rect 5956 4340 5962 4374
rect 5910 4299 5962 4340
rect 5910 4265 5922 4299
rect 5956 4265 5962 4299
rect 5910 4249 5962 4265
rect 6064 8522 6266 11362
tri 6266 11341 6287 11362 nw
rect 6647 11431 6849 12951
rect 6923 13740 7125 14080
rect 7204 14063 7376 14093
tri 7376 14063 7406 14093 sw
rect 7204 13980 7406 14063
rect 7204 13946 7216 13980
rect 7250 13946 7288 13980
rect 7322 13946 7360 13980
rect 7394 13946 7406 13980
rect 7204 13940 7406 13946
rect 6923 13706 6929 13740
rect 6963 13706 7125 13740
rect 6923 13652 7125 13706
rect 6923 13618 6929 13652
rect 6963 13618 7125 13652
rect 6923 13485 7125 13618
rect 6923 13451 6929 13485
rect 6963 13451 7125 13485
rect 6923 13397 7125 13451
rect 6923 13363 6929 13397
rect 6963 13363 7125 13397
rect 6923 13228 7125 13363
rect 6923 13194 6929 13228
rect 6963 13194 7125 13228
rect 6923 13140 7125 13194
rect 6923 13106 6929 13140
rect 6963 13106 7125 13140
rect 6923 13003 7125 13106
rect 6923 12972 6930 13003
rect 6923 12938 6929 12972
rect 6982 12951 6994 13003
rect 7046 12951 7058 13003
rect 7110 12951 7125 13003
rect 6963 12938 7125 12951
rect 6923 12884 7125 12938
rect 6923 12850 6929 12884
rect 6963 12850 7125 12884
rect 6923 12528 7125 12850
rect 7204 13835 7406 13841
rect 7256 13783 7279 13835
rect 7331 13783 7354 13835
rect 7204 13767 7406 13783
rect 7256 13715 7279 13767
rect 7331 13715 7354 13767
rect 7204 13699 7406 13715
rect 7256 13647 7279 13699
rect 7331 13647 7354 13699
rect 7204 13631 7406 13647
rect 7256 13579 7279 13631
rect 7331 13579 7354 13631
rect 7204 13563 7406 13579
rect 7256 13511 7279 13563
rect 7331 13511 7354 13563
rect 7204 13312 7406 13511
rect 7204 13278 7216 13312
rect 7250 13278 7288 13312
rect 7322 13278 7360 13312
rect 7394 13278 7406 13312
rect 7204 12800 7406 13278
rect 7204 12766 7216 12800
rect 7250 12766 7288 12800
rect 7322 12766 7360 12800
rect 7394 12766 7406 12800
rect 7204 12644 7406 12766
rect 7204 12610 7216 12644
rect 7250 12610 7288 12644
rect 7322 12610 7360 12644
rect 7394 12610 7406 12644
rect 7204 12528 7406 12610
rect 7485 13568 7687 14144
rect 8003 14132 9110 14138
rect 7485 13534 7497 13568
rect 7531 13534 7569 13568
rect 7603 13534 7641 13568
rect 7675 13534 7687 13568
rect 7485 13056 7687 13534
rect 7485 13022 7497 13056
rect 7531 13022 7569 13056
rect 7603 13022 7641 13056
rect 7675 13022 7687 13056
rect 7485 12600 7687 13022
tri 7485 12567 7518 12600 ne
rect 7518 12567 7687 12600
tri 7518 12553 7532 12567 ne
rect 7532 12553 7687 12567
tri 7532 12528 7557 12553 ne
rect 6887 12386 7504 12392
rect 6887 12352 6899 12386
rect 6933 12352 6978 12386
rect 7012 12352 7058 12386
rect 7092 12352 7138 12386
rect 7172 12352 7218 12386
rect 7252 12352 7298 12386
rect 7332 12352 7378 12386
rect 7412 12352 7458 12386
rect 7492 12352 7504 12386
rect 6887 12346 7504 12352
tri 7433 12321 7458 12346 ne
rect 6877 12175 7430 12181
rect 6877 12141 6889 12175
rect 6923 12141 6971 12175
rect 7005 12141 7053 12175
rect 7087 12141 7135 12175
rect 7169 12141 7218 12175
rect 7252 12141 7301 12175
rect 7335 12141 7384 12175
rect 7418 12141 7430 12175
rect 6877 12120 7430 12141
rect 6877 12103 7263 12120
rect 7379 12103 7430 12120
rect 6877 12069 6889 12103
rect 6923 12069 6971 12103
rect 7005 12069 7053 12103
rect 7087 12069 7135 12103
rect 7169 12069 7218 12103
rect 7252 12069 7263 12103
rect 7379 12069 7384 12103
rect 7418 12069 7430 12103
rect 6877 12031 7263 12069
rect 7379 12031 7430 12069
rect 6877 11997 6889 12031
rect 6923 11997 6971 12031
rect 7005 11997 7053 12031
rect 7087 11997 7135 12031
rect 7169 11997 7218 12031
rect 7252 12004 7263 12031
rect 7379 12004 7384 12031
rect 7252 11997 7301 12004
rect 7335 11997 7384 12004
rect 7418 11997 7430 12031
rect 6877 11991 7430 11997
tri 7417 11842 7458 11883 se
rect 7458 11842 7504 12346
rect 7417 11836 7504 11842
rect 7469 11833 7504 11836
tri 7469 11798 7504 11833 nw
rect 7417 11763 7469 11784
tri 7392 11729 7417 11754 se
rect 6889 11723 7417 11729
rect 6889 11689 6901 11723
rect 6935 11689 6976 11723
rect 7010 11689 7051 11723
rect 7085 11689 7126 11723
rect 7160 11689 7201 11723
rect 7235 11689 7276 11723
rect 7310 11689 7351 11723
rect 7385 11711 7417 11723
rect 7385 11689 7423 11711
rect 7457 11689 7469 11711
rect 6889 11683 7417 11689
tri 7392 11658 7417 11683 ne
rect 7557 11723 7687 12553
rect 7755 14093 7801 14105
rect 7755 14059 7761 14093
rect 7795 14059 7801 14093
rect 7755 14018 7801 14059
rect 8003 14098 8015 14132
rect 8049 14098 8089 14132
rect 8123 14098 8164 14132
rect 8198 14098 8239 14132
rect 8273 14098 8314 14132
rect 8348 14098 8389 14132
rect 8423 14098 8464 14132
rect 8498 14098 8539 14132
rect 8573 14098 8614 14132
rect 8648 14098 8689 14132
rect 8723 14098 8764 14132
rect 8798 14098 8839 14132
rect 8873 14098 8914 14132
rect 8948 14098 8989 14132
rect 9023 14098 9064 14132
rect 9098 14098 9110 14132
rect 9359 14126 9909 14194
tri 9909 14169 9934 14194 nw
tri 11046 14169 11071 14194 ne
tri 7801 14018 7822 14039 sw
tri 7982 14018 8003 14039 se
rect 8003 14018 9110 14098
rect 7755 13984 7761 14018
rect 7795 14014 7822 14018
tri 7822 14014 7826 14018 sw
tri 7978 14014 7982 14018 se
rect 7982 14014 9110 14018
rect 7795 13984 7861 14014
rect 7863 14013 7899 14014
rect 7755 13962 7861 13984
rect 7862 13963 7900 14013
rect 7863 13962 7899 13963
rect 7901 13962 9110 14014
rect 7755 13946 7810 13962
tri 7810 13946 7826 13962 nw
tri 7978 13946 7994 13962 ne
rect 7994 13946 9110 13962
rect 7755 13943 7807 13946
tri 7807 13943 7810 13946 nw
tri 7994 13943 7997 13946 ne
rect 7997 13943 9110 13946
rect 7755 13909 7761 13943
rect 7795 13909 7801 13943
tri 7801 13937 7807 13943 nw
tri 7997 13937 8003 13943 ne
rect 7755 13868 7801 13909
rect 7755 13834 7761 13868
rect 7795 13834 7801 13868
rect 7755 13793 7801 13834
rect 7755 13759 7761 13793
rect 7795 13759 7801 13793
rect 7755 13718 7801 13759
rect 7755 13684 7761 13718
rect 7795 13684 7801 13718
rect 7755 13643 7801 13684
rect 7755 13609 7761 13643
rect 7795 13609 7801 13643
rect 7755 13568 7801 13609
rect 7755 13534 7761 13568
rect 7795 13534 7801 13568
rect 7755 13493 7801 13534
rect 7755 13459 7761 13493
rect 7795 13459 7801 13493
rect 7755 13418 7801 13459
rect 7755 13384 7761 13418
rect 7795 13384 7801 13418
rect 7755 13343 7801 13384
rect 7755 13309 7761 13343
rect 7795 13309 7801 13343
rect 7755 13268 7801 13309
rect 7755 13234 7761 13268
rect 7795 13234 7801 13268
rect 7755 13193 7801 13234
rect 7755 13159 7761 13193
rect 7795 13159 7801 13193
rect 7755 13119 7801 13159
rect 7755 13085 7761 13119
rect 7795 13085 7801 13119
rect 7755 13045 7801 13085
rect 8003 13835 9110 13943
rect 8003 13783 8053 13835
rect 8105 13783 8130 13835
rect 8182 13783 8207 13835
rect 8259 13783 8284 13835
rect 8336 13783 8361 13835
rect 8413 13783 8441 13835
rect 8493 13783 8518 13835
rect 8570 13783 8595 13835
rect 8647 13783 8672 13835
rect 8724 13783 8749 13835
rect 8801 13783 8826 13835
rect 8878 13783 8900 13835
rect 8952 13783 8975 13835
rect 9027 13783 9050 13835
rect 9102 13783 9110 13835
rect 8003 13767 9110 13783
rect 8003 13715 8053 13767
rect 8105 13715 8130 13767
rect 8182 13715 8207 13767
rect 8259 13715 8284 13767
rect 8336 13715 8361 13767
rect 8413 13715 8441 13767
rect 8493 13715 8518 13767
rect 8570 13715 8595 13767
rect 8647 13715 8672 13767
rect 8724 13715 8749 13767
rect 8801 13715 8826 13767
rect 8878 13715 8900 13767
rect 8952 13715 8975 13767
rect 9027 13715 9050 13767
rect 9102 13715 9110 13767
rect 8003 13699 9110 13715
rect 8003 13647 8053 13699
rect 8105 13647 8130 13699
rect 8182 13647 8207 13699
rect 8259 13647 8284 13699
rect 8336 13647 8361 13699
rect 8413 13647 8441 13699
rect 8493 13647 8518 13699
rect 8570 13647 8595 13699
rect 8647 13647 8672 13699
rect 8724 13647 8749 13699
rect 8801 13647 8826 13699
rect 8878 13647 8900 13699
rect 8952 13647 8975 13699
rect 9027 13647 9050 13699
rect 9102 13647 9110 13699
rect 8003 13631 9110 13647
rect 8003 13579 8053 13631
rect 8105 13579 8130 13631
rect 8182 13579 8207 13631
rect 8259 13579 8284 13631
rect 8336 13579 8361 13631
rect 8413 13579 8441 13631
rect 8493 13579 8518 13631
rect 8570 13579 8595 13631
rect 8647 13579 8672 13631
rect 8724 13579 8749 13631
rect 8801 13579 8826 13631
rect 8878 13579 8900 13631
rect 8952 13579 8975 13631
rect 9027 13579 9050 13631
rect 9102 13579 9110 13631
rect 8003 13563 9110 13579
rect 8003 13511 8053 13563
rect 8105 13511 8130 13563
rect 8182 13511 8207 13563
rect 8259 13511 8284 13563
rect 8336 13511 8361 13563
rect 8413 13511 8441 13563
rect 8493 13511 8518 13563
rect 8570 13511 8595 13563
rect 8647 13511 8672 13563
rect 8724 13511 8749 13563
rect 8801 13511 8826 13563
rect 8878 13511 8900 13563
rect 8952 13511 8975 13563
rect 9027 13511 9050 13563
rect 9102 13511 9110 13563
rect 7755 13011 7761 13045
rect 7795 13011 7801 13045
rect 7895 13073 7947 13079
tri 7801 13011 7818 13028 sw
tri 7878 13011 7895 13028 se
rect 7895 13011 7947 13021
rect 7755 13003 7818 13011
tri 7818 13003 7826 13011 sw
tri 7870 13003 7878 13011 se
rect 7878 13009 7947 13011
rect 7878 13003 7895 13009
rect 7755 12971 7829 13003
rect 7755 12937 7761 12971
rect 7795 12951 7829 12971
rect 7830 12952 7831 13002
rect 7867 12952 7868 13002
rect 7869 12957 7895 13003
rect 7869 12951 7947 12957
rect 7795 12937 7812 12951
tri 7812 12937 7826 12951 nw
rect 7755 12929 7804 12937
tri 7804 12929 7812 12937 nw
rect 7755 12897 7801 12929
tri 7801 12926 7804 12929 nw
rect 7755 12863 7761 12897
rect 7795 12863 7801 12897
rect 7755 12823 7801 12863
rect 7755 12789 7761 12823
rect 7795 12789 7801 12823
rect 7755 12749 7801 12789
rect 7755 12715 7761 12749
rect 7795 12715 7801 12749
rect 7755 12675 7801 12715
rect 7755 12641 7761 12675
rect 7795 12641 7801 12675
rect 7755 12601 7801 12641
rect 7755 12567 7761 12601
rect 7795 12567 7801 12601
rect 7755 12527 7801 12567
rect 7755 12493 7761 12527
rect 7795 12493 7801 12527
rect 7755 12481 7801 12493
rect 8003 12482 9110 13511
rect 8003 12448 8015 12482
rect 8049 12448 8089 12482
rect 8123 12448 8164 12482
rect 8198 12448 8239 12482
rect 8273 12448 8314 12482
rect 8348 12448 8389 12482
rect 8423 12448 8464 12482
rect 8498 12448 8539 12482
rect 8573 12448 8614 12482
rect 8648 12448 8689 12482
rect 8723 12448 8764 12482
rect 8798 12448 8839 12482
rect 8873 12448 8914 12482
rect 8948 12448 8989 12482
rect 9023 12448 9064 12482
rect 9098 12448 9110 12482
rect 9285 14093 9331 14105
rect 9285 14059 9291 14093
rect 9325 14059 9331 14093
rect 9285 14018 9331 14059
rect 9285 13984 9291 14018
rect 9325 13984 9331 14018
rect 9285 13943 9331 13984
rect 9285 13909 9291 13943
rect 9325 13909 9331 13943
rect 9285 13868 9331 13909
rect 9285 13834 9291 13868
rect 9325 13834 9331 13868
rect 9285 13793 9331 13834
rect 9285 13759 9291 13793
rect 9325 13759 9331 13793
rect 9285 13718 9331 13759
rect 9285 13684 9291 13718
rect 9325 13684 9331 13718
rect 9285 13643 9331 13684
rect 9285 13609 9291 13643
rect 9325 13609 9331 13643
rect 9285 13568 9331 13609
rect 9285 13534 9291 13568
rect 9325 13534 9331 13568
rect 9285 13493 9331 13534
rect 9285 13459 9291 13493
rect 9325 13459 9331 13493
rect 9285 13418 9331 13459
rect 9285 13384 9291 13418
rect 9325 13384 9331 13418
rect 9285 13343 9331 13384
rect 9285 13309 9291 13343
rect 9325 13309 9331 13343
rect 9285 13268 9331 13309
rect 9285 13234 9291 13268
rect 9325 13234 9331 13268
rect 9285 13193 9331 13234
rect 9285 13159 9291 13193
rect 9325 13159 9331 13193
rect 9285 13119 9331 13159
rect 9285 13085 9291 13119
rect 9325 13085 9331 13119
rect 9285 13045 9331 13085
rect 9285 13011 9291 13045
rect 9325 13011 9331 13045
rect 9285 12971 9331 13011
rect 9285 12937 9291 12971
rect 9325 12937 9331 12971
rect 9285 12897 9331 12937
rect 9285 12863 9291 12897
rect 9325 12863 9331 12897
rect 9285 12823 9331 12863
rect 9285 12789 9291 12823
rect 9325 12789 9331 12823
rect 9285 12749 9331 12789
rect 9285 12715 9291 12749
rect 9325 12715 9331 12749
rect 9285 12675 9331 12715
rect 9285 12641 9291 12675
rect 9325 12641 9331 12675
rect 9285 12601 9331 12641
rect 9285 12567 9291 12601
rect 9325 12567 9331 12601
rect 9285 12527 9331 12567
rect 9285 12493 9291 12527
rect 9325 12493 9331 12527
rect 9285 12481 9331 12493
rect 9359 14092 9380 14126
rect 9414 14092 9459 14126
rect 9493 14092 9538 14126
rect 9572 14092 9617 14126
rect 9651 14092 9696 14126
rect 9730 14092 9775 14126
rect 9809 14092 9854 14126
rect 9888 14092 9909 14126
rect 9359 14012 9909 14092
rect 9359 13978 9397 14012
rect 9431 13978 9471 14012
rect 9505 13978 9544 14012
rect 9578 13978 9617 14012
rect 9651 13978 9690 14012
rect 9724 13978 9763 14012
rect 9797 13980 9909 14012
rect 9797 13978 9869 13980
rect 9359 13972 9869 13978
rect 9359 13908 9411 13972
tri 9411 13947 9436 13972 nw
tri 9832 13947 9857 13972 ne
rect 9857 13946 9869 13972
rect 9903 13946 9909 13980
rect 9359 13874 9365 13908
rect 9399 13874 9411 13908
rect 9510 13881 9516 13933
rect 9568 13881 9608 13933
rect 9660 13881 9700 13933
rect 9752 13881 9758 13933
rect 9857 13907 9909 13946
rect 9359 13836 9411 13874
rect 9857 13873 9869 13907
rect 9903 13873 9909 13907
rect 9359 13802 9365 13836
rect 9399 13802 9411 13836
rect 9359 13764 9411 13802
rect 9359 13730 9365 13764
rect 9399 13730 9411 13764
rect 9359 13692 9411 13730
rect 9359 13658 9365 13692
rect 9399 13658 9411 13692
rect 9359 13620 9411 13658
rect 9359 13586 9365 13620
rect 9399 13586 9411 13620
rect 9359 13547 9411 13586
rect 9359 13513 9365 13547
rect 9399 13513 9411 13547
rect 9359 13474 9411 13513
rect 9359 13440 9365 13474
rect 9399 13440 9411 13474
rect 9359 13401 9411 13440
rect 9359 13367 9365 13401
rect 9399 13367 9411 13401
rect 9359 13328 9411 13367
rect 9359 13294 9365 13328
rect 9399 13294 9411 13328
rect 9359 13255 9411 13294
rect 9359 13221 9365 13255
rect 9399 13221 9411 13255
rect 9359 13182 9411 13221
rect 9359 13148 9365 13182
rect 9399 13148 9411 13182
rect 9359 13109 9411 13148
rect 9359 13075 9365 13109
rect 9399 13075 9411 13109
rect 9359 13036 9411 13075
rect 9359 13002 9365 13036
rect 9399 13002 9411 13036
rect 9359 12963 9411 13002
rect 9359 12929 9365 12963
rect 9399 12929 9411 12963
rect 9359 12890 9411 12929
rect 9452 13827 9504 13839
rect 9452 13793 9461 13827
rect 9495 13793 9504 13827
rect 9452 13754 9504 13793
rect 9452 13720 9461 13754
rect 9495 13720 9504 13754
rect 9452 13681 9504 13720
rect 9452 13647 9461 13681
rect 9495 13647 9504 13681
rect 9452 13608 9504 13647
rect 9452 13574 9461 13608
rect 9495 13574 9504 13608
rect 9452 13535 9504 13574
rect 9452 13501 9461 13535
rect 9495 13501 9504 13535
rect 9452 13461 9504 13501
rect 9452 13449 9461 13461
rect 9495 13449 9504 13461
rect 9452 13387 9504 13397
rect 9452 13385 9461 13387
rect 9495 13385 9504 13387
rect 9452 13321 9504 13333
rect 9452 13257 9504 13269
rect 9452 13193 9504 13205
rect 9452 13131 9461 13141
rect 9495 13131 9504 13141
rect 9452 13091 9504 13131
rect 9452 13057 9461 13091
rect 9495 13057 9504 13091
rect 9452 13017 9504 13057
rect 9452 12983 9461 13017
rect 9495 12983 9504 13017
rect 9452 12943 9504 12983
rect 9452 12909 9461 12943
rect 9495 12909 9504 12943
rect 9452 12897 9504 12909
rect 9606 13827 9658 13842
rect 9606 13793 9618 13827
rect 9652 13793 9658 13827
rect 9606 13754 9658 13793
rect 9606 13720 9618 13754
rect 9652 13720 9658 13754
rect 9606 13681 9658 13720
rect 9606 13647 9618 13681
rect 9652 13647 9658 13681
rect 9606 13608 9658 13647
rect 9606 13574 9618 13608
rect 9652 13574 9658 13608
rect 9606 13535 9658 13574
rect 9606 13501 9618 13535
rect 9652 13501 9658 13535
rect 9606 13461 9658 13501
rect 9606 13427 9618 13461
rect 9652 13427 9658 13461
rect 9606 13387 9658 13427
rect 9606 13353 9618 13387
rect 9652 13353 9658 13387
rect 9606 13313 9658 13353
rect 9606 13279 9618 13313
rect 9652 13279 9658 13313
rect 9606 13239 9658 13279
rect 9606 13205 9618 13239
rect 9652 13205 9658 13239
rect 9606 13165 9658 13205
rect 9606 13131 9618 13165
rect 9652 13131 9658 13165
rect 9606 13091 9658 13131
rect 9606 13057 9618 13091
rect 9652 13057 9658 13091
rect 9606 13017 9658 13057
rect 9606 12983 9618 13017
rect 9652 12983 9658 13017
rect 9606 12943 9658 12983
rect 9606 12909 9618 12943
rect 9652 12909 9658 12943
rect 9359 12856 9365 12890
rect 9399 12856 9411 12890
rect 9359 12817 9411 12856
rect 9359 12783 9365 12817
rect 9399 12791 9411 12817
tri 9411 12791 9436 12816 sw
rect 9399 12785 9529 12791
rect 9399 12783 9483 12785
rect 9359 12751 9483 12783
rect 9517 12751 9529 12785
rect 9359 12709 9529 12751
rect 9359 12675 9453 12709
rect 9487 12675 9529 12709
rect 9359 12631 9529 12675
rect 9359 12597 9453 12631
rect 9487 12597 9529 12631
rect 9359 12553 9529 12597
rect 9359 12519 9453 12553
rect 9487 12519 9529 12553
rect 9606 12643 9658 12909
rect 9764 13827 9816 13839
rect 9764 13793 9773 13827
rect 9807 13793 9816 13827
rect 9764 13754 9816 13793
rect 9764 13720 9773 13754
rect 9807 13720 9816 13754
rect 9764 13681 9816 13720
rect 9764 13647 9773 13681
rect 9807 13647 9816 13681
rect 9764 13608 9816 13647
rect 9764 13574 9773 13608
rect 9807 13574 9816 13608
rect 9764 13535 9816 13574
rect 9764 13501 9773 13535
rect 9807 13501 9816 13535
rect 9764 13461 9816 13501
rect 9764 13449 9773 13461
rect 9807 13449 9816 13461
rect 9764 13387 9816 13397
rect 9764 13385 9773 13387
rect 9807 13385 9816 13387
rect 9764 13321 9816 13333
rect 9764 13257 9816 13269
rect 9764 13193 9816 13205
rect 9764 13131 9773 13141
rect 9807 13131 9816 13141
rect 9764 13091 9816 13131
rect 9764 13057 9773 13091
rect 9807 13057 9816 13091
rect 9764 13017 9816 13057
rect 9764 12983 9773 13017
rect 9807 12983 9816 13017
rect 9764 12943 9816 12983
rect 9764 12909 9773 12943
rect 9807 12909 9816 12943
rect 9764 12897 9816 12909
rect 9857 13834 9909 13873
rect 9857 13800 9869 13834
rect 9903 13800 9909 13834
rect 9857 13761 9909 13800
rect 9857 13727 9869 13761
rect 9903 13727 9909 13761
rect 9857 13688 9909 13727
rect 9857 13654 9869 13688
rect 9903 13654 9909 13688
rect 9857 13615 9909 13654
rect 9857 13581 9869 13615
rect 9903 13581 9909 13615
rect 9857 13542 9909 13581
rect 9857 13508 9869 13542
rect 9903 13508 9909 13542
rect 9857 13469 9909 13508
rect 9857 13435 9869 13469
rect 9903 13435 9909 13469
rect 9857 13396 9909 13435
rect 9857 13362 9869 13396
rect 9903 13362 9909 13396
rect 9857 13323 9909 13362
rect 9857 13289 9869 13323
rect 9903 13289 9909 13323
rect 9857 13250 9909 13289
rect 9857 13216 9869 13250
rect 9903 13216 9909 13250
rect 9857 13177 9909 13216
rect 9857 13143 9869 13177
rect 9903 13143 9909 13177
rect 9857 13105 9909 13143
rect 9857 13071 9869 13105
rect 9903 13071 9909 13105
rect 9857 13033 9909 13071
rect 9857 12999 9869 13033
rect 9903 12999 9909 13033
rect 9857 12961 9909 12999
rect 9857 12927 9869 12961
rect 9903 12927 9909 12961
rect 9857 12889 9909 12927
rect 9857 12855 9869 12889
rect 9903 12855 9909 12889
tri 9832 12791 9857 12816 se
rect 9857 12791 9909 12855
rect 9606 12579 9658 12591
rect 9606 12521 9658 12527
rect 9730 12785 9909 12791
rect 9730 12751 9742 12785
rect 9776 12751 9837 12785
rect 9871 12751 9909 12785
rect 9730 12709 9909 12751
rect 9730 12675 9783 12709
rect 9817 12675 9909 12709
rect 9730 12631 9909 12675
rect 9730 12597 9783 12631
rect 9817 12597 9909 12631
rect 9730 12553 9909 12597
rect 8003 12442 9110 12448
rect 9359 12475 9529 12519
rect 9359 12441 9453 12475
rect 9487 12441 9529 12475
tri 9334 12386 9359 12411 se
rect 9359 12386 9529 12441
rect 9730 12519 9783 12553
rect 9817 12519 9909 12553
rect 9730 12475 9909 12519
rect 9730 12441 9783 12475
rect 9817 12441 9909 12475
tri 9529 12386 9554 12411 sw
tri 9705 12386 9730 12411 se
rect 9730 12386 9909 12441
rect 11071 14162 11077 14194
rect 11111 14162 11117 14196
rect 11071 14122 11117 14162
rect 11071 14088 11077 14122
rect 11111 14088 11117 14122
rect 11071 14048 11117 14088
rect 11071 14014 11077 14048
rect 11111 14014 11117 14048
rect 11071 13974 11117 14014
rect 11071 13940 11077 13974
rect 11111 13940 11117 13974
rect 11071 13900 11117 13940
rect 11071 13866 11077 13900
rect 11111 13866 11117 13900
rect 11071 13826 11117 13866
rect 11071 13792 11077 13826
rect 11111 13792 11117 13826
rect 11071 13752 11117 13792
rect 11071 13718 11077 13752
rect 11111 13718 11117 13752
rect 11071 13678 11117 13718
rect 11071 13644 11077 13678
rect 11111 13644 11117 13678
rect 11071 13604 11117 13644
rect 11071 13570 11077 13604
rect 11111 13570 11117 13604
rect 11071 13530 11117 13570
rect 11071 13496 11077 13530
rect 11111 13496 11117 13530
rect 11071 13456 11117 13496
rect 11071 13422 11077 13456
rect 11111 13422 11117 13456
rect 11071 13382 11117 13422
rect 11071 13348 11077 13382
rect 11111 13348 11117 13382
rect 11071 13308 11117 13348
rect 11071 13274 11077 13308
rect 11111 13274 11117 13308
rect 11071 13234 11117 13274
rect 11071 13200 11077 13234
rect 11111 13200 11117 13234
rect 11071 13160 11117 13200
rect 11071 13126 11077 13160
rect 11111 13126 11117 13160
rect 11071 13086 11117 13126
rect 11071 13052 11077 13086
rect 11111 13052 11117 13086
rect 11071 13012 11117 13052
rect 11071 12978 11077 13012
rect 11111 12978 11117 13012
rect 11071 12938 11117 12978
rect 11071 12904 11077 12938
rect 11111 12904 11117 12938
rect 11071 12864 11117 12904
rect 11071 12830 11077 12864
rect 11111 12830 11117 12864
rect 11071 12790 11117 12830
rect 11071 12756 11077 12790
rect 11111 12756 11117 12790
rect 11071 12716 11117 12756
rect 11071 12682 11077 12716
rect 11111 12682 11117 12716
rect 11071 12642 11117 12682
rect 11071 12608 11077 12642
rect 11111 12608 11117 12642
rect 11071 12568 11117 12608
rect 11071 12534 11077 12568
rect 11111 12534 11117 12568
rect 11071 12494 11117 12534
rect 11071 12460 11077 12494
rect 11111 12460 11117 12494
rect 11071 12420 11117 12460
tri 9909 12386 9934 12411 sw
rect 11071 12386 11077 12420
rect 11111 12386 11117 12420
rect 7790 12380 10954 12386
rect 7790 12346 7802 12380
rect 7836 12346 7874 12380
rect 7908 12346 7946 12380
rect 7980 12346 8018 12380
rect 8052 12346 8090 12380
rect 8124 12346 8162 12380
rect 8196 12346 8234 12380
rect 8268 12346 8306 12380
rect 8340 12346 8378 12380
rect 8412 12346 8450 12380
rect 8484 12346 8522 12380
rect 8556 12346 8594 12380
rect 8628 12346 8666 12380
rect 8700 12346 8738 12380
rect 8772 12346 8810 12380
rect 8844 12346 8882 12380
rect 8916 12346 8954 12380
rect 8988 12346 9026 12380
rect 9060 12346 9098 12380
rect 9132 12346 9170 12380
rect 9204 12346 9242 12380
rect 9276 12346 9314 12380
rect 9348 12346 9386 12380
rect 9420 12346 9458 12380
rect 9492 12346 9530 12380
rect 9564 12346 9602 12380
rect 9636 12346 9674 12380
rect 9708 12346 9747 12380
rect 9781 12346 9820 12380
rect 9854 12346 9893 12380
rect 9927 12346 9966 12380
rect 10000 12346 10065 12380
rect 10099 12346 10141 12380
rect 10175 12346 10217 12380
rect 10251 12346 10293 12380
rect 10327 12346 10369 12380
rect 10403 12346 10446 12380
rect 10480 12346 10523 12380
rect 10557 12346 10600 12380
rect 10634 12346 10677 12380
rect 10711 12346 10754 12380
rect 10788 12346 10831 12380
rect 10865 12346 10908 12380
rect 10942 12346 10954 12380
rect 11071 12352 11117 12386
rect 7790 12340 10954 12346
tri 9868 12315 9893 12340 ne
rect 8970 12270 9100 12276
rect 7791 12175 8874 12181
rect 7791 12141 7803 12175
rect 7837 12141 7876 12175
rect 7910 12141 7949 12175
rect 7983 12141 8022 12175
rect 8056 12141 8095 12175
rect 8129 12141 8168 12175
rect 8202 12141 8241 12175
rect 8275 12141 8314 12175
rect 8348 12141 8387 12175
rect 8421 12141 8460 12175
rect 8494 12141 8533 12175
rect 8567 12141 8606 12175
rect 8640 12141 8680 12175
rect 8714 12141 8754 12175
rect 8788 12141 8828 12175
rect 8862 12141 8874 12175
rect 7791 12120 8874 12141
rect 7791 12103 8277 12120
rect 8393 12103 8874 12120
rect 7791 12069 7803 12103
rect 7837 12069 7876 12103
rect 7910 12069 7949 12103
rect 7983 12069 8022 12103
rect 8056 12069 8095 12103
rect 8129 12069 8168 12103
rect 8202 12069 8241 12103
rect 8275 12069 8277 12103
rect 8421 12069 8460 12103
rect 8494 12069 8533 12103
rect 8567 12069 8606 12103
rect 8640 12069 8680 12103
rect 8714 12069 8754 12103
rect 8788 12069 8828 12103
rect 8862 12069 8874 12103
rect 7791 12031 8277 12069
rect 8393 12031 8874 12069
rect 7791 11997 7803 12031
rect 7837 11997 7876 12031
rect 7910 11997 7949 12031
rect 7983 11997 8022 12031
rect 8056 11997 8095 12031
rect 8129 11997 8168 12031
rect 8202 11997 8241 12031
rect 8275 12004 8277 12031
rect 8275 11997 8314 12004
rect 8348 11997 8387 12004
rect 8421 11997 8460 12031
rect 8494 11997 8533 12031
rect 8567 11997 8606 12031
rect 8640 11997 8680 12031
rect 8714 11997 8754 12031
rect 8788 11997 8828 12031
rect 8862 11997 8874 12031
rect 7791 11991 8874 11997
rect 9086 12154 9100 12270
tri 7687 11723 7701 11737 sw
rect 7557 11689 7701 11723
tri 7701 11689 7735 11723 sw
rect 7557 11683 7735 11689
tri 7557 11650 7590 11683 ne
rect 7590 11650 7735 11683
tri 7735 11650 7774 11689 sw
rect 7814 11680 7820 11732
rect 7872 11680 7886 11732
rect 7938 11680 7952 11732
rect 8004 11723 8018 11732
rect 8070 11723 8084 11732
rect 8136 11723 8150 11732
rect 8202 11723 8216 11732
rect 8268 11723 8282 11732
rect 8010 11689 8018 11723
rect 8268 11689 8276 11723
rect 8004 11680 8018 11689
rect 8070 11680 8084 11689
rect 8136 11680 8150 11689
rect 8202 11680 8216 11689
rect 8268 11680 8282 11689
rect 8334 11680 8348 11732
rect 8400 11680 8414 11732
rect 8466 11680 8480 11732
rect 8532 11723 8546 11732
rect 8598 11723 8612 11732
rect 8664 11723 8677 11732
rect 8729 11723 8742 11732
rect 8538 11689 8546 11723
rect 8729 11689 8732 11723
rect 8532 11680 8546 11689
rect 8598 11680 8612 11689
rect 8664 11680 8677 11689
rect 8729 11680 8742 11689
rect 8794 11680 8807 11732
rect 8859 11680 8872 11732
rect 8924 11680 8930 11732
rect 7417 11616 7423 11637
rect 7457 11616 7469 11637
tri 7590 11616 7624 11650 ne
rect 7624 11616 7774 11650
tri 7774 11616 7808 11650 sw
rect 7417 11615 7469 11616
tri 7624 11577 7663 11616 ne
rect 7663 11610 7808 11616
tri 7808 11610 7814 11616 sw
rect 7663 11577 7814 11610
rect 7417 11543 7423 11563
rect 7457 11543 7469 11563
tri 7663 11556 7684 11577 ne
rect 7417 11541 7469 11543
rect 7417 11470 7423 11489
rect 7457 11470 7469 11489
rect 7417 11467 7469 11470
tri 6849 11431 6864 11446 sw
rect 6647 11425 6864 11431
tri 6864 11425 6870 11431 sw
rect 6647 11362 6870 11425
rect 7417 11397 7423 11415
rect 7457 11409 7469 11415
rect 7457 11397 7463 11409
tri 6647 11341 6668 11362 ne
rect 6064 8488 6076 8522
rect 6110 8488 6148 8522
rect 6182 8488 6220 8522
rect 6254 8488 6266 8522
rect 6064 5098 6266 8488
rect 6064 5064 6076 5098
rect 6110 5064 6148 5098
rect 6182 5064 6220 5098
rect 6254 5064 6266 5098
rect 5828 4193 5840 4227
rect 5874 4193 5880 4227
rect 5828 4154 5880 4193
rect 5828 4120 5840 4154
rect 5874 4120 5880 4154
rect 5828 4081 5880 4120
rect 5828 4047 5840 4081
rect 5874 4047 5880 4081
rect 6064 4052 6266 5064
rect 6366 11248 6568 11254
rect 6366 11214 6378 11248
rect 6412 11214 6450 11248
rect 6484 11214 6522 11248
rect 6556 11214 6568 11248
rect 6366 11090 6568 11214
rect 6366 11056 6378 11090
rect 6412 11056 6450 11090
rect 6484 11056 6522 11090
rect 6556 11056 6568 11090
rect 6366 9378 6568 11056
rect 6366 9344 6378 9378
rect 6412 9344 6450 9378
rect 6484 9344 6522 9378
rect 6556 9344 6568 9378
rect 6366 7666 6568 9344
rect 6366 7632 6378 7666
rect 6412 7632 6450 7666
rect 6484 7632 6522 7666
rect 6556 7632 6568 7666
rect 6366 5954 6568 7632
rect 6366 5920 6378 5954
rect 6412 5920 6450 5954
rect 6484 5920 6522 5954
rect 6556 5920 6568 5954
rect 6366 4242 6568 5920
rect 6366 4208 6378 4242
rect 6412 4208 6450 4242
rect 6484 4208 6522 4242
rect 6556 4208 6568 4242
rect 6366 4084 6568 4208
rect 5828 4008 5880 4047
rect 5828 3974 5840 4008
rect 5874 3981 5880 4008
rect 6366 4050 6378 4084
rect 6412 4050 6450 4084
rect 6484 4050 6522 4084
rect 6556 4050 6568 4084
rect 6668 10234 6870 11362
rect 6898 11362 7181 11368
rect 7183 11367 7219 11368
rect 6898 11328 6910 11362
rect 6944 11328 6990 11362
rect 7024 11328 7181 11362
rect 6898 11324 7181 11328
rect 6898 11322 7114 11324
tri 7083 11297 7108 11322 ne
rect 7108 11290 7114 11322
rect 7148 11290 7181 11324
rect 7108 11251 7181 11290
rect 7108 11217 7114 11251
rect 7148 11217 7181 11251
rect 7108 11178 7181 11217
rect 7108 11144 7114 11178
rect 7148 11144 7181 11178
rect 7108 11105 7181 11144
rect 7108 11071 7114 11105
rect 7148 11071 7181 11105
rect 6668 10200 6680 10234
rect 6714 10200 6752 10234
rect 6786 10200 6824 10234
rect 6858 10200 6870 10234
rect 6668 9849 6870 10200
rect 6668 9797 6703 9849
rect 6755 9797 6783 9849
rect 6835 9797 6870 9849
rect 6668 9783 6870 9797
rect 6668 9731 6703 9783
rect 6755 9731 6783 9783
rect 6835 9731 6870 9783
rect 6668 6810 6870 9731
rect 6668 6776 6680 6810
rect 6714 6776 6752 6810
rect 6786 6776 6824 6810
rect 6858 6776 6870 6810
rect 6668 4052 6870 6776
rect 7026 11033 7078 11045
rect 7026 10999 7032 11033
rect 7066 10999 7078 11033
rect 7026 10967 7078 10999
rect 7026 10901 7078 10915
rect 7026 10811 7078 10849
rect 7026 10777 7032 10811
rect 7066 10777 7078 10811
rect 7026 10737 7078 10777
rect 7026 10703 7032 10737
rect 7066 10703 7078 10737
rect 7026 10663 7078 10703
rect 7026 10629 7032 10663
rect 7066 10629 7078 10663
rect 7026 10589 7078 10629
rect 7026 10555 7032 10589
rect 7066 10555 7078 10589
rect 7026 10515 7078 10555
rect 7026 10481 7032 10515
rect 7066 10481 7078 10515
rect 7026 10441 7078 10481
rect 7026 10407 7032 10441
rect 7066 10407 7078 10441
rect 7026 10366 7078 10407
rect 7026 10332 7032 10366
rect 7066 10332 7078 10366
rect 7026 10291 7078 10332
rect 7026 10257 7032 10291
rect 7066 10257 7078 10291
rect 7026 10177 7078 10257
rect 7026 10143 7032 10177
rect 7066 10143 7078 10177
rect 7026 10103 7078 10143
rect 7026 10069 7032 10103
rect 7066 10069 7078 10103
rect 7026 10029 7078 10069
rect 7026 9995 7032 10029
rect 7066 9995 7078 10029
rect 7026 9955 7078 9995
rect 7026 9921 7032 9955
rect 7066 9921 7078 9955
rect 7026 9881 7078 9921
rect 7026 9847 7032 9881
rect 7066 9847 7078 9881
rect 7026 9807 7078 9847
rect 7026 9773 7032 9807
rect 7066 9773 7078 9807
rect 7026 9733 7078 9773
rect 7026 9699 7032 9733
rect 7066 9699 7078 9733
rect 7026 9659 7078 9699
rect 7026 9625 7032 9659
rect 7066 9625 7078 9659
rect 7026 9585 7078 9625
rect 7026 9551 7032 9585
rect 7066 9551 7078 9585
rect 7026 9510 7078 9551
rect 7026 9476 7032 9510
rect 7066 9476 7078 9510
rect 7026 9435 7078 9476
rect 7026 9401 7032 9435
rect 7066 9401 7078 9435
rect 7026 7609 7078 9401
rect 7026 7575 7032 7609
rect 7066 7575 7078 7609
rect 7026 7535 7078 7575
rect 7026 7501 7032 7535
rect 7066 7501 7078 7535
rect 7026 7461 7078 7501
rect 7026 7427 7032 7461
rect 7066 7427 7078 7461
rect 7026 7387 7078 7427
rect 7026 7353 7032 7387
rect 7066 7353 7078 7387
rect 7026 7313 7078 7353
rect 7026 7279 7032 7313
rect 7066 7279 7078 7313
rect 7026 7239 7078 7279
rect 7026 7205 7032 7239
rect 7066 7205 7078 7239
rect 7026 7165 7078 7205
rect 7026 7131 7032 7165
rect 7066 7131 7078 7165
rect 7026 7091 7078 7131
rect 7026 7057 7032 7091
rect 7066 7057 7078 7091
rect 7026 7043 7078 7057
rect 7026 6983 7032 6991
rect 7066 6983 7078 6991
rect 7026 6977 7078 6983
rect 7026 6908 7032 6925
rect 7066 6908 7078 6925
rect 7026 6867 7078 6908
rect 7026 6833 7032 6867
rect 7066 6833 7078 6867
rect 7026 6753 7078 6833
rect 7026 6719 7032 6753
rect 7066 6719 7078 6753
rect 7026 6679 7078 6719
rect 7026 6645 7032 6679
rect 7066 6645 7078 6679
rect 7026 6605 7078 6645
rect 7026 6571 7032 6605
rect 7066 6571 7078 6605
rect 7026 6531 7078 6571
rect 7026 6497 7032 6531
rect 7066 6497 7078 6531
rect 7026 6457 7078 6497
rect 7026 6423 7032 6457
rect 7066 6423 7078 6457
rect 7026 6383 7078 6423
rect 7026 6349 7032 6383
rect 7066 6349 7078 6383
rect 7026 6309 7078 6349
rect 7026 6275 7032 6309
rect 7066 6275 7078 6309
rect 7026 6235 7078 6275
rect 7026 6201 7032 6235
rect 7066 6201 7078 6235
rect 7026 6161 7078 6201
rect 7026 6127 7032 6161
rect 7066 6127 7078 6161
rect 7026 6086 7078 6127
rect 7026 6052 7032 6086
rect 7066 6052 7078 6086
rect 7026 6011 7078 6052
rect 7026 5977 7032 6011
rect 7066 5977 7078 6011
rect 7026 4249 7078 5977
rect 7108 11032 7181 11071
rect 7108 10998 7114 11032
rect 7148 10998 7181 11032
rect 7108 10959 7181 10998
rect 7108 10925 7114 10959
rect 7148 10925 7181 10959
rect 7108 10886 7181 10925
rect 7108 10852 7114 10886
rect 7148 10852 7181 10886
rect 7108 10813 7181 10852
rect 7108 10779 7114 10813
rect 7148 10779 7181 10813
rect 7108 10740 7181 10779
rect 7108 10706 7114 10740
rect 7148 10706 7181 10740
rect 7108 10667 7181 10706
rect 7108 10633 7114 10667
rect 7148 10633 7181 10667
rect 7108 10594 7181 10633
rect 7108 10560 7114 10594
rect 7148 10560 7181 10594
rect 7108 10521 7181 10560
rect 7108 10487 7114 10521
rect 7148 10487 7181 10521
rect 7108 10448 7181 10487
rect 7108 10414 7114 10448
rect 7148 10414 7181 10448
rect 7108 10375 7181 10414
rect 7108 10341 7114 10375
rect 7148 10341 7181 10375
rect 7108 10302 7181 10341
rect 7108 10268 7114 10302
rect 7148 10268 7181 10302
rect 7108 10229 7181 10268
rect 7108 10195 7114 10229
rect 7148 10195 7181 10229
rect 7108 10156 7181 10195
rect 7108 10122 7114 10156
rect 7148 10122 7181 10156
rect 7108 10083 7181 10122
rect 7108 10049 7114 10083
rect 7148 10049 7181 10083
rect 7108 10010 7181 10049
rect 7108 9976 7114 10010
rect 7148 9976 7181 10010
rect 7108 9937 7181 9976
rect 7108 9903 7114 9937
rect 7148 9903 7181 9937
rect 7108 9864 7181 9903
rect 7108 9830 7114 9864
rect 7148 9830 7181 9864
rect 7108 9791 7181 9830
rect 7108 9757 7114 9791
rect 7148 9757 7181 9791
rect 7108 9718 7181 9757
rect 7108 9684 7114 9718
rect 7148 9684 7181 9718
rect 7108 9645 7181 9684
rect 7108 9611 7114 9645
rect 7148 9611 7181 9645
rect 7108 9572 7181 9611
rect 7108 9538 7114 9572
rect 7148 9538 7181 9572
rect 7108 9499 7181 9538
rect 7108 9465 7114 9499
rect 7148 9465 7181 9499
rect 7108 9426 7181 9465
rect 7108 9392 7114 9426
rect 7148 9392 7181 9426
rect 7108 9353 7181 9392
rect 7108 9319 7114 9353
rect 7148 9319 7181 9353
rect 7108 9280 7181 9319
rect 7108 9246 7114 9280
rect 7148 9246 7181 9280
rect 7108 9207 7181 9246
rect 7108 9173 7114 9207
rect 7148 9173 7181 9207
rect 7108 9134 7181 9173
rect 7108 9100 7114 9134
rect 7148 9100 7181 9134
rect 7108 9061 7181 9100
rect 7108 9027 7114 9061
rect 7148 9027 7181 9061
rect 7108 8988 7181 9027
rect 7108 8954 7114 8988
rect 7148 8954 7181 8988
rect 7108 8915 7181 8954
rect 7108 8881 7114 8915
rect 7148 8881 7181 8915
rect 7108 8842 7181 8881
rect 7108 8808 7114 8842
rect 7148 8808 7181 8842
rect 7108 8769 7181 8808
rect 7108 8735 7114 8769
rect 7148 8735 7181 8769
rect 7108 8696 7181 8735
rect 7108 8662 7114 8696
rect 7148 8662 7181 8696
rect 7108 8623 7181 8662
rect 7108 8589 7114 8623
rect 7148 8589 7181 8623
rect 7108 8550 7181 8589
rect 7108 8516 7114 8550
rect 7148 8516 7181 8550
rect 7108 8477 7181 8516
rect 7108 8443 7114 8477
rect 7148 8443 7181 8477
rect 7108 8404 7181 8443
rect 7108 8370 7114 8404
rect 7148 8370 7181 8404
rect 7108 8331 7181 8370
rect 7108 8297 7114 8331
rect 7148 8297 7181 8331
rect 7108 8258 7181 8297
rect 7108 8224 7114 8258
rect 7148 8224 7181 8258
rect 7108 8185 7181 8224
rect 7108 8151 7114 8185
rect 7148 8151 7181 8185
rect 7108 8112 7181 8151
rect 7108 8078 7114 8112
rect 7148 8078 7181 8112
rect 7108 8040 7181 8078
rect 7108 8006 7114 8040
rect 7148 8006 7181 8040
rect 7108 7968 7181 8006
rect 7108 7934 7114 7968
rect 7148 7934 7181 7968
rect 7108 7896 7181 7934
rect 7108 7862 7114 7896
rect 7148 7862 7181 7896
rect 7108 7824 7181 7862
rect 7108 7790 7114 7824
rect 7148 7790 7181 7824
rect 7108 7752 7181 7790
rect 7108 7718 7114 7752
rect 7148 7718 7181 7752
rect 7108 7680 7181 7718
rect 7108 7646 7114 7680
rect 7148 7646 7181 7680
rect 7108 7608 7181 7646
rect 7108 7574 7114 7608
rect 7148 7574 7181 7608
rect 7108 7536 7181 7574
rect 7108 7502 7114 7536
rect 7148 7502 7181 7536
rect 7108 7464 7181 7502
rect 7108 7430 7114 7464
rect 7148 7430 7181 7464
rect 7108 7392 7181 7430
rect 7108 7358 7114 7392
rect 7148 7358 7181 7392
rect 7108 7320 7181 7358
rect 7108 7286 7114 7320
rect 7148 7286 7181 7320
rect 7108 7248 7181 7286
rect 7108 7214 7114 7248
rect 7148 7214 7181 7248
rect 7108 7176 7181 7214
rect 7108 7142 7114 7176
rect 7148 7142 7181 7176
rect 7108 7104 7181 7142
rect 7108 7070 7114 7104
rect 7148 7070 7181 7104
rect 7108 7032 7181 7070
rect 7108 6998 7114 7032
rect 7148 6998 7181 7032
rect 7108 6960 7181 6998
rect 7108 6926 7114 6960
rect 7148 6926 7181 6960
rect 7108 6888 7181 6926
rect 7108 6854 7114 6888
rect 7148 6854 7181 6888
rect 7108 6816 7181 6854
rect 7108 6782 7114 6816
rect 7148 6782 7181 6816
rect 7108 6744 7181 6782
rect 7108 6710 7114 6744
rect 7148 6710 7181 6744
rect 7108 6672 7181 6710
rect 7108 6638 7114 6672
rect 7148 6638 7181 6672
rect 7108 6600 7181 6638
rect 7108 6566 7114 6600
rect 7148 6566 7181 6600
rect 7108 6528 7181 6566
rect 7108 6494 7114 6528
rect 7148 6494 7181 6528
rect 7108 6456 7181 6494
rect 7108 6422 7114 6456
rect 7148 6422 7181 6456
rect 7108 6384 7181 6422
rect 7108 6350 7114 6384
rect 7148 6350 7181 6384
rect 7108 6312 7181 6350
rect 7108 6278 7114 6312
rect 7148 6278 7181 6312
rect 7108 6240 7181 6278
rect 7108 6206 7114 6240
rect 7148 6206 7181 6240
rect 7108 6168 7181 6206
rect 7108 6134 7114 6168
rect 7148 6134 7181 6168
rect 7108 6096 7181 6134
rect 7108 6062 7114 6096
rect 7148 6062 7181 6096
rect 7108 6024 7181 6062
rect 7108 5990 7114 6024
rect 7148 5990 7181 6024
rect 7108 5952 7181 5990
rect 7108 5918 7114 5952
rect 7148 5918 7181 5952
rect 7108 5880 7181 5918
rect 7108 5846 7114 5880
rect 7148 5846 7181 5880
rect 7108 5808 7181 5846
rect 7108 5774 7114 5808
rect 7148 5774 7181 5808
rect 7108 5736 7181 5774
rect 7108 5702 7114 5736
rect 7148 5702 7181 5736
rect 7108 5664 7181 5702
rect 7108 5630 7114 5664
rect 7148 5630 7181 5664
rect 7108 5592 7181 5630
rect 7108 5558 7114 5592
rect 7148 5558 7181 5592
rect 7108 5520 7181 5558
rect 7108 5486 7114 5520
rect 7148 5486 7181 5520
rect 7108 5448 7181 5486
rect 7108 5414 7114 5448
rect 7148 5414 7181 5448
rect 7108 5376 7181 5414
rect 7108 5342 7114 5376
rect 7148 5342 7181 5376
rect 7108 5304 7181 5342
rect 7108 5270 7114 5304
rect 7148 5270 7181 5304
rect 7108 5232 7181 5270
rect 7108 5198 7114 5232
rect 7148 5198 7181 5232
rect 7108 5160 7181 5198
rect 7108 5126 7114 5160
rect 7148 5126 7181 5160
rect 7108 5088 7181 5126
rect 7108 5054 7114 5088
rect 7148 5054 7181 5088
rect 7108 5016 7181 5054
rect 7108 4982 7114 5016
rect 7148 4982 7181 5016
rect 7108 4944 7181 4982
rect 7108 4910 7114 4944
rect 7148 4910 7181 4944
rect 7108 4872 7181 4910
rect 7108 4838 7114 4872
rect 7148 4838 7181 4872
rect 7108 4800 7181 4838
rect 7108 4766 7114 4800
rect 7148 4766 7181 4800
rect 7108 4728 7181 4766
rect 7108 4694 7114 4728
rect 7148 4694 7181 4728
rect 7108 4656 7181 4694
rect 7108 4622 7114 4656
rect 7148 4622 7181 4656
rect 7108 4584 7181 4622
rect 7108 4550 7114 4584
rect 7148 4550 7181 4584
rect 7108 4512 7181 4550
rect 7108 4478 7114 4512
rect 7148 4478 7181 4512
rect 7108 4440 7181 4478
rect 7108 4406 7114 4440
rect 7148 4406 7181 4440
rect 7108 4368 7181 4406
rect 7108 4334 7114 4368
rect 7148 4334 7181 4368
rect 7108 4296 7181 4334
rect 7108 4262 7114 4296
rect 7148 4262 7181 4296
rect 7108 4224 7181 4262
rect 7108 4190 7114 4224
rect 7148 4190 7181 4224
rect 7108 4152 7181 4190
rect 7108 4118 7114 4152
rect 7148 4118 7181 4152
rect 7108 4080 7181 4118
tri 5880 3981 5900 4001 sw
tri 6346 3981 6366 4001 se
rect 6366 3981 6568 4050
rect 7108 4046 7114 4080
rect 7148 4046 7181 4080
tri 6568 3981 6588 4001 sw
tri 7088 3981 7108 4001 se
rect 7108 3981 7181 4046
rect 5874 3976 5900 3981
tri 5900 3976 5905 3981 sw
tri 6341 3976 6346 3981 se
rect 6346 3976 6588 3981
tri 6588 3976 6593 3981 sw
tri 7083 3976 7088 3981 se
rect 7088 3976 7181 3981
rect 5874 3974 6299 3976
rect 5828 3970 6299 3974
rect 5828 3936 5978 3970
rect 6012 3936 6064 3970
rect 6098 3936 6150 3970
rect 6184 3936 6237 3970
rect 6271 3936 6299 3970
rect 5790 3930 5826 3931
rect 5828 3930 6299 3936
rect 6300 3931 6301 3975
rect 6337 3931 6338 3975
rect 6339 3930 6606 3976
rect 6607 3931 6608 3975
rect 6644 3931 6645 3975
rect 6646 3970 7181 3976
rect 6646 3936 6671 3970
rect 6705 3936 6752 3970
rect 6786 3936 6833 3970
rect 6867 3936 6914 3970
rect 6948 3936 6995 3970
rect 7029 3936 7076 3970
rect 7110 3936 7181 3970
rect 6646 3930 7181 3936
rect 7182 3931 7220 11367
rect 7221 7341 7389 11368
rect 7221 7161 7266 7341
rect 7382 7161 7389 7341
rect 7221 6819 7389 7161
rect 7221 6639 7266 6819
rect 7382 6639 7389 6819
rect 7221 5638 7389 6639
rect 7221 5458 7266 5638
rect 7382 5458 7389 5638
rect 7221 4203 7389 5458
rect 7221 4023 7266 4203
rect 7382 4023 7389 4203
rect 7183 3930 7219 3931
rect 7221 3930 7389 4023
tri 6341 3909 6362 3930 ne
rect 6362 3909 6572 3930
tri 6572 3909 6593 3930 nw
tri 7234 3909 7255 3930 ne
rect 7255 3909 7389 3930
rect 3761 2060 3891 3906
tri 3891 3905 3892 3906 nw
tri 4525 3905 4526 3906 ne
tri 4503 3799 4526 3822 se
rect 4526 3799 4728 3906
tri 4728 3905 4729 3906 nw
tri 4469 3765 4503 3799 se
rect 4503 3765 4728 3799
tri 4464 3760 4469 3765 se
rect 4469 3760 4728 3765
tri 4430 3726 4464 3760 se
rect 4464 3738 4728 3760
rect 4464 3726 4716 3738
tri 4716 3726 4728 3738 nw
rect 5548 3872 5557 3906
rect 5591 3872 5600 3906
tri 6362 3905 6366 3909 ne
rect 5548 3833 5600 3872
rect 5548 3799 5557 3833
rect 5591 3799 5600 3833
tri 6343 3799 6366 3822 se
rect 6366 3799 6568 3909
tri 6568 3905 6572 3909 nw
tri 7255 3905 7259 3909 ne
rect 5548 3760 5600 3799
tri 6309 3765 6343 3799 se
rect 6343 3765 6568 3799
rect 5548 3726 5557 3760
rect 5591 3726 5600 3760
tri 6294 3750 6309 3765 se
rect 6309 3750 6568 3765
tri 6271 3727 6294 3750 se
rect 6294 3738 6568 3750
rect 6294 3727 6557 3738
tri 6557 3727 6568 3738 nw
tri 4397 3693 4430 3726 se
rect 4430 3693 4683 3726
tri 4683 3693 4716 3726 nw
tri 4391 3687 4397 3693 se
rect 4397 3687 4677 3693
tri 4677 3687 4683 3693 nw
rect 5548 3687 5600 3726
tri 6237 3693 6271 3727 se
rect 6271 3693 6523 3727
tri 6523 3693 6557 3727 nw
tri 4357 3653 4391 3687 se
rect 4391 3653 4643 3687
tri 4643 3653 4677 3687 nw
rect 5548 3653 5557 3687
rect 5591 3653 5600 3687
tri 6199 3655 6237 3693 se
rect 6237 3655 6485 3693
tri 6485 3655 6523 3693 nw
tri 4325 3621 4357 3653 se
rect 4357 3621 4611 3653
tri 4611 3621 4643 3653 nw
rect 5548 3641 5600 3653
tri 6185 3641 6199 3655 se
rect 6199 3641 6451 3655
tri 6165 3621 6185 3641 se
rect 6185 3621 6451 3641
tri 6451 3621 6485 3655 nw
tri 4295 3591 4325 3621 se
rect 4325 3591 4581 3621
tri 4581 3591 4611 3621 nw
tri 6135 3591 6165 3621 se
rect 6165 3591 6421 3621
tri 6421 3591 6451 3621 nw
tri 4287 3583 4295 3591 se
rect 4295 3583 4573 3591
tri 4573 3583 4581 3591 nw
tri 6127 3583 6135 3591 se
rect 6135 3583 6413 3591
tri 6413 3583 6421 3591 nw
tri 4253 3549 4287 3583 se
rect 4287 3549 4539 3583
tri 4539 3549 4573 3583 nw
tri 6093 3549 6127 3583 se
rect 6127 3549 6379 3583
tri 6379 3549 6413 3583 nw
tri 4240 3536 4253 3549 se
rect 4253 3536 4526 3549
tri 4526 3536 4539 3549 nw
tri 6080 3536 6093 3549 se
rect 6093 3536 6366 3549
tri 6366 3536 6379 3549 nw
tri 4238 3534 4240 3536 se
rect 4240 3534 4524 3536
tri 4524 3534 4526 3536 nw
tri 6078 3534 6080 3536 se
rect 6080 3534 6364 3536
tri 6364 3534 6366 3536 nw
tri 4231 3527 4238 3534 se
rect 4238 3527 4517 3534
tri 4517 3527 4524 3534 nw
tri 6071 3527 6078 3534 se
rect 6078 3527 6357 3534
tri 6357 3527 6364 3534 nw
tri 4215 3511 4231 3527 se
rect 4231 3511 4501 3527
tri 4501 3511 4517 3527 nw
tri 6055 3511 6071 3527 se
rect 6071 3511 6341 3527
tri 6341 3511 6357 3527 nw
tri 4181 3477 4215 3511 se
rect 4215 3477 4467 3511
tri 4467 3477 4501 3511 nw
tri 6021 3477 6055 3511 se
rect 6055 3477 6307 3511
tri 6307 3477 6341 3511 nw
tri 4166 3462 4181 3477 se
rect 4181 3462 4452 3477
tri 4452 3462 4467 3477 nw
tri 6006 3462 6021 3477 se
rect 6021 3462 6292 3477
tri 6292 3462 6307 3477 nw
tri 4144 3440 4166 3462 se
rect 4166 3440 4430 3462
tri 4430 3440 4452 3462 nw
tri 5984 3440 6006 3462 se
rect 6006 3440 6270 3462
tri 6270 3440 6292 3462 nw
tri 4143 3439 4144 3440 se
rect 4144 3439 4429 3440
tri 4429 3439 4430 3440 nw
tri 5983 3439 5984 3440 se
rect 5984 3439 6269 3440
tri 6269 3439 6270 3440 nw
tri 4133 3429 4143 3439 se
rect 4143 3429 4395 3439
rect 4133 3405 4395 3429
tri 4395 3405 4429 3439 nw
tri 5973 3429 5983 3439 se
rect 5983 3429 6235 3439
rect 5973 3405 6235 3429
tri 6235 3405 6269 3439 nw
rect 4133 3390 4380 3405
tri 4380 3390 4395 3405 nw
rect 5973 3390 6220 3405
tri 6220 3390 6235 3405 nw
rect 4133 3367 4357 3390
tri 4357 3367 4380 3390 nw
rect 4133 2864 4332 3367
tri 4332 3342 4357 3367 nw
rect 4904 3324 4910 3376
rect 4962 3324 4974 3376
rect 5026 3324 5038 3376
rect 5090 3324 5096 3376
rect 5973 3367 6197 3390
tri 6197 3367 6220 3390 nw
rect 6788 3376 6980 3382
rect 5363 3132 5619 3138
rect 4948 3069 5140 3127
tri 4923 3048 4944 3069 ne
rect 4944 3048 5140 3069
rect 5363 3098 5413 3132
rect 5447 3098 5493 3132
rect 5527 3098 5573 3132
rect 5607 3098 5619 3132
rect 5363 3092 5619 3098
rect 5363 3079 5503 3092
tri 5503 3079 5516 3092 nw
tri 4944 3044 4948 3048 ne
tri 4332 2864 4357 2889 sw
rect 4133 2604 4191 2864
tri 4191 2793 4216 2818 nw
tri 4936 2627 4948 2639 se
rect 4948 2627 5140 3048
rect 4134 2602 4190 2603
tri 4923 2614 4936 2627 se
rect 4936 2614 5140 2627
rect 3761 2026 3773 2060
rect 3807 2026 3845 2060
rect 3879 2026 3891 2060
rect 3761 1985 3891 2026
rect 3761 1951 3773 1985
rect 3807 1951 3845 1985
rect 3879 1951 3891 1985
rect 3761 1910 3891 1951
rect 3761 1876 3773 1910
rect 3807 1876 3845 1910
rect 3879 1876 3891 1910
rect 3761 1835 3891 1876
rect 3761 1801 3773 1835
rect 3807 1801 3845 1835
rect 3879 1801 3891 1835
rect 3761 1760 3891 1801
rect 3334 955 3340 1007
rect 3392 955 3404 1007
rect 3456 955 3464 1007
rect 3500 1747 3552 1759
rect 3500 1713 3506 1747
rect 3540 1713 3552 1747
rect 3500 1673 3552 1713
rect 3500 1639 3506 1673
rect 3540 1639 3552 1673
rect 3500 1599 3552 1639
rect 3500 1565 3506 1599
rect 3540 1565 3552 1599
rect 3500 1525 3552 1565
rect 3500 1491 3506 1525
rect 3540 1491 3552 1525
rect 3500 1451 3552 1491
rect 3500 1417 3506 1451
rect 3540 1417 3552 1451
rect 3500 1377 3552 1417
rect 3500 1343 3506 1377
rect 3540 1343 3552 1377
rect 3500 1303 3552 1343
rect 3500 1269 3506 1303
rect 3540 1269 3552 1303
rect 3500 1229 3552 1269
rect 3500 1195 3506 1229
rect 3540 1195 3552 1229
rect 3500 1185 3552 1195
rect 3500 1121 3506 1133
rect 3540 1121 3552 1133
rect 3500 1046 3506 1069
rect 3540 1046 3552 1069
rect 3500 1005 3552 1046
rect 3500 971 3506 1005
rect 3540 971 3552 1005
rect 3500 959 3552 971
rect 3761 1726 3773 1760
rect 3807 1726 3845 1760
rect 3879 1726 3891 1760
rect 3761 1685 3891 1726
rect 3761 1651 3773 1685
rect 3807 1651 3845 1685
rect 3879 1651 3891 1685
rect 3761 1610 3891 1651
rect 3761 1576 3773 1610
rect 3807 1576 3845 1610
rect 3879 1576 3891 1610
rect 3761 1535 3891 1576
rect 3761 1501 3773 1535
rect 3807 1501 3845 1535
rect 3879 1501 3891 1535
rect 3761 1460 3891 1501
rect 3761 1426 3773 1460
rect 3807 1426 3845 1460
rect 3879 1426 3891 1460
rect 3761 1385 3891 1426
rect 3761 1351 3773 1385
rect 3807 1351 3845 1385
rect 3879 1351 3891 1385
rect 3761 1310 3891 1351
rect 3761 1276 3773 1310
rect 3807 1276 3845 1310
rect 3879 1276 3891 1310
rect 4134 2565 4190 2566
rect 4133 2358 4191 2564
rect 4923 2556 5140 2614
tri 4923 2544 4935 2556 ne
rect 4935 2544 5140 2556
tri 4935 2532 4947 2544 ne
rect 4947 2532 5140 2544
tri 4947 2531 4948 2532 ne
tri 4191 2358 4216 2383 sw
rect 4133 2300 4291 2358
rect 4133 2279 4195 2300
tri 4195 2279 4216 2300 nw
rect 4133 1846 4191 2279
tri 4191 2275 4195 2279 nw
tri 4942 2121 4948 2127 se
rect 4948 2121 5140 2532
tri 4933 2112 4942 2121 se
rect 4942 2112 5140 2121
tri 4927 2106 4933 2112 se
rect 4933 2106 5140 2112
tri 4922 2101 4927 2106 se
rect 4927 2101 5140 2106
rect 4922 2045 5140 2101
tri 4922 2033 4934 2045 ne
rect 4934 2033 5140 2045
tri 4934 2021 4946 2033 ne
rect 4946 2021 5140 2033
tri 4946 2019 4948 2021 ne
tri 4191 1846 4216 1871 sw
rect 4133 1788 4291 1846
rect 4133 1768 4196 1788
tri 4196 1768 4216 1788 nw
rect 4133 1334 4191 1768
tri 4191 1763 4196 1768 nw
tri 4943 1610 4948 1615 se
rect 4948 1610 5140 2021
tri 4925 1592 4943 1610 se
rect 4943 1592 5140 1610
tri 4922 1589 4925 1592 se
rect 4925 1589 5140 1592
rect 4922 1533 5140 1589
tri 4922 1518 4937 1533 ne
rect 4937 1518 5140 1533
tri 4937 1510 4945 1518 ne
rect 4945 1510 5140 1518
tri 4945 1507 4948 1510 ne
tri 4191 1334 4216 1359 sw
rect 4133 1276 4291 1334
rect 3761 1235 3891 1276
rect 3761 1201 3773 1235
rect 3807 1201 3845 1235
rect 3879 1201 3891 1235
rect 3761 1160 3891 1201
rect 3761 1126 3773 1160
rect 3807 1126 3845 1160
rect 3879 1126 3891 1160
rect 3761 1085 3891 1126
rect 3761 1051 3773 1085
rect 3807 1051 3845 1085
rect 3879 1051 3891 1085
rect 3761 1010 3891 1051
rect 3761 976 3773 1010
rect 3807 976 3845 1010
rect 3879 976 3891 1010
rect 2303 892 2385 899
tri 2385 892 2392 899 nw
tri 2790 892 2797 899 ne
rect 2797 892 2897 899
tri 2897 892 2904 899 nw
rect 2303 708 2367 892
tri 2367 874 2385 892 nw
tri 2797 874 2815 892 ne
rect 2303 674 2316 708
rect 2350 674 2367 708
rect 2048 671 2167 674
tri 2167 671 2170 674 nw
rect 2048 658 2154 671
tri 2154 658 2167 671 nw
rect 2048 656 2132 658
rect 2048 622 2060 656
rect 2094 636 2132 656
tri 2132 636 2154 658 nw
rect 2303 636 2367 674
rect 2094 622 2102 636
rect 2048 606 2102 622
tri 2102 606 2132 636 nw
rect 2303 624 2316 636
rect 2350 624 2367 636
rect 2303 572 2309 624
rect 2361 572 2367 624
rect 2303 564 2367 572
rect 2303 560 2316 564
rect 2350 560 2367 564
rect 2303 508 2309 560
rect 2361 508 2367 560
rect 2559 716 2565 768
rect 2617 716 2623 768
rect 2559 704 2572 716
rect 2606 704 2623 716
rect 2559 652 2565 704
rect 2617 652 2623 704
rect 2559 624 2572 652
rect 2606 624 2623 652
rect 2559 586 2623 624
rect 2559 552 2572 586
rect 2606 552 2623 586
rect 2559 546 2623 552
rect 2815 708 2879 892
tri 2879 874 2897 892 nw
rect 3169 800 3287 812
rect 2815 674 2828 708
rect 2862 674 2879 708
rect 2815 636 2879 674
rect 2815 624 2828 636
rect 2862 624 2879 636
rect 2815 572 2821 624
rect 2873 572 2879 624
rect 2815 564 2879 572
rect 2815 560 2828 564
rect 2862 560 2879 564
rect 2815 508 2821 560
rect 2873 508 2879 560
rect 3071 716 3077 768
rect 3129 716 3135 768
rect 3169 766 3175 800
rect 3209 766 3247 800
rect 3281 766 3287 800
rect 3169 754 3287 766
tri 3219 751 3222 754 ne
rect 3222 751 3287 754
tri 3222 744 3229 751 ne
rect 3229 744 3287 751
tri 3229 730 3243 744 ne
rect 3243 730 3287 744
tri 3243 729 3244 730 ne
rect 3071 704 3084 716
rect 3118 704 3135 716
rect 3071 652 3077 704
rect 3129 652 3135 704
rect 3071 624 3084 652
rect 3118 624 3135 652
rect 3244 646 3287 730
rect 3334 771 3464 955
rect 3761 935 3891 976
rect 3761 901 3773 935
rect 3807 901 3845 935
rect 3879 901 3891 935
rect 3334 768 3462 771
tri 3462 769 3464 771 nw
rect 3500 871 3546 875
tri 3546 871 3550 875 sw
rect 3500 870 3550 871
tri 3550 870 3551 871 sw
rect 3500 863 3551 870
rect 3500 796 3506 863
rect 3540 860 3551 863
tri 3551 860 3561 870 sw
rect 3761 860 3891 901
rect 3540 848 3561 860
tri 3561 848 3573 860 sw
rect 3558 796 3570 848
rect 3622 796 3628 848
rect 3761 826 3773 860
rect 3807 826 3845 860
rect 3879 826 3891 860
rect 3500 791 3563 796
tri 3244 636 3254 646 ne
rect 3254 636 3287 646
tri 3287 636 3306 655 sw
rect 3334 652 3340 768
rect 3456 652 3462 768
rect 3500 757 3506 791
rect 3540 788 3563 791
tri 3563 788 3571 796 nw
rect 3540 785 3560 788
tri 3560 785 3563 788 nw
rect 3761 785 3891 826
rect 3931 944 4047 1247
tri 4935 1090 4948 1103 se
rect 4948 1090 5140 1510
tri 4931 1086 4935 1090 se
rect 4935 1086 5140 1090
tri 4930 1085 4931 1086 se
rect 4931 1085 5140 1086
tri 4923 1078 4930 1085 se
rect 4930 1078 5140 1085
rect 4948 1020 5140 1078
rect 5188 3036 5240 3048
rect 5188 3002 5194 3036
rect 5228 3002 5240 3036
rect 5188 2964 5240 3002
rect 5188 2930 5194 2964
rect 5228 2930 5240 2964
rect 5188 2892 5240 2930
rect 5188 2858 5194 2892
rect 5228 2858 5240 2892
rect 5188 2820 5240 2858
rect 5188 2786 5194 2820
rect 5228 2786 5240 2820
rect 5188 2748 5240 2786
rect 5188 2714 5194 2748
rect 5228 2714 5240 2748
rect 5188 2676 5240 2714
rect 5188 2642 5194 2676
rect 5228 2642 5240 2676
rect 5188 2604 5240 2642
rect 5188 2570 5194 2604
rect 5228 2570 5240 2604
rect 5188 2532 5240 2570
rect 5188 2498 5194 2532
rect 5228 2498 5240 2532
rect 5188 2459 5240 2498
rect 5188 2425 5194 2459
rect 5228 2425 5240 2459
rect 5188 2386 5240 2425
rect 5188 2352 5194 2386
rect 5228 2352 5240 2386
rect 5188 2313 5240 2352
rect 5188 2279 5194 2313
rect 5228 2279 5240 2313
rect 5188 2240 5240 2279
rect 5188 2206 5194 2240
rect 5228 2206 5240 2240
rect 5188 2167 5240 2206
rect 5188 2133 5194 2167
rect 5228 2133 5240 2167
rect 5188 2094 5240 2133
rect 5188 2060 5194 2094
rect 5228 2060 5240 2094
rect 5188 2021 5240 2060
rect 5188 1987 5194 2021
rect 5228 1987 5240 2021
rect 5188 1948 5240 1987
rect 5188 1914 5194 1948
rect 5228 1914 5240 1948
rect 5188 1875 5240 1914
rect 5188 1841 5194 1875
rect 5228 1841 5240 1875
rect 5188 1802 5240 1841
rect 5188 1768 5194 1802
rect 5228 1768 5240 1802
rect 5188 1729 5240 1768
rect 5188 1695 5194 1729
rect 5228 1695 5240 1729
rect 5188 1656 5240 1695
rect 5188 1622 5194 1656
rect 5228 1622 5240 1656
rect 5188 1583 5240 1622
rect 5188 1549 5194 1583
rect 5228 1549 5240 1583
rect 5188 1510 5240 1549
rect 5188 1476 5194 1510
rect 5228 1476 5240 1510
rect 5188 1437 5240 1476
rect 5188 1403 5194 1437
rect 5228 1403 5240 1437
rect 5188 1364 5240 1403
rect 5188 1330 5194 1364
rect 5228 1330 5240 1364
rect 5188 1291 5240 1330
rect 5188 1257 5194 1291
rect 5228 1257 5240 1291
rect 5188 1218 5240 1257
rect 5188 1185 5194 1218
rect 5228 1185 5240 1218
rect 5188 1121 5194 1133
rect 5228 1121 5240 1133
rect 5188 1055 5240 1069
rect 5363 2685 5491 3079
tri 5491 3067 5503 3079 nw
rect 5706 3048 5752 3060
rect 5706 3014 5712 3048
rect 5746 3014 5752 3048
rect 5706 3002 5752 3014
tri 5752 3002 5757 3007 sw
rect 5706 2982 5757 3002
tri 5757 2982 5777 3002 sw
rect 5706 2976 5823 2982
rect 5706 2942 5712 2976
rect 5746 2973 5823 2976
tri 5823 2973 5832 2982 sw
rect 5746 2964 5832 2973
tri 5832 2964 5841 2973 sw
rect 5746 2942 5841 2964
rect 5706 2930 5841 2942
tri 5841 2930 5875 2964 sw
tri 5801 2908 5823 2930 ne
rect 5823 2920 5875 2930
tri 5875 2920 5885 2930 sw
rect 5823 2908 5885 2920
tri 5823 2902 5829 2908 ne
rect 5829 2902 5885 2908
rect 5541 2901 5766 2902
tri 5766 2901 5767 2902 sw
tri 5829 2901 5830 2902 ne
rect 5830 2901 5885 2902
rect 5541 2896 5767 2901
rect 5541 2862 5553 2896
rect 5587 2862 5627 2896
rect 5661 2862 5701 2896
rect 5735 2892 5767 2896
tri 5767 2892 5776 2901 sw
tri 5830 2898 5833 2901 ne
rect 5735 2871 5776 2892
tri 5776 2871 5797 2892 sw
rect 5735 2862 5797 2871
rect 5541 2856 5797 2862
tri 5644 2831 5669 2856 ne
tri 5491 2685 5498 2692 sw
rect 5363 2676 5498 2685
tri 5498 2676 5507 2685 sw
rect 5363 2667 5507 2676
tri 5507 2667 5516 2676 sw
rect 5363 2661 5619 2667
rect 5363 2627 5413 2661
rect 5447 2627 5493 2661
rect 5527 2627 5573 2661
rect 5607 2627 5619 2661
rect 5363 2621 5619 2627
rect 5363 2613 5508 2621
tri 5508 2613 5516 2621 nw
rect 5363 2604 5499 2613
tri 5499 2604 5508 2613 nw
tri 4923 1017 4926 1020 ne
rect 4926 1017 5140 1020
tri 4926 1014 4929 1017 ne
rect 4929 1014 5140 1017
tri 4929 1010 4933 1014 ne
rect 4933 1010 5140 1014
tri 4933 1000 4943 1010 ne
rect 4943 1000 5140 1010
tri 4943 995 4948 1000 ne
tri 4047 944 4050 947 sw
rect 3931 942 4050 944
tri 4050 942 4052 944 sw
rect 3931 935 4052 942
tri 4052 935 4059 942 sw
rect 3931 926 4059 935
tri 4059 926 4068 935 sw
rect 3931 922 4068 926
tri 4068 922 4072 926 sw
rect 3931 864 4160 922
rect 3931 812 4854 864
rect 3931 797 4160 812
tri 4135 788 4144 797 ne
rect 4144 788 4160 797
tri 4144 785 4147 788 ne
rect 4147 785 4160 788
rect 3540 757 3546 785
tri 3546 771 3560 785 nw
rect 3500 745 3546 757
rect 3761 751 3773 785
rect 3807 751 3845 785
rect 3879 751 3891 785
tri 4147 778 4154 785 ne
rect 4154 778 4160 785
tri 4154 772 4160 778 ne
rect 3500 705 3546 717
rect 3500 671 3506 705
rect 3540 671 3546 705
tri 3487 636 3500 649 se
rect 3500 636 3546 671
tri 3254 634 3256 636 ne
rect 3256 634 3306 636
tri 3306 634 3308 636 sw
tri 3485 634 3487 636 se
rect 3487 634 3546 636
tri 3256 633 3257 634 ne
rect 3257 633 3308 634
tri 3308 633 3309 634 sw
tri 3484 633 3485 634 se
rect 3485 633 3546 634
rect 3071 586 3135 624
tri 3257 603 3287 633 ne
rect 3287 624 3309 633
tri 3309 624 3318 633 sw
tri 3475 624 3484 633 se
rect 3484 624 3506 633
rect 3287 603 3506 624
tri 3287 599 3291 603 ne
rect 3291 599 3506 603
rect 3540 599 3546 633
tri 3291 588 3302 599 ne
rect 3302 588 3546 599
tri 3490 587 3491 588 ne
rect 3491 587 3546 588
rect 3761 710 3891 751
rect 3761 676 3773 710
rect 3807 676 3845 710
rect 3879 676 3891 710
rect 3761 634 3891 676
rect 3761 600 3773 634
rect 3807 600 3845 634
rect 3879 600 3891 634
rect 3071 552 3084 586
rect 3118 552 3135 586
rect 3071 546 3135 552
rect 3256 508 3264 560
rect 3316 508 3328 560
rect 3380 508 3386 560
rect 3761 558 3891 600
rect 3761 524 3773 558
rect 3807 524 3845 558
rect 3879 524 3891 558
tri 1658 482 1681 505 sw
rect 3761 482 3891 524
rect 1612 480 1681 482
tri 1681 480 1683 482 sw
rect 1612 428 1618 480
rect 1670 428 1682 480
rect 1734 428 1740 480
rect 3761 448 3773 482
rect 3807 448 3845 482
rect 3879 448 3891 482
rect 4160 754 4443 771
rect 4160 744 4458 754
tri 4458 744 4468 754 nw
tri 4944 744 4948 748 se
rect 4948 744 5140 1000
rect 5363 899 5491 2604
tri 5491 2596 5499 2604 nw
rect 5363 783 5369 899
rect 5485 783 5491 899
rect 5522 2544 5638 2556
rect 5522 2510 5563 2544
rect 5597 2510 5638 2544
rect 5522 2471 5638 2510
rect 5522 2437 5563 2471
rect 5597 2437 5638 2471
rect 5522 2398 5638 2437
rect 5522 2364 5563 2398
rect 5597 2364 5638 2398
rect 5522 2325 5638 2364
rect 5522 2291 5563 2325
rect 5597 2291 5638 2325
rect 5522 2252 5638 2291
rect 5522 2218 5563 2252
rect 5597 2218 5638 2252
rect 5522 2179 5638 2218
rect 5522 2145 5563 2179
rect 5597 2145 5638 2179
rect 5522 2106 5638 2145
rect 5522 2072 5563 2106
rect 5597 2072 5638 2106
rect 5522 2033 5638 2072
rect 5522 1999 5563 2033
rect 5597 1999 5638 2033
rect 5522 1960 5638 1999
rect 5522 1926 5563 1960
rect 5597 1926 5638 1960
rect 5522 1887 5638 1926
rect 5522 1853 5563 1887
rect 5597 1853 5638 1887
rect 5522 1814 5638 1853
rect 5522 1780 5563 1814
rect 5597 1780 5638 1814
rect 5522 1740 5638 1780
rect 5522 1706 5563 1740
rect 5597 1706 5638 1740
rect 5522 1666 5638 1706
rect 5522 1632 5563 1666
rect 5597 1632 5638 1666
rect 5522 1592 5638 1632
rect 5522 1558 5563 1592
rect 5597 1558 5638 1592
rect 5522 1518 5638 1558
rect 5522 1484 5563 1518
rect 5597 1484 5638 1518
rect 5522 1444 5638 1484
rect 5522 1410 5563 1444
rect 5597 1410 5638 1444
rect 5522 1370 5638 1410
rect 5522 1336 5563 1370
rect 5597 1336 5638 1370
rect 5522 1296 5638 1336
rect 5522 1262 5563 1296
rect 5597 1262 5638 1296
rect 5522 1222 5638 1262
rect 5522 1188 5563 1222
rect 5597 1188 5638 1222
rect 5522 1148 5638 1188
rect 5522 1114 5563 1148
rect 5597 1114 5638 1148
rect 5522 1074 5638 1114
rect 5522 1040 5563 1074
rect 5597 1040 5638 1074
rect 5522 1000 5638 1040
rect 5522 966 5563 1000
rect 5597 966 5638 1000
rect 5522 926 5638 966
rect 5522 892 5563 926
rect 5597 892 5638 926
rect 5522 852 5638 892
rect 5522 818 5563 852
rect 5597 818 5638 852
rect 4160 730 4444 744
tri 4444 730 4458 744 nw
tri 4930 730 4944 744 se
rect 4944 730 5140 744
rect 4160 522 4443 730
tri 4443 729 4444 730 nw
tri 4929 729 4930 730 se
rect 4930 729 5140 730
tri 4923 723 4929 729 se
rect 4929 723 5140 729
tri 4538 710 4551 723 se
rect 4551 710 5140 723
tri 4532 704 4538 710 se
rect 4538 704 5140 710
rect 5522 778 5638 818
rect 5669 899 5797 2856
rect 5669 783 5675 899
rect 5791 783 5797 899
rect 5522 744 5563 778
rect 5597 744 5638 778
rect 5522 704 5638 744
tri 4520 692 4532 704 se
rect 4532 692 5140 704
tri 4486 658 4520 692 se
rect 4520 658 5140 692
tri 4484 656 4486 658 se
rect 4486 656 5140 658
rect 4484 628 5140 656
rect 4484 600 5112 628
tri 5112 600 5140 628 nw
rect 5180 692 5232 704
rect 5180 658 5192 692
rect 5226 658 5232 692
rect 5180 600 5232 658
rect 4484 598 5078 600
tri 4484 566 4516 598 ne
rect 4516 566 5078 598
tri 5078 566 5112 600 nw
rect 5180 566 5192 600
rect 5226 566 5232 600
tri 4516 558 4524 566 ne
rect 4524 558 5070 566
tri 5070 558 5078 566 nw
tri 4524 556 4526 558 ne
rect 4526 556 5068 558
tri 5068 556 5070 558 nw
tri 4526 531 4551 556 ne
rect 4551 531 5043 556
tri 5043 531 5068 556 nw
tri 4443 522 4446 525 sw
rect 4160 513 4446 522
tri 4446 513 4455 522 sw
rect 4160 510 4455 513
tri 4455 510 4458 513 sw
rect 4160 500 4458 510
tri 4458 500 4468 510 sw
rect 4160 466 4443 500
rect 5180 482 5232 566
rect 5522 670 5563 704
rect 5597 670 5638 704
rect 5522 630 5638 670
rect 5522 596 5563 630
rect 5597 596 5638 630
rect 5522 556 5638 596
rect 5522 522 5563 556
rect 5597 522 5638 556
tri 5232 482 5255 505 sw
rect 5522 482 5638 522
tri 5810 482 5833 505 se
rect 5833 482 5885 2901
rect 5973 2864 6172 3367
tri 6172 3342 6197 3367 nw
rect 6786 3324 6792 3376
rect 6844 3324 6856 3376
rect 6908 3324 6920 3376
rect 6972 3324 6980 3376
tri 6763 3318 6769 3324 ne
rect 6769 3318 6980 3324
tri 6769 3299 6788 3318 ne
tri 6763 3126 6788 3151 se
rect 6788 3068 6980 3318
tri 6763 3045 6786 3068 ne
rect 6786 3045 6980 3068
tri 6786 3043 6788 3045 ne
tri 6172 2864 6197 2889 sw
rect 5973 2605 6031 2864
tri 6031 2793 6056 2818 nw
rect 5974 2603 6030 2604
tri 6763 2614 6788 2639 se
rect 6788 2614 6980 3045
rect 5974 2566 6030 2567
rect 5973 2358 6031 2565
rect 6763 2556 6980 2614
tri 6763 2541 6778 2556 ne
rect 6778 2541 6980 2556
tri 6778 2532 6787 2541 ne
rect 6787 2532 6980 2541
tri 6787 2531 6788 2532 ne
tri 6031 2358 6056 2383 sw
rect 5973 2300 6131 2358
rect 5973 2279 6035 2300
tri 6035 2279 6056 2300 nw
rect 5973 1846 6031 2279
tri 6031 2275 6035 2279 nw
tri 6782 2121 6788 2127 se
rect 6788 2121 6980 2532
tri 6773 2112 6782 2121 se
rect 6782 2112 6980 2121
tri 6762 2101 6773 2112 se
rect 6773 2101 6980 2112
rect 6762 2045 6980 2101
tri 6762 2026 6781 2045 ne
rect 6781 2026 6980 2045
tri 6781 2022 6785 2026 ne
rect 6785 2022 6980 2026
tri 6785 2021 6786 2022 ne
rect 6786 2021 6980 2022
tri 6786 2019 6788 2021 ne
tri 6031 1846 6056 1871 sw
rect 5973 1788 6131 1846
rect 5973 1768 6036 1788
tri 6036 1768 6056 1788 nw
rect 5973 1334 6031 1768
tri 6031 1763 6036 1768 nw
tri 6783 1610 6788 1615 se
rect 6788 1610 6980 2021
tri 6762 1589 6783 1610 se
rect 6783 1589 6980 1610
rect 6762 1588 6980 1589
rect 6762 1533 6794 1588
tri 6762 1510 6785 1533 ne
rect 6785 1510 6794 1533
tri 6785 1507 6788 1510 ne
tri 6031 1334 6056 1359 sw
rect 5973 1276 6131 1334
rect 6788 1280 6794 1510
rect 6974 1280 6980 1588
tri 6775 1090 6788 1103 se
rect 6788 1090 6980 1280
tri 6771 1086 6775 1090 se
rect 6775 1086 6980 1090
tri 6770 1085 6771 1086 se
rect 6771 1085 6980 1086
tri 6763 1078 6770 1085 se
rect 6770 1078 6980 1085
rect 6788 1020 6980 1078
rect 7020 3036 7072 3048
rect 7020 3002 7032 3036
rect 7066 3002 7072 3036
rect 7020 2964 7072 3002
rect 7020 2930 7032 2964
rect 7066 2930 7072 2964
rect 7020 2892 7072 2930
rect 7020 2858 7032 2892
rect 7066 2858 7072 2892
rect 7020 2820 7072 2858
rect 7020 2786 7032 2820
rect 7066 2786 7072 2820
rect 7020 2748 7072 2786
rect 7020 2714 7032 2748
rect 7066 2714 7072 2748
rect 7020 2676 7072 2714
rect 7020 2642 7032 2676
rect 7066 2642 7072 2676
rect 7020 2604 7072 2642
rect 7020 2570 7032 2604
rect 7066 2570 7072 2604
rect 7020 2532 7072 2570
rect 7020 2498 7032 2532
rect 7066 2498 7072 2532
rect 7020 2459 7072 2498
rect 7020 2425 7032 2459
rect 7066 2425 7072 2459
rect 7020 2386 7072 2425
rect 7020 2352 7032 2386
rect 7066 2352 7072 2386
rect 7020 2313 7072 2352
rect 7020 2279 7032 2313
rect 7066 2279 7072 2313
rect 7020 2240 7072 2279
rect 7020 2206 7032 2240
rect 7066 2206 7072 2240
rect 7020 2167 7072 2206
rect 7020 2133 7032 2167
rect 7066 2133 7072 2167
rect 7020 2094 7072 2133
rect 7020 2060 7032 2094
rect 7066 2060 7072 2094
rect 7020 2021 7072 2060
rect 7020 1987 7032 2021
rect 7066 1987 7072 2021
rect 7020 1948 7072 1987
rect 7020 1914 7032 1948
rect 7066 1914 7072 1948
rect 7020 1875 7072 1914
rect 7020 1841 7032 1875
rect 7066 1841 7072 1875
rect 7020 1802 7072 1841
rect 7020 1768 7032 1802
rect 7066 1768 7072 1802
rect 7020 1729 7072 1768
rect 7020 1695 7032 1729
rect 7066 1695 7072 1729
rect 7020 1656 7072 1695
rect 7020 1622 7032 1656
rect 7066 1622 7072 1656
rect 7020 1583 7072 1622
rect 7020 1549 7032 1583
rect 7066 1549 7072 1583
rect 7020 1510 7072 1549
rect 7020 1476 7032 1510
rect 7066 1476 7072 1510
rect 7020 1437 7072 1476
rect 7020 1403 7032 1437
rect 7066 1403 7072 1437
rect 7020 1364 7072 1403
rect 7020 1330 7032 1364
rect 7066 1330 7072 1364
rect 7020 1291 7072 1330
rect 7020 1257 7032 1291
rect 7066 1257 7072 1291
rect 7020 1218 7072 1257
rect 7020 1185 7032 1218
rect 7066 1185 7072 1218
rect 7020 1121 7032 1133
rect 7066 1121 7072 1133
rect 7020 1055 7072 1069
rect 7259 2060 7389 3909
rect 7417 11359 7463 11397
rect 7417 11325 7423 11359
rect 7457 11325 7463 11359
rect 7417 11287 7463 11325
rect 7417 11253 7423 11287
rect 7457 11253 7463 11287
rect 7417 11215 7463 11253
rect 7417 11181 7423 11215
rect 7457 11181 7463 11215
rect 7417 11143 7463 11181
rect 7417 11109 7423 11143
rect 7457 11109 7463 11143
rect 7417 11071 7463 11109
rect 7417 11037 7423 11071
rect 7457 11037 7463 11071
rect 7417 10999 7463 11037
rect 7417 10965 7423 10999
rect 7457 10965 7463 10999
rect 7417 10927 7463 10965
rect 7417 10893 7423 10927
rect 7457 10893 7463 10927
rect 7417 10855 7463 10893
rect 7417 10821 7423 10855
rect 7457 10821 7463 10855
rect 7417 10783 7463 10821
rect 7417 10749 7423 10783
rect 7457 10749 7463 10783
rect 7417 10711 7463 10749
rect 7417 10677 7423 10711
rect 7457 10677 7463 10711
rect 7417 10639 7463 10677
rect 7417 10605 7423 10639
rect 7457 10605 7463 10639
rect 7417 10567 7463 10605
rect 7417 10533 7423 10567
rect 7457 10533 7463 10567
rect 7417 10495 7463 10533
rect 7417 10461 7423 10495
rect 7457 10461 7463 10495
rect 7417 10423 7463 10461
rect 7417 10389 7423 10423
rect 7457 10389 7463 10423
rect 7417 10351 7463 10389
rect 7417 10317 7423 10351
rect 7457 10317 7463 10351
rect 7417 10279 7463 10317
rect 7417 10245 7423 10279
rect 7457 10249 7463 10279
rect 7491 11279 7568 11285
rect 7491 11227 7516 11279
rect 7491 11215 7568 11227
rect 7491 11163 7516 11215
rect 7491 11151 7568 11163
rect 7491 11099 7516 11151
rect 7491 11087 7568 11099
rect 7491 11035 7516 11087
rect 7491 10274 7568 11035
tri 7491 10268 7497 10274 ne
tri 7463 10249 7469 10255 sw
rect 7457 10245 7469 10249
rect 7417 10243 7469 10245
rect 7417 10179 7423 10191
rect 7457 10179 7469 10191
rect 7417 10114 7423 10127
rect 7457 10114 7469 10127
rect 7417 10029 7423 10062
rect 7457 10056 7469 10062
rect 7457 10029 7463 10056
tri 7463 10050 7469 10056 nw
tri 7494 10034 7497 10037 se
rect 7497 10034 7568 10274
rect 7417 9991 7463 10029
rect 7417 9957 7423 9991
rect 7457 9957 7463 9991
rect 7417 9919 7463 9957
rect 7417 9885 7423 9919
rect 7457 9885 7463 9919
rect 7417 9847 7463 9885
rect 7417 9813 7423 9847
rect 7457 9813 7463 9847
rect 7417 9775 7463 9813
rect 7417 9741 7423 9775
rect 7457 9741 7463 9775
rect 7417 9703 7463 9741
rect 7417 9669 7423 9703
rect 7457 9669 7463 9703
rect 7417 9631 7463 9669
rect 7417 9597 7423 9631
rect 7457 9597 7463 9631
rect 7417 9559 7463 9597
rect 7417 9525 7423 9559
rect 7457 9525 7463 9559
rect 7417 9487 7463 9525
rect 7417 9453 7423 9487
rect 7457 9453 7463 9487
rect 7417 9415 7463 9453
rect 7417 9381 7423 9415
rect 7457 9381 7463 9415
rect 7417 9343 7463 9381
rect 7417 9309 7423 9343
rect 7457 9309 7463 9343
rect 7417 9271 7463 9309
rect 7417 9237 7423 9271
rect 7457 9237 7463 9271
rect 7417 9199 7463 9237
rect 7417 9165 7423 9199
rect 7457 9165 7463 9199
rect 7417 9127 7463 9165
rect 7417 9093 7423 9127
rect 7457 9093 7463 9127
rect 7417 9055 7463 9093
rect 7417 9021 7423 9055
rect 7457 9021 7463 9055
rect 7417 8983 7463 9021
rect 7417 8949 7423 8983
rect 7457 8949 7463 8983
rect 7417 8911 7463 8949
rect 7417 8877 7423 8911
rect 7457 8877 7463 8911
rect 7417 8839 7463 8877
rect 7417 8805 7423 8839
rect 7457 8805 7463 8839
rect 7417 8767 7463 8805
rect 7417 8733 7423 8767
rect 7457 8733 7463 8767
rect 7417 8695 7463 8733
rect 7417 8661 7423 8695
rect 7457 8661 7463 8695
rect 7417 8623 7463 8661
rect 7417 8589 7423 8623
rect 7457 8589 7463 8623
rect 7417 8551 7463 8589
rect 7417 8517 7423 8551
rect 7457 8517 7463 8551
rect 7417 8479 7463 8517
rect 7417 8445 7423 8479
rect 7457 8445 7463 8479
rect 7417 8407 7463 8445
rect 7417 8373 7423 8407
rect 7457 8373 7463 8407
rect 7417 8335 7463 8373
rect 7417 8301 7423 8335
rect 7457 8301 7463 8335
rect 7417 8263 7463 8301
rect 7417 8229 7423 8263
rect 7457 8229 7463 8263
rect 7417 8191 7463 8229
rect 7417 8157 7423 8191
rect 7457 8157 7463 8191
tri 7491 10031 7494 10034 se
rect 7494 10031 7568 10034
rect 7491 8179 7568 10031
tri 7491 8173 7497 8179 ne
rect 7417 8152 7463 8157
tri 7463 8152 7469 8158 sw
rect 7417 8146 7469 8152
rect 7417 8085 7423 8094
rect 7457 8085 7469 8094
rect 7417 8082 7469 8085
rect 7417 8017 7423 8030
rect 7457 8017 7469 8030
rect 7417 7941 7423 7965
rect 7457 7959 7469 7965
rect 7457 7941 7463 7959
tri 7463 7953 7469 7959 nw
rect 7417 7903 7463 7941
rect 7417 7869 7423 7903
rect 7457 7869 7463 7903
rect 7417 7831 7463 7869
rect 7417 7797 7423 7831
rect 7457 7797 7463 7831
rect 7417 7759 7463 7797
rect 7417 7725 7423 7759
rect 7457 7725 7463 7759
rect 7417 7687 7463 7725
rect 7417 7653 7423 7687
rect 7457 7653 7463 7687
rect 7417 7615 7463 7653
rect 7417 7581 7423 7615
rect 7457 7581 7463 7615
rect 7417 7543 7463 7581
rect 7417 7509 7423 7543
rect 7457 7509 7463 7543
rect 7417 7471 7463 7509
rect 7417 7437 7423 7471
rect 7457 7437 7463 7471
rect 7417 7399 7463 7437
rect 7417 7365 7423 7399
rect 7457 7365 7463 7399
rect 7417 7327 7463 7365
rect 7417 7293 7423 7327
rect 7457 7293 7463 7327
rect 7417 7255 7463 7293
rect 7417 7221 7423 7255
rect 7457 7221 7463 7255
rect 7417 7183 7463 7221
rect 7417 7149 7423 7183
rect 7457 7149 7463 7183
rect 7417 7111 7463 7149
rect 7417 7077 7423 7111
rect 7457 7077 7463 7111
rect 7417 7039 7463 7077
rect 7417 7005 7423 7039
rect 7457 7005 7463 7039
rect 7417 6967 7463 7005
rect 7417 6933 7423 6967
rect 7457 6933 7463 6967
rect 7417 6895 7463 6933
rect 7417 6861 7423 6895
rect 7457 6861 7463 6895
rect 7417 6823 7463 6861
rect 7417 6789 7423 6823
rect 7457 6789 7463 6823
rect 7417 6751 7463 6789
rect 7417 6717 7423 6751
rect 7457 6717 7463 6751
rect 7417 6679 7463 6717
rect 7417 6645 7423 6679
rect 7457 6645 7463 6679
rect 7417 6607 7463 6645
rect 7417 6573 7423 6607
rect 7457 6573 7463 6607
rect 7417 6535 7463 6573
rect 7417 6501 7423 6535
rect 7457 6501 7463 6535
rect 7417 6463 7463 6501
rect 7417 6429 7423 6463
rect 7457 6429 7463 6463
rect 7417 6391 7463 6429
rect 7417 6357 7423 6391
rect 7457 6357 7463 6391
rect 7417 6319 7463 6357
rect 7417 6285 7423 6319
rect 7457 6285 7463 6319
rect 7417 6247 7463 6285
rect 7417 6213 7423 6247
rect 7457 6213 7463 6247
rect 7417 6175 7463 6213
rect 7417 6141 7423 6175
rect 7457 6141 7463 6175
rect 7417 6103 7463 6141
rect 7417 6069 7423 6103
rect 7457 6069 7463 6103
rect 7417 6031 7463 6069
rect 7417 5997 7423 6031
rect 7457 5997 7463 6031
rect 7417 5959 7463 5997
rect 7417 5925 7423 5959
rect 7457 5925 7463 5959
rect 7417 5887 7463 5925
rect 7417 5853 7423 5887
rect 7457 5853 7463 5887
rect 7417 5815 7463 5853
rect 7417 5781 7423 5815
rect 7457 5781 7463 5815
rect 7417 5743 7463 5781
rect 7417 5709 7423 5743
rect 7457 5709 7463 5743
rect 7417 5671 7463 5709
rect 7417 5637 7423 5671
rect 7457 5637 7463 5671
rect 7417 5599 7463 5637
rect 7417 5565 7423 5599
rect 7457 5565 7463 5599
rect 7417 5527 7463 5565
rect 7417 5493 7423 5527
rect 7457 5493 7463 5527
rect 7417 5455 7463 5493
rect 7417 5421 7423 5455
rect 7457 5421 7463 5455
rect 7417 5383 7463 5421
rect 7417 5349 7423 5383
rect 7457 5349 7463 5383
rect 7417 5311 7463 5349
rect 7417 5277 7423 5311
rect 7457 5277 7463 5311
rect 7417 5239 7463 5277
rect 7417 5205 7423 5239
rect 7457 5205 7463 5239
rect 7417 5167 7463 5205
rect 7417 5133 7423 5167
rect 7457 5133 7463 5167
rect 7417 5095 7463 5133
rect 7417 5061 7423 5095
rect 7457 5061 7463 5095
rect 7417 5023 7463 5061
rect 7417 4989 7423 5023
rect 7457 4989 7463 5023
rect 7417 4951 7463 4989
rect 7417 4917 7423 4951
rect 7457 4917 7463 4951
rect 7417 4886 7463 4917
tri 7491 7934 7497 7940 se
rect 7497 7934 7568 8179
rect 7491 4914 7568 7934
rect 7596 11228 7648 11240
rect 7596 11194 7608 11228
rect 7642 11194 7648 11228
rect 7596 11154 7648 11194
rect 7596 11120 7608 11154
rect 7642 11120 7648 11154
rect 7596 11080 7648 11120
rect 7596 11046 7608 11080
rect 7642 11046 7648 11080
rect 7596 11006 7648 11046
rect 7596 10972 7608 11006
rect 7642 10972 7648 11006
rect 7596 10932 7648 10972
rect 7596 10898 7608 10932
rect 7642 10898 7648 10932
rect 7596 10858 7648 10898
rect 7596 10824 7608 10858
rect 7642 10824 7648 10858
rect 7596 10784 7648 10824
rect 7596 10750 7608 10784
rect 7642 10750 7648 10784
rect 7596 10710 7648 10750
rect 7596 10676 7608 10710
rect 7642 10676 7648 10710
rect 7596 10636 7648 10676
rect 7596 10602 7608 10636
rect 7642 10602 7648 10636
rect 7596 10561 7648 10602
rect 7596 10527 7608 10561
rect 7642 10527 7648 10561
rect 7596 10486 7648 10527
rect 7596 10452 7608 10486
rect 7642 10452 7648 10486
rect 7596 10142 7648 10452
rect 7596 10108 7608 10142
rect 7642 10108 7648 10142
rect 7596 10068 7648 10108
rect 7596 10034 7608 10068
rect 7642 10034 7648 10068
rect 7596 9994 7648 10034
rect 7596 9960 7608 9994
rect 7642 9960 7648 9994
rect 7596 9920 7648 9960
rect 7596 9886 7608 9920
rect 7642 9886 7648 9920
rect 7596 9849 7648 9886
rect 7596 9783 7648 9797
rect 7596 9698 7648 9731
rect 7596 9664 7608 9698
rect 7642 9664 7648 9698
rect 7596 9624 7648 9664
rect 7596 9590 7608 9624
rect 7642 9590 7648 9624
rect 7596 9550 7648 9590
rect 7596 9516 7608 9550
rect 7642 9516 7648 9550
rect 7596 9475 7648 9516
rect 7596 9441 7608 9475
rect 7642 9441 7648 9475
rect 7596 9400 7648 9441
rect 7596 9366 7608 9400
rect 7642 9366 7648 9400
rect 7596 9286 7648 9366
rect 7596 9252 7608 9286
rect 7642 9252 7648 9286
rect 7596 9212 7648 9252
rect 7596 9178 7608 9212
rect 7642 9178 7648 9212
rect 7596 9138 7648 9178
rect 7596 9104 7608 9138
rect 7642 9104 7648 9138
rect 7596 9064 7648 9104
rect 7596 9030 7608 9064
rect 7642 9030 7648 9064
rect 7596 8990 7648 9030
rect 7596 8956 7608 8990
rect 7642 8956 7648 8990
rect 7596 8916 7648 8956
rect 7596 8882 7608 8916
rect 7642 8882 7648 8916
rect 7596 8842 7648 8882
rect 7596 8808 7608 8842
rect 7642 8808 7648 8842
rect 7596 8768 7648 8808
rect 7596 8734 7608 8768
rect 7642 8734 7648 8768
rect 7596 8694 7648 8734
rect 7596 8660 7608 8694
rect 7642 8660 7648 8694
rect 7596 8619 7648 8660
rect 7596 8585 7608 8619
rect 7642 8585 7648 8619
rect 7596 8544 7648 8585
rect 7596 8510 7608 8544
rect 7642 8510 7648 8544
rect 7596 8200 7648 8510
rect 7596 8166 7608 8200
rect 7642 8166 7648 8200
rect 7596 8126 7648 8166
rect 7596 8092 7608 8126
rect 7642 8092 7648 8126
rect 7596 8052 7648 8092
rect 7596 8018 7608 8052
rect 7642 8018 7648 8052
rect 7596 7978 7648 8018
rect 7596 7944 7608 7978
rect 7642 7944 7648 7978
rect 7596 7904 7648 7944
rect 7596 7870 7608 7904
rect 7642 7870 7648 7904
rect 7596 7830 7648 7870
rect 7596 7796 7608 7830
rect 7642 7796 7648 7830
rect 7596 7756 7648 7796
rect 7596 7722 7608 7756
rect 7642 7722 7648 7756
rect 7596 7682 7648 7722
rect 7596 7648 7608 7682
rect 7642 7648 7648 7682
rect 7596 7608 7648 7648
rect 7596 7574 7608 7608
rect 7642 7574 7648 7608
rect 7596 7533 7648 7574
rect 7596 7499 7608 7533
rect 7642 7499 7648 7533
rect 7596 7458 7648 7499
rect 7596 7424 7608 7458
rect 7642 7424 7648 7458
rect 7596 7412 7648 7424
rect 7684 7763 7814 11577
rect 7684 7647 7698 7763
tri 7491 4908 7497 4914 ne
tri 7463 4886 7469 4892 sw
rect 7417 4880 7469 4886
rect 7417 4814 7469 4828
rect 7417 4756 7469 4762
rect 7417 4735 7463 4756
tri 7463 4750 7469 4756 nw
rect 7417 4701 7423 4735
rect 7457 4701 7463 4735
rect 7417 4663 7463 4701
rect 7417 4629 7423 4663
rect 7457 4629 7463 4663
rect 7417 4591 7463 4629
rect 7417 4557 7423 4591
rect 7457 4557 7463 4591
rect 7417 4519 7463 4557
rect 7417 4485 7423 4519
rect 7457 4485 7463 4519
rect 7417 4447 7463 4485
rect 7417 4413 7423 4447
rect 7457 4413 7463 4447
rect 7417 4375 7463 4413
rect 7417 4341 7423 4375
rect 7457 4341 7463 4375
rect 7417 4303 7463 4341
rect 7417 4269 7423 4303
rect 7457 4269 7463 4303
rect 7417 4231 7463 4269
rect 7417 4197 7423 4231
rect 7457 4197 7463 4231
rect 7417 4159 7463 4197
rect 7417 4125 7423 4159
rect 7457 4125 7463 4159
rect 7417 4087 7463 4125
rect 7417 4053 7423 4087
rect 7457 4053 7463 4087
rect 7417 4015 7463 4053
rect 7417 3981 7423 4015
rect 7457 3981 7463 4015
rect 7417 3943 7463 3981
rect 7417 3909 7423 3943
rect 7457 3909 7463 3943
rect 7417 3871 7463 3909
rect 7417 3837 7423 3871
rect 7457 3837 7463 3871
rect 7417 3799 7463 3837
rect 7417 3765 7423 3799
rect 7457 3765 7463 3799
rect 7417 3727 7463 3765
rect 7417 3693 7423 3727
rect 7457 3693 7463 3727
rect 7417 3655 7463 3693
rect 7417 3621 7423 3655
rect 7457 3621 7463 3655
rect 7417 3583 7463 3621
rect 7417 3549 7423 3583
rect 7457 3549 7463 3583
rect 7417 3511 7463 3549
rect 7417 3477 7423 3511
rect 7457 3477 7463 3511
rect 7417 3439 7463 3477
rect 7417 3405 7423 3439
rect 7457 3405 7463 3439
rect 7417 3367 7463 3405
rect 7417 3333 7423 3367
rect 7457 3333 7463 3367
rect 7417 3295 7463 3333
rect 7417 3261 7423 3295
rect 7457 3261 7463 3295
rect 7417 3223 7463 3261
rect 7417 3189 7423 3223
rect 7457 3189 7463 3223
rect 7417 3151 7463 3189
rect 7417 3117 7423 3151
rect 7457 3117 7463 3151
rect 7417 3079 7463 3117
rect 7417 3045 7423 3079
rect 7457 3045 7463 3079
rect 7417 3007 7463 3045
rect 7417 2973 7423 3007
rect 7457 2973 7463 3007
rect 7417 2935 7463 2973
rect 7417 2901 7423 2935
rect 7457 2901 7463 2935
rect 7417 2863 7463 2901
rect 7417 2829 7423 2863
rect 7457 2829 7463 2863
rect 7417 2791 7463 2829
rect 7417 2757 7423 2791
rect 7457 2757 7463 2791
rect 7417 2719 7463 2757
rect 7417 2685 7423 2719
rect 7457 2685 7463 2719
rect 7417 2647 7463 2685
rect 7417 2613 7423 2647
rect 7457 2613 7463 2647
rect 7417 2575 7463 2613
rect 7417 2541 7423 2575
rect 7457 2541 7463 2575
rect 7417 2503 7463 2541
rect 7417 2469 7423 2503
rect 7457 2469 7463 2503
rect 7417 2431 7463 2469
rect 7417 2397 7423 2431
rect 7457 2397 7463 2431
rect 7417 2359 7463 2397
rect 7417 2325 7423 2359
rect 7457 2325 7463 2359
rect 7417 2287 7463 2325
rect 7417 2253 7423 2287
rect 7457 2253 7463 2287
rect 7417 2215 7463 2253
rect 7417 2181 7423 2215
rect 7457 2181 7463 2215
rect 7417 2169 7463 2181
tri 7491 4729 7497 4735 se
rect 7497 4729 7568 4914
rect 7259 2026 7271 2060
rect 7305 2026 7343 2060
rect 7377 2026 7389 2060
rect 7259 1985 7389 2026
rect 7259 1951 7271 1985
rect 7305 1951 7343 1985
rect 7377 1951 7389 1985
rect 7259 1910 7389 1951
rect 7259 1876 7271 1910
rect 7305 1876 7343 1910
rect 7377 1876 7389 1910
rect 7259 1835 7389 1876
rect 7259 1801 7271 1835
rect 7305 1801 7343 1835
rect 7377 1801 7389 1835
rect 7259 1760 7389 1801
rect 7259 1726 7271 1760
rect 7305 1726 7343 1760
rect 7377 1726 7389 1760
rect 7259 1685 7389 1726
rect 7259 1651 7271 1685
rect 7305 1651 7343 1685
rect 7377 1651 7389 1685
rect 7259 1610 7389 1651
rect 7259 1588 7271 1610
rect 7305 1588 7343 1610
rect 7377 1588 7389 1610
rect 7259 1280 7266 1588
rect 7382 1280 7389 1588
rect 7259 1276 7271 1280
rect 7305 1276 7343 1280
rect 7377 1276 7389 1280
rect 7259 1235 7389 1276
rect 7259 1201 7271 1235
rect 7305 1201 7343 1235
rect 7377 1201 7389 1235
tri 7490 1229 7491 1230 se
rect 7491 1229 7568 4729
rect 7596 6468 7648 6480
rect 7596 6434 7608 6468
rect 7642 6434 7648 6468
rect 7596 6392 7648 6434
rect 7596 6358 7608 6392
rect 7642 6358 7648 6392
rect 7596 6316 7648 6358
rect 7596 6282 7608 6316
rect 7642 6282 7648 6316
rect 7596 6258 7648 6282
rect 7596 6205 7608 6206
rect 7642 6205 7648 6206
rect 7596 6192 7648 6205
rect 7596 6128 7608 6140
rect 7642 6128 7648 6140
rect 7596 6085 7648 6128
rect 7596 6051 7608 6085
rect 7642 6051 7648 6085
rect 7596 6008 7648 6051
rect 7596 5974 7608 6008
rect 7642 5974 7648 6008
rect 7596 5931 7648 5974
rect 7596 5897 7608 5931
rect 7642 5897 7648 5931
rect 7596 5854 7648 5897
rect 7596 5820 7608 5854
rect 7642 5820 7648 5854
rect 7596 5777 7648 5820
rect 7596 5743 7608 5777
rect 7642 5743 7648 5777
rect 7596 5700 7648 5743
rect 7596 5666 7608 5700
rect 7642 5666 7648 5700
rect 7596 5382 7648 5666
rect 7596 5348 7608 5382
rect 7642 5348 7648 5382
rect 7596 5308 7648 5348
rect 7596 5274 7608 5308
rect 7642 5274 7648 5308
rect 7596 5234 7648 5274
rect 7596 5200 7608 5234
rect 7642 5200 7648 5234
rect 7596 5160 7648 5200
rect 7596 5126 7608 5160
rect 7642 5126 7648 5160
rect 7596 5086 7648 5126
rect 7596 5052 7608 5086
rect 7642 5052 7648 5086
rect 7596 5012 7648 5052
rect 7596 4978 7608 5012
rect 7642 4978 7648 5012
rect 7596 4938 7648 4978
rect 7596 4904 7608 4938
rect 7642 4904 7648 4938
rect 7596 4864 7648 4904
rect 7596 4830 7608 4864
rect 7642 4830 7648 4864
rect 7596 4790 7648 4830
rect 7596 4756 7608 4790
rect 7642 4756 7648 4790
rect 7596 4715 7648 4756
rect 7596 4681 7608 4715
rect 7642 4681 7648 4715
rect 7596 4640 7648 4681
rect 7596 4606 7608 4640
rect 7642 4606 7648 4640
rect 7596 4526 7648 4606
rect 7596 4492 7608 4526
rect 7642 4492 7648 4526
rect 7596 4452 7648 4492
rect 7596 4418 7608 4452
rect 7642 4418 7648 4452
rect 7596 4378 7648 4418
rect 7596 4344 7608 4378
rect 7642 4344 7648 4378
rect 7596 4304 7648 4344
rect 7596 4270 7608 4304
rect 7642 4270 7648 4304
rect 7596 4230 7648 4270
rect 7596 4196 7608 4230
rect 7642 4196 7648 4230
rect 7596 4156 7648 4196
rect 7596 4122 7608 4156
rect 7642 4122 7648 4156
rect 7596 4082 7648 4122
rect 7596 4048 7608 4082
rect 7642 4048 7648 4082
rect 7596 4008 7648 4048
rect 7596 3974 7608 4008
rect 7642 3974 7648 4008
rect 7596 3934 7648 3974
rect 7596 3900 7608 3934
rect 7642 3900 7648 3934
rect 7596 3859 7648 3900
rect 7596 3825 7608 3859
rect 7642 3825 7648 3859
rect 7596 3784 7648 3825
rect 7596 3750 7608 3784
rect 7642 3750 7648 3784
rect 7596 3440 7648 3750
rect 7596 3406 7608 3440
rect 7642 3406 7648 3440
rect 7596 3366 7648 3406
rect 7596 3332 7608 3366
rect 7642 3332 7648 3366
rect 7596 3292 7648 3332
rect 7596 3258 7608 3292
rect 7642 3258 7648 3292
rect 7596 3218 7648 3258
rect 7596 3184 7608 3218
rect 7642 3184 7648 3218
rect 7596 3144 7648 3184
rect 7596 3110 7608 3144
rect 7642 3110 7648 3144
rect 7596 3070 7648 3110
rect 7596 3036 7608 3070
rect 7642 3036 7648 3070
rect 7596 2996 7648 3036
rect 7596 2962 7608 2996
rect 7642 2962 7648 2996
rect 7596 2922 7648 2962
rect 7596 2888 7608 2922
rect 7642 2888 7648 2922
rect 7596 2848 7648 2888
rect 7596 2814 7608 2848
rect 7642 2814 7648 2848
rect 7596 2773 7648 2814
rect 7596 2739 7608 2773
rect 7642 2739 7648 2773
rect 7596 2698 7648 2739
rect 7596 2664 7608 2698
rect 7642 2664 7648 2698
rect 7596 2652 7648 2664
rect 7684 4288 7814 7647
rect 7915 11429 8914 11435
rect 7915 11251 7927 11429
rect 8537 11395 8576 11429
rect 8610 11395 8649 11429
rect 8683 11395 8722 11429
rect 8756 11395 8795 11429
rect 8829 11395 8868 11429
rect 8902 11395 8914 11429
rect 8537 11357 8914 11395
rect 8537 11323 8576 11357
rect 8610 11323 8649 11357
rect 8683 11323 8722 11357
rect 8756 11323 8795 11357
rect 8829 11323 8868 11357
rect 8902 11323 8914 11357
rect 8537 11285 8914 11323
rect 8537 11251 8576 11285
rect 8610 11251 8649 11285
rect 8683 11251 8722 11285
rect 8756 11251 8795 11285
rect 8829 11251 8868 11285
rect 8902 11251 8914 11285
rect 7915 10396 8914 11251
rect 7915 10218 7927 10396
rect 8537 10362 8576 10396
rect 8610 10362 8649 10396
rect 8683 10362 8722 10396
rect 8756 10362 8795 10396
rect 8829 10362 8868 10396
rect 8902 10362 8914 10396
rect 8537 10324 8914 10362
rect 8537 10290 8576 10324
rect 8610 10290 8649 10324
rect 8683 10290 8722 10324
rect 8756 10290 8795 10324
rect 8829 10290 8868 10324
rect 8902 10290 8914 10324
rect 8537 10252 8914 10290
rect 8537 10218 8576 10252
rect 8610 10218 8649 10252
rect 8683 10218 8722 10252
rect 8756 10218 8795 10252
rect 8829 10218 8868 10252
rect 8902 10218 8914 10252
rect 7915 9343 8914 10218
rect 7915 9309 7927 9343
rect 7961 9309 7999 9343
rect 8033 9309 8071 9343
rect 8105 9309 8143 9343
rect 8177 9309 8215 9343
rect 8249 9309 8287 9343
rect 8321 9309 8359 9343
rect 8393 9309 8431 9343
rect 8465 9309 8503 9343
rect 8537 9309 8576 9343
rect 8610 9309 8649 9343
rect 8683 9309 8722 9343
rect 8756 9309 8795 9343
rect 8829 9309 8868 9343
rect 8902 9309 8914 9343
rect 7915 8483 8914 9309
rect 7915 8449 7927 8483
rect 7961 8449 7999 8483
rect 8033 8449 8071 8483
rect 8105 8449 8143 8483
rect 8177 8449 8215 8483
rect 8249 8449 8287 8483
rect 8321 8449 8359 8483
rect 8393 8449 8431 8483
rect 8465 8449 8503 8483
rect 8537 8449 8576 8483
rect 8610 8449 8649 8483
rect 8683 8449 8722 8483
rect 8756 8449 8795 8483
rect 8829 8449 8868 8483
rect 8902 8449 8914 8483
rect 7915 8359 8914 8449
rect 7915 8253 7927 8359
rect 8537 8325 8576 8359
rect 8610 8325 8649 8359
rect 8683 8325 8722 8359
rect 8756 8325 8795 8359
rect 8829 8325 8868 8359
rect 8902 8325 8914 8359
rect 8537 8287 8914 8325
rect 8537 8253 8576 8287
rect 8610 8253 8649 8287
rect 8683 8253 8722 8287
rect 8756 8253 8795 8287
rect 8829 8253 8868 8287
rect 8902 8253 8914 8287
rect 7915 7476 8914 8253
rect 7915 7424 8664 7476
rect 8716 7424 8728 7476
rect 8780 7424 8792 7476
rect 8844 7424 8856 7476
rect 8908 7424 8914 7476
rect 7915 7401 8914 7424
rect 7915 7223 7927 7401
rect 8537 7367 8576 7401
rect 8610 7367 8649 7401
rect 8683 7367 8722 7401
rect 8756 7367 8795 7401
rect 8829 7367 8868 7401
rect 8902 7367 8914 7401
rect 8537 7329 8914 7367
rect 8537 7295 8576 7329
rect 8610 7295 8649 7329
rect 8683 7295 8722 7329
rect 8756 7295 8795 7329
rect 8829 7295 8868 7329
rect 8902 7295 8914 7329
rect 8537 7257 8914 7295
rect 8537 7223 8576 7257
rect 8610 7223 8649 7257
rect 8683 7223 8722 7257
rect 8756 7223 8795 7257
rect 8829 7223 8868 7257
rect 8902 7223 8914 7257
rect 7915 7207 8914 7223
tri 8945 6675 8970 6700 se
rect 8970 6675 9100 12154
rect 9410 12175 9865 12181
rect 9410 12141 9422 12175
rect 9456 12141 9501 12175
rect 9535 12141 9580 12175
rect 9614 12141 9659 12175
rect 9693 12141 9739 12175
rect 9773 12141 9819 12175
rect 9853 12141 9865 12175
rect 9410 12103 9865 12141
rect 9410 12069 9422 12103
rect 9456 12069 9501 12103
rect 9535 12069 9580 12103
rect 9614 12069 9659 12103
rect 9693 12069 9739 12103
rect 9773 12069 9819 12103
rect 9853 12069 9865 12103
rect 9410 12031 9865 12069
rect 9410 11997 9422 12031
rect 9456 11997 9501 12031
rect 9535 11997 9580 12031
rect 9614 11997 9659 12031
rect 9693 11997 9739 12031
rect 9773 11997 9819 12031
rect 9853 11997 9865 12031
rect 9410 11991 9865 11997
tri 9866 11920 9893 11947 se
rect 9893 11920 9939 12340
tri 9939 12315 9964 12340 nw
rect 9995 12175 10279 12181
rect 9995 12141 10007 12175
rect 10041 12141 10082 12175
rect 10116 12141 10157 12175
rect 10191 12141 10233 12175
rect 10267 12141 10279 12175
rect 9995 12103 10279 12141
rect 9995 12069 10007 12103
rect 10041 12069 10082 12103
rect 10116 12069 10157 12103
rect 10191 12069 10233 12103
rect 10267 12069 10279 12103
rect 9995 12031 10279 12069
rect 9995 11997 10007 12031
rect 10041 11997 10082 12031
rect 10116 11997 10157 12031
rect 10191 11997 10233 12031
rect 10267 11997 10279 12031
rect 9995 11991 10279 11997
rect 10471 12175 11211 12181
rect 10471 12141 10483 12175
rect 10517 12141 10558 12175
rect 10592 12141 10633 12175
rect 10667 12141 10709 12175
rect 10743 12141 10785 12175
rect 10819 12141 10861 12175
rect 10895 12141 10937 12175
rect 10971 12141 11013 12175
rect 11047 12141 11089 12175
rect 11123 12141 11165 12175
rect 11199 12141 11211 12175
rect 10471 12103 11211 12141
rect 10471 12069 10483 12103
rect 10517 12069 10558 12103
rect 10592 12069 10633 12103
rect 10667 12069 10709 12103
rect 10743 12069 10785 12103
rect 10819 12069 10861 12103
rect 10895 12069 10937 12103
rect 10971 12069 11013 12103
rect 11047 12069 11089 12103
rect 11123 12069 11165 12103
rect 11199 12069 11211 12103
rect 10471 12031 11211 12069
rect 10471 11997 10483 12031
rect 10517 11997 10558 12031
rect 10592 11997 10633 12031
rect 10667 11997 10709 12031
rect 10743 11997 10785 12031
rect 10819 11997 10861 12031
rect 10895 11997 10937 12031
rect 10971 11997 11013 12031
rect 11047 11997 11089 12031
rect 11123 11997 11165 12031
rect 11199 11997 11211 12031
rect 10471 11991 11211 11997
tri 9939 11920 9966 11947 sw
tri 9804 11858 9866 11920 se
rect 9866 11868 9890 11920
rect 9942 11868 9966 11920
rect 9866 11858 9966 11868
rect 9804 11847 9966 11858
rect 9804 11795 9890 11847
rect 9942 11836 9966 11847
tri 9966 11836 10050 11920 sw
rect 9942 11795 10050 11836
rect 9804 11773 10050 11795
tri 9779 11729 9804 11754 se
rect 9804 11729 9890 11773
rect 9335 11723 9890 11729
rect 9335 11689 9347 11723
rect 9381 11689 9427 11723
rect 9461 11689 9507 11723
rect 9541 11689 9587 11723
rect 9621 11689 9667 11723
rect 9701 11689 9747 11723
rect 9781 11689 9827 11723
rect 9861 11721 9890 11723
rect 9942 11721 10050 11773
rect 9861 11699 9899 11721
rect 9933 11699 10050 11721
rect 9861 11689 9890 11699
rect 9335 11683 9890 11689
tri 9779 11658 9804 11683 ne
rect 9804 11647 9890 11683
rect 9942 11647 10050 11699
rect 9804 11625 9899 11647
rect 9933 11625 10050 11647
rect 9804 11573 9890 11625
rect 9942 11573 10050 11625
rect 9804 11551 9899 11573
rect 9933 11551 10050 11573
rect 9804 11499 9890 11551
rect 9942 11499 10050 11551
rect 9804 11470 9899 11499
rect 9933 11470 10050 11499
rect 9804 11431 10050 11470
rect 9804 11397 9899 11431
rect 9933 11397 10050 11431
rect 9804 11358 10050 11397
rect 9804 11324 9899 11358
rect 9933 11324 10050 11358
rect 9804 11285 10050 11324
rect 9804 11251 9899 11285
rect 9933 11251 10050 11285
rect 9712 11228 9764 11240
rect 9712 11194 9718 11228
rect 9752 11194 9764 11228
rect 9712 11154 9764 11194
rect 9712 11120 9718 11154
rect 9752 11120 9764 11154
rect 9712 11080 9764 11120
rect 9712 11046 9718 11080
rect 9752 11046 9764 11080
rect 9712 11006 9764 11046
rect 9712 10972 9718 11006
rect 9752 10972 9764 11006
rect 9712 10932 9764 10972
rect 9712 10898 9718 10932
rect 9752 10898 9764 10932
rect 9712 10858 9764 10898
rect 9712 10824 9718 10858
rect 9752 10824 9764 10858
rect 9712 10784 9764 10824
rect 9712 10750 9718 10784
rect 9752 10750 9764 10784
rect 9712 10710 9764 10750
rect 9712 10676 9718 10710
rect 9752 10676 9764 10710
rect 9712 10636 9764 10676
rect 9712 10602 9718 10636
rect 9752 10602 9764 10636
rect 9712 10561 9764 10602
rect 9712 10527 9718 10561
rect 9752 10527 9764 10561
rect 9712 10486 9764 10527
rect 9712 10452 9718 10486
rect 9752 10452 9764 10486
rect 9712 10142 9764 10452
rect 9712 10108 9718 10142
rect 9752 10108 9764 10142
rect 9712 10068 9764 10108
rect 9712 10034 9718 10068
rect 9752 10034 9764 10068
rect 9712 9994 9764 10034
rect 9712 9960 9718 9994
rect 9752 9960 9764 9994
rect 9712 9920 9764 9960
rect 9712 9886 9718 9920
rect 9752 9886 9764 9920
rect 9712 9849 9764 9886
rect 9712 9783 9764 9797
rect 9712 9698 9764 9731
rect 9712 9664 9718 9698
rect 9752 9664 9764 9698
rect 9712 9624 9764 9664
rect 9712 9590 9718 9624
rect 9752 9590 9764 9624
rect 9712 9550 9764 9590
rect 9712 9516 9718 9550
rect 9752 9516 9764 9550
rect 9712 9475 9764 9516
rect 9712 9441 9718 9475
rect 9752 9441 9764 9475
rect 9712 9400 9764 9441
rect 9712 9366 9718 9400
rect 9752 9366 9764 9400
rect 9712 9286 9764 9366
rect 9712 9252 9718 9286
rect 9752 9252 9764 9286
rect 9712 9212 9764 9252
rect 9712 9178 9718 9212
rect 9752 9178 9764 9212
rect 9712 9138 9764 9178
rect 9712 9104 9718 9138
rect 9752 9104 9764 9138
rect 9712 9064 9764 9104
rect 9712 9030 9718 9064
rect 9752 9030 9764 9064
rect 9712 8990 9764 9030
rect 9712 8956 9718 8990
rect 9752 8956 9764 8990
rect 9712 8916 9764 8956
rect 9712 8882 9718 8916
rect 9752 8882 9764 8916
rect 9712 8842 9764 8882
rect 9712 8808 9718 8842
rect 9752 8808 9764 8842
rect 9712 8768 9764 8808
rect 9712 8734 9718 8768
rect 9752 8734 9764 8768
rect 9712 8694 9764 8734
rect 9712 8660 9718 8694
rect 9752 8660 9764 8694
rect 9712 8619 9764 8660
rect 9712 8585 9718 8619
rect 9752 8585 9764 8619
rect 9712 8544 9764 8585
rect 9712 8510 9718 8544
rect 9752 8510 9764 8544
rect 9712 8200 9764 8510
rect 9712 8166 9718 8200
rect 9752 8166 9764 8200
rect 9712 8126 9764 8166
rect 9712 8092 9718 8126
rect 9752 8092 9764 8126
rect 9712 8052 9764 8092
rect 9712 8018 9718 8052
rect 9752 8018 9764 8052
rect 9712 7978 9764 8018
rect 9712 7944 9718 7978
rect 9752 7944 9764 7978
rect 9712 7904 9764 7944
rect 9712 7870 9718 7904
rect 9752 7870 9764 7904
rect 9712 7830 9764 7870
rect 9712 7796 9718 7830
rect 9752 7796 9764 7830
rect 9712 7756 9764 7796
rect 9712 7722 9718 7756
rect 9752 7722 9764 7756
rect 9712 7682 9764 7722
rect 9712 7648 9718 7682
rect 9752 7648 9764 7682
rect 9712 7608 9764 7648
rect 9712 7574 9718 7608
rect 9752 7574 9764 7608
rect 9712 7533 9764 7574
rect 9712 7499 9718 7533
rect 9752 7499 9764 7533
rect 9712 7458 9764 7499
rect 9712 7424 9718 7458
rect 9752 7424 9764 7458
rect 9712 7412 9764 7424
rect 9804 11212 10050 11251
rect 9804 11178 9899 11212
rect 9933 11178 10050 11212
rect 9804 11139 10050 11178
rect 9804 11105 9899 11139
rect 9933 11105 10050 11139
rect 9804 11066 10050 11105
rect 9804 11032 9899 11066
rect 9933 11032 10050 11066
rect 9804 10993 10050 11032
rect 9804 10959 9899 10993
rect 9933 10959 10050 10993
rect 9804 10920 10050 10959
rect 9804 10886 9899 10920
rect 9933 10886 10050 10920
rect 9804 10847 10050 10886
rect 9804 10813 9899 10847
rect 9933 10813 10050 10847
rect 9804 10774 10050 10813
rect 9804 10740 9899 10774
rect 9933 10740 10050 10774
rect 9804 10701 10050 10740
rect 9804 10667 9899 10701
rect 9933 10667 10050 10701
rect 9804 10628 10050 10667
rect 9804 10594 9899 10628
rect 9933 10594 10050 10628
rect 9804 10555 10050 10594
rect 9804 10521 9899 10555
rect 9933 10521 10050 10555
rect 9804 10482 10050 10521
rect 9804 10448 9899 10482
rect 9933 10448 10050 10482
rect 9804 10409 10050 10448
rect 9804 10375 9899 10409
rect 9933 10375 10050 10409
rect 9804 10336 10050 10375
rect 9804 10302 9899 10336
rect 9933 10302 10050 10336
rect 9804 10263 10050 10302
rect 9804 10243 9899 10263
rect 9933 10243 10050 10263
rect 10048 10127 10050 10243
rect 9804 10117 10050 10127
rect 9804 10114 9899 10117
rect 9933 10114 10050 10117
rect 9856 10062 9868 10114
rect 9920 10062 9932 10083
rect 9984 10062 9996 10114
rect 10048 10062 10050 10114
rect 9804 10044 10050 10062
rect 9804 10010 9899 10044
rect 9933 10010 10050 10044
rect 9804 9971 10050 10010
rect 9804 9937 9899 9971
rect 9933 9937 10050 9971
rect 9804 9898 10050 9937
rect 9804 9864 9899 9898
rect 9933 9864 10050 9898
rect 9804 9825 10050 9864
rect 9804 9791 9899 9825
rect 9933 9791 10050 9825
rect 9804 9752 10050 9791
rect 9804 9718 9899 9752
rect 9933 9718 10050 9752
rect 9804 9679 10050 9718
rect 9804 9645 9899 9679
rect 9933 9645 10050 9679
rect 9804 9606 10050 9645
rect 9804 9572 9899 9606
rect 9933 9572 10050 9606
rect 9804 9533 10050 9572
rect 9804 9499 9899 9533
rect 9933 9499 10050 9533
rect 9804 9460 10050 9499
rect 9804 9426 9899 9460
rect 9933 9426 10050 9460
rect 9804 9387 10050 9426
rect 9804 9353 9899 9387
rect 9933 9353 10050 9387
rect 9804 9314 10050 9353
tri 10078 9620 10090 9632 se
rect 10090 9620 10194 9632
rect 10078 9614 10194 9620
rect 10078 9485 10194 9498
rect 10130 9433 10142 9485
rect 10078 9420 10194 9433
rect 10130 9368 10142 9420
rect 10078 9362 10194 9368
tri 10078 9350 10090 9362 ne
rect 10090 9350 10194 9362
rect 9804 9280 9899 9314
rect 9933 9280 10050 9314
rect 9804 9241 10050 9280
rect 9804 9207 9899 9241
rect 9933 9207 10050 9241
rect 9804 9168 10050 9207
rect 9804 9134 9899 9168
rect 9933 9134 10050 9168
rect 9804 9095 10050 9134
rect 9804 9061 9899 9095
rect 9933 9061 10050 9095
rect 9804 9022 10050 9061
rect 9804 8988 9899 9022
rect 9933 8988 10050 9022
rect 9804 8949 10050 8988
rect 9804 8915 9899 8949
rect 9933 8915 10050 8949
rect 9804 8876 10050 8915
rect 9804 8842 9899 8876
rect 9933 8842 10050 8876
rect 9804 8803 10050 8842
rect 9804 8769 9899 8803
rect 9933 8769 10050 8803
rect 9804 8730 10050 8769
rect 9804 8696 9899 8730
rect 9933 8696 10050 8730
rect 9804 8657 10050 8696
rect 9804 8623 9899 8657
rect 9933 8623 10050 8657
rect 9804 8584 10050 8623
rect 9804 8550 9899 8584
rect 9933 8550 10050 8584
rect 9804 8511 10050 8550
rect 9804 8477 9899 8511
rect 9933 8477 10050 8511
rect 9804 8438 10050 8477
rect 9804 8404 9899 8438
rect 9933 8404 10050 8438
rect 9804 8365 10050 8404
rect 9804 8331 9899 8365
rect 9933 8331 10050 8365
rect 9804 8292 10050 8331
rect 9804 8258 9899 8292
rect 9933 8258 10050 8292
tri 10078 8546 10090 8558 se
rect 10090 8546 10194 8558
rect 10078 8540 10194 8546
rect 10130 8488 10142 8540
rect 10078 8473 10194 8488
rect 10130 8421 10142 8473
rect 10078 8406 10194 8421
rect 10130 8354 10142 8406
rect 10078 8338 10194 8354
rect 10130 8286 10142 8338
rect 10078 8280 10194 8286
tri 10078 8268 10090 8280 ne
rect 10090 8268 10194 8280
rect 9804 8219 10050 8258
rect 9804 8185 9899 8219
rect 9933 8185 10050 8219
rect 9804 8146 10050 8185
rect 10048 8030 10050 8146
rect 9804 8017 10050 8030
rect 9856 7965 9868 8017
rect 9920 8000 9932 8017
rect 9920 7965 9932 7966
rect 9984 7965 9996 8017
rect 10048 7965 10050 8017
rect 10305 7997 10311 8049
rect 10363 7997 10376 8049
rect 10428 7997 10441 8049
rect 10493 8040 10506 8049
rect 10558 8040 10571 8049
rect 10623 8040 10636 8049
rect 10688 8040 10701 8049
rect 10753 8040 10766 8049
rect 10818 8040 10831 8049
rect 10883 8040 10896 8049
rect 10495 8006 10506 8040
rect 10567 8006 10571 8040
rect 10818 8006 10821 8040
rect 10883 8006 10893 8040
rect 10493 7997 10506 8006
rect 10558 7997 10571 8006
rect 10623 7997 10636 8006
rect 10688 7997 10701 8006
rect 10753 7997 10766 8006
rect 10818 7997 10831 8006
rect 10883 7997 10896 8006
rect 10948 7997 10961 8049
rect 11013 7997 11026 8049
rect 11078 7997 11091 8049
rect 11143 7997 11156 8049
rect 11208 8040 11221 8049
rect 11273 8040 11286 8049
rect 11338 8040 11350 8049
rect 11402 8040 11414 8049
rect 11466 8040 11478 8049
rect 11530 8040 11542 8049
rect 11215 8006 11221 8040
rect 11466 8006 11469 8040
rect 11530 8006 11541 8040
rect 11208 7997 11221 8006
rect 11273 7997 11286 8006
rect 11338 7997 11350 8006
rect 11402 7997 11414 8006
rect 11466 7997 11478 8006
rect 11530 7997 11542 8006
rect 11594 7997 11606 8049
rect 11658 7997 11670 8049
rect 11722 7997 11734 8049
rect 11786 8040 11798 8049
rect 11850 8040 11862 8049
rect 11914 8040 11926 8049
rect 11978 8040 11990 8049
rect 12042 8040 12054 8049
rect 12106 8040 12118 8049
rect 11791 8006 11798 8040
rect 12042 8006 12045 8040
rect 12106 8006 12117 8040
rect 11786 7997 11798 8006
rect 11850 7997 11862 8006
rect 11914 7997 11926 8006
rect 11978 7997 11990 8006
rect 12042 7997 12054 8006
rect 12106 7997 12118 8006
rect 12170 7997 12182 8049
rect 12234 7997 12246 8049
rect 12298 7997 12310 8049
rect 12362 8040 12374 8049
rect 12426 8040 12438 8049
rect 12490 8040 12502 8049
rect 12554 8040 12566 8049
rect 12618 8040 12630 8049
rect 12367 8006 12374 8040
rect 12618 8006 12624 8040
rect 12362 7997 12374 8006
rect 12426 7997 12438 8006
rect 12490 7997 12502 8006
rect 12554 7997 12566 8006
rect 12618 7997 12630 8006
rect 12682 7997 12694 8049
rect 12746 7997 12758 8049
rect 12810 8023 12816 8049
tri 12816 8023 12842 8049 sw
rect 12810 7997 12842 8023
tri 12793 7974 12816 7997 ne
rect 12816 7974 12842 7997
rect 9804 7927 10050 7965
tri 12816 7948 12842 7974 ne
tri 12842 7948 12917 8023 sw
rect 9804 7893 9899 7927
rect 9933 7893 10050 7927
rect 9804 7854 10050 7893
tri 12842 7873 12917 7948 ne
tri 12917 7873 12992 7948 sw
rect 9804 7820 9899 7854
rect 9933 7820 10050 7854
rect 9804 7782 10050 7820
tri 12917 7798 12992 7873 ne
tri 12992 7798 13067 7873 sw
rect 9804 7748 9899 7782
rect 9933 7748 10050 7782
tri 12992 7775 13015 7798 ne
rect 9804 7710 10050 7748
rect 9804 7676 9899 7710
rect 9933 7676 10050 7710
rect 9804 7638 10050 7676
rect 9804 7604 9899 7638
rect 9933 7604 10050 7638
rect 9804 7566 10050 7604
rect 9804 7532 9899 7566
rect 9933 7532 10050 7566
rect 9804 7494 10050 7532
rect 9804 7460 9899 7494
rect 9933 7460 10050 7494
rect 9804 7422 10050 7460
rect 9804 7388 9899 7422
rect 9933 7388 10050 7422
rect 9804 7350 10050 7388
rect 9804 7316 9899 7350
rect 9933 7316 10050 7350
rect 9804 7278 10050 7316
rect 9804 7244 9899 7278
rect 9933 7244 10050 7278
rect 9804 7206 10050 7244
rect 9804 7172 9899 7206
rect 9933 7172 10050 7206
rect 9804 7134 10050 7172
rect 9804 7100 9899 7134
rect 9933 7100 10050 7134
rect 9804 7062 10050 7100
rect 9804 7028 9899 7062
rect 9933 7028 10050 7062
rect 9804 6990 10050 7028
rect 9804 6956 9899 6990
rect 9933 6956 10050 6990
rect 9804 6918 10050 6956
rect 9804 6884 9899 6918
rect 9933 6884 10050 6918
rect 9804 6846 10050 6884
rect 9804 6812 9899 6846
rect 9933 6812 10050 6846
rect 9804 6774 10050 6812
rect 9804 6740 9899 6774
rect 9933 6740 10050 6774
rect 9804 6702 10050 6740
tri 9100 6675 9125 6700 sw
rect 7684 4236 7692 4288
rect 7744 4236 7756 4288
rect 7808 4236 7814 4288
rect 7259 1160 7389 1201
tri 7456 1195 7490 1229 se
rect 7490 1195 7568 1229
rect 7259 1126 7271 1160
rect 7305 1126 7343 1160
rect 7377 1126 7389 1160
rect 7259 1085 7389 1126
tri 6763 1017 6766 1020 ne
rect 6766 1017 6980 1020
tri 6766 1014 6769 1017 ne
rect 6769 1014 6980 1017
tri 6769 1010 6773 1014 ne
rect 6773 1010 6980 1014
tri 6773 995 6788 1010 ne
tri 6785 944 6788 947 se
rect 6788 944 6980 1010
tri 6783 942 6785 944 se
rect 6785 942 6980 944
tri 6776 935 6783 942 se
rect 6783 935 6980 942
tri 6763 922 6776 935 se
rect 6776 922 6980 935
rect 6788 864 6980 922
rect 6059 812 6980 864
rect 6788 754 6980 812
tri 6763 751 6766 754 ne
rect 6766 751 6980 754
tri 6766 750 6767 751 ne
rect 6767 750 6980 751
tri 6767 730 6787 750 ne
rect 6787 730 6980 750
tri 6787 729 6788 730 ne
tri 6256 710 6271 725 se
rect 6271 710 6623 725
tri 6623 710 6638 725 sw
tri 6238 692 6256 710 se
rect 6256 692 6638 710
tri 6638 692 6656 710 sw
tri 6204 658 6238 692 se
rect 6238 658 6656 692
tri 6656 658 6690 692 sw
tri 6202 656 6204 658 se
rect 6204 656 6690 658
tri 6690 656 6692 658 sw
rect 6202 598 6692 656
tri 6202 586 6214 598 ne
rect 6214 586 6680 598
tri 6680 586 6692 598 nw
tri 6214 578 6222 586 ne
rect 6222 578 6672 586
tri 6672 578 6680 586 nw
tri 6222 558 6242 578 ne
rect 6242 558 6652 578
tri 6652 558 6672 578 nw
tri 6242 547 6253 558 ne
rect 6253 547 6641 558
tri 6641 547 6652 558 nw
tri 6253 533 6267 547 ne
rect 6267 533 6627 547
tri 6627 533 6641 547 nw
tri 6776 513 6788 525 se
rect 6788 513 6980 730
rect 7259 1051 7271 1085
rect 7305 1051 7343 1085
rect 7377 1051 7389 1085
tri 7452 1191 7456 1195 se
rect 7456 1191 7568 1195
rect 7452 1185 7568 1191
rect 7452 1063 7568 1069
rect 7596 1747 7648 1759
rect 7596 1713 7608 1747
rect 7642 1713 7648 1747
rect 7596 1673 7648 1713
rect 7596 1639 7608 1673
rect 7642 1639 7648 1673
rect 7596 1599 7648 1639
rect 7596 1565 7608 1599
rect 7642 1565 7648 1599
rect 7596 1525 7648 1565
rect 7596 1491 7608 1525
rect 7642 1491 7648 1525
rect 7596 1451 7648 1491
rect 7596 1417 7608 1451
rect 7642 1417 7648 1451
rect 7596 1377 7648 1417
rect 7596 1343 7608 1377
rect 7642 1343 7648 1377
rect 7596 1303 7648 1343
rect 7596 1269 7608 1303
rect 7642 1269 7648 1303
rect 7596 1229 7648 1269
rect 7596 1195 7608 1229
rect 7642 1195 7648 1229
rect 7596 1185 7648 1195
rect 7596 1121 7608 1133
rect 7642 1121 7648 1133
rect 7259 1010 7389 1051
rect 7259 976 7271 1010
rect 7305 976 7343 1010
rect 7377 976 7389 1010
rect 7259 935 7389 976
rect 7596 1046 7608 1069
rect 7642 1046 7648 1069
rect 7596 1005 7648 1046
rect 7596 971 7608 1005
rect 7642 971 7648 1005
rect 7596 959 7648 971
rect 7259 901 7271 935
rect 7305 901 7343 935
rect 7377 901 7389 935
rect 7259 860 7389 901
rect 7259 826 7271 860
rect 7305 826 7343 860
rect 7377 826 7389 860
rect 7259 785 7389 826
rect 7259 751 7271 785
rect 7305 751 7343 785
rect 7377 751 7389 785
rect 7259 710 7389 751
rect 7575 860 7633 866
rect 7575 826 7587 860
rect 7621 826 7633 860
rect 7575 788 7633 826
rect 7575 754 7587 788
rect 7621 754 7633 788
rect 7684 768 7814 4236
rect 8139 6669 9138 6675
rect 8139 6491 8151 6669
rect 8761 6635 8800 6669
rect 8834 6635 8873 6669
rect 8907 6635 8946 6669
rect 8980 6635 9019 6669
rect 9053 6635 9092 6669
rect 9126 6635 9138 6669
rect 8761 6597 9138 6635
rect 8761 6563 8800 6597
rect 8834 6563 8873 6597
rect 8907 6563 8946 6597
rect 8980 6563 9019 6597
rect 9053 6563 9092 6597
rect 9126 6563 9138 6597
rect 8761 6525 9138 6563
rect 8761 6491 8800 6525
rect 8834 6491 8873 6525
rect 8907 6491 8946 6525
rect 8980 6491 9019 6525
rect 9053 6491 9092 6525
rect 9126 6491 9138 6525
rect 8139 5610 9138 6491
rect 9804 6668 9899 6702
rect 9933 6668 10050 6702
rect 9804 6630 10050 6668
rect 9804 6596 9899 6630
rect 9933 6596 10050 6630
rect 9804 6558 10050 6596
rect 9804 6524 9899 6558
rect 9933 6540 10050 6558
rect 9933 6524 10023 6540
rect 9804 6513 10023 6524
tri 10023 6513 10050 6540 nw
rect 10193 7705 12837 7711
rect 10193 7699 10277 7705
rect 10193 7665 10205 7699
rect 10239 7671 10277 7699
rect 10311 7671 10349 7705
rect 10383 7671 10421 7705
rect 10455 7671 10493 7705
rect 10527 7671 10565 7705
rect 10599 7671 10637 7705
rect 10671 7671 10709 7705
rect 10743 7671 10782 7705
rect 10816 7671 10855 7705
rect 10889 7671 10928 7705
rect 10962 7671 11001 7705
rect 11035 7671 11074 7705
rect 11108 7671 11147 7705
rect 11181 7671 11220 7705
rect 11254 7671 11293 7705
rect 11327 7671 11366 7705
rect 11400 7671 11439 7705
rect 11473 7671 11512 7705
rect 11546 7671 11585 7705
rect 11619 7671 11658 7705
rect 11692 7671 11731 7705
rect 11765 7671 11804 7705
rect 11838 7671 11877 7705
rect 11911 7671 11950 7705
rect 11984 7671 12023 7705
rect 12057 7671 12096 7705
rect 12130 7671 12169 7705
rect 12203 7671 12242 7705
rect 12276 7671 12315 7705
rect 12349 7671 12388 7705
rect 12422 7671 12461 7705
rect 12495 7671 12534 7705
rect 12568 7671 12607 7705
rect 12641 7671 12680 7705
rect 12714 7671 12753 7705
rect 12787 7672 12837 7705
tri 12837 7672 12876 7711 sw
rect 12787 7671 12876 7672
rect 10239 7665 12876 7671
rect 10193 7627 10245 7665
tri 10245 7640 10270 7665 nw
tri 12808 7640 12833 7665 ne
rect 12833 7640 12876 7665
rect 10193 7593 10205 7627
rect 10239 7593 10245 7627
tri 12833 7597 12876 7640 ne
tri 12876 7597 12951 7672 sw
rect 10193 7555 10245 7593
rect 10193 7521 10205 7555
rect 10239 7521 10245 7555
rect 10193 7483 10245 7521
rect 10193 7449 10205 7483
rect 10239 7449 10245 7483
rect 10193 7411 10245 7449
rect 10193 7377 10205 7411
rect 10239 7377 10245 7411
rect 10193 7341 10245 7377
rect 10193 7277 10245 7289
rect 10193 7213 10245 7225
rect 10193 7123 10245 7161
rect 10193 7089 10205 7123
rect 10239 7089 10245 7123
rect 10193 7051 10245 7089
rect 10193 7017 10205 7051
rect 10239 7017 10245 7051
rect 10193 6979 10245 7017
rect 10193 6945 10205 6979
rect 10239 6945 10245 6979
rect 10193 6907 10245 6945
rect 10193 6873 10205 6907
rect 10239 6873 10245 6907
rect 10193 6835 10245 6873
rect 10193 6819 10205 6835
rect 10239 6819 10245 6835
rect 10193 6763 10245 6767
rect 10193 6755 10205 6763
rect 10239 6755 10245 6763
rect 10193 6691 10245 6703
rect 10193 6619 10245 6639
rect 10193 6585 10205 6619
rect 10239 6585 10245 6619
rect 10193 6547 10245 6585
rect 10193 6513 10205 6547
rect 10239 6513 10245 6547
rect 9804 6512 10022 6513
tri 10022 6512 10023 6513 nw
rect 9804 6486 9990 6512
rect 8139 5432 8151 5610
rect 8761 5576 8800 5610
rect 8834 5576 8873 5610
rect 8907 5576 8946 5610
rect 8980 5576 9019 5610
rect 9053 5576 9092 5610
rect 9126 5576 9138 5610
rect 8761 5538 9138 5576
rect 8761 5504 8800 5538
rect 8834 5504 8873 5538
rect 8907 5504 8946 5538
rect 8980 5504 9019 5538
rect 9053 5504 9092 5538
rect 9126 5504 9138 5538
rect 8761 5466 9138 5504
rect 8761 5432 8800 5466
rect 8834 5432 8873 5466
rect 8907 5432 8946 5466
rect 8980 5432 9019 5466
rect 9053 5432 9092 5466
rect 9126 5432 9138 5466
rect 8139 4583 9138 5432
rect 8139 4549 8151 4583
rect 8185 4549 8223 4583
rect 8257 4549 8295 4583
rect 8329 4549 8367 4583
rect 8401 4549 8439 4583
rect 8473 4549 8511 4583
rect 8545 4549 8583 4583
rect 8617 4549 8655 4583
rect 8689 4549 8727 4583
rect 8761 4549 8800 4583
rect 8834 4549 8873 4583
rect 8907 4549 8946 4583
rect 8980 4549 9019 4583
rect 9053 4549 9092 4583
rect 9126 4549 9138 4583
rect 8139 3697 9138 4549
rect 8139 3591 8151 3697
rect 8761 3663 8800 3697
rect 8834 3663 8873 3697
rect 8907 3663 8946 3697
rect 8980 3663 9019 3697
rect 9053 3663 9092 3697
rect 9126 3663 9138 3697
rect 8761 3625 9138 3663
rect 8761 3591 8800 3625
rect 8834 3591 8873 3625
rect 8907 3591 8946 3625
rect 8980 3591 9019 3625
rect 9053 3591 9092 3625
rect 9126 3591 9138 3625
rect 8139 3527 9138 3591
rect 8139 3493 8151 3527
rect 8185 3493 8223 3527
rect 8257 3493 8295 3527
rect 8329 3493 8367 3527
rect 8401 3493 8439 3527
rect 8473 3493 8511 3527
rect 8545 3493 8583 3527
rect 8617 3493 8655 3527
rect 8689 3493 8727 3527
rect 8761 3493 8800 3527
rect 8834 3493 8873 3527
rect 8907 3493 8946 3527
rect 8980 3493 9019 3527
rect 9053 3493 9092 3527
rect 9126 3493 9138 3527
rect 8139 2641 9138 3493
rect 9712 6468 9764 6480
rect 9712 6434 9718 6468
rect 9752 6434 9764 6468
rect 9712 6392 9764 6434
rect 9712 6358 9718 6392
rect 9752 6358 9764 6392
rect 9712 6316 9764 6358
rect 9712 6282 9718 6316
rect 9752 6282 9764 6316
rect 9712 6258 9764 6282
rect 9712 6205 9718 6206
rect 9752 6205 9764 6206
rect 9712 6192 9764 6205
rect 9712 6128 9718 6140
rect 9752 6128 9764 6140
rect 9712 6085 9764 6128
rect 9712 6051 9718 6085
rect 9752 6051 9764 6085
rect 9712 6008 9764 6051
rect 9712 5974 9718 6008
rect 9752 5974 9764 6008
rect 9712 5931 9764 5974
rect 9712 5897 9718 5931
rect 9752 5897 9764 5931
rect 9712 5854 9764 5897
rect 9712 5820 9718 5854
rect 9752 5820 9764 5854
rect 9712 5777 9764 5820
rect 9712 5743 9718 5777
rect 9752 5743 9764 5777
rect 9712 5700 9764 5743
rect 9712 5666 9718 5700
rect 9752 5666 9764 5700
rect 9712 5382 9764 5666
rect 9712 5348 9718 5382
rect 9752 5348 9764 5382
rect 9712 5308 9764 5348
rect 9712 5274 9718 5308
rect 9752 5274 9764 5308
rect 9712 5234 9764 5274
rect 9712 5200 9718 5234
rect 9752 5200 9764 5234
rect 9712 5160 9764 5200
rect 9712 5126 9718 5160
rect 9752 5126 9764 5160
rect 9712 5086 9764 5126
rect 9712 5052 9718 5086
rect 9752 5052 9764 5086
rect 9712 5012 9764 5052
rect 9712 4978 9718 5012
rect 9752 4978 9764 5012
rect 9712 4938 9764 4978
rect 9712 4904 9718 4938
rect 9752 4904 9764 4938
rect 9712 4864 9764 4904
rect 9712 4830 9718 4864
rect 9752 4830 9764 4864
rect 9712 4790 9764 4830
rect 9712 4756 9718 4790
rect 9752 4756 9764 4790
rect 9712 4715 9764 4756
rect 9712 4681 9718 4715
rect 9752 4681 9764 4715
rect 9712 4640 9764 4681
rect 9712 4606 9718 4640
rect 9752 4606 9764 4640
rect 9712 4526 9764 4606
rect 9712 4492 9718 4526
rect 9752 4492 9764 4526
rect 9712 4452 9764 4492
rect 9712 4418 9718 4452
rect 9752 4418 9764 4452
rect 9712 4378 9764 4418
rect 9712 4344 9718 4378
rect 9752 4344 9764 4378
rect 9712 4304 9764 4344
rect 9712 4270 9718 4304
rect 9752 4270 9764 4304
rect 9712 4230 9764 4270
rect 9712 4196 9718 4230
rect 9752 4196 9764 4230
rect 9712 4156 9764 4196
rect 9712 4122 9718 4156
rect 9752 4122 9764 4156
rect 9712 4082 9764 4122
rect 9712 4048 9718 4082
rect 9752 4048 9764 4082
rect 9712 4008 9764 4048
rect 9712 3974 9718 4008
rect 9752 3974 9764 4008
rect 9712 3934 9764 3974
rect 9712 3900 9718 3934
rect 9752 3900 9764 3934
rect 9712 3859 9764 3900
rect 9712 3825 9718 3859
rect 9752 3825 9764 3859
rect 9712 3784 9764 3825
rect 9712 3750 9718 3784
rect 9752 3750 9764 3784
rect 9712 3440 9764 3750
rect 9712 3406 9718 3440
rect 9752 3406 9764 3440
rect 9712 3366 9764 3406
rect 9712 3332 9718 3366
rect 9752 3332 9764 3366
rect 9712 3292 9764 3332
rect 9712 3258 9718 3292
rect 9752 3258 9764 3292
rect 9712 3218 9764 3258
rect 9712 3184 9718 3218
rect 9752 3184 9764 3218
rect 9712 3144 9764 3184
rect 9712 3110 9718 3144
rect 9752 3110 9764 3144
rect 9712 3070 9764 3110
rect 9712 3036 9718 3070
rect 9752 3036 9764 3070
rect 9712 2996 9764 3036
rect 9712 2962 9718 2996
rect 9752 2962 9764 2996
rect 9712 2922 9764 2962
rect 9712 2888 9718 2922
rect 9752 2888 9764 2922
rect 9712 2848 9764 2888
rect 9712 2814 9718 2848
rect 9752 2814 9764 2848
rect 9712 2773 9764 2814
rect 9712 2739 9718 2773
rect 9752 2739 9764 2773
rect 9712 2698 9764 2739
rect 9712 2664 9718 2698
rect 9752 2664 9764 2698
rect 9712 2652 9764 2664
rect 9804 6452 9899 6486
rect 9933 6480 9990 6486
tri 9990 6480 10022 6512 nw
rect 9933 6478 9988 6480
tri 9988 6478 9990 6480 nw
rect 9933 6475 9985 6478
tri 9985 6475 9988 6478 nw
rect 9933 6452 9951 6475
rect 9804 6441 9951 6452
tri 9951 6441 9985 6475 nw
rect 10047 6474 10099 6480
rect 9804 6440 9950 6441
tri 9950 6440 9951 6441 nw
rect 9804 6414 9939 6440
tri 9939 6429 9950 6440 nw
rect 9804 6380 9899 6414
rect 9933 6380 9939 6414
rect 9804 6342 9939 6380
rect 9804 6308 9899 6342
rect 9933 6308 9939 6342
rect 9804 6270 9939 6308
rect 9804 6236 9899 6270
rect 9933 6236 9939 6270
rect 10047 6408 10099 6422
rect 9804 6198 9939 6236
rect 9804 6164 9899 6198
rect 9933 6164 9939 6198
rect 9804 6126 9939 6164
rect 9804 6092 9899 6126
rect 9933 6092 9939 6126
rect 9804 6054 9939 6092
rect 9804 6020 9899 6054
rect 9933 6020 9939 6054
rect 9804 5982 9939 6020
rect 9804 5948 9899 5982
rect 9933 5948 9939 5982
rect 9804 5910 9939 5948
rect 9804 5876 9899 5910
rect 9933 5876 9939 5910
rect 9804 5838 9939 5876
rect 9804 5804 9899 5838
rect 9933 5804 9939 5838
rect 9804 5766 9939 5804
rect 9804 5732 9899 5766
rect 9933 5732 9939 5766
rect 9804 5694 9939 5732
rect 9804 5660 9899 5694
rect 9933 5660 9939 5694
rect 9804 5622 9939 5660
rect 9804 5588 9899 5622
rect 9933 5588 9939 5622
rect 9804 5550 9939 5588
rect 9804 5516 9899 5550
rect 9933 5516 9939 5550
rect 9804 5478 9939 5516
rect 9804 5444 9899 5478
rect 9933 5444 9939 5478
rect 9804 5406 9939 5444
rect 9804 5372 9899 5406
rect 9933 5372 9939 5406
rect 9804 5334 9939 5372
rect 9804 5300 9899 5334
rect 9933 5300 9939 5334
rect 9804 5262 9939 5300
rect 9804 5228 9899 5262
rect 9933 5228 9939 5262
rect 9804 5190 9939 5228
rect 9804 5156 9899 5190
rect 9933 5156 9939 5190
rect 9804 5118 9939 5156
rect 9804 5084 9899 5118
rect 9933 5084 9939 5118
rect 9804 5046 9939 5084
rect 9804 5012 9899 5046
rect 9933 5012 9939 5046
rect 9804 4974 9939 5012
rect 9804 4940 9899 4974
rect 9933 4940 9939 4974
rect 9804 4902 9939 4940
rect 9804 4880 9899 4902
rect 9804 4828 9817 4880
rect 9869 4828 9881 4880
rect 9804 4814 9899 4828
rect 9804 4762 9817 4814
rect 9869 4762 9881 4814
rect 9933 4762 9939 4902
rect 9804 4758 9939 4762
rect 9804 4724 9899 4758
rect 9933 4724 9939 4758
rect 9804 4686 9939 4724
rect 9804 4652 9899 4686
rect 9933 4652 9939 4686
rect 9804 4614 9939 4652
rect 9804 4580 9899 4614
rect 9933 4580 9939 4614
rect 9804 4542 9939 4580
rect 9804 4508 9899 4542
rect 9933 4508 9939 4542
rect 9804 4470 9939 4508
rect 9804 4436 9899 4470
rect 9933 4436 9939 4470
rect 9804 4398 9939 4436
rect 9804 4364 9899 4398
rect 9933 4364 9939 4398
rect 9804 4326 9939 4364
rect 9804 4292 9899 4326
rect 9933 4292 9939 4326
rect 9804 4254 9939 4292
rect 9804 4220 9899 4254
rect 9933 4220 9939 4254
rect 9804 4182 9939 4220
rect 9804 4148 9899 4182
rect 9933 4148 9939 4182
rect 9804 4110 9939 4148
rect 9804 4076 9899 4110
rect 9933 4076 9939 4110
rect 9804 4038 9939 4076
rect 9804 4004 9899 4038
rect 9933 4004 9939 4038
rect 9804 3966 9939 4004
rect 9804 3932 9899 3966
rect 9933 3932 9939 3966
rect 9804 3894 9939 3932
rect 9967 6258 10019 6264
rect 9967 6192 10019 6206
rect 9967 4022 10019 6140
rect 10047 4065 10099 6356
rect 10193 6475 10245 6513
rect 10193 6441 10205 6475
rect 10239 6441 10245 6475
rect 10193 6403 10245 6441
rect 10193 6369 10205 6403
rect 10239 6369 10245 6403
rect 10193 6331 10245 6369
rect 10193 6297 10205 6331
rect 10239 6297 10245 6331
rect 10193 6259 10245 6297
rect 10193 6225 10205 6259
rect 10239 6225 10245 6259
rect 10193 6187 10245 6225
rect 10193 6153 10205 6187
rect 10239 6153 10245 6187
rect 10193 6115 10245 6153
rect 10193 6081 10205 6115
rect 10239 6081 10245 6115
rect 10193 6043 10245 6081
rect 10193 6009 10205 6043
rect 10239 6009 10245 6043
rect 10193 5971 10245 6009
rect 10193 5937 10205 5971
rect 10239 5937 10245 5971
rect 10193 5899 10245 5937
rect 10193 5865 10205 5899
rect 10239 5865 10245 5899
rect 10193 5827 10245 5865
rect 10193 5793 10205 5827
rect 10239 5793 10245 5827
rect 10193 5755 10245 5793
rect 10193 5721 10205 5755
rect 10239 5721 10245 5755
rect 10193 5683 10245 5721
rect 10193 5649 10205 5683
rect 10239 5649 10245 5683
rect 10193 5638 10245 5649
rect 10193 5577 10205 5586
rect 10239 5577 10245 5586
rect 10193 5574 10245 5577
rect 10193 5510 10205 5522
rect 10239 5510 10245 5522
rect 10193 5433 10205 5458
rect 10239 5433 10245 5458
rect 10193 5395 10245 5433
rect 10193 5361 10205 5395
rect 10239 5361 10245 5395
rect 10193 5323 10245 5361
rect 10193 5289 10205 5323
rect 10239 5289 10245 5323
rect 10193 5251 10245 5289
rect 10193 5217 10205 5251
rect 10239 5217 10245 5251
rect 10193 5179 10245 5217
rect 10193 5145 10205 5179
rect 10239 5145 10245 5179
rect 10193 5107 10245 5145
rect 10193 5073 10205 5107
rect 10239 5073 10245 5107
rect 10193 5035 10245 5073
rect 10193 5001 10205 5035
rect 10239 5001 10245 5035
rect 10193 4963 10245 5001
rect 10193 4929 10205 4963
rect 10239 4929 10245 4963
rect 10193 4891 10245 4929
rect 10193 4857 10205 4891
rect 10239 4857 10245 4891
rect 10193 4819 10245 4857
rect 10193 4785 10205 4819
rect 10239 4785 10245 4819
rect 10193 4747 10245 4785
rect 10193 4713 10205 4747
rect 10239 4713 10245 4747
rect 10193 4675 10245 4713
rect 10193 4641 10205 4675
rect 10239 4641 10245 4675
rect 10193 4603 10245 4641
rect 10193 4569 10205 4603
rect 10239 4569 10245 4603
rect 10193 4531 10245 4569
rect 10193 4497 10205 4531
rect 10239 4497 10245 4531
rect 10193 4459 10245 4497
rect 10193 4425 10205 4459
rect 10239 4425 10245 4459
rect 10193 4387 10245 4425
rect 10193 4353 10205 4387
rect 10239 4353 10245 4387
rect 10193 4315 10245 4353
rect 10193 4281 10205 4315
rect 10239 4281 10245 4315
rect 10193 4243 10245 4281
rect 10193 4209 10205 4243
rect 10239 4209 10245 4243
rect 10193 4171 10245 4209
rect 10193 4137 10205 4171
rect 10239 4137 10245 4171
rect 10193 4099 10245 4137
tri 10099 4065 10111 4077 sw
rect 10193 4065 10205 4099
rect 10239 4065 10245 4099
rect 10047 4064 10111 4065
tri 10111 4064 10112 4065 sw
rect 10047 4052 10112 4064
tri 10112 4052 10124 4064 sw
rect 10047 4046 10163 4052
rect 10099 3994 10111 4046
rect 10047 3988 10163 3994
rect 10193 4027 10245 4065
rect 10193 3993 10205 4027
rect 10239 3993 10245 4027
rect 9967 3956 10019 3970
rect 9967 3898 10019 3904
rect 10193 3955 10245 3993
rect 10193 3921 10205 3955
rect 10239 3921 10245 3955
rect 9804 3860 9899 3894
rect 9933 3860 9939 3894
rect 10193 3883 10245 3921
rect 9804 3849 9939 3860
tri 9939 3849 9959 3869 sw
rect 10193 3849 10205 3883
rect 10239 3849 10245 3883
rect 9804 3848 9959 3849
tri 9959 3848 9960 3849 sw
rect 9804 3822 9960 3848
rect 9804 3788 9899 3822
rect 9933 3814 9960 3822
tri 9960 3814 9994 3848 sw
rect 9933 3811 9994 3814
tri 9994 3811 9997 3814 sw
rect 10193 3811 10245 3849
rect 9933 3788 9997 3811
rect 9804 3777 9997 3788
tri 9997 3777 10031 3811 sw
rect 10193 3777 10205 3811
rect 10239 3777 10245 3811
rect 9804 3776 10031 3777
tri 10031 3776 10032 3777 sw
rect 9804 3758 10032 3776
tri 10032 3758 10050 3776 sw
rect 9804 3750 10050 3758
rect 9804 3716 9899 3750
rect 9933 3716 10050 3750
rect 9804 3678 10050 3716
rect 9804 3644 9899 3678
rect 9933 3644 10050 3678
rect 9804 3606 10050 3644
rect 9804 3572 9899 3606
rect 9933 3572 10050 3606
rect 9804 3534 10050 3572
rect 9804 3500 9899 3534
rect 9933 3500 10050 3534
rect 9804 3462 10050 3500
rect 9804 3428 9899 3462
rect 9933 3428 10050 3462
rect 9804 3390 10050 3428
rect 9804 3356 9899 3390
rect 9933 3356 10050 3390
rect 9804 3318 10050 3356
rect 9804 3284 9899 3318
rect 9933 3284 10050 3318
rect 9804 3246 10050 3284
rect 9804 3212 9899 3246
rect 9933 3212 10050 3246
rect 9804 3174 10050 3212
rect 9804 3140 9899 3174
rect 9933 3140 10050 3174
rect 9804 3102 10050 3140
rect 9804 3068 9899 3102
rect 9933 3068 10050 3102
rect 9804 3030 10050 3068
rect 9804 2996 9899 3030
rect 9933 2996 10050 3030
rect 9804 2958 10050 2996
rect 9804 2924 9899 2958
rect 9933 2924 10050 2958
rect 9804 2886 10050 2924
rect 9804 2852 9899 2886
rect 9933 2852 10050 2886
rect 9804 2814 10050 2852
rect 9804 2780 9899 2814
rect 9933 2780 10050 2814
rect 9804 2742 10050 2780
rect 9804 2708 9899 2742
rect 9933 2708 10050 2742
rect 9804 2670 10050 2708
rect 8139 2463 8151 2641
rect 8761 2607 8800 2641
rect 8834 2607 8873 2641
rect 8907 2607 8946 2641
rect 8980 2607 9019 2641
rect 9053 2607 9092 2641
rect 9126 2607 9138 2641
rect 8761 2569 9138 2607
rect 8761 2535 8800 2569
rect 8834 2535 8873 2569
rect 8907 2535 8946 2569
rect 8980 2535 9019 2569
rect 9053 2535 9092 2569
rect 9126 2535 9138 2569
rect 8761 2497 9138 2535
rect 8761 2463 8800 2497
rect 8834 2463 8873 2497
rect 8907 2463 8946 2497
rect 8980 2463 9019 2497
rect 9053 2463 9092 2497
rect 9126 2463 9138 2497
rect 8139 2447 9138 2463
rect 9804 2636 9899 2670
rect 9933 2636 10050 2670
rect 9804 2598 10050 2636
rect 9804 2564 9899 2598
rect 9933 2564 10050 2598
rect 9804 2526 10050 2564
rect 9804 2492 9899 2526
rect 9933 2492 10050 2526
rect 9804 2454 10050 2492
tri 8945 2422 8970 2447 ne
rect 8139 1588 8845 1838
rect 8139 1536 8151 1588
rect 8203 1536 8217 1588
rect 8269 1536 8283 1588
rect 8335 1536 8349 1588
rect 8401 1536 8415 1588
rect 8467 1536 8481 1588
rect 8533 1536 8546 1588
rect 8598 1536 8611 1588
rect 8663 1536 8676 1588
rect 8728 1536 8741 1588
rect 8793 1536 8845 1588
rect 8139 1524 8845 1536
rect 8139 1472 8151 1524
rect 8203 1472 8217 1524
rect 8269 1472 8283 1524
rect 8335 1472 8349 1524
rect 8401 1472 8415 1524
rect 8467 1472 8481 1524
rect 8533 1472 8546 1524
rect 8598 1472 8611 1524
rect 8663 1472 8676 1524
rect 8728 1472 8741 1524
rect 8793 1472 8845 1524
rect 8139 1460 8845 1472
rect 8139 1408 8151 1460
rect 8203 1408 8217 1460
rect 8269 1408 8283 1460
rect 8335 1408 8349 1460
rect 8401 1408 8415 1460
rect 8467 1408 8481 1460
rect 8533 1408 8546 1460
rect 8598 1408 8611 1460
rect 8663 1408 8676 1460
rect 8728 1408 8741 1460
rect 8793 1408 8845 1460
rect 8139 1396 8845 1408
rect 8139 1344 8151 1396
rect 8203 1344 8217 1396
rect 8269 1344 8283 1396
rect 8335 1344 8349 1396
rect 8401 1344 8415 1396
rect 8467 1344 8481 1396
rect 8533 1344 8546 1396
rect 8598 1344 8611 1396
rect 8663 1344 8676 1396
rect 8728 1344 8741 1396
rect 8793 1344 8845 1396
rect 8139 1332 8845 1344
rect 8139 1280 8151 1332
rect 8203 1280 8217 1332
rect 8269 1280 8283 1332
rect 8335 1280 8349 1332
rect 8401 1280 8415 1332
rect 8467 1280 8481 1332
rect 8533 1280 8546 1332
rect 8598 1280 8611 1332
rect 8663 1280 8676 1332
rect 8728 1280 8741 1332
rect 8793 1280 8845 1332
tri 8118 1195 8139 1216 se
rect 8139 1195 8845 1280
tri 8114 1191 8118 1195 se
rect 8118 1191 8845 1195
rect 8023 1185 8075 1191
rect 8077 1190 8113 1191
rect 8023 1121 8075 1133
rect 8023 1063 8075 1069
rect 8076 1064 8114 1190
rect 8077 1063 8113 1064
rect 8115 1063 8845 1191
tri 8114 1046 8131 1063 ne
rect 8131 1046 8845 1063
tri 8131 1041 8136 1046 ne
rect 8136 1041 8845 1046
tri 8136 1038 8139 1041 ne
rect 8139 899 8845 1041
tri 8244 896 8247 899 ne
rect 8247 896 8355 899
tri 8355 896 8358 899 nw
tri 8756 896 8759 899 ne
rect 8759 896 8845 899
tri 8247 874 8269 896 ne
rect 7575 748 7633 754
tri 7675 750 7684 759 se
rect 7684 750 7692 768
tri 7673 748 7675 750 se
rect 7675 748 7692 750
tri 7655 730 7673 748 se
rect 7673 730 7692 748
tri 7645 720 7655 730 se
rect 7655 720 7692 730
tri 6773 510 6776 513 se
rect 6776 510 6980 513
tri 6763 500 6773 510 se
rect 6773 500 6980 510
rect 5180 480 5255 482
tri 5255 480 5257 482 sw
rect 3761 436 3891 448
rect 5180 428 5186 480
rect 5238 428 5250 480
rect 5302 428 5308 480
rect 5522 448 5563 482
rect 5597 448 5638 482
tri 5808 480 5810 482 se
rect 5810 480 5885 482
rect 5522 436 5638 448
rect 5757 428 5763 480
rect 5815 428 5827 480
rect 5879 428 5885 480
rect 6788 442 6980 500
rect 7026 692 7078 704
rect 7026 658 7032 692
rect 7066 658 7078 692
rect 7026 620 7078 658
rect 7026 586 7032 620
rect 7066 586 7078 620
rect 7026 550 7078 586
rect 7026 486 7078 498
rect 7259 676 7271 710
rect 7305 676 7343 710
rect 7377 676 7389 710
rect 7259 634 7389 676
rect 7259 600 7271 634
rect 7305 600 7343 634
rect 7377 600 7389 634
rect 7259 558 7389 600
rect 7612 708 7692 720
rect 7612 674 7618 708
rect 7652 674 7692 708
rect 7612 652 7692 674
rect 7808 652 7814 768
rect 8013 716 8019 768
rect 8071 716 8077 768
rect 8013 704 8030 716
rect 8064 704 8077 716
rect 8013 652 8019 704
rect 8071 652 8077 704
rect 7612 636 7698 652
rect 7612 602 7618 636
rect 7652 624 7698 636
tri 7698 624 7726 652 nw
rect 8013 624 8030 652
rect 8064 624 8077 652
rect 7652 602 7676 624
tri 7676 602 7698 624 nw
rect 7612 590 7664 602
tri 7664 590 7676 602 nw
rect 7259 524 7271 558
rect 7305 524 7343 558
rect 7377 524 7389 558
rect 7762 585 7892 591
rect 7814 533 7826 585
rect 7878 578 7892 585
rect 7880 544 7892 578
rect 8013 586 8077 624
rect 8013 552 8030 586
rect 8064 552 8077 586
rect 8013 546 8077 552
rect 8269 708 8333 896
tri 8333 874 8355 896 nw
tri 8759 874 8781 896 ne
rect 8269 674 8286 708
rect 8320 674 8333 708
rect 8269 636 8333 674
rect 8269 624 8286 636
rect 8320 624 8333 636
rect 8269 572 8275 624
rect 8327 572 8333 624
rect 8269 564 8333 572
rect 8269 560 8286 564
rect 8320 560 8333 564
rect 7878 533 7892 544
rect 7762 527 7892 533
rect 7259 482 7389 524
rect 8269 508 8275 560
rect 8327 508 8333 560
rect 8525 716 8531 768
rect 8583 716 8589 768
rect 8525 704 8542 716
rect 8576 704 8589 716
rect 8525 652 8531 704
rect 8583 652 8589 704
rect 8525 624 8542 652
rect 8576 624 8589 652
rect 8525 586 8589 624
rect 8525 552 8542 586
rect 8576 552 8589 586
rect 8525 546 8589 552
rect 8781 708 8845 896
rect 8781 674 8798 708
rect 8832 674 8845 708
rect 8970 1195 9100 2447
tri 9100 2422 9125 2447 nw
rect 9804 2420 9899 2454
rect 9933 2420 10050 2454
rect 9804 2382 10050 2420
rect 9804 2348 9899 2382
rect 9933 2348 10050 2382
rect 9804 2310 10050 2348
rect 9804 2276 9899 2310
rect 9933 2276 10050 2310
rect 9804 2238 10050 2276
rect 9804 2204 9899 2238
rect 9933 2204 10050 2238
rect 9804 2166 10050 2204
rect 9804 2132 9899 2166
rect 9933 2132 10050 2166
rect 9804 2094 10050 2132
rect 9804 2060 9899 2094
rect 9933 2060 10050 2094
rect 9804 2022 10050 2060
rect 9804 1988 9899 2022
rect 9933 1988 10050 2022
rect 9804 1950 10050 1988
rect 9804 1916 9899 1950
rect 9933 1916 10050 1950
rect 9804 1878 10050 1916
rect 9804 1844 9899 1878
rect 9933 1844 10050 1878
rect 9804 1806 10050 1844
rect 9804 1772 9899 1806
rect 9933 1772 10050 1806
rect 9712 1747 9764 1759
rect 9712 1713 9718 1747
rect 9752 1713 9764 1747
rect 9712 1673 9764 1713
rect 9712 1639 9718 1673
rect 9752 1639 9764 1673
rect 9712 1599 9764 1639
rect 9712 1565 9718 1599
rect 9752 1565 9764 1599
rect 9712 1525 9764 1565
rect 9712 1491 9718 1525
rect 9752 1491 9764 1525
rect 9712 1451 9764 1491
rect 9712 1417 9718 1451
rect 9752 1417 9764 1451
rect 9712 1377 9764 1417
rect 9712 1343 9718 1377
rect 9752 1343 9764 1377
rect 9712 1303 9764 1343
rect 9712 1269 9718 1303
rect 9752 1269 9764 1303
rect 9712 1229 9764 1269
tri 9100 1195 9121 1216 sw
rect 9712 1195 9718 1229
rect 9752 1195 9764 1229
rect 8970 1191 9121 1195
tri 9121 1191 9125 1195 sw
rect 8970 1063 9123 1191
rect 9124 1064 9125 1190
rect 9161 1064 9162 1190
rect 9163 1185 9215 1191
rect 9163 1121 9215 1133
rect 9163 1063 9215 1069
rect 9712 1185 9764 1195
rect 9712 1121 9718 1133
rect 9752 1121 9764 1133
rect 8970 1046 9108 1063
tri 9108 1046 9125 1063 nw
rect 9712 1046 9718 1069
rect 9752 1046 9764 1069
rect 8970 1041 9103 1046
tri 9103 1041 9108 1046 nw
rect 8970 800 9100 1041
tri 9100 1038 9103 1041 nw
rect 9712 1005 9764 1046
rect 9712 971 9718 1005
rect 9752 971 9764 1005
rect 9712 959 9764 971
rect 9804 1734 10050 1772
rect 9804 1700 9899 1734
rect 9933 1700 10050 1734
rect 9804 1662 10050 1700
rect 9804 1628 9899 1662
rect 9933 1628 10050 1662
rect 9804 1590 10050 1628
rect 9804 1556 9899 1590
rect 9933 1556 10050 1590
rect 9804 1518 10050 1556
rect 9804 1484 9899 1518
rect 9933 1484 10050 1518
rect 9804 1446 10050 1484
rect 9804 1412 9899 1446
rect 9933 1412 10050 1446
rect 9804 1374 10050 1412
rect 9804 1340 9899 1374
rect 9933 1340 10050 1374
rect 9804 1302 10050 1340
rect 9804 1268 9899 1302
rect 9933 1268 10050 1302
rect 9804 1230 10050 1268
rect 9804 1196 9899 1230
rect 9933 1196 10050 1230
rect 9804 1158 10050 1196
rect 9804 1124 9899 1158
rect 9933 1124 10050 1158
rect 9804 1086 10050 1124
rect 9804 1052 9899 1086
rect 9933 1052 10050 1086
rect 9804 1014 10050 1052
rect 9804 980 9899 1014
rect 9933 980 10050 1014
rect 8970 766 9054 800
rect 9088 766 9100 800
rect 8970 728 9100 766
rect 8970 694 9054 728
rect 9088 694 9100 728
rect 9804 942 10050 980
rect 9804 908 9899 942
rect 9933 908 10050 942
rect 9804 870 10050 908
rect 9804 836 9899 870
rect 9933 836 10050 870
rect 9804 798 10050 836
rect 9804 764 9899 798
rect 9933 764 10050 798
rect 9804 726 10050 764
rect 8970 682 9100 694
tri 8970 674 8978 682 ne
rect 8978 674 9100 682
rect 8781 636 8845 674
tri 8978 656 8996 674 ne
rect 8996 656 9100 674
rect 8781 624 8798 636
rect 8832 624 8845 636
rect 8781 572 8787 624
rect 8839 572 8845 624
tri 8996 622 9030 656 ne
rect 9030 622 9054 656
rect 9088 622 9100 656
tri 9030 606 9046 622 ne
rect 9046 606 9100 622
rect 9193 708 9257 714
rect 9193 674 9210 708
rect 9244 674 9257 708
rect 9193 636 9257 674
rect 9193 624 9210 636
rect 9244 624 9257 636
rect 8781 564 8845 572
rect 8781 560 8798 564
rect 8832 560 8845 564
rect 8781 508 8787 560
rect 8839 508 8845 560
rect 9193 572 9199 624
rect 9251 572 9257 624
rect 9193 564 9257 572
rect 9193 560 9210 564
rect 9244 560 9257 564
rect 9193 508 9199 560
rect 9251 508 9257 560
rect 9804 692 9899 726
rect 9933 692 10050 726
rect 9804 654 10050 692
rect 9804 620 9899 654
rect 9933 620 10050 654
rect 9804 582 10050 620
rect 9804 548 9899 582
rect 9933 548 10050 582
rect 9804 510 10050 548
rect 7259 448 7271 482
rect 7305 448 7343 482
rect 7377 448 7389 482
rect 7259 436 7389 448
rect 9804 476 9899 510
rect 9933 476 10050 510
rect 9804 438 10050 476
rect 7026 428 7078 434
rect 1117 379 1185 413
rect 1219 379 1225 413
rect 1117 341 1225 379
rect 1117 307 1185 341
rect 1219 307 1225 341
rect 9804 404 9899 438
rect 9933 404 10050 438
rect 9804 366 10050 404
rect 9804 332 9899 366
rect 9933 332 10050 366
rect 1117 269 1225 307
tri 9791 294 9804 307 se
rect 9804 294 10050 332
rect 10193 3739 10245 3777
rect 10193 3705 10205 3739
rect 10239 3705 10245 3739
rect 10193 3667 10245 3705
rect 10193 3633 10205 3667
rect 10239 3633 10245 3667
rect 10193 3595 10245 3633
rect 10193 3561 10205 3595
rect 10239 3561 10245 3595
rect 10193 3523 10245 3561
rect 10193 3489 10205 3523
rect 10239 3489 10245 3523
rect 10193 3451 10245 3489
rect 10193 3417 10205 3451
rect 10239 3417 10245 3451
rect 10193 3379 10245 3417
rect 10193 3345 10205 3379
rect 10239 3345 10245 3379
rect 10193 3307 10245 3345
rect 10193 3273 10205 3307
rect 10239 3273 10245 3307
rect 10193 3235 10245 3273
rect 10193 3201 10205 3235
rect 10239 3201 10245 3235
rect 10193 3163 10245 3201
rect 10193 3129 10205 3163
rect 10239 3129 10245 3163
rect 10193 3091 10245 3129
rect 10193 3057 10205 3091
rect 10239 3057 10245 3091
rect 10193 3019 10245 3057
rect 10193 2985 10205 3019
rect 10239 2985 10245 3019
rect 10193 2947 10245 2985
rect 10193 2913 10205 2947
rect 10239 2913 10245 2947
rect 10193 2875 10245 2913
rect 10193 2841 10205 2875
rect 10239 2841 10245 2875
rect 10193 2803 10245 2841
rect 10193 2769 10205 2803
rect 10239 2769 10245 2803
rect 10193 2731 10245 2769
rect 10193 2697 10205 2731
rect 10239 2697 10245 2731
rect 10193 2659 10245 2697
rect 10193 2625 10205 2659
rect 10239 2625 10245 2659
rect 10193 2587 10245 2625
rect 10193 2553 10205 2587
rect 10239 2553 10245 2587
rect 10193 2515 10245 2553
rect 10193 2481 10205 2515
rect 10239 2481 10245 2515
rect 10193 2443 10245 2481
rect 10193 2409 10205 2443
rect 10239 2409 10245 2443
rect 10193 2371 10245 2409
rect 10193 2337 10205 2371
rect 10239 2337 10245 2371
rect 10193 2299 10245 2337
rect 10193 2265 10205 2299
rect 10239 2265 10245 2299
rect 10193 2227 10245 2265
rect 10193 2193 10205 2227
rect 10239 2193 10245 2227
rect 10193 2155 10245 2193
rect 10193 2121 10205 2155
rect 10239 2121 10245 2155
rect 10193 2083 10245 2121
rect 10193 2060 10205 2083
rect 10239 2060 10245 2083
rect 10193 1996 10205 2008
rect 10239 1996 10245 2008
rect 10193 1939 10245 1944
rect 10193 1932 10205 1939
rect 10239 1932 10245 1939
rect 10193 1868 10245 1880
rect 10193 1804 10245 1816
rect 10193 1723 10245 1752
rect 10193 1689 10205 1723
rect 10239 1689 10245 1723
rect 10193 1651 10245 1689
rect 10193 1617 10205 1651
rect 10239 1617 10245 1651
rect 10193 1579 10245 1617
rect 10193 1545 10205 1579
rect 10239 1545 10245 1579
rect 10193 1507 10245 1545
rect 10193 1473 10205 1507
rect 10239 1473 10245 1507
rect 10193 1435 10245 1473
rect 10193 1401 10205 1435
rect 10239 1401 10245 1435
rect 10193 1363 10245 1401
rect 10193 1329 10205 1363
rect 10239 1329 10245 1363
rect 10193 1291 10245 1329
rect 10193 1257 10205 1291
rect 10239 1257 10245 1291
rect 10193 1219 10245 1257
rect 10193 1185 10205 1219
rect 10239 1185 10245 1219
rect 10193 1147 10245 1185
rect 10193 1113 10205 1147
rect 10239 1113 10245 1147
rect 10193 1075 10245 1113
rect 10193 1041 10205 1075
rect 10239 1041 10245 1075
rect 10193 1003 10245 1041
rect 10193 969 10205 1003
rect 10239 969 10245 1003
rect 10193 930 10245 969
rect 10193 896 10205 930
rect 10239 896 10245 930
rect 10193 857 10245 896
rect 10193 823 10205 857
rect 10239 823 10245 857
rect 10193 784 10245 823
rect 10193 750 10205 784
rect 10239 750 10245 784
rect 10193 711 10245 750
rect 10193 677 10205 711
rect 10239 677 10245 711
rect 10193 638 10245 677
rect 10193 604 10205 638
rect 10239 604 10245 638
rect 10193 565 10245 604
rect 10193 531 10205 565
rect 10239 531 10245 565
rect 10193 506 10245 531
rect 12876 7589 12951 7597
tri 12951 7589 12959 7597 sw
rect 12876 7016 12959 7589
rect 13015 7172 13067 7798
tri 13067 7172 13109 7214 sw
rect 13015 7160 13109 7172
rect 13015 7126 13069 7160
rect 13103 7126 13109 7160
rect 13015 7088 13109 7126
rect 13015 7054 13069 7088
rect 13103 7054 13109 7088
rect 13015 7045 13109 7054
tri 13015 7027 13033 7045 ne
rect 13033 7027 13109 7045
tri 12959 7016 12970 7027 sw
tri 13033 7016 13044 7027 ne
rect 13044 7016 13109 7027
rect 12876 6982 12970 7016
tri 12970 6982 13004 7016 sw
tri 13044 6997 13063 7016 ne
rect 13063 6982 13069 7016
rect 13103 6982 13109 7016
rect 12876 6979 13004 6982
tri 13004 6979 13007 6982 sw
rect 12876 6819 13007 6979
rect 12876 6639 12891 6819
rect 12876 5638 13007 6639
rect 12876 5586 12891 5638
rect 12943 5586 12955 5638
rect 12876 5564 13007 5586
rect 12876 5512 12891 5564
rect 12943 5512 12955 5564
rect 12876 5490 13007 5512
rect 12876 5438 12891 5490
rect 12943 5438 12955 5490
rect 12876 5416 13007 5438
rect 12876 5364 12891 5416
rect 12943 5364 12955 5416
rect 12876 5341 13007 5364
rect 12876 5289 12891 5341
rect 12943 5289 12955 5341
rect 12876 5266 13007 5289
rect 12876 5214 12891 5266
rect 12943 5214 12955 5266
rect 12876 5191 13007 5214
rect 12876 5139 12891 5191
rect 12943 5139 12955 5191
rect 12876 2066 13007 5139
rect 12876 2014 12891 2066
rect 12943 2014 12955 2066
rect 12876 2001 13007 2014
rect 12876 1949 12891 2001
rect 12943 1949 12955 2001
rect 12876 1936 13007 1949
rect 12876 1884 12891 1936
rect 12943 1884 12955 1936
rect 12876 1870 13007 1884
rect 12876 1818 12891 1870
rect 12943 1818 12955 1870
rect 12876 1804 13007 1818
rect 12876 1752 12891 1804
rect 12943 1752 12955 1804
tri 10245 506 10250 511 sw
tri 12871 506 12876 511 se
rect 12876 506 13007 1752
rect 10193 492 10250 506
rect 10193 458 10205 492
rect 10239 486 10250 492
tri 10250 486 10270 506 sw
tri 12851 486 12871 506 se
rect 12871 486 13007 506
rect 10239 480 13007 486
rect 10239 458 10277 480
rect 10193 446 10277 458
rect 10311 446 10350 480
rect 10384 446 10423 480
rect 10457 446 10496 480
rect 10530 446 10569 480
rect 10603 446 10642 480
rect 10676 446 10715 480
rect 10749 446 10788 480
rect 10822 446 10861 480
rect 10895 446 10934 480
rect 10968 446 11007 480
rect 11041 446 11080 480
rect 11114 446 11153 480
rect 11187 446 11226 480
rect 11260 446 11299 480
rect 11333 446 11372 480
rect 11406 446 11445 480
rect 11479 446 11518 480
rect 11552 446 11591 480
rect 11625 446 11664 480
rect 11698 446 11737 480
rect 11771 446 11810 480
rect 11844 446 11883 480
rect 11917 446 11956 480
rect 11990 446 12029 480
rect 12063 446 12102 480
rect 12136 446 12175 480
rect 12209 446 12248 480
rect 12282 446 12321 480
rect 12355 446 12393 480
rect 12427 446 12465 480
rect 12499 446 12537 480
rect 12571 446 12609 480
rect 12643 446 12681 480
rect 12715 446 12753 480
rect 12787 446 13007 480
rect 10193 409 13007 446
rect 10193 399 12997 409
tri 12997 399 13007 409 nw
rect 13063 6944 13109 6982
rect 13063 6910 13069 6944
rect 13103 6910 13109 6944
rect 13063 6872 13109 6910
rect 13063 6838 13069 6872
rect 13103 6838 13109 6872
rect 13063 6800 13109 6838
rect 13063 6766 13069 6800
rect 13103 6766 13109 6800
rect 13063 6728 13109 6766
rect 13063 6694 13069 6728
rect 13103 6694 13109 6728
rect 13063 6656 13109 6694
rect 13063 6622 13069 6656
rect 13103 6622 13109 6656
rect 13063 6584 13109 6622
rect 13063 6550 13069 6584
rect 13103 6550 13109 6584
rect 13063 6512 13109 6550
rect 13063 6478 13069 6512
rect 13103 6478 13109 6512
rect 13063 6440 13109 6478
rect 13063 6406 13069 6440
rect 13103 6406 13109 6440
rect 13063 6368 13109 6406
rect 13063 6334 13069 6368
rect 13103 6334 13109 6368
rect 13063 6296 13109 6334
rect 13063 6262 13069 6296
rect 13103 6262 13109 6296
rect 13063 6224 13109 6262
rect 13063 6190 13069 6224
rect 13103 6190 13109 6224
rect 13063 6152 13109 6190
rect 13063 6118 13069 6152
rect 13103 6118 13109 6152
rect 13063 6080 13109 6118
rect 13063 6046 13069 6080
rect 13103 6046 13109 6080
rect 13063 6008 13109 6046
rect 13063 5974 13069 6008
rect 13103 5974 13109 6008
rect 13063 5936 13109 5974
rect 13063 5902 13069 5936
rect 13103 5902 13109 5936
rect 13063 5864 13109 5902
rect 13063 5830 13069 5864
rect 13103 5830 13109 5864
rect 13063 5792 13109 5830
rect 13063 5758 13069 5792
rect 13103 5758 13109 5792
rect 13063 5720 13109 5758
rect 13063 5686 13069 5720
rect 13103 5686 13109 5720
rect 13063 5648 13109 5686
rect 13063 5614 13069 5648
rect 13103 5614 13109 5648
rect 13063 5576 13109 5614
rect 13063 5542 13069 5576
rect 13103 5542 13109 5576
rect 13063 5504 13109 5542
rect 13063 5470 13069 5504
rect 13103 5470 13109 5504
rect 13063 5432 13109 5470
rect 13063 5398 13069 5432
rect 13103 5398 13109 5432
rect 13063 5360 13109 5398
rect 13063 5326 13069 5360
rect 13103 5326 13109 5360
rect 13063 5288 13109 5326
rect 13063 5254 13069 5288
rect 13103 5254 13109 5288
rect 13063 5216 13109 5254
rect 13063 5182 13069 5216
rect 13103 5182 13109 5216
rect 13063 5144 13109 5182
rect 13063 5110 13069 5144
rect 13103 5110 13109 5144
rect 13063 5072 13109 5110
rect 13063 5038 13069 5072
rect 13103 5038 13109 5072
rect 13063 5000 13109 5038
rect 13063 4966 13069 5000
rect 13103 4966 13109 5000
rect 13063 4928 13109 4966
rect 13063 4894 13069 4928
rect 13103 4894 13109 4928
rect 13063 4886 13109 4894
tri 13109 4886 13115 4892 sw
rect 13063 4880 13115 4886
rect 13063 4822 13069 4828
rect 13103 4822 13115 4828
rect 13063 4814 13115 4822
rect 13063 4750 13069 4762
rect 13103 4756 13115 4762
rect 13103 4750 13109 4756
tri 13109 4750 13115 4756 nw
rect 13063 4712 13109 4750
rect 13063 4678 13069 4712
rect 13103 4678 13109 4712
rect 13063 4640 13109 4678
rect 13063 4606 13069 4640
rect 13103 4606 13109 4640
rect 13063 4568 13109 4606
rect 13063 4534 13069 4568
rect 13103 4534 13109 4568
rect 13063 4496 13109 4534
rect 13063 4462 13069 4496
rect 13103 4462 13109 4496
rect 13063 4424 13109 4462
rect 13063 4390 13069 4424
rect 13103 4390 13109 4424
rect 13063 4352 13109 4390
rect 13063 4318 13069 4352
rect 13103 4318 13109 4352
rect 13063 4280 13109 4318
rect 13063 4246 13069 4280
rect 13103 4246 13109 4280
rect 13063 4208 13109 4246
rect 13063 4174 13069 4208
rect 13103 4174 13109 4208
rect 13063 4136 13109 4174
rect 13063 4102 13069 4136
rect 13103 4102 13109 4136
rect 13063 4064 13109 4102
rect 13063 4030 13069 4064
rect 13103 4030 13109 4064
rect 13063 3992 13109 4030
rect 13063 3958 13069 3992
rect 13103 3958 13109 3992
rect 13063 3920 13109 3958
rect 13063 3886 13069 3920
rect 13103 3886 13109 3920
rect 13063 3848 13109 3886
rect 13063 3814 13069 3848
rect 13103 3814 13109 3848
rect 13063 3776 13109 3814
rect 13063 3742 13069 3776
rect 13103 3742 13109 3776
rect 13063 3704 13109 3742
rect 13063 3670 13069 3704
rect 13103 3670 13109 3704
rect 13063 3632 13109 3670
rect 13063 3598 13069 3632
rect 13103 3598 13109 3632
rect 13063 3560 13109 3598
rect 13063 3526 13069 3560
rect 13103 3526 13109 3560
rect 13063 3488 13109 3526
rect 13063 3454 13069 3488
rect 13103 3454 13109 3488
rect 13063 3416 13109 3454
rect 13063 3382 13069 3416
rect 13103 3382 13109 3416
rect 13063 3344 13109 3382
rect 13063 3310 13069 3344
rect 13103 3310 13109 3344
rect 13063 3272 13109 3310
rect 13063 3238 13069 3272
rect 13103 3238 13109 3272
rect 13063 3200 13109 3238
rect 13063 3166 13069 3200
rect 13103 3166 13109 3200
rect 13063 3128 13109 3166
rect 13063 3094 13069 3128
rect 13103 3094 13109 3128
rect 13063 3056 13109 3094
rect 13063 3022 13069 3056
rect 13103 3022 13109 3056
rect 13063 2984 13109 3022
rect 13063 2950 13069 2984
rect 13103 2950 13109 2984
rect 13063 2912 13109 2950
rect 13063 2878 13069 2912
rect 13103 2878 13109 2912
rect 13063 2840 13109 2878
rect 13063 2806 13069 2840
rect 13103 2806 13109 2840
rect 13063 2768 13109 2806
rect 13063 2734 13069 2768
rect 13103 2734 13109 2768
rect 13063 2696 13109 2734
rect 13063 2662 13069 2696
rect 13103 2662 13109 2696
rect 13063 2623 13109 2662
rect 13063 2589 13069 2623
rect 13103 2589 13109 2623
rect 13063 2550 13109 2589
rect 13063 2516 13069 2550
rect 13103 2516 13109 2550
rect 13063 2477 13109 2516
rect 13063 2443 13069 2477
rect 13103 2443 13109 2477
rect 13063 2404 13109 2443
rect 13063 2370 13069 2404
rect 13103 2370 13109 2404
rect 13063 2331 13109 2370
rect 13063 2297 13069 2331
rect 13103 2297 13109 2331
rect 13063 2258 13109 2297
rect 13063 2224 13069 2258
rect 13103 2224 13109 2258
rect 13063 2185 13109 2224
rect 13063 2151 13069 2185
rect 13103 2151 13109 2185
rect 13063 2112 13109 2151
rect 13063 2078 13069 2112
rect 13103 2078 13109 2112
rect 13063 2039 13109 2078
rect 13063 2005 13069 2039
rect 13103 2005 13109 2039
rect 13063 1966 13109 2005
rect 13063 1932 13069 1966
rect 13103 1932 13109 1966
rect 13063 1893 13109 1932
rect 13063 1859 13069 1893
rect 13103 1859 13109 1893
rect 13063 1820 13109 1859
rect 13063 1786 13069 1820
rect 13103 1786 13109 1820
rect 13063 1747 13109 1786
rect 13063 1713 13069 1747
rect 13103 1713 13109 1747
rect 13063 1674 13109 1713
rect 13063 1640 13069 1674
rect 13103 1640 13109 1674
rect 13063 1601 13109 1640
rect 13063 1567 13069 1601
rect 13103 1567 13109 1601
rect 13063 1528 13109 1567
rect 13063 1494 13069 1528
rect 13103 1494 13109 1528
rect 13063 1455 13109 1494
rect 13063 1421 13069 1455
rect 13103 1421 13109 1455
rect 13063 1382 13109 1421
rect 13063 1348 13069 1382
rect 13103 1348 13109 1382
rect 13063 1309 13109 1348
rect 13063 1275 13069 1309
rect 13103 1275 13109 1309
rect 13063 1236 13109 1275
rect 13063 1202 13069 1236
rect 13103 1202 13109 1236
rect 13063 1163 13109 1202
rect 13063 1129 13069 1163
rect 13103 1129 13109 1163
rect 13063 1090 13109 1129
rect 13063 1056 13069 1090
rect 13103 1056 13109 1090
rect 13063 1017 13109 1056
rect 13063 983 13069 1017
rect 13103 983 13109 1017
rect 13063 944 13109 983
rect 13063 910 13069 944
rect 13103 910 13109 944
rect 13063 871 13109 910
rect 13063 837 13069 871
rect 13103 837 13109 871
rect 13063 798 13109 837
rect 13063 764 13069 798
rect 13103 764 13109 798
rect 13063 725 13109 764
rect 13063 691 13069 725
rect 13103 691 13109 725
rect 13063 652 13109 691
rect 13063 618 13069 652
rect 13103 618 13109 652
rect 13063 579 13109 618
rect 13063 545 13069 579
rect 13103 545 13109 579
rect 13063 506 13109 545
rect 13063 472 13069 506
rect 13103 472 13109 506
rect 13063 433 13109 472
rect 13063 399 13069 433
rect 13103 399 13109 433
rect 10193 360 12958 399
tri 12958 360 12997 399 nw
tri 13045 360 13063 378 se
rect 13063 360 13109 399
rect 10193 347 12945 360
tri 12945 347 12958 360 nw
tri 13032 347 13045 360 se
rect 13045 347 13069 360
rect 10193 326 12924 347
tri 12924 326 12945 347 nw
tri 13011 326 13032 347 se
rect 13032 326 13069 347
rect 13103 326 13109 360
rect 10193 316 12914 326
tri 12914 316 12924 326 nw
tri 13001 316 13011 326 se
rect 13011 316 13109 326
tri 12992 307 13001 316 se
rect 13001 307 13109 316
tri 9782 285 9791 294 se
rect 9791 285 9899 294
rect 1117 235 1185 269
rect 1219 260 1225 269
tri 1225 260 1250 285 sw
tri 9757 260 9782 285 se
rect 9782 260 9899 285
rect 9933 287 10050 294
tri 10050 287 10070 307 sw
tri 12972 287 12992 307 se
rect 12992 287 13109 307
rect 9933 260 10070 287
tri 10070 260 10097 287 sw
tri 12945 260 12972 287 se
rect 12972 260 13069 287
rect 1219 253 13069 260
rect 13103 253 13109 287
rect 1219 235 13109 253
rect 1117 222 13109 235
rect 1117 197 9899 222
rect 1117 163 1185 197
rect 1219 163 1257 197
rect 1291 163 1329 197
rect 1363 163 1401 197
rect 1435 163 1473 197
rect 1507 163 1545 197
rect 1579 163 1617 197
rect 1651 163 1689 197
rect 1723 163 1761 197
rect 1795 163 1833 197
rect 1867 163 1905 197
rect 1939 163 1977 197
rect 2011 163 2049 197
rect 2083 163 2121 197
rect 2155 163 2193 197
rect 2227 163 2265 197
rect 2299 163 2337 197
rect 2371 163 2409 197
rect 2443 163 2481 197
rect 2515 163 2553 197
rect 2587 163 2625 197
rect 2659 163 2697 197
rect 2731 163 2769 197
rect 2803 163 2841 197
rect 2875 163 2913 197
rect 2947 163 2985 197
rect 3019 163 3057 197
rect 3091 163 3129 197
rect 3163 163 3201 197
rect 3235 163 3273 197
rect 3307 163 3345 197
rect 3379 163 3417 197
rect 3451 163 3489 197
rect 3523 163 3561 197
rect 3595 163 3633 197
rect 3667 163 3705 197
rect 3739 163 3777 197
rect 3811 163 3849 197
rect 3883 163 3921 197
rect 3955 163 3993 197
rect 4027 163 4065 197
rect 4099 163 4137 197
rect 4171 163 4209 197
rect 4243 163 4281 197
rect 4315 163 4353 197
rect 4387 163 4425 197
rect 4459 163 4497 197
rect 4531 163 4569 197
rect 4603 163 4641 197
rect 4675 163 4713 197
rect 4747 163 4785 197
rect 4819 163 4857 197
rect 4891 163 4929 197
rect 4963 163 5001 197
rect 5035 163 5073 197
rect 5107 163 5145 197
rect 5179 163 5217 197
rect 5251 163 5289 197
rect 5323 163 5361 197
rect 5395 163 5433 197
rect 5467 163 5505 197
rect 5539 163 5577 197
rect 5611 163 5649 197
rect 5683 163 5721 197
rect 5755 163 5793 197
rect 5827 163 5865 197
rect 5899 163 5937 197
rect 5971 163 6009 197
rect 6043 163 6081 197
rect 6115 163 6153 197
rect 6187 163 6225 197
rect 6259 163 6297 197
rect 6331 163 6369 197
rect 6403 163 6441 197
rect 6475 163 6513 197
rect 6547 163 6585 197
rect 6619 163 6657 197
rect 6691 163 6729 197
rect 6763 163 6801 197
rect 6835 163 6873 197
rect 6907 163 6945 197
rect 6979 163 7017 197
rect 7051 163 7089 197
rect 7123 163 7161 197
rect 7195 163 7233 197
rect 7267 163 7305 197
rect 7339 163 7377 197
rect 7411 163 7449 197
rect 7483 163 7521 197
rect 7555 163 7593 197
rect 7627 163 7665 197
rect 7699 163 7737 197
rect 7771 163 7809 197
rect 7843 163 7881 197
rect 7915 163 7953 197
rect 7987 163 8025 197
rect 8059 163 8097 197
rect 8131 163 8169 197
rect 8203 163 8241 197
rect 8275 163 8313 197
rect 8347 163 8385 197
rect 8419 163 8457 197
rect 8491 163 8529 197
rect 8563 163 8601 197
rect 8635 163 8673 197
rect 8707 163 8745 197
rect 8779 163 8817 197
rect 8851 163 8889 197
rect 8923 163 8961 197
rect 8995 163 9033 197
rect 9067 163 9105 197
rect 9139 163 9177 197
rect 9211 163 9249 197
rect 9283 163 9321 197
rect 9355 163 9393 197
rect 9427 163 9465 197
rect 9499 163 9537 197
rect 9571 163 9609 197
rect 9643 163 9681 197
rect 9715 163 9754 197
rect 9788 163 9827 197
rect 9861 188 9899 197
rect 9933 214 13109 222
rect 9933 197 13069 214
rect 9933 188 9971 197
rect 9861 163 9971 188
rect 10005 163 10044 197
rect 10078 163 10117 197
rect 10151 163 10189 197
rect 10223 163 10261 197
rect 10295 163 10333 197
rect 10367 163 10405 197
rect 10439 163 10477 197
rect 10511 163 10549 197
rect 10583 163 10621 197
rect 10655 163 10693 197
rect 10727 163 10765 197
rect 10799 163 10837 197
rect 10871 163 10909 197
rect 10943 163 10981 197
rect 11015 163 11053 197
rect 11087 163 11125 197
rect 11159 163 11197 197
rect 11231 163 11269 197
rect 11303 163 11341 197
rect 11375 163 11413 197
rect 11447 163 11485 197
rect 11519 163 11557 197
rect 11591 163 11629 197
rect 11663 163 11701 197
rect 11735 163 11773 197
rect 11807 163 11845 197
rect 11879 163 11917 197
rect 11951 163 11989 197
rect 12023 163 12061 197
rect 12095 163 12133 197
rect 12167 163 12205 197
rect 12239 163 12277 197
rect 12311 163 12349 197
rect 12383 163 12421 197
rect 12455 163 12493 197
rect 12527 163 12565 197
rect 12599 163 12637 197
rect 12671 163 12709 197
rect 12743 163 12781 197
rect 12815 163 12853 197
rect 12887 163 12925 197
rect 12959 163 12997 197
rect 13031 180 13069 197
rect 13103 180 13109 214
rect 13031 166 13109 180
rect 13031 163 13080 166
rect 1117 137 13080 163
tri 13080 137 13109 166 nw
<< rmetal1 >>
rect 3212 14013 3214 14014
rect 3250 14013 3252 14014
rect 3212 13963 3213 14013
rect 3251 13963 3252 14013
rect 3212 13962 3214 13963
rect 3250 13962 3252 13963
rect 3214 13002 3216 13003
rect 3214 12952 3215 13002
rect 3214 12951 3216 12952
rect 3252 13002 3254 13003
rect 3253 12952 3254 13002
rect 3252 12951 3254 12952
rect 1984 1190 1986 1191
rect 1984 1185 1985 1190
rect 1984 1121 1985 1133
rect 1984 1064 1985 1069
rect 1984 1063 1986 1064
rect 2022 1190 2024 1191
rect 2023 1064 2024 1190
rect 2022 1063 2024 1064
rect 3033 1190 3035 1191
rect 3071 1190 3073 1191
rect 3033 1064 3034 1190
rect 3072 1064 3073 1190
rect 3033 1063 3035 1064
rect 3071 1063 3073 1064
rect 3928 11367 3930 11368
rect 3966 11367 3968 11368
rect 3928 3931 3929 11367
rect 3967 3931 3968 11367
rect 5320 11367 5322 11368
rect 5358 11367 5360 11368
rect 4453 3975 4455 3976
rect 3928 3930 3930 3931
rect 3966 3930 3968 3931
rect 4453 3931 4454 3975
rect 4453 3930 4455 3931
rect 4491 3975 4493 3976
rect 4492 3931 4493 3975
rect 4491 3930 4493 3931
rect 4769 3975 4771 3976
rect 4769 3931 4770 3975
rect 4769 3930 4771 3931
rect 4807 3975 4809 3976
rect 4808 3931 4809 3975
rect 4807 3930 4809 3931
rect 5320 3931 5321 11367
rect 5359 3931 5360 11367
rect 5320 3930 5322 3931
rect 5358 3930 5360 3931
rect 5788 11367 5790 11368
rect 5826 11367 5828 11368
rect 5788 7341 5789 11367
rect 5788 6819 5789 7161
rect 5788 5638 5789 6639
rect 5788 4203 5789 5458
rect 5788 3931 5789 4023
rect 5827 3931 5828 11367
rect 7861 14013 7863 14014
rect 7899 14013 7901 14014
rect 7861 13963 7862 14013
rect 7900 13963 7901 14013
rect 7861 13962 7863 13963
rect 7899 13962 7901 13963
rect 7829 13002 7831 13003
rect 7829 12952 7830 13002
rect 7829 12951 7831 12952
rect 7867 13002 7869 13003
rect 7868 12952 7869 13002
rect 7867 12951 7869 12952
rect 7181 11367 7183 11368
rect 7219 11367 7221 11368
rect 6299 3975 6301 3976
rect 5788 3930 5790 3931
rect 5826 3930 5828 3931
rect 6299 3931 6300 3975
rect 6299 3930 6301 3931
rect 6337 3975 6339 3976
rect 6338 3931 6339 3975
rect 6337 3930 6339 3931
rect 6606 3975 6608 3976
rect 6606 3931 6607 3975
rect 6606 3930 6608 3931
rect 6644 3975 6646 3976
rect 6645 3931 6646 3975
rect 6644 3930 6646 3931
rect 7181 3931 7182 11367
rect 7220 3931 7221 11367
rect 7181 3930 7183 3931
rect 7219 3930 7221 3931
rect 4133 2603 4191 2604
rect 4133 2602 4134 2603
rect 4190 2602 4191 2603
rect 4133 2565 4134 2566
rect 4190 2565 4191 2566
rect 4133 2564 4191 2565
rect 5973 2604 6031 2605
rect 5973 2603 5974 2604
rect 6030 2603 6031 2604
rect 5973 2566 5974 2567
rect 6030 2566 6031 2567
rect 5973 2565 6031 2566
rect 8075 1190 8077 1191
rect 8113 1190 8115 1191
rect 8075 1064 8076 1190
rect 8114 1064 8115 1190
rect 8075 1063 8077 1064
rect 8113 1063 8115 1064
rect 9123 1190 9125 1191
rect 9123 1064 9124 1190
rect 9123 1063 9125 1064
rect 9161 1190 9163 1191
rect 9162 1064 9163 1190
rect 9161 1063 9163 1064
<< via1 >>
rect 1348 13881 1400 13933
rect 1413 13881 1465 13933
rect 1176 11784 1228 11836
rect 1176 11723 1228 11763
rect 1176 11711 1185 11723
rect 1185 11711 1219 11723
rect 1219 11711 1228 11723
rect 1176 11689 1185 11690
rect 1185 11689 1219 11690
rect 1219 11689 1228 11690
rect 1176 11650 1228 11689
rect 1176 11638 1185 11650
rect 1185 11638 1219 11650
rect 1219 11638 1228 11650
rect 1176 11616 1185 11617
rect 1185 11616 1219 11617
rect 1219 11616 1228 11617
rect 1176 11577 1228 11616
rect 1604 13783 1656 13835
rect 1604 13715 1656 13767
rect 1604 13647 1656 13699
rect 1604 13579 1656 13631
rect 1604 13511 1656 13563
rect 1996 13309 2048 13361
rect 2073 13309 2125 13361
rect 2150 13309 2202 13361
rect 2227 13309 2279 13361
rect 2304 13309 2356 13361
rect 2384 13309 2436 13361
rect 2461 13309 2513 13361
rect 2538 13309 2590 13361
rect 2615 13309 2667 13361
rect 2692 13309 2744 13361
rect 2769 13309 2821 13361
rect 2843 13309 2895 13361
rect 2918 13309 2970 13361
rect 2993 13309 3045 13361
rect 1996 13241 2048 13293
rect 2073 13241 2125 13293
rect 2150 13241 2202 13293
rect 2227 13241 2279 13293
rect 2304 13241 2356 13293
rect 2384 13241 2436 13293
rect 2461 13241 2513 13293
rect 2538 13241 2590 13293
rect 2615 13241 2667 13293
rect 2692 13241 2744 13293
rect 2769 13241 2821 13293
rect 2843 13241 2895 13293
rect 2918 13241 2970 13293
rect 2993 13241 3045 13293
rect 1996 13173 2048 13225
rect 2073 13173 2125 13225
rect 2150 13173 2202 13225
rect 2227 13173 2279 13225
rect 2304 13173 2356 13225
rect 2384 13173 2436 13225
rect 2461 13173 2513 13225
rect 2538 13173 2590 13225
rect 2615 13173 2667 13225
rect 2692 13173 2744 13225
rect 2769 13173 2821 13225
rect 2843 13173 2895 13225
rect 2918 13173 2970 13225
rect 2993 13173 3045 13225
rect 1996 13105 2048 13157
rect 2073 13105 2125 13157
rect 2150 13105 2202 13157
rect 2227 13105 2279 13157
rect 2304 13105 2356 13157
rect 2384 13105 2436 13157
rect 2461 13105 2513 13157
rect 2538 13105 2590 13157
rect 2615 13105 2667 13157
rect 2692 13105 2744 13157
rect 2769 13105 2821 13157
rect 2843 13105 2895 13157
rect 2918 13105 2970 13157
rect 2993 13105 3045 13157
rect 1996 13037 2048 13089
rect 2073 13037 2125 13089
rect 2150 13037 2202 13089
rect 2227 13037 2279 13089
rect 2304 13037 2356 13089
rect 2384 13037 2436 13089
rect 2461 13037 2513 13089
rect 2538 13037 2590 13089
rect 2615 13037 2667 13089
rect 2692 13037 2744 13089
rect 2769 13037 2821 13089
rect 2843 13037 2895 13089
rect 2918 13037 2970 13089
rect 2993 13037 3045 13089
rect 3135 12945 3187 12997
rect 3135 12881 3187 12933
rect 1447 12458 1499 12467
rect 1447 12424 1474 12458
rect 1474 12424 1499 12458
rect 1447 12415 1499 12424
rect 1511 12458 1563 12467
rect 1511 12424 1529 12458
rect 1529 12424 1563 12458
rect 1511 12415 1563 12424
rect 3477 12591 3529 12643
rect 3477 12527 3529 12579
rect 3688 13312 3740 13361
rect 3688 13309 3700 13312
rect 3700 13309 3734 13312
rect 3734 13309 3740 13312
rect 3762 13312 3814 13361
rect 3762 13309 3772 13312
rect 3772 13309 3806 13312
rect 3806 13309 3814 13312
rect 3838 13312 3890 13361
rect 3838 13309 3844 13312
rect 3844 13309 3878 13312
rect 3878 13309 3890 13312
rect 3688 13278 3700 13293
rect 3700 13278 3734 13293
rect 3734 13278 3740 13293
rect 3688 13241 3740 13278
rect 3762 13278 3772 13293
rect 3772 13278 3806 13293
rect 3806 13278 3814 13293
rect 3762 13241 3814 13278
rect 3838 13278 3844 13293
rect 3844 13278 3878 13293
rect 3878 13278 3890 13293
rect 3838 13241 3890 13278
rect 3688 13173 3740 13225
rect 3762 13173 3814 13225
rect 3838 13173 3890 13225
rect 3688 13105 3740 13157
rect 3762 13105 3814 13157
rect 3838 13105 3890 13157
rect 3688 13037 3740 13089
rect 3762 13037 3814 13089
rect 3838 13037 3890 13089
rect 3975 12951 4027 13003
rect 4039 12951 4091 13003
rect 4103 12972 4155 13003
rect 4103 12951 4131 12972
rect 4131 12951 4155 12972
rect 1176 11565 1185 11577
rect 1185 11565 1219 11577
rect 1219 11565 1228 11577
rect 1176 11543 1185 11544
rect 1185 11543 1219 11544
rect 1219 11543 1228 11544
rect 1176 11504 1228 11543
rect 1176 11492 1185 11504
rect 1185 11492 1219 11504
rect 1219 11492 1228 11504
rect 1176 11431 1228 11470
rect 1176 11418 1185 11431
rect 1185 11418 1219 11431
rect 1219 11418 1228 11431
rect 1117 10189 1169 10241
rect 1181 10205 1233 10241
rect 1181 10189 1185 10205
rect 1185 10189 1219 10205
rect 1219 10189 1233 10205
rect 1117 10062 1169 10114
rect 1181 10099 1185 10114
rect 1185 10099 1219 10114
rect 1219 10099 1233 10114
rect 1181 10062 1233 10099
rect 1117 8117 1233 8146
rect 1117 8083 1185 8117
rect 1185 8083 1219 8117
rect 1219 8083 1233 8117
rect 1117 8045 1233 8083
rect 1117 8030 1185 8045
rect 1185 8030 1219 8045
rect 1219 8030 1233 8045
rect 1117 7965 1169 8017
rect 1181 8011 1185 8017
rect 1185 8011 1219 8017
rect 1219 8011 1233 8017
rect 1181 7973 1233 8011
rect 1181 7965 1185 7973
rect 1185 7965 1219 7973
rect 1219 7965 1233 7973
rect 1117 4828 1169 4880
rect 1181 4877 1233 4880
rect 1181 4843 1185 4877
rect 1185 4843 1219 4877
rect 1219 4843 1233 4877
rect 1181 4828 1233 4843
rect 1117 4762 1169 4814
rect 1181 4805 1233 4814
rect 1181 4771 1185 4805
rect 1185 4771 1219 4805
rect 1219 4771 1233 4805
rect 1181 4762 1233 4771
rect 1758 12103 1874 12120
rect 1758 12069 1777 12103
rect 1777 12069 1836 12103
rect 1836 12069 1870 12103
rect 1870 12069 1874 12103
rect 1758 12031 1874 12069
rect 1758 12004 1777 12031
rect 1777 12004 1836 12031
rect 1836 12004 1870 12031
rect 1870 12004 1874 12031
rect 2048 12154 2164 12270
rect 1624 11723 1676 11732
rect 1624 11689 1630 11723
rect 1630 11689 1664 11723
rect 1664 11689 1676 11723
rect 1624 11680 1676 11689
rect 1689 11723 1741 11732
rect 1754 11723 1806 11732
rect 1819 11723 1871 11732
rect 1884 11723 1936 11732
rect 1689 11689 1713 11723
rect 1713 11689 1741 11723
rect 1754 11689 1796 11723
rect 1796 11689 1806 11723
rect 1819 11689 1830 11723
rect 1830 11689 1871 11723
rect 1884 11689 1913 11723
rect 1913 11689 1936 11723
rect 1689 11680 1741 11689
rect 1754 11680 1806 11689
rect 1819 11680 1871 11689
rect 1884 11680 1936 11689
rect 1950 11723 2002 11732
rect 1950 11689 1962 11723
rect 1962 11689 1996 11723
rect 1996 11689 2002 11723
rect 1950 11680 2002 11689
rect 1384 9846 1436 9849
rect 1384 9812 1396 9846
rect 1396 9812 1430 9846
rect 1430 9812 1436 9846
rect 1384 9797 1436 9812
rect 1384 9772 1436 9783
rect 1384 9738 1396 9772
rect 1396 9738 1430 9772
rect 1430 9738 1436 9772
rect 1384 9731 1436 9738
rect 1384 6468 1436 6474
rect 1384 6434 1396 6468
rect 1396 6434 1430 6468
rect 1430 6434 1436 6468
rect 1384 6422 1436 6434
rect 1384 6394 1436 6408
rect 1384 6360 1396 6394
rect 1396 6360 1430 6394
rect 1430 6360 1436 6394
rect 1384 6356 1436 6360
rect 1384 1155 1436 1185
rect 1384 1133 1396 1155
rect 1396 1133 1430 1155
rect 1430 1133 1436 1155
rect 1384 1080 1436 1121
rect 1384 1069 1396 1080
rect 1396 1069 1430 1080
rect 1430 1069 1436 1080
rect 1532 866 1584 918
rect 1532 802 1584 854
rect 2720 12103 2836 12120
rect 2720 12069 2746 12103
rect 2746 12069 2780 12103
rect 2780 12069 2823 12103
rect 2823 12069 2836 12103
rect 2720 12031 2836 12069
rect 2720 12004 2746 12031
rect 2746 12004 2780 12031
rect 2780 12004 2823 12031
rect 2823 12004 2836 12031
rect 2224 11723 2276 11732
rect 2224 11689 2230 11723
rect 2230 11689 2264 11723
rect 2264 11689 2276 11723
rect 2224 11680 2276 11689
rect 2292 11723 2344 11732
rect 2292 11689 2302 11723
rect 2302 11689 2336 11723
rect 2336 11689 2344 11723
rect 2292 11680 2344 11689
rect 2360 11723 2412 11732
rect 2360 11689 2374 11723
rect 2374 11689 2408 11723
rect 2408 11689 2412 11723
rect 2360 11680 2412 11689
rect 2428 11723 2480 11732
rect 2428 11689 2446 11723
rect 2446 11689 2480 11723
rect 2428 11680 2480 11689
rect 2496 11723 2548 11732
rect 2564 11723 2616 11732
rect 2632 11723 2684 11732
rect 2700 11723 2752 11732
rect 2768 11723 2820 11732
rect 2836 11723 2888 11732
rect 2904 11723 2956 11732
rect 2972 11723 3024 11732
rect 3040 11723 3092 11732
rect 3108 11723 3160 11732
rect 2496 11689 2518 11723
rect 2518 11689 2548 11723
rect 2564 11689 2591 11723
rect 2591 11689 2616 11723
rect 2632 11689 2664 11723
rect 2664 11689 2684 11723
rect 2700 11689 2737 11723
rect 2737 11689 2752 11723
rect 2768 11689 2771 11723
rect 2771 11689 2810 11723
rect 2810 11689 2820 11723
rect 2836 11689 2844 11723
rect 2844 11689 2883 11723
rect 2883 11689 2888 11723
rect 2904 11689 2917 11723
rect 2917 11689 2956 11723
rect 2972 11689 2990 11723
rect 2990 11689 3024 11723
rect 3040 11689 3063 11723
rect 3063 11689 3092 11723
rect 3108 11689 3136 11723
rect 3136 11689 3160 11723
rect 2496 11680 2548 11689
rect 2564 11680 2616 11689
rect 2632 11680 2684 11689
rect 2700 11680 2752 11689
rect 2768 11680 2820 11689
rect 2836 11680 2888 11689
rect 2904 11680 2956 11689
rect 2972 11680 3024 11689
rect 3040 11680 3092 11689
rect 3108 11680 3160 11689
rect 3175 11723 3227 11732
rect 3175 11689 3209 11723
rect 3209 11689 3227 11723
rect 3175 11680 3227 11689
rect 3242 11723 3294 11732
rect 3242 11689 3248 11723
rect 3248 11689 3282 11723
rect 3282 11689 3294 11723
rect 3242 11680 3294 11689
rect 3309 11723 3361 11732
rect 3309 11689 3321 11723
rect 3321 11689 3355 11723
rect 3355 11689 3361 11723
rect 3309 11680 3361 11689
rect 3767 12004 3883 12120
rect 3681 11784 3733 11836
rect 3681 11723 3733 11762
rect 3681 11710 3693 11723
rect 3693 11710 3727 11723
rect 3727 11710 3733 11723
rect 3681 11650 3733 11688
rect 3681 11636 3693 11650
rect 3693 11636 3727 11650
rect 3727 11636 3733 11650
rect 3681 11577 3733 11614
rect 3681 11562 3693 11577
rect 3693 11562 3727 11577
rect 3727 11562 3733 11577
rect 2983 7532 3035 7584
rect 3047 7532 3099 7584
rect 3111 7532 3163 7584
rect 3175 7532 3227 7584
rect 3681 11504 3733 11540
rect 3681 11488 3693 11504
rect 3693 11488 3727 11504
rect 3727 11488 3733 11504
rect 3681 11431 3733 11467
rect 4526 13309 4578 13361
rect 4601 13309 4653 13361
rect 4676 13309 4728 13361
rect 4526 13241 4578 13293
rect 4601 13241 4653 13293
rect 4676 13241 4728 13293
rect 4526 13173 4578 13225
rect 4601 13173 4653 13225
rect 4676 13173 4728 13225
rect 4526 13105 4578 13157
rect 4601 13105 4653 13157
rect 4676 13105 4728 13157
rect 4526 13037 4578 13089
rect 4601 13037 4653 13089
rect 4676 13037 4728 13089
rect 5262 13921 5314 13933
rect 5262 13887 5268 13921
rect 5268 13887 5302 13921
rect 5302 13887 5314 13921
rect 5262 13881 5314 13887
rect 5326 13921 5378 13933
rect 5326 13887 5342 13921
rect 5342 13887 5376 13921
rect 5376 13887 5378 13921
rect 5326 13881 5378 13887
rect 5390 13921 5442 13933
rect 5454 13921 5506 13933
rect 5518 13921 5570 13933
rect 5582 13921 5634 13933
rect 5646 13921 5698 13933
rect 5390 13887 5416 13921
rect 5416 13887 5442 13921
rect 5454 13887 5490 13921
rect 5490 13887 5506 13921
rect 5518 13887 5524 13921
rect 5524 13887 5564 13921
rect 5564 13887 5570 13921
rect 5582 13887 5598 13921
rect 5598 13887 5634 13921
rect 5646 13887 5672 13921
rect 5672 13887 5698 13921
rect 5390 13881 5442 13887
rect 5454 13881 5506 13887
rect 5518 13881 5570 13887
rect 5582 13881 5634 13887
rect 5646 13881 5698 13887
rect 5710 13921 5762 13933
rect 5710 13887 5712 13921
rect 5712 13887 5746 13921
rect 5746 13887 5762 13921
rect 5710 13881 5762 13887
rect 5774 13921 5826 13933
rect 5774 13887 5786 13921
rect 5786 13887 5820 13921
rect 5820 13887 5826 13921
rect 5774 13881 5826 13887
rect 4813 12951 4865 13003
rect 4877 12951 4929 13003
rect 4941 12951 4993 13003
rect 4475 12218 4527 12270
rect 4475 12154 4527 12206
rect 4493 11723 4545 11732
rect 4493 11689 4499 11723
rect 4499 11689 4533 11723
rect 4533 11689 4545 11723
rect 4493 11680 4545 11689
rect 4565 11723 4617 11732
rect 4565 11689 4573 11723
rect 4573 11689 4607 11723
rect 4607 11689 4617 11723
rect 4565 11680 4617 11689
rect 4637 11723 4689 11732
rect 4637 11689 4647 11723
rect 4647 11689 4681 11723
rect 4681 11689 4689 11723
rect 4637 11680 4689 11689
rect 4709 11723 4761 11732
rect 4709 11689 4721 11723
rect 4721 11689 4755 11723
rect 4755 11689 4761 11723
rect 4709 11680 4761 11689
rect 3681 11415 3693 11431
rect 3693 11415 3727 11431
rect 3727 11415 3733 11431
rect 3681 10207 3733 10243
rect 3681 10191 3693 10207
rect 3693 10191 3727 10207
rect 3727 10191 3733 10207
rect 3681 10173 3693 10179
rect 3693 10173 3727 10179
rect 3727 10173 3733 10179
rect 3681 10135 3733 10173
rect 3681 10127 3693 10135
rect 3693 10127 3727 10135
rect 3727 10127 3733 10135
rect 3681 10101 3693 10114
rect 3693 10101 3727 10114
rect 3727 10101 3733 10114
rect 3681 10063 3733 10101
rect 3681 10062 3693 10063
rect 3693 10062 3727 10063
rect 3727 10062 3733 10063
rect 3500 9846 3552 9849
rect 3500 9812 3506 9846
rect 3506 9812 3540 9846
rect 3540 9812 3552 9846
rect 3500 9797 3552 9812
rect 3500 9772 3552 9783
rect 3500 9738 3506 9772
rect 3506 9738 3540 9772
rect 3540 9738 3552 9772
rect 3500 9731 3552 9738
rect 3681 8119 3733 8146
rect 3681 8094 3693 8119
rect 3693 8094 3727 8119
rect 3727 8094 3733 8119
rect 3681 8047 3733 8082
rect 3681 8030 3693 8047
rect 3693 8030 3727 8047
rect 3727 8030 3733 8047
rect 3681 8013 3693 8017
rect 3693 8013 3727 8017
rect 3727 8013 3733 8017
rect 3681 7975 3733 8013
rect 3681 7965 3693 7975
rect 3693 7965 3727 7975
rect 3727 7965 3733 7975
rect 3340 3909 3392 3961
rect 3404 3909 3456 3961
rect 1933 1133 1985 1185
rect 1933 1069 1985 1121
rect 1833 602 1904 624
rect 1904 602 1938 624
rect 1938 602 1949 624
rect 1833 564 1949 602
rect 1833 530 1904 564
rect 1904 530 1938 564
rect 1938 530 1949 564
rect 1833 508 1949 530
rect 2354 1536 2406 1588
rect 2420 1536 2472 1588
rect 2486 1536 2538 1588
rect 2552 1536 2604 1588
rect 2618 1536 2670 1588
rect 2684 1536 2736 1588
rect 2749 1536 2801 1588
rect 2814 1536 2866 1588
rect 2879 1536 2931 1588
rect 2944 1536 2996 1588
rect 2354 1472 2406 1524
rect 2420 1472 2472 1524
rect 2486 1472 2538 1524
rect 2552 1472 2604 1524
rect 2618 1472 2670 1524
rect 2684 1472 2736 1524
rect 2749 1472 2801 1524
rect 2814 1472 2866 1524
rect 2879 1472 2931 1524
rect 2944 1472 2996 1524
rect 2354 1408 2406 1460
rect 2420 1408 2472 1460
rect 2486 1408 2538 1460
rect 2552 1408 2604 1460
rect 2618 1408 2670 1460
rect 2684 1408 2736 1460
rect 2749 1408 2801 1460
rect 2814 1408 2866 1460
rect 2879 1408 2931 1460
rect 2944 1408 2996 1460
rect 2354 1344 2406 1396
rect 2420 1344 2472 1396
rect 2486 1344 2538 1396
rect 2552 1344 2604 1396
rect 2618 1344 2670 1396
rect 2684 1344 2736 1396
rect 2749 1344 2801 1396
rect 2814 1344 2866 1396
rect 2879 1344 2931 1396
rect 2944 1344 2996 1396
rect 2354 1280 2406 1332
rect 2420 1280 2472 1332
rect 2486 1280 2538 1332
rect 2552 1280 2604 1332
rect 2618 1280 2670 1332
rect 2684 1280 2736 1332
rect 2749 1280 2801 1332
rect 2814 1280 2866 1332
rect 2879 1280 2931 1332
rect 2944 1280 2996 1332
rect 3073 1133 3125 1185
rect 3073 1069 3125 1121
rect 3500 6468 3552 6474
rect 3500 6434 3506 6468
rect 3506 6434 3540 6468
rect 3540 6434 3552 6468
rect 3500 6422 3552 6434
rect 3500 6394 3552 6408
rect 3500 6360 3506 6394
rect 3506 6360 3540 6394
rect 3540 6360 3552 6394
rect 3500 6356 3552 6360
rect 3681 4879 3733 4880
rect 3681 4845 3693 4879
rect 3693 4845 3727 4879
rect 3727 4845 3733 4879
rect 3681 4828 3733 4845
rect 3681 4807 3733 4814
rect 3681 4773 3693 4807
rect 3693 4773 3727 4807
rect 3727 4773 3733 4807
rect 3681 4762 3733 4773
rect 3768 7161 3884 7341
rect 3768 6639 3884 6819
rect 3768 5458 3884 5638
rect 3768 4023 3884 4203
rect 4070 8951 4122 8983
rect 4070 8931 4082 8951
rect 4082 8931 4116 8951
rect 4116 8931 4122 8951
rect 4070 8877 4122 8917
rect 4070 8865 4082 8877
rect 4082 8865 4116 8877
rect 4116 8865 4122 8877
rect 4070 5271 4082 5282
rect 4082 5271 4116 5282
rect 4116 5271 4122 5282
rect 4070 5230 4122 5271
rect 4070 5196 4082 5216
rect 4082 5196 4116 5216
rect 4116 5196 4122 5216
rect 4070 5164 4122 5196
rect 5215 13829 5267 13835
rect 5215 13795 5224 13829
rect 5224 13795 5258 13829
rect 5258 13795 5267 13829
rect 5215 13783 5267 13795
rect 5215 13753 5267 13767
rect 5215 13719 5224 13753
rect 5224 13719 5258 13753
rect 5258 13719 5267 13753
rect 5215 13715 5267 13719
rect 5215 13677 5267 13699
rect 5215 13647 5224 13677
rect 5224 13647 5258 13677
rect 5258 13647 5267 13677
rect 5215 13602 5267 13631
rect 5215 13579 5224 13602
rect 5224 13579 5258 13602
rect 5258 13579 5267 13602
rect 5215 13527 5267 13563
rect 5215 13511 5224 13527
rect 5224 13511 5258 13527
rect 5258 13511 5267 13527
rect 5371 13343 5380 13361
rect 5380 13343 5414 13361
rect 5414 13343 5423 13361
rect 5371 13309 5423 13343
rect 5371 13268 5380 13293
rect 5380 13268 5414 13293
rect 5414 13268 5423 13293
rect 5371 13241 5423 13268
rect 5371 13193 5380 13225
rect 5380 13193 5414 13225
rect 5414 13193 5423 13225
rect 5371 13173 5423 13193
rect 5371 13152 5423 13157
rect 5371 13118 5380 13152
rect 5380 13118 5414 13152
rect 5414 13118 5423 13152
rect 5371 13105 5423 13118
rect 5371 13077 5423 13089
rect 5371 13043 5380 13077
rect 5380 13043 5414 13077
rect 5414 13043 5423 13077
rect 5371 13037 5423 13043
rect 5527 13829 5579 13835
rect 5527 13795 5536 13829
rect 5536 13795 5570 13829
rect 5570 13795 5579 13829
rect 5527 13783 5579 13795
rect 5527 13753 5579 13767
rect 5527 13719 5536 13753
rect 5536 13719 5570 13753
rect 5570 13719 5579 13753
rect 5527 13715 5579 13719
rect 5527 13677 5579 13699
rect 5527 13647 5536 13677
rect 5536 13647 5570 13677
rect 5570 13647 5579 13677
rect 5527 13602 5579 13631
rect 5527 13579 5536 13602
rect 5536 13579 5570 13602
rect 5570 13579 5579 13602
rect 5527 13527 5579 13563
rect 5527 13511 5536 13527
rect 5536 13511 5570 13527
rect 5570 13511 5579 13527
rect 5683 13343 5692 13361
rect 5692 13343 5726 13361
rect 5726 13343 5735 13361
rect 5683 13309 5735 13343
rect 5683 13268 5692 13293
rect 5692 13268 5726 13293
rect 5726 13268 5735 13293
rect 5683 13241 5735 13268
rect 5683 13193 5692 13225
rect 5692 13193 5726 13225
rect 5726 13193 5735 13225
rect 5683 13173 5735 13193
rect 5683 13152 5735 13157
rect 5683 13118 5692 13152
rect 5692 13118 5726 13152
rect 5726 13118 5735 13152
rect 5683 13105 5735 13118
rect 5683 13077 5735 13089
rect 5683 13043 5692 13077
rect 5692 13043 5726 13077
rect 5726 13043 5735 13077
rect 5683 13037 5735 13043
rect 5839 13829 5891 13835
rect 5839 13795 5848 13829
rect 5848 13795 5882 13829
rect 5882 13795 5891 13829
rect 5839 13783 5891 13795
rect 5839 13753 5891 13767
rect 5839 13719 5848 13753
rect 5848 13719 5882 13753
rect 5882 13719 5891 13753
rect 5839 13715 5891 13719
rect 5839 13677 5891 13699
rect 5839 13647 5848 13677
rect 5848 13647 5882 13677
rect 5882 13647 5891 13677
rect 5839 13602 5891 13631
rect 5839 13579 5848 13602
rect 5848 13579 5882 13602
rect 5882 13579 5891 13602
rect 5839 13527 5891 13563
rect 5839 13511 5848 13527
rect 5848 13511 5882 13527
rect 5882 13511 5891 13527
rect 5447 12626 5457 12643
rect 5457 12626 5491 12643
rect 5491 12626 5499 12643
rect 5447 12591 5499 12626
rect 5447 12560 5499 12579
rect 5447 12527 5457 12560
rect 5457 12527 5491 12560
rect 5491 12527 5499 12560
rect 5495 12458 5547 12467
rect 5495 12424 5500 12458
rect 5500 12424 5534 12458
rect 5534 12424 5547 12458
rect 5495 12415 5547 12424
rect 5559 12458 5611 12467
rect 5559 12424 5572 12458
rect 5572 12424 5606 12458
rect 5606 12424 5611 12458
rect 5559 12415 5611 12424
rect 5478 12103 5594 12120
rect 5478 12069 5497 12103
rect 5497 12069 5541 12103
rect 5541 12069 5575 12103
rect 5575 12069 5594 12103
rect 5478 12031 5594 12069
rect 5478 12004 5497 12031
rect 5497 12004 5541 12031
rect 5541 12004 5575 12031
rect 5575 12004 5594 12031
rect 5055 11723 5107 11732
rect 5055 11689 5061 11723
rect 5061 11689 5095 11723
rect 5095 11689 5107 11723
rect 5055 11680 5107 11689
rect 5122 11723 5174 11732
rect 5189 11723 5241 11732
rect 5256 11723 5308 11732
rect 5323 11723 5375 11732
rect 5122 11689 5145 11723
rect 5145 11689 5174 11723
rect 5189 11689 5230 11723
rect 5230 11689 5241 11723
rect 5256 11689 5264 11723
rect 5264 11689 5308 11723
rect 5323 11689 5349 11723
rect 5349 11689 5375 11723
rect 5122 11680 5174 11689
rect 5189 11680 5241 11689
rect 5256 11680 5308 11689
rect 5323 11680 5375 11689
rect 5390 11723 5442 11732
rect 5390 11689 5400 11723
rect 5400 11689 5434 11723
rect 5434 11689 5442 11723
rect 5390 11680 5442 11689
rect 5457 11723 5509 11732
rect 5524 11723 5576 11732
rect 5591 11723 5643 11732
rect 5657 11723 5709 11732
rect 5723 11723 5775 11732
rect 5789 11723 5841 11732
rect 5855 11723 5907 11732
rect 5457 11689 5485 11723
rect 5485 11689 5509 11723
rect 5524 11689 5557 11723
rect 5557 11689 5576 11723
rect 5591 11689 5629 11723
rect 5629 11689 5643 11723
rect 5657 11689 5663 11723
rect 5663 11689 5703 11723
rect 5703 11689 5709 11723
rect 5723 11689 5737 11723
rect 5737 11689 5775 11723
rect 5789 11689 5811 11723
rect 5811 11689 5841 11723
rect 5855 11689 5885 11723
rect 5885 11689 5907 11723
rect 5457 11680 5509 11689
rect 5524 11680 5576 11689
rect 5591 11680 5643 11689
rect 5657 11680 5709 11689
rect 5723 11680 5775 11689
rect 5789 11680 5841 11689
rect 5855 11680 5907 11689
rect 5921 11723 5973 11732
rect 5921 11689 5925 11723
rect 5925 11689 5959 11723
rect 5959 11689 5973 11723
rect 5921 11680 5973 11689
rect 5987 11723 6039 11732
rect 5987 11689 5999 11723
rect 5999 11689 6033 11723
rect 6033 11689 6039 11723
rect 5987 11680 6039 11689
rect 6366 13783 6418 13835
rect 6442 13783 6494 13835
rect 6516 13783 6568 13835
rect 6366 13715 6418 13767
rect 6442 13715 6494 13767
rect 6516 13715 6568 13767
rect 6366 13647 6418 13699
rect 6442 13647 6494 13699
rect 6516 13647 6568 13699
rect 6366 13579 6418 13631
rect 6442 13579 6494 13631
rect 6516 13579 6568 13631
rect 6366 13511 6418 13563
rect 6442 13511 6494 13563
rect 6516 13511 6568 13563
rect 6653 12951 6705 13003
rect 6717 12951 6769 13003
rect 6781 12951 6833 13003
rect 6315 12218 6367 12270
rect 6315 12154 6367 12206
rect 6333 11723 6385 11732
rect 6333 11689 6339 11723
rect 6339 11689 6373 11723
rect 6373 11689 6385 11723
rect 6333 11680 6385 11689
rect 6405 11723 6457 11732
rect 6405 11689 6413 11723
rect 6413 11689 6447 11723
rect 6447 11689 6457 11723
rect 6405 11680 6457 11689
rect 6477 11723 6529 11732
rect 6477 11689 6487 11723
rect 6487 11689 6521 11723
rect 6521 11689 6529 11723
rect 6477 11680 6529 11689
rect 6549 11723 6601 11732
rect 6549 11689 6561 11723
rect 6561 11689 6595 11723
rect 6595 11689 6601 11723
rect 6549 11680 6601 11689
rect 4850 9797 4902 9849
rect 4930 9797 4982 9849
rect 4850 9731 4902 9783
rect 4930 9731 4982 9783
rect 5186 10959 5238 10967
rect 5186 10925 5192 10959
rect 5192 10925 5226 10959
rect 5226 10925 5238 10959
rect 5186 10915 5238 10925
rect 5186 10885 5238 10901
rect 5186 10851 5192 10885
rect 5192 10851 5226 10885
rect 5226 10851 5238 10885
rect 5186 10849 5238 10851
rect 5186 7017 5238 7043
rect 5186 6991 5192 7017
rect 5192 6991 5226 7017
rect 5226 6991 5238 7017
rect 5186 6942 5238 6977
rect 5186 6925 5192 6942
rect 5192 6925 5226 6942
rect 5226 6925 5238 6942
rect 5367 4023 5483 4203
rect 5548 10211 5600 10243
rect 5548 10191 5557 10211
rect 5557 10191 5591 10211
rect 5591 10191 5600 10211
rect 5548 10177 5557 10179
rect 5557 10177 5591 10179
rect 5591 10177 5600 10179
rect 5548 10139 5600 10177
rect 5548 10127 5557 10139
rect 5557 10127 5591 10139
rect 5591 10127 5600 10139
rect 5548 10105 5557 10114
rect 5557 10105 5591 10114
rect 5591 10105 5600 10114
rect 5548 10067 5600 10105
rect 5548 10062 5557 10067
rect 5557 10062 5591 10067
rect 5591 10062 5600 10067
rect 5548 8123 5600 8146
rect 5548 8094 5557 8123
rect 5557 8094 5591 8123
rect 5591 8094 5600 8123
rect 5548 8051 5600 8082
rect 5548 8030 5557 8051
rect 5557 8030 5591 8051
rect 5591 8030 5600 8051
rect 5548 7979 5600 8017
rect 5548 7965 5557 7979
rect 5557 7965 5591 7979
rect 5591 7965 5600 7979
rect 5548 4855 5600 4880
rect 5548 4828 5557 4855
rect 5557 4828 5591 4855
rect 5591 4828 5600 4855
rect 5548 4782 5600 4814
rect 5548 4762 5557 4782
rect 5557 4762 5591 4782
rect 5591 4762 5600 4782
rect 5678 7161 5794 7341
rect 5678 6639 5794 6819
rect 5678 5458 5794 5638
rect 5678 4023 5794 4203
rect 5910 8951 5962 8983
rect 5910 8931 5922 8951
rect 5922 8931 5956 8951
rect 5956 8931 5962 8951
rect 5910 8877 5962 8917
rect 5910 8865 5922 8877
rect 5922 8865 5956 8877
rect 5956 8865 5962 8877
rect 5910 5271 5922 5282
rect 5922 5271 5956 5282
rect 5956 5271 5962 5282
rect 5910 5230 5962 5271
rect 5910 5196 5922 5216
rect 5922 5196 5956 5216
rect 5956 5196 5962 5216
rect 5910 5164 5962 5196
rect 6930 12972 6982 13003
rect 6930 12951 6963 12972
rect 6963 12951 6982 12972
rect 6994 12951 7046 13003
rect 7058 12951 7110 13003
rect 7204 13824 7256 13835
rect 7204 13790 7216 13824
rect 7216 13790 7250 13824
rect 7250 13790 7256 13824
rect 7204 13783 7256 13790
rect 7279 13824 7331 13835
rect 7279 13790 7288 13824
rect 7288 13790 7322 13824
rect 7322 13790 7331 13824
rect 7279 13783 7331 13790
rect 7354 13824 7406 13835
rect 7354 13790 7360 13824
rect 7360 13790 7394 13824
rect 7394 13790 7406 13824
rect 7354 13783 7406 13790
rect 7204 13715 7256 13767
rect 7279 13715 7331 13767
rect 7354 13715 7406 13767
rect 7204 13647 7256 13699
rect 7279 13647 7331 13699
rect 7354 13647 7406 13699
rect 7204 13579 7256 13631
rect 7279 13579 7331 13631
rect 7354 13579 7406 13631
rect 7204 13511 7256 13563
rect 7279 13511 7331 13563
rect 7354 13511 7406 13563
rect 7263 12103 7379 12120
rect 7263 12069 7301 12103
rect 7301 12069 7335 12103
rect 7335 12069 7379 12103
rect 7263 12031 7379 12069
rect 7263 12004 7301 12031
rect 7301 12004 7335 12031
rect 7335 12004 7379 12031
rect 7417 11784 7469 11836
rect 7417 11723 7469 11763
rect 7417 11711 7423 11723
rect 7423 11711 7457 11723
rect 7457 11711 7469 11723
rect 7417 11650 7469 11689
rect 8053 13783 8105 13835
rect 8130 13783 8182 13835
rect 8207 13783 8259 13835
rect 8284 13783 8336 13835
rect 8361 13783 8413 13835
rect 8441 13783 8493 13835
rect 8518 13783 8570 13835
rect 8595 13783 8647 13835
rect 8672 13783 8724 13835
rect 8749 13783 8801 13835
rect 8826 13783 8878 13835
rect 8900 13783 8952 13835
rect 8975 13783 9027 13835
rect 9050 13783 9102 13835
rect 8053 13715 8105 13767
rect 8130 13715 8182 13767
rect 8207 13715 8259 13767
rect 8284 13715 8336 13767
rect 8361 13715 8413 13767
rect 8441 13715 8493 13767
rect 8518 13715 8570 13767
rect 8595 13715 8647 13767
rect 8672 13715 8724 13767
rect 8749 13715 8801 13767
rect 8826 13715 8878 13767
rect 8900 13715 8952 13767
rect 8975 13715 9027 13767
rect 9050 13715 9102 13767
rect 8053 13647 8105 13699
rect 8130 13647 8182 13699
rect 8207 13647 8259 13699
rect 8284 13647 8336 13699
rect 8361 13647 8413 13699
rect 8441 13647 8493 13699
rect 8518 13647 8570 13699
rect 8595 13647 8647 13699
rect 8672 13647 8724 13699
rect 8749 13647 8801 13699
rect 8826 13647 8878 13699
rect 8900 13647 8952 13699
rect 8975 13647 9027 13699
rect 9050 13647 9102 13699
rect 8053 13579 8105 13631
rect 8130 13579 8182 13631
rect 8207 13579 8259 13631
rect 8284 13579 8336 13631
rect 8361 13579 8413 13631
rect 8441 13579 8493 13631
rect 8518 13579 8570 13631
rect 8595 13579 8647 13631
rect 8672 13579 8724 13631
rect 8749 13579 8801 13631
rect 8826 13579 8878 13631
rect 8900 13579 8952 13631
rect 8975 13579 9027 13631
rect 9050 13579 9102 13631
rect 8053 13511 8105 13563
rect 8130 13511 8182 13563
rect 8207 13511 8259 13563
rect 8284 13511 8336 13563
rect 8361 13511 8413 13563
rect 8441 13511 8493 13563
rect 8518 13511 8570 13563
rect 8595 13511 8647 13563
rect 8672 13511 8724 13563
rect 8749 13511 8801 13563
rect 8826 13511 8878 13563
rect 8900 13511 8952 13563
rect 8975 13511 9027 13563
rect 9050 13511 9102 13563
rect 7895 13021 7947 13073
rect 7895 12957 7947 13009
rect 9516 13921 9568 13933
rect 9516 13887 9522 13921
rect 9522 13887 9556 13921
rect 9556 13887 9568 13921
rect 9516 13881 9568 13887
rect 9608 13921 9660 13933
rect 9608 13887 9617 13921
rect 9617 13887 9651 13921
rect 9651 13887 9660 13921
rect 9608 13881 9660 13887
rect 9700 13921 9752 13933
rect 9700 13887 9712 13921
rect 9712 13887 9746 13921
rect 9746 13887 9752 13921
rect 9700 13881 9752 13887
rect 9452 13427 9461 13449
rect 9461 13427 9495 13449
rect 9495 13427 9504 13449
rect 9452 13397 9504 13427
rect 9452 13353 9461 13385
rect 9461 13353 9495 13385
rect 9495 13353 9504 13385
rect 9452 13333 9504 13353
rect 9452 13313 9504 13321
rect 9452 13279 9461 13313
rect 9461 13279 9495 13313
rect 9495 13279 9504 13313
rect 9452 13269 9504 13279
rect 9452 13239 9504 13257
rect 9452 13205 9461 13239
rect 9461 13205 9495 13239
rect 9495 13205 9504 13239
rect 9452 13165 9504 13193
rect 9452 13141 9461 13165
rect 9461 13141 9495 13165
rect 9495 13141 9504 13165
rect 9764 13427 9773 13449
rect 9773 13427 9807 13449
rect 9807 13427 9816 13449
rect 9764 13397 9816 13427
rect 9764 13353 9773 13385
rect 9773 13353 9807 13385
rect 9807 13353 9816 13385
rect 9764 13333 9816 13353
rect 9764 13313 9816 13321
rect 9764 13279 9773 13313
rect 9773 13279 9807 13313
rect 9807 13279 9816 13313
rect 9764 13269 9816 13279
rect 9764 13239 9816 13257
rect 9764 13205 9773 13239
rect 9773 13205 9807 13239
rect 9807 13205 9816 13239
rect 9764 13165 9816 13193
rect 9764 13141 9773 13165
rect 9773 13141 9807 13165
rect 9807 13141 9816 13165
rect 9606 12591 9658 12643
rect 9606 12527 9658 12579
rect 8277 12103 8393 12120
rect 8277 12069 8314 12103
rect 8314 12069 8348 12103
rect 8348 12069 8387 12103
rect 8387 12069 8393 12103
rect 8277 12031 8393 12069
rect 8277 12004 8314 12031
rect 8314 12004 8348 12031
rect 8348 12004 8387 12031
rect 8387 12004 8393 12031
rect 8970 12154 9086 12270
rect 7820 11723 7872 11732
rect 7820 11689 7826 11723
rect 7826 11689 7860 11723
rect 7860 11689 7872 11723
rect 7820 11680 7872 11689
rect 7886 11723 7938 11732
rect 7886 11689 7901 11723
rect 7901 11689 7935 11723
rect 7935 11689 7938 11723
rect 7886 11680 7938 11689
rect 7952 11723 8004 11732
rect 8018 11723 8070 11732
rect 8084 11723 8136 11732
rect 8150 11723 8202 11732
rect 8216 11723 8268 11732
rect 8282 11723 8334 11732
rect 7952 11689 7976 11723
rect 7976 11689 8004 11723
rect 8018 11689 8051 11723
rect 8051 11689 8070 11723
rect 8084 11689 8085 11723
rect 8085 11689 8126 11723
rect 8126 11689 8136 11723
rect 8150 11689 8160 11723
rect 8160 11689 8201 11723
rect 8201 11689 8202 11723
rect 8216 11689 8235 11723
rect 8235 11689 8268 11723
rect 8282 11689 8310 11723
rect 8310 11689 8334 11723
rect 7952 11680 8004 11689
rect 8018 11680 8070 11689
rect 8084 11680 8136 11689
rect 8150 11680 8202 11689
rect 8216 11680 8268 11689
rect 8282 11680 8334 11689
rect 8348 11723 8400 11732
rect 8348 11689 8352 11723
rect 8352 11689 8386 11723
rect 8386 11689 8400 11723
rect 8348 11680 8400 11689
rect 8414 11723 8466 11732
rect 8414 11689 8428 11723
rect 8428 11689 8462 11723
rect 8462 11689 8466 11723
rect 8414 11680 8466 11689
rect 8480 11723 8532 11732
rect 8546 11723 8598 11732
rect 8612 11723 8664 11732
rect 8677 11723 8729 11732
rect 8742 11723 8794 11732
rect 8480 11689 8504 11723
rect 8504 11689 8532 11723
rect 8546 11689 8580 11723
rect 8580 11689 8598 11723
rect 8612 11689 8614 11723
rect 8614 11689 8656 11723
rect 8656 11689 8664 11723
rect 8677 11689 8690 11723
rect 8690 11689 8729 11723
rect 8742 11689 8766 11723
rect 8766 11689 8794 11723
rect 8480 11680 8532 11689
rect 8546 11680 8598 11689
rect 8612 11680 8664 11689
rect 8677 11680 8729 11689
rect 8742 11680 8794 11689
rect 8807 11723 8859 11732
rect 8807 11689 8808 11723
rect 8808 11689 8842 11723
rect 8842 11689 8859 11723
rect 8807 11680 8859 11689
rect 8872 11723 8924 11732
rect 8872 11689 8884 11723
rect 8884 11689 8918 11723
rect 8918 11689 8924 11723
rect 8872 11680 8924 11689
rect 7417 11637 7423 11650
rect 7423 11637 7457 11650
rect 7457 11637 7469 11650
rect 7417 11577 7469 11615
rect 7417 11563 7423 11577
rect 7423 11563 7457 11577
rect 7457 11563 7469 11577
rect 7417 11504 7469 11541
rect 7417 11489 7423 11504
rect 7423 11489 7457 11504
rect 7457 11489 7469 11504
rect 7417 11431 7469 11467
rect 7417 11415 7423 11431
rect 7423 11415 7457 11431
rect 7457 11415 7469 11431
rect 6703 9797 6755 9849
rect 6783 9797 6835 9849
rect 6703 9731 6755 9783
rect 6783 9731 6835 9783
rect 7026 10959 7078 10967
rect 7026 10925 7032 10959
rect 7032 10925 7066 10959
rect 7066 10925 7078 10959
rect 7026 10915 7078 10925
rect 7026 10885 7078 10901
rect 7026 10851 7032 10885
rect 7032 10851 7066 10885
rect 7066 10851 7078 10885
rect 7026 10849 7078 10851
rect 7026 7017 7078 7043
rect 7026 6991 7032 7017
rect 7032 6991 7066 7017
rect 7066 6991 7078 7017
rect 7026 6942 7078 6977
rect 7026 6925 7032 6942
rect 7032 6925 7066 6942
rect 7066 6925 7078 6942
rect 7266 7161 7382 7341
rect 7266 6639 7382 6819
rect 7266 5458 7382 5638
rect 7266 4023 7382 4203
rect 4910 3324 4962 3376
rect 4974 3324 5026 3376
rect 5038 3324 5090 3376
rect 3340 955 3392 1007
rect 3404 955 3456 1007
rect 3500 1155 3552 1185
rect 3500 1133 3506 1155
rect 3506 1133 3540 1155
rect 3540 1133 3552 1155
rect 3500 1080 3552 1121
rect 3500 1069 3506 1080
rect 3506 1069 3540 1080
rect 3540 1069 3552 1080
rect 2309 602 2316 624
rect 2316 602 2350 624
rect 2350 602 2361 624
rect 2309 572 2361 602
rect 2309 530 2316 560
rect 2316 530 2350 560
rect 2350 530 2361 560
rect 2309 508 2361 530
rect 2565 730 2617 768
rect 2565 716 2572 730
rect 2572 716 2606 730
rect 2606 716 2617 730
rect 2565 696 2572 704
rect 2572 696 2606 704
rect 2606 696 2617 704
rect 2565 658 2617 696
rect 2565 652 2572 658
rect 2572 652 2606 658
rect 2606 652 2617 658
rect 2821 602 2828 624
rect 2828 602 2862 624
rect 2862 602 2873 624
rect 2821 572 2873 602
rect 2821 530 2828 560
rect 2828 530 2862 560
rect 2862 530 2873 560
rect 2821 508 2873 530
rect 3077 730 3129 768
rect 3077 716 3084 730
rect 3084 716 3118 730
rect 3118 716 3129 730
rect 3077 696 3084 704
rect 3084 696 3118 704
rect 3118 696 3129 704
rect 3077 658 3129 696
rect 3077 652 3084 658
rect 3084 652 3118 658
rect 3118 652 3129 658
rect 3506 829 3540 848
rect 3540 829 3558 848
rect 3506 796 3558 829
rect 3570 796 3622 848
rect 3340 652 3456 768
rect 5188 1184 5194 1185
rect 5194 1184 5228 1185
rect 5228 1184 5240 1185
rect 5188 1145 5240 1184
rect 5188 1133 5194 1145
rect 5194 1133 5228 1145
rect 5228 1133 5240 1145
rect 5188 1111 5194 1121
rect 5194 1111 5228 1121
rect 5228 1111 5240 1121
rect 5188 1069 5240 1111
rect 3264 553 3316 560
rect 3264 519 3268 553
rect 3268 519 3302 553
rect 3302 519 3316 553
rect 3264 508 3316 519
rect 3328 553 3380 560
rect 3328 519 3340 553
rect 3340 519 3374 553
rect 3374 519 3380 553
rect 3328 508 3380 519
rect 1618 428 1670 480
rect 1682 428 1734 480
rect 5369 783 5485 899
rect 5675 783 5791 899
rect 6792 3324 6844 3376
rect 6856 3324 6908 3376
rect 6920 3324 6972 3376
rect 6794 1280 6974 1588
rect 7020 1184 7032 1185
rect 7032 1184 7066 1185
rect 7066 1184 7072 1185
rect 7020 1145 7072 1184
rect 7020 1133 7032 1145
rect 7032 1133 7066 1145
rect 7066 1133 7072 1145
rect 7020 1111 7032 1121
rect 7032 1111 7066 1121
rect 7066 1111 7072 1121
rect 7020 1069 7072 1111
rect 7516 11227 7568 11279
rect 7516 11163 7568 11215
rect 7516 11099 7568 11151
rect 7516 11035 7568 11087
rect 7417 10207 7469 10243
rect 7417 10191 7423 10207
rect 7423 10191 7457 10207
rect 7457 10191 7469 10207
rect 7417 10173 7423 10179
rect 7423 10173 7457 10179
rect 7457 10173 7469 10179
rect 7417 10135 7469 10173
rect 7417 10127 7423 10135
rect 7423 10127 7457 10135
rect 7457 10127 7469 10135
rect 7417 10101 7423 10114
rect 7423 10101 7457 10114
rect 7457 10101 7469 10114
rect 7417 10063 7469 10101
rect 7417 10062 7423 10063
rect 7423 10062 7457 10063
rect 7457 10062 7469 10063
rect 7417 8119 7469 8146
rect 7417 8094 7423 8119
rect 7423 8094 7457 8119
rect 7457 8094 7469 8119
rect 7417 8047 7469 8082
rect 7417 8030 7423 8047
rect 7423 8030 7457 8047
rect 7457 8030 7469 8047
rect 7417 8013 7423 8017
rect 7423 8013 7457 8017
rect 7457 8013 7469 8017
rect 7417 7975 7469 8013
rect 7417 7965 7423 7975
rect 7423 7965 7457 7975
rect 7457 7965 7469 7975
rect 7596 9846 7648 9849
rect 7596 9812 7608 9846
rect 7608 9812 7642 9846
rect 7642 9812 7648 9846
rect 7596 9797 7648 9812
rect 7596 9772 7648 9783
rect 7596 9738 7608 9772
rect 7608 9738 7642 9772
rect 7642 9738 7648 9772
rect 7596 9731 7648 9738
rect 7698 7647 7814 7763
rect 7417 4879 7469 4880
rect 7417 4845 7423 4879
rect 7423 4845 7457 4879
rect 7457 4845 7469 4879
rect 7417 4828 7469 4845
rect 7417 4807 7469 4814
rect 7417 4773 7423 4807
rect 7423 4773 7457 4807
rect 7457 4773 7469 4807
rect 7417 4762 7469 4773
rect 7266 1576 7271 1588
rect 7271 1576 7305 1588
rect 7305 1576 7343 1588
rect 7343 1576 7377 1588
rect 7377 1576 7382 1588
rect 7266 1535 7382 1576
rect 7266 1501 7271 1535
rect 7271 1501 7305 1535
rect 7305 1501 7343 1535
rect 7343 1501 7377 1535
rect 7377 1501 7382 1535
rect 7266 1460 7382 1501
rect 7266 1426 7271 1460
rect 7271 1426 7305 1460
rect 7305 1426 7343 1460
rect 7343 1426 7377 1460
rect 7377 1426 7382 1460
rect 7266 1385 7382 1426
rect 7266 1351 7271 1385
rect 7271 1351 7305 1385
rect 7305 1351 7343 1385
rect 7343 1351 7377 1385
rect 7377 1351 7382 1385
rect 7266 1310 7382 1351
rect 7266 1280 7271 1310
rect 7271 1280 7305 1310
rect 7305 1280 7343 1310
rect 7343 1280 7377 1310
rect 7377 1280 7382 1310
rect 7596 6239 7648 6258
rect 7596 6206 7608 6239
rect 7608 6206 7642 6239
rect 7642 6206 7648 6239
rect 7596 6162 7648 6192
rect 7596 6140 7608 6162
rect 7608 6140 7642 6162
rect 7642 6140 7648 6162
rect 8664 7424 8716 7476
rect 8728 7424 8780 7476
rect 8792 7424 8844 7476
rect 8856 7424 8908 7476
rect 9890 11868 9942 11920
rect 9890 11795 9942 11847
rect 9890 11723 9942 11773
rect 9890 11721 9899 11723
rect 9899 11721 9933 11723
rect 9933 11721 9942 11723
rect 9890 11689 9899 11699
rect 9899 11689 9933 11699
rect 9933 11689 9942 11699
rect 9890 11650 9942 11689
rect 9890 11647 9899 11650
rect 9899 11647 9933 11650
rect 9933 11647 9942 11650
rect 9890 11616 9899 11625
rect 9899 11616 9933 11625
rect 9933 11616 9942 11625
rect 9890 11577 9942 11616
rect 9890 11573 9899 11577
rect 9899 11573 9933 11577
rect 9933 11573 9942 11577
rect 9890 11543 9899 11551
rect 9899 11543 9933 11551
rect 9933 11543 9942 11551
rect 9890 11504 9942 11543
rect 9890 11499 9899 11504
rect 9899 11499 9933 11504
rect 9933 11499 9942 11504
rect 9712 9846 9764 9849
rect 9712 9812 9718 9846
rect 9718 9812 9752 9846
rect 9752 9812 9764 9846
rect 9712 9797 9764 9812
rect 9712 9772 9764 9783
rect 9712 9738 9718 9772
rect 9718 9738 9752 9772
rect 9752 9738 9764 9772
rect 9712 9731 9764 9738
rect 9804 10229 9899 10243
rect 9899 10229 9933 10243
rect 9933 10229 10048 10243
rect 9804 10190 10048 10229
rect 9804 10156 9899 10190
rect 9899 10156 9933 10190
rect 9933 10156 10048 10190
rect 9804 10127 10048 10156
rect 9804 10062 9856 10114
rect 9868 10083 9899 10114
rect 9899 10083 9920 10114
rect 9932 10083 9933 10114
rect 9933 10083 9984 10114
rect 9868 10062 9920 10083
rect 9932 10062 9984 10083
rect 9996 10062 10048 10114
rect 10078 9498 10194 9614
rect 10078 9433 10130 9485
rect 10142 9433 10194 9485
rect 10078 9368 10130 9420
rect 10142 9368 10194 9420
rect 10078 8488 10130 8540
rect 10142 8488 10194 8540
rect 10078 8421 10130 8473
rect 10142 8421 10194 8473
rect 10078 8354 10130 8406
rect 10142 8354 10194 8406
rect 10078 8286 10130 8338
rect 10142 8286 10194 8338
rect 9804 8112 9899 8146
rect 9899 8112 9933 8146
rect 9933 8112 10048 8146
rect 9804 8073 10048 8112
rect 9804 8039 9899 8073
rect 9899 8039 9933 8073
rect 9933 8039 10048 8073
rect 9804 8030 10048 8039
rect 9804 7965 9856 8017
rect 9868 8000 9920 8017
rect 9932 8000 9984 8017
rect 9868 7966 9899 8000
rect 9899 7966 9920 8000
rect 9932 7966 9933 8000
rect 9933 7966 9984 8000
rect 9868 7965 9920 7966
rect 9932 7965 9984 7966
rect 9996 7965 10048 8017
rect 10311 8040 10363 8049
rect 10311 8006 10317 8040
rect 10317 8006 10351 8040
rect 10351 8006 10363 8040
rect 10311 7997 10363 8006
rect 10376 8040 10428 8049
rect 10376 8006 10389 8040
rect 10389 8006 10423 8040
rect 10423 8006 10428 8040
rect 10376 7997 10428 8006
rect 10441 8040 10493 8049
rect 10506 8040 10558 8049
rect 10571 8040 10623 8049
rect 10636 8040 10688 8049
rect 10701 8040 10753 8049
rect 10766 8040 10818 8049
rect 10831 8040 10883 8049
rect 10896 8040 10948 8049
rect 10441 8006 10461 8040
rect 10461 8006 10493 8040
rect 10506 8006 10533 8040
rect 10533 8006 10558 8040
rect 10571 8006 10605 8040
rect 10605 8006 10623 8040
rect 10636 8006 10639 8040
rect 10639 8006 10677 8040
rect 10677 8006 10688 8040
rect 10701 8006 10711 8040
rect 10711 8006 10749 8040
rect 10749 8006 10753 8040
rect 10766 8006 10783 8040
rect 10783 8006 10818 8040
rect 10831 8006 10855 8040
rect 10855 8006 10883 8040
rect 10896 8006 10927 8040
rect 10927 8006 10948 8040
rect 10441 7997 10493 8006
rect 10506 7997 10558 8006
rect 10571 7997 10623 8006
rect 10636 7997 10688 8006
rect 10701 7997 10753 8006
rect 10766 7997 10818 8006
rect 10831 7997 10883 8006
rect 10896 7997 10948 8006
rect 10961 8040 11013 8049
rect 10961 8006 10965 8040
rect 10965 8006 10999 8040
rect 10999 8006 11013 8040
rect 10961 7997 11013 8006
rect 11026 8040 11078 8049
rect 11026 8006 11037 8040
rect 11037 8006 11071 8040
rect 11071 8006 11078 8040
rect 11026 7997 11078 8006
rect 11091 8040 11143 8049
rect 11091 8006 11109 8040
rect 11109 8006 11143 8040
rect 11091 7997 11143 8006
rect 11156 8040 11208 8049
rect 11221 8040 11273 8049
rect 11286 8040 11338 8049
rect 11350 8040 11402 8049
rect 11414 8040 11466 8049
rect 11478 8040 11530 8049
rect 11542 8040 11594 8049
rect 11156 8006 11181 8040
rect 11181 8006 11208 8040
rect 11221 8006 11253 8040
rect 11253 8006 11273 8040
rect 11286 8006 11287 8040
rect 11287 8006 11325 8040
rect 11325 8006 11338 8040
rect 11350 8006 11359 8040
rect 11359 8006 11397 8040
rect 11397 8006 11402 8040
rect 11414 8006 11431 8040
rect 11431 8006 11466 8040
rect 11478 8006 11503 8040
rect 11503 8006 11530 8040
rect 11542 8006 11575 8040
rect 11575 8006 11594 8040
rect 11156 7997 11208 8006
rect 11221 7997 11273 8006
rect 11286 7997 11338 8006
rect 11350 7997 11402 8006
rect 11414 7997 11466 8006
rect 11478 7997 11530 8006
rect 11542 7997 11594 8006
rect 11606 8040 11658 8049
rect 11606 8006 11613 8040
rect 11613 8006 11647 8040
rect 11647 8006 11658 8040
rect 11606 7997 11658 8006
rect 11670 8040 11722 8049
rect 11670 8006 11685 8040
rect 11685 8006 11719 8040
rect 11719 8006 11722 8040
rect 11670 7997 11722 8006
rect 11734 8040 11786 8049
rect 11798 8040 11850 8049
rect 11862 8040 11914 8049
rect 11926 8040 11978 8049
rect 11990 8040 12042 8049
rect 12054 8040 12106 8049
rect 12118 8040 12170 8049
rect 11734 8006 11757 8040
rect 11757 8006 11786 8040
rect 11798 8006 11829 8040
rect 11829 8006 11850 8040
rect 11862 8006 11863 8040
rect 11863 8006 11901 8040
rect 11901 8006 11914 8040
rect 11926 8006 11935 8040
rect 11935 8006 11973 8040
rect 11973 8006 11978 8040
rect 11990 8006 12007 8040
rect 12007 8006 12042 8040
rect 12054 8006 12079 8040
rect 12079 8006 12106 8040
rect 12118 8006 12151 8040
rect 12151 8006 12170 8040
rect 11734 7997 11786 8006
rect 11798 7997 11850 8006
rect 11862 7997 11914 8006
rect 11926 7997 11978 8006
rect 11990 7997 12042 8006
rect 12054 7997 12106 8006
rect 12118 7997 12170 8006
rect 12182 8040 12234 8049
rect 12182 8006 12189 8040
rect 12189 8006 12223 8040
rect 12223 8006 12234 8040
rect 12182 7997 12234 8006
rect 12246 8040 12298 8049
rect 12246 8006 12261 8040
rect 12261 8006 12295 8040
rect 12295 8006 12298 8040
rect 12246 7997 12298 8006
rect 12310 8040 12362 8049
rect 12374 8040 12426 8049
rect 12438 8040 12490 8049
rect 12502 8040 12554 8049
rect 12566 8040 12618 8049
rect 12630 8040 12682 8049
rect 12310 8006 12333 8040
rect 12333 8006 12362 8040
rect 12374 8006 12405 8040
rect 12405 8006 12426 8040
rect 12438 8006 12439 8040
rect 12439 8006 12478 8040
rect 12478 8006 12490 8040
rect 12502 8006 12512 8040
rect 12512 8006 12551 8040
rect 12551 8006 12554 8040
rect 12566 8006 12585 8040
rect 12585 8006 12618 8040
rect 12630 8006 12658 8040
rect 12658 8006 12682 8040
rect 12310 7997 12362 8006
rect 12374 7997 12426 8006
rect 12438 7997 12490 8006
rect 12502 7997 12554 8006
rect 12566 7997 12618 8006
rect 12630 7997 12682 8006
rect 12694 8040 12746 8049
rect 12694 8006 12697 8040
rect 12697 8006 12731 8040
rect 12731 8006 12746 8040
rect 12694 7997 12746 8006
rect 12758 8040 12810 8049
rect 12758 8006 12770 8040
rect 12770 8006 12804 8040
rect 12804 8006 12810 8040
rect 12758 7997 12810 8006
rect 7692 4236 7744 4288
rect 7756 4236 7808 4288
rect 7452 1069 7568 1185
rect 7596 1155 7648 1185
rect 7596 1133 7608 1155
rect 7608 1133 7642 1155
rect 7642 1133 7648 1155
rect 7596 1080 7648 1121
rect 7596 1069 7608 1080
rect 7608 1069 7642 1080
rect 7642 1069 7648 1080
rect 10193 7339 10245 7341
rect 10193 7305 10205 7339
rect 10205 7305 10239 7339
rect 10239 7305 10245 7339
rect 10193 7289 10245 7305
rect 10193 7267 10245 7277
rect 10193 7233 10205 7267
rect 10205 7233 10239 7267
rect 10239 7233 10245 7267
rect 10193 7225 10245 7233
rect 10193 7195 10245 7213
rect 10193 7161 10205 7195
rect 10205 7161 10239 7195
rect 10239 7161 10245 7195
rect 10193 6801 10205 6819
rect 10205 6801 10239 6819
rect 10239 6801 10245 6819
rect 10193 6767 10245 6801
rect 10193 6729 10205 6755
rect 10205 6729 10239 6755
rect 10239 6729 10245 6755
rect 10193 6703 10245 6729
rect 10193 6657 10205 6691
rect 10205 6657 10239 6691
rect 10239 6657 10245 6691
rect 10193 6639 10245 6657
rect 9712 6239 9764 6258
rect 9712 6206 9718 6239
rect 9718 6206 9752 6239
rect 9752 6206 9764 6239
rect 9712 6162 9764 6192
rect 9712 6140 9718 6162
rect 9718 6140 9752 6162
rect 9752 6140 9764 6162
rect 10047 6422 10099 6474
rect 10047 6356 10099 6408
rect 9817 4828 9869 4880
rect 9881 4868 9899 4880
rect 9899 4868 9933 4880
rect 9881 4830 9933 4868
rect 9881 4828 9899 4830
rect 9899 4828 9933 4830
rect 9817 4762 9869 4814
rect 9881 4796 9899 4814
rect 9899 4796 9933 4814
rect 9881 4762 9933 4796
rect 9967 6206 10019 6258
rect 9967 6140 10019 6192
rect 9967 3970 10019 4022
rect 10193 5611 10245 5638
rect 10193 5586 10205 5611
rect 10205 5586 10239 5611
rect 10239 5586 10245 5611
rect 10193 5539 10245 5574
rect 10193 5522 10205 5539
rect 10205 5522 10239 5539
rect 10239 5522 10245 5539
rect 10193 5505 10205 5510
rect 10205 5505 10239 5510
rect 10239 5505 10245 5510
rect 10193 5467 10245 5505
rect 10193 5458 10205 5467
rect 10205 5458 10239 5467
rect 10239 5458 10245 5467
rect 10047 3994 10099 4046
rect 10111 3994 10163 4046
rect 9967 3904 10019 3956
rect 8151 1536 8203 1588
rect 8217 1536 8269 1588
rect 8283 1536 8335 1588
rect 8349 1536 8401 1588
rect 8415 1536 8467 1588
rect 8481 1536 8533 1588
rect 8546 1536 8598 1588
rect 8611 1536 8663 1588
rect 8676 1536 8728 1588
rect 8741 1536 8793 1588
rect 8151 1472 8203 1524
rect 8217 1472 8269 1524
rect 8283 1472 8335 1524
rect 8349 1472 8401 1524
rect 8415 1472 8467 1524
rect 8481 1472 8533 1524
rect 8546 1472 8598 1524
rect 8611 1472 8663 1524
rect 8676 1472 8728 1524
rect 8741 1472 8793 1524
rect 8151 1408 8203 1460
rect 8217 1408 8269 1460
rect 8283 1408 8335 1460
rect 8349 1408 8401 1460
rect 8415 1408 8467 1460
rect 8481 1408 8533 1460
rect 8546 1408 8598 1460
rect 8611 1408 8663 1460
rect 8676 1408 8728 1460
rect 8741 1408 8793 1460
rect 8151 1344 8203 1396
rect 8217 1344 8269 1396
rect 8283 1344 8335 1396
rect 8349 1344 8401 1396
rect 8415 1344 8467 1396
rect 8481 1344 8533 1396
rect 8546 1344 8598 1396
rect 8611 1344 8663 1396
rect 8676 1344 8728 1396
rect 8741 1344 8793 1396
rect 8151 1280 8203 1332
rect 8217 1280 8269 1332
rect 8283 1280 8335 1332
rect 8349 1280 8401 1332
rect 8415 1280 8467 1332
rect 8481 1280 8533 1332
rect 8546 1280 8598 1332
rect 8611 1280 8663 1332
rect 8676 1280 8728 1332
rect 8741 1280 8793 1332
rect 8023 1133 8075 1185
rect 8023 1069 8075 1121
rect 5186 428 5238 480
rect 5250 428 5302 480
rect 5763 428 5815 480
rect 5827 428 5879 480
rect 7026 547 7078 550
rect 7026 513 7032 547
rect 7032 513 7066 547
rect 7066 513 7078 547
rect 7026 498 7078 513
rect 7026 434 7078 486
rect 7692 652 7808 768
rect 8019 730 8071 768
rect 8019 716 8030 730
rect 8030 716 8064 730
rect 8064 716 8071 730
rect 8019 696 8030 704
rect 8030 696 8064 704
rect 8064 696 8071 704
rect 8019 658 8071 696
rect 8019 652 8030 658
rect 8030 652 8064 658
rect 8064 652 8071 658
rect 7762 578 7814 585
rect 7762 544 7774 578
rect 7774 544 7808 578
rect 7808 544 7814 578
rect 7762 533 7814 544
rect 7826 578 7878 585
rect 7826 544 7846 578
rect 7846 544 7878 578
rect 8275 602 8286 624
rect 8286 602 8320 624
rect 8320 602 8327 624
rect 8275 572 8327 602
rect 7826 533 7878 544
rect 8275 530 8286 560
rect 8286 530 8320 560
rect 8320 530 8327 560
rect 8275 508 8327 530
rect 8531 730 8583 768
rect 8531 716 8542 730
rect 8542 716 8576 730
rect 8576 716 8583 730
rect 8531 696 8542 704
rect 8542 696 8576 704
rect 8576 696 8583 704
rect 8531 658 8583 696
rect 8531 652 8542 658
rect 8542 652 8576 658
rect 8576 652 8583 658
rect 9163 1133 9215 1185
rect 9163 1069 9215 1121
rect 9712 1155 9764 1185
rect 9712 1133 9718 1155
rect 9718 1133 9752 1155
rect 9752 1133 9764 1155
rect 9712 1080 9764 1121
rect 9712 1069 9718 1080
rect 9718 1069 9752 1080
rect 9752 1069 9764 1080
rect 8787 602 8798 624
rect 8798 602 8832 624
rect 8832 602 8839 624
rect 8787 572 8839 602
rect 8787 530 8798 560
rect 8798 530 8832 560
rect 8832 530 8839 560
rect 8787 508 8839 530
rect 9199 602 9210 624
rect 9210 602 9244 624
rect 9244 602 9251 624
rect 9199 572 9251 602
rect 9199 530 9210 560
rect 9210 530 9244 560
rect 9244 530 9251 560
rect 9199 508 9251 530
rect 10193 2049 10205 2060
rect 10205 2049 10239 2060
rect 10239 2049 10245 2060
rect 10193 2011 10245 2049
rect 10193 2008 10205 2011
rect 10205 2008 10239 2011
rect 10239 2008 10245 2011
rect 10193 1977 10205 1996
rect 10205 1977 10239 1996
rect 10239 1977 10245 1996
rect 10193 1944 10245 1977
rect 10193 1905 10205 1932
rect 10205 1905 10239 1932
rect 10239 1905 10245 1932
rect 10193 1880 10245 1905
rect 10193 1867 10245 1868
rect 10193 1833 10205 1867
rect 10205 1833 10239 1867
rect 10239 1833 10245 1867
rect 10193 1816 10245 1833
rect 10193 1795 10245 1804
rect 10193 1761 10205 1795
rect 10205 1761 10239 1795
rect 10239 1761 10245 1795
rect 10193 1752 10245 1761
rect 12891 6639 13007 6819
rect 12891 5586 12943 5638
rect 12955 5586 13007 5638
rect 12891 5512 12943 5564
rect 12955 5512 13007 5564
rect 12891 5438 12943 5490
rect 12955 5438 13007 5490
rect 12891 5364 12943 5416
rect 12955 5364 13007 5416
rect 12891 5289 12943 5341
rect 12955 5289 13007 5341
rect 12891 5214 12943 5266
rect 12955 5214 13007 5266
rect 12891 5139 12943 5191
rect 12955 5139 13007 5191
rect 12891 2014 12943 2066
rect 12955 2014 13007 2066
rect 12891 1949 12943 2001
rect 12955 1949 13007 2001
rect 12891 1884 12943 1936
rect 12955 1884 13007 1936
rect 12891 1818 12943 1870
rect 12955 1818 13007 1870
rect 12891 1752 12943 1804
rect 12955 1752 13007 1804
rect 13063 4856 13115 4880
rect 13063 4828 13069 4856
rect 13069 4828 13103 4856
rect 13103 4828 13115 4856
rect 13063 4784 13115 4814
rect 13063 4762 13069 4784
rect 13069 4762 13103 4784
rect 13103 4762 13115 4784
<< metal2 >>
rect 1202 13989 11178 14527
rect 1342 13881 1348 13933
rect 1400 13881 1413 13933
rect 1465 13881 5262 13933
rect 5314 13881 5326 13933
rect 5378 13881 5390 13933
rect 5442 13881 5454 13933
rect 5506 13881 5518 13933
rect 5570 13881 5582 13933
rect 5634 13881 5646 13933
rect 5698 13881 5710 13933
rect 5762 13881 5774 13933
rect 5826 13881 9516 13933
rect 9568 13881 9608 13933
rect 9660 13881 9700 13933
rect 9752 13881 9758 13933
rect 1604 13835 10127 13841
rect 1656 13783 5215 13835
rect 5267 13783 5527 13835
rect 5579 13783 5839 13835
rect 5891 13783 6366 13835
rect 6418 13783 6442 13835
rect 6494 13783 6516 13835
rect 6568 13783 7204 13835
rect 7256 13783 7279 13835
rect 7331 13783 7354 13835
rect 7406 13783 8053 13835
rect 8105 13783 8130 13835
rect 8182 13783 8207 13835
rect 8259 13783 8284 13835
rect 8336 13783 8361 13835
rect 8413 13783 8441 13835
rect 8493 13783 8518 13835
rect 8570 13783 8595 13835
rect 8647 13783 8672 13835
rect 8724 13783 8749 13835
rect 8801 13783 8826 13835
rect 8878 13783 8900 13835
rect 8952 13783 8975 13835
rect 9027 13783 9050 13835
rect 9102 13783 10127 13835
rect 1604 13767 10127 13783
rect 1656 13715 5215 13767
rect 5267 13715 5527 13767
rect 5579 13715 5839 13767
rect 5891 13715 6366 13767
rect 6418 13715 6442 13767
rect 6494 13715 6516 13767
rect 6568 13715 7204 13767
rect 7256 13715 7279 13767
rect 7331 13715 7354 13767
rect 7406 13715 8053 13767
rect 8105 13715 8130 13767
rect 8182 13715 8207 13767
rect 8259 13715 8284 13767
rect 8336 13715 8361 13767
rect 8413 13715 8441 13767
rect 8493 13715 8518 13767
rect 8570 13715 8595 13767
rect 8647 13715 8672 13767
rect 8724 13715 8749 13767
rect 8801 13715 8826 13767
rect 8878 13715 8900 13767
rect 8952 13715 8975 13767
rect 9027 13715 9050 13767
rect 9102 13715 10127 13767
rect 1604 13699 10127 13715
rect 1656 13647 5215 13699
rect 5267 13647 5527 13699
rect 5579 13647 5839 13699
rect 5891 13647 6366 13699
rect 6418 13647 6442 13699
rect 6494 13647 6516 13699
rect 6568 13647 7204 13699
rect 7256 13647 7279 13699
rect 7331 13647 7354 13699
rect 7406 13647 8053 13699
rect 8105 13647 8130 13699
rect 8182 13647 8207 13699
rect 8259 13647 8284 13699
rect 8336 13647 8361 13699
rect 8413 13647 8441 13699
rect 8493 13647 8518 13699
rect 8570 13647 8595 13699
rect 8647 13647 8672 13699
rect 8724 13647 8749 13699
rect 8801 13647 8826 13699
rect 8878 13647 8900 13699
rect 8952 13647 8975 13699
rect 9027 13647 9050 13699
rect 9102 13647 10127 13699
rect 1604 13631 10127 13647
rect 1656 13579 5215 13631
rect 5267 13579 5527 13631
rect 5579 13579 5839 13631
rect 5891 13579 6366 13631
rect 6418 13579 6442 13631
rect 6494 13579 6516 13631
rect 6568 13579 7204 13631
rect 7256 13579 7279 13631
rect 7331 13579 7354 13631
rect 7406 13579 8053 13631
rect 8105 13579 8130 13631
rect 8182 13579 8207 13631
rect 8259 13579 8284 13631
rect 8336 13579 8361 13631
rect 8413 13579 8441 13631
rect 8493 13579 8518 13631
rect 8570 13579 8595 13631
rect 8647 13579 8672 13631
rect 8724 13579 8749 13631
rect 8801 13579 8826 13631
rect 8878 13579 8900 13631
rect 8952 13579 8975 13631
rect 9027 13579 9050 13631
rect 9102 13579 10127 13631
rect 1604 13563 10127 13579
rect 1656 13511 5215 13563
rect 5267 13511 5527 13563
rect 5579 13511 5839 13563
rect 5891 13511 6366 13563
rect 6418 13511 6442 13563
rect 6494 13511 6516 13563
rect 6568 13511 7204 13563
rect 7256 13511 7279 13563
rect 7331 13511 7354 13563
rect 7406 13511 8053 13563
rect 8105 13511 8130 13563
rect 8182 13511 8207 13563
rect 8259 13511 8284 13563
rect 8336 13511 8361 13563
rect 8413 13511 8441 13563
rect 8493 13511 8518 13563
rect 8570 13511 8595 13563
rect 8647 13511 8672 13563
rect 8724 13511 8749 13563
rect 8801 13511 8826 13563
rect 8878 13511 8900 13563
rect 8952 13511 8975 13563
rect 9027 13511 9050 13563
rect 9102 13511 10127 13563
rect 1604 13505 10127 13511
rect 7621 13449 9816 13455
rect 7621 13397 9452 13449
rect 9504 13397 9764 13449
rect 7621 13385 9816 13397
rect 1983 13361 7423 13367
rect 1983 13309 1996 13361
rect 2048 13309 2073 13361
rect 2125 13309 2150 13361
rect 2202 13309 2227 13361
rect 2279 13309 2304 13361
rect 2356 13309 2384 13361
rect 2436 13309 2461 13361
rect 2513 13309 2538 13361
rect 2590 13309 2615 13361
rect 2667 13309 2692 13361
rect 2744 13309 2769 13361
rect 2821 13309 2843 13361
rect 2895 13309 2918 13361
rect 2970 13309 2993 13361
rect 3045 13309 3688 13361
rect 3740 13309 3762 13361
rect 3814 13309 3838 13361
rect 3890 13309 4526 13361
rect 4578 13309 4601 13361
rect 4653 13309 4676 13361
rect 4728 13309 5371 13361
rect 5423 13309 5683 13361
rect 5735 13309 7423 13361
rect 1983 13293 7423 13309
rect 1983 13241 1996 13293
rect 2048 13241 2073 13293
rect 2125 13241 2150 13293
rect 2202 13241 2227 13293
rect 2279 13241 2304 13293
rect 2356 13241 2384 13293
rect 2436 13241 2461 13293
rect 2513 13241 2538 13293
rect 2590 13241 2615 13293
rect 2667 13241 2692 13293
rect 2744 13241 2769 13293
rect 2821 13241 2843 13293
rect 2895 13241 2918 13293
rect 2970 13241 2993 13293
rect 3045 13241 3688 13293
rect 3740 13241 3762 13293
rect 3814 13241 3838 13293
rect 3890 13241 4526 13293
rect 4578 13241 4601 13293
rect 4653 13241 4676 13293
rect 4728 13241 5371 13293
rect 5423 13241 5683 13293
rect 5735 13241 7423 13293
rect 1983 13225 7423 13241
rect 1983 13173 1996 13225
rect 2048 13173 2073 13225
rect 2125 13173 2150 13225
rect 2202 13173 2227 13225
rect 2279 13173 2304 13225
rect 2356 13173 2384 13225
rect 2436 13173 2461 13225
rect 2513 13173 2538 13225
rect 2590 13173 2615 13225
rect 2667 13173 2692 13225
rect 2744 13173 2769 13225
rect 2821 13173 2843 13225
rect 2895 13173 2918 13225
rect 2970 13173 2993 13225
rect 3045 13173 3688 13225
rect 3740 13173 3762 13225
rect 3814 13173 3838 13225
rect 3890 13173 4526 13225
rect 4578 13173 4601 13225
rect 4653 13173 4676 13225
rect 4728 13173 5371 13225
rect 5423 13173 5683 13225
rect 5735 13173 7423 13225
rect 1983 13157 7423 13173
rect 1983 13105 1996 13157
rect 2048 13105 2073 13157
rect 2125 13105 2150 13157
rect 2202 13105 2227 13157
rect 2279 13105 2304 13157
rect 2356 13105 2384 13157
rect 2436 13105 2461 13157
rect 2513 13105 2538 13157
rect 2590 13105 2615 13157
rect 2667 13105 2692 13157
rect 2744 13105 2769 13157
rect 2821 13105 2843 13157
rect 2895 13105 2918 13157
rect 2970 13105 2993 13157
rect 3045 13105 3688 13157
rect 3740 13105 3762 13157
rect 3814 13105 3838 13157
rect 3890 13105 4526 13157
rect 4578 13105 4601 13157
rect 4653 13105 4676 13157
rect 4728 13105 5371 13157
rect 5423 13105 5683 13157
rect 5735 13105 7423 13157
rect 7621 13333 9452 13385
rect 9504 13333 9764 13385
rect 7621 13321 9816 13333
rect 7621 13269 9452 13321
rect 9504 13269 9764 13321
rect 7621 13257 9816 13269
rect 7621 13205 9452 13257
rect 9504 13205 9764 13257
rect 7621 13193 9816 13205
rect 7621 13141 9452 13193
rect 9504 13141 9764 13193
rect 7621 13135 9816 13141
rect 1983 13089 7423 13105
rect 1983 13037 1996 13089
rect 2048 13037 2073 13089
rect 2125 13037 2150 13089
rect 2202 13037 2227 13089
rect 2279 13037 2304 13089
rect 2356 13037 2384 13089
rect 2436 13037 2461 13089
rect 2513 13037 2538 13089
rect 2590 13037 2615 13089
rect 2667 13037 2692 13089
rect 2744 13037 2769 13089
rect 2821 13037 2843 13089
rect 2895 13037 2918 13089
rect 2970 13037 2993 13089
rect 3045 13037 3688 13089
rect 3740 13037 3762 13089
rect 3814 13037 3838 13089
rect 3890 13037 4526 13089
rect 4578 13037 4601 13089
rect 4653 13037 4676 13089
rect 4728 13037 5371 13089
rect 5423 13037 5683 13089
rect 5735 13037 7423 13089
rect 1983 13031 7423 13037
rect 7895 13073 7947 13079
tri 7888 13021 7895 13028 se
tri 7876 13009 7888 13021 se
rect 7888 13009 7947 13021
tri 7870 13003 7876 13009 se
rect 7876 13003 7895 13009
rect 3135 12997 3975 13003
rect 3187 12951 3975 12997
rect 4027 12951 4039 13003
rect 4091 12951 4103 13003
rect 4155 12951 4813 13003
rect 4865 12951 4877 13003
rect 4929 12951 4941 13003
rect 4993 12951 4999 13003
rect 6647 12951 6653 13003
rect 6705 12951 6717 13003
rect 6769 12951 6781 13003
rect 6833 12951 6930 13003
rect 6982 12951 6994 13003
rect 7046 12951 7058 13003
rect 7110 12957 7895 13003
rect 7110 12951 7947 12957
rect 3135 12933 3187 12945
tri 3187 12926 3212 12951 nw
rect 3135 12875 3187 12881
rect 1202 12847 3087 12872
tri 3087 12847 3112 12872 sw
tri 3210 12847 3235 12872 se
rect 3235 12847 11178 12872
rect 1202 12820 11178 12847
tri 3062 12795 3087 12820 ne
rect 3087 12795 3235 12820
tri 3235 12795 3260 12820 nw
tri 12181 12649 12296 12764 se
rect 12296 12649 13266 12764
rect 3477 12643 9658 12649
rect 3529 12591 5447 12643
rect 5499 12591 9606 12643
rect 3477 12579 9658 12591
rect 3529 12527 5447 12579
rect 5499 12527 9606 12579
rect 3477 12521 9658 12527
tri 12053 12521 12181 12649 se
rect 12181 12542 13266 12649
rect 12181 12521 12296 12542
tri 11999 12467 12053 12521 se
rect 12053 12467 12296 12521
rect 1441 12415 1447 12467
rect 1499 12415 1511 12467
rect 1563 12415 5495 12467
rect 5547 12415 5559 12467
rect 5611 12415 5617 12467
tri 11982 12450 11999 12467 se
rect 11999 12450 12296 12467
tri 12296 12450 12388 12542 nw
tri 12516 12450 12552 12486 se
rect 12552 12450 13266 12486
tri 11947 12415 11982 12450 se
rect 11982 12415 12076 12450
tri 11808 12276 11947 12415 se
rect 11947 12276 12076 12415
rect 2048 12270 4527 12276
rect 2164 12218 4475 12270
rect 2164 12206 4527 12218
rect 2164 12154 4475 12206
rect 2048 12148 4527 12154
rect 6315 12270 9086 12276
rect 6367 12218 8970 12270
rect 6315 12206 8970 12218
rect 6367 12154 8970 12206
tri 11736 12204 11808 12276 se
rect 11808 12230 12076 12276
tri 12076 12230 12296 12450 nw
tri 12378 12312 12516 12450 se
rect 12516 12356 13266 12450
rect 12516 12312 12552 12356
tri 12552 12312 12596 12356 nw
tri 12296 12230 12378 12312 se
rect 12378 12300 12540 12312
tri 12540 12300 12552 12312 nw
rect 12378 12260 12500 12300
tri 12500 12260 12540 12300 nw
tri 12540 12260 12580 12300 se
rect 12580 12260 13266 12300
rect 12378 12230 12460 12260
rect 11808 12204 12050 12230
tri 12050 12204 12076 12230 nw
tri 12270 12204 12296 12230 se
rect 12296 12220 12460 12230
tri 12460 12220 12500 12260 nw
tri 12500 12220 12540 12260 se
rect 12540 12220 13266 12260
rect 12296 12206 12446 12220
tri 12446 12206 12460 12220 nw
tri 12486 12206 12500 12220 se
rect 12500 12206 13266 12220
rect 12296 12204 12406 12206
rect 6315 12148 9086 12154
tri 9142 12148 9198 12204 se
rect 9198 12148 11830 12204
tri 9114 12120 9142 12148 se
rect 9142 12120 11830 12148
rect 1202 12004 1758 12120
rect 1874 12004 2720 12120
rect 2836 12004 3767 12120
rect 3883 12004 5478 12120
rect 5594 12004 7263 12120
rect 7379 12004 8277 12120
rect 8393 12004 11830 12120
rect 1202 11984 11830 12004
tri 11830 11984 12050 12204 nw
tri 12204 12138 12270 12204 se
rect 12270 12166 12406 12204
tri 12406 12166 12446 12206 nw
tri 12446 12166 12486 12206 se
rect 12486 12170 13266 12206
rect 12486 12166 12580 12170
rect 12270 12138 12378 12166
tri 12378 12138 12406 12166 nw
tri 12418 12138 12446 12166 se
rect 12446 12138 12580 12166
tri 12050 11984 12204 12138 se
rect 12204 12126 12366 12138
tri 12366 12126 12378 12138 nw
tri 12406 12126 12418 12138 se
rect 12418 12126 12580 12138
tri 12580 12126 12624 12170 nw
rect 12204 12086 12326 12126
tri 12326 12086 12366 12126 nw
tri 12366 12086 12406 12126 se
rect 12204 12046 12286 12086
tri 12286 12046 12326 12086 nw
tri 12326 12046 12366 12086 se
rect 12366 12046 12406 12086
rect 12204 12032 12272 12046
tri 12272 12032 12286 12046 nw
tri 12312 12032 12326 12046 se
rect 12326 12032 12406 12046
rect 12204 11992 12232 12032
tri 12232 11992 12272 12032 nw
tri 12272 11992 12312 12032 se
rect 12312 11992 12406 12032
rect 1202 11982 11828 11984
tri 11828 11982 11830 11984 nw
tri 12048 11982 12050 11984 se
rect 12050 11982 12204 11984
rect 1202 11920 9228 11982
tri 9228 11920 9290 11982 nw
tri 12030 11964 12048 11982 se
rect 12048 11964 12204 11982
tri 12204 11964 12232 11992 nw
tri 12244 11964 12272 11992 se
rect 12272 11964 12406 11992
tri 11992 11926 12030 11964 se
rect 12030 11952 12192 11964
tri 12192 11952 12204 11964 nw
tri 12232 11952 12244 11964 se
rect 12244 11952 12406 11964
tri 12406 11952 12580 12126 nw
rect 12030 11926 12152 11952
tri 9743 11920 9749 11926 se
rect 9749 11920 11505 11926
rect 1202 11898 9206 11920
tri 9206 11898 9228 11920 nw
tri 9721 11898 9743 11920 se
rect 9743 11898 9890 11920
tri 9691 11868 9721 11898 se
rect 9721 11868 9890 11898
rect 9942 11868 11505 11920
tri 9670 11847 9691 11868 se
rect 9691 11847 11505 11868
tri 9665 11842 9670 11847 se
rect 9670 11842 9890 11847
rect 1176 11836 9890 11842
rect 1228 11784 3681 11836
rect 3733 11784 7417 11836
rect 7469 11795 9890 11836
rect 9942 11795 11505 11847
rect 7469 11784 11505 11795
tri 11856 11790 11992 11926 se
rect 11992 11912 12152 11926
tri 12152 11912 12192 11952 nw
tri 12192 11912 12232 11952 se
rect 11992 11872 12112 11912
tri 12112 11872 12152 11912 nw
tri 12152 11872 12192 11912 se
rect 12192 11872 12232 11912
rect 11992 11858 12098 11872
tri 12098 11858 12112 11872 nw
tri 12138 11858 12152 11872 se
rect 12152 11858 12232 11872
rect 11992 11818 12058 11858
tri 12058 11818 12098 11858 nw
tri 12098 11818 12138 11858 se
rect 12138 11818 12232 11858
rect 11992 11790 12030 11818
tri 12030 11790 12058 11818 nw
tri 12070 11790 12098 11818 se
rect 12098 11790 12232 11818
rect 1176 11773 11505 11784
rect 1176 11763 9890 11773
rect 1228 11762 7417 11763
rect 1228 11732 3681 11762
rect 1228 11711 1624 11732
rect 1176 11690 1624 11711
rect 1228 11680 1624 11690
rect 1676 11680 1689 11732
rect 1741 11680 1754 11732
rect 1806 11680 1819 11732
rect 1871 11680 1884 11732
rect 1936 11680 1950 11732
rect 2002 11680 2224 11732
rect 2276 11680 2292 11732
rect 2344 11680 2360 11732
rect 2412 11680 2428 11732
rect 2480 11680 2496 11732
rect 2548 11680 2564 11732
rect 2616 11680 2632 11732
rect 2684 11680 2700 11732
rect 2752 11680 2768 11732
rect 2820 11680 2836 11732
rect 2888 11680 2904 11732
rect 2956 11680 2972 11732
rect 3024 11680 3040 11732
rect 3092 11680 3108 11732
rect 3160 11680 3175 11732
rect 3227 11680 3242 11732
rect 3294 11680 3309 11732
rect 3361 11710 3681 11732
rect 3733 11732 7417 11762
rect 3733 11710 4493 11732
rect 3361 11688 4493 11710
rect 3361 11680 3681 11688
rect 1228 11638 3681 11680
rect 1176 11636 3681 11638
rect 3733 11680 4493 11688
rect 4545 11680 4565 11732
rect 4617 11680 4637 11732
rect 4689 11680 4709 11732
rect 4761 11680 5055 11732
rect 5107 11680 5122 11732
rect 5174 11680 5189 11732
rect 5241 11680 5256 11732
rect 5308 11680 5323 11732
rect 5375 11680 5390 11732
rect 5442 11680 5457 11732
rect 5509 11680 5524 11732
rect 5576 11680 5591 11732
rect 5643 11680 5657 11732
rect 5709 11680 5723 11732
rect 5775 11680 5789 11732
rect 5841 11680 5855 11732
rect 5907 11680 5921 11732
rect 5973 11680 5987 11732
rect 6039 11680 6333 11732
rect 6385 11680 6405 11732
rect 6457 11680 6477 11732
rect 6529 11680 6549 11732
rect 6601 11711 7417 11732
rect 7469 11732 9890 11763
rect 7469 11711 7820 11732
rect 6601 11689 7820 11711
rect 6601 11680 7417 11689
rect 3733 11637 7417 11680
rect 7469 11680 7820 11689
rect 7872 11680 7886 11732
rect 7938 11680 7952 11732
rect 8004 11680 8018 11732
rect 8070 11680 8084 11732
rect 8136 11680 8150 11732
rect 8202 11680 8216 11732
rect 8268 11680 8282 11732
rect 8334 11680 8348 11732
rect 8400 11680 8414 11732
rect 8466 11680 8480 11732
rect 8532 11680 8546 11732
rect 8598 11680 8612 11732
rect 8664 11680 8677 11732
rect 8729 11680 8742 11732
rect 8794 11680 8807 11732
rect 8859 11680 8872 11732
rect 8924 11721 9890 11732
rect 9942 11721 11505 11773
rect 8924 11699 11505 11721
rect 8924 11680 9890 11699
rect 7469 11647 9890 11680
rect 9942 11647 11505 11699
rect 7469 11637 11505 11647
rect 3733 11636 11505 11637
rect 1176 11625 11505 11636
rect 1176 11617 9890 11625
rect 1228 11615 9890 11617
rect 1228 11614 7417 11615
rect 1228 11565 3681 11614
rect 1176 11562 3681 11565
rect 3733 11563 7417 11614
rect 7469 11573 9890 11615
rect 9942 11573 11505 11625
tri 11682 11616 11856 11790 se
rect 11856 11778 12018 11790
tri 12018 11778 12030 11790 nw
tri 12058 11778 12070 11790 se
rect 12070 11778 12232 11790
tri 12232 11778 12406 11952 nw
rect 11856 11738 11978 11778
tri 11978 11738 12018 11778 nw
tri 12018 11738 12058 11778 se
rect 11856 11698 11938 11738
tri 11938 11698 11978 11738 nw
tri 11978 11698 12018 11738 se
rect 12018 11698 12058 11738
rect 11856 11684 11924 11698
tri 11924 11684 11938 11698 nw
tri 11964 11684 11978 11698 se
rect 11978 11684 12058 11698
rect 11856 11644 11884 11684
tri 11884 11644 11924 11684 nw
tri 11924 11644 11964 11684 se
rect 11964 11644 12058 11684
tri 11856 11616 11884 11644 nw
tri 11896 11616 11924 11644 se
rect 11924 11616 12058 11644
rect 7469 11563 11505 11573
rect 3733 11562 11505 11563
rect 1176 11551 11505 11562
rect 1176 11544 9890 11551
rect 1228 11541 9890 11544
rect 1228 11540 7417 11541
rect 1228 11492 3681 11540
rect 1176 11488 3681 11492
rect 3733 11489 7417 11540
rect 7469 11499 9890 11541
rect 9942 11499 11505 11551
rect 7469 11493 11505 11499
tri 11559 11493 11682 11616 se
rect 11682 11604 11844 11616
tri 11844 11604 11856 11616 nw
tri 11884 11604 11896 11616 se
rect 11896 11604 12058 11616
tri 12058 11604 12232 11778 nw
rect 11682 11564 11804 11604
tri 11804 11564 11844 11604 nw
tri 11844 11564 11884 11604 se
rect 11682 11524 11764 11564
tri 11764 11524 11804 11564 nw
tri 11804 11524 11844 11564 se
rect 11844 11524 11884 11564
rect 11682 11510 11750 11524
tri 11750 11510 11764 11524 nw
tri 11790 11510 11804 11524 se
rect 11804 11510 11884 11524
rect 11682 11493 11710 11510
rect 7469 11489 9845 11493
rect 3733 11488 9845 11489
rect 1176 11470 9845 11488
rect 1228 11467 9845 11470
rect 1228 11418 3681 11467
rect 1176 11415 3681 11418
rect 3733 11415 7417 11467
rect 7469 11415 9845 11467
rect 1176 11412 9845 11415
rect 1179 11409 9845 11412
tri 9845 11409 9929 11493 nw
tri 11508 11442 11559 11493 se
rect 11559 11470 11710 11493
tri 11710 11470 11750 11510 nw
tri 11750 11470 11790 11510 se
rect 11790 11470 11884 11510
rect 11559 11442 11682 11470
tri 11682 11442 11710 11470 nw
tri 11722 11442 11750 11470 se
rect 11750 11442 11884 11470
tri 11475 11409 11508 11442 se
rect 11508 11430 11670 11442
tri 11670 11430 11682 11442 nw
tri 11710 11430 11722 11442 se
rect 11722 11430 11884 11442
tri 11884 11430 12058 11604 nw
rect 11508 11409 11630 11430
tri 11351 11285 11475 11409 se
rect 11475 11390 11630 11409
tri 11630 11390 11670 11430 nw
tri 11670 11390 11710 11430 se
rect 11475 11350 11590 11390
tri 11590 11350 11630 11390 nw
tri 11630 11350 11670 11390 se
rect 11670 11350 11710 11390
rect 11475 11336 11576 11350
tri 11576 11336 11590 11350 nw
tri 11616 11336 11630 11350 se
rect 11630 11336 11710 11350
rect 11475 11296 11536 11336
tri 11536 11296 11576 11336 nw
tri 11576 11296 11616 11336 se
rect 11616 11296 11710 11336
rect 11475 11285 11508 11296
rect 7516 11279 7568 11285
rect 7516 11215 7568 11227
rect 7516 11157 7568 11163
tri 7568 11157 7696 11285 sw
tri 11334 11268 11351 11285 se
rect 11351 11268 11508 11285
tri 11508 11268 11536 11296 nw
tri 11548 11268 11576 11296 se
rect 11576 11268 11710 11296
tri 11223 11157 11334 11268 se
rect 11334 11256 11496 11268
tri 11496 11256 11508 11268 nw
tri 11536 11256 11548 11268 se
rect 11548 11256 11710 11268
tri 11710 11256 11884 11430 nw
rect 11334 11216 11456 11256
tri 11456 11216 11496 11256 nw
tri 11496 11216 11536 11256 se
rect 11334 11197 11437 11216
tri 11437 11197 11456 11216 nw
tri 11477 11197 11496 11216 se
rect 11496 11197 11536 11216
rect 11334 11157 11397 11197
tri 11397 11157 11437 11197 nw
tri 11437 11157 11477 11197 se
rect 11477 11157 11536 11197
rect 7516 11151 11362 11157
rect 7568 11122 11362 11151
tri 11362 11122 11397 11157 nw
tri 11402 11122 11437 11157 se
rect 11437 11122 11536 11157
rect 7568 11099 11322 11122
rect 7516 11087 11322 11099
rect 7568 11082 11322 11087
tri 11322 11082 11362 11122 nw
tri 11362 11082 11402 11122 se
rect 11402 11082 11536 11122
tri 11536 11082 11710 11256 nw
rect 7568 11042 11282 11082
tri 11282 11042 11322 11082 nw
tri 11322 11042 11362 11082 se
rect 11362 11042 11427 11082
rect 7568 11035 11269 11042
rect 7516 11029 11269 11035
tri 11269 11029 11282 11042 nw
tri 11309 11029 11322 11042 se
rect 11322 11029 11427 11042
tri 11253 10973 11309 11029 se
rect 11309 10973 11427 11029
tri 11427 10973 11536 11082 nw
rect 5186 10967 11297 10973
rect 5238 10915 7026 10967
rect 7078 10915 11297 10967
rect 5186 10901 11297 10915
rect 5238 10849 7026 10901
rect 7078 10849 11297 10901
rect 5186 10843 11297 10849
tri 11297 10843 11427 10973 nw
rect 1202 10735 9539 10787
tri 9517 10713 9539 10735 ne
tri 9539 10713 9613 10787 sw
tri 9539 10648 9604 10713 ne
rect 9604 10648 9613 10713
tri 9613 10648 9678 10713 sw
tri 9604 10596 9656 10648 ne
rect 9656 10596 9846 10648
rect 1117 10243 12868 10249
rect 1117 10241 3681 10243
rect 1169 10189 1181 10241
rect 1233 10191 3681 10241
rect 3733 10191 5548 10243
rect 5600 10191 7417 10243
rect 7469 10191 9804 10243
rect 1233 10189 9804 10191
rect 1117 10179 9804 10189
rect 1117 10127 3681 10179
rect 3733 10127 5548 10179
rect 5600 10127 7417 10179
rect 7469 10127 9804 10179
rect 10048 10127 12868 10243
rect 1117 10114 12868 10127
rect 1169 10062 1181 10114
rect 1233 10062 3681 10114
rect 3733 10062 5548 10114
rect 5600 10062 7417 10114
rect 7469 10062 9804 10114
rect 9856 10062 9868 10114
rect 9920 10062 9932 10114
rect 9984 10062 9996 10114
rect 10048 10062 12868 10114
rect 1117 10056 12868 10062
rect 1384 9849 5320 9855
rect 1436 9797 3500 9849
rect 3552 9797 4850 9849
rect 4902 9797 4930 9849
rect 4982 9797 5320 9849
rect 1384 9783 5320 9797
rect 1436 9731 3500 9783
rect 3552 9731 4850 9783
rect 4902 9731 4930 9783
rect 4982 9731 5320 9783
rect 1384 9725 5320 9731
rect 5840 9849 9764 9855
rect 5840 9797 6703 9849
rect 6755 9797 6783 9849
rect 6835 9797 7596 9849
rect 7648 9797 9712 9849
rect 5840 9783 9764 9797
rect 5840 9731 6703 9783
rect 6755 9731 6783 9783
rect 6835 9731 7596 9783
rect 7648 9731 9712 9783
rect 5840 9725 9764 9731
tri 1245 9614 1251 9620 se
rect 1251 9614 10206 9620
tri 1145 9514 1245 9614 se
rect 1245 9514 10078 9614
rect 1117 9498 10078 9514
rect 10194 9498 10206 9614
rect 1117 9485 10206 9498
rect 1117 9433 10078 9485
rect 10130 9433 10142 9485
rect 10194 9433 10206 9485
rect 1117 9420 10206 9433
rect 1117 9368 10078 9420
rect 10130 9368 10142 9420
rect 10194 9368 10206 9420
rect 1117 9362 10206 9368
rect 1117 9230 1226 9362
tri 1226 9230 1358 9362 nw
rect 1202 9124 9846 9176
rect 4070 8983 5962 8989
rect 4122 8931 5910 8983
rect 4070 8917 5962 8931
rect 4122 8865 5910 8917
rect 4070 8859 5962 8865
rect 1117 8540 10206 8546
rect 1117 8488 10078 8540
rect 10130 8488 10142 8540
rect 10194 8488 10206 8540
rect 1117 8473 10206 8488
rect 1117 8421 10078 8473
rect 10130 8421 10142 8473
rect 10194 8421 10206 8473
rect 1117 8406 10206 8421
rect 1117 8354 10078 8406
rect 10130 8354 10142 8406
rect 10194 8354 10206 8406
rect 1117 8338 10206 8354
rect 1117 8286 10078 8338
rect 10130 8286 10142 8338
rect 10194 8286 10206 8338
rect 1117 8280 10206 8286
rect 1117 8146 12868 8152
rect 1233 8094 3681 8146
rect 3733 8094 5548 8146
rect 5600 8094 7417 8146
rect 7469 8094 9804 8146
rect 1233 8082 9804 8094
rect 1233 8030 3681 8082
rect 3733 8030 5548 8082
rect 5600 8030 7417 8082
rect 7469 8030 9804 8082
rect 10048 8049 12868 8146
rect 10048 8030 10311 8049
rect 1117 8017 10311 8030
rect 1169 7965 1181 8017
rect 1233 7965 3681 8017
rect 3733 7965 5548 8017
rect 5600 7965 7417 8017
rect 7469 7965 9804 8017
rect 9856 7965 9868 8017
rect 9920 7965 9932 8017
rect 9984 7965 9996 8017
rect 10048 7997 10311 8017
rect 10363 7997 10376 8049
rect 10428 7997 10441 8049
rect 10493 7997 10506 8049
rect 10558 7997 10571 8049
rect 10623 7997 10636 8049
rect 10688 7997 10701 8049
rect 10753 7997 10766 8049
rect 10818 7997 10831 8049
rect 10883 7997 10896 8049
rect 10948 7997 10961 8049
rect 11013 7997 11026 8049
rect 11078 7997 11091 8049
rect 11143 7997 11156 8049
rect 11208 7997 11221 8049
rect 11273 7997 11286 8049
rect 11338 7997 11350 8049
rect 11402 7997 11414 8049
rect 11466 7997 11478 8049
rect 11530 7997 11542 8049
rect 11594 7997 11606 8049
rect 11658 7997 11670 8049
rect 11722 7997 11734 8049
rect 11786 7997 11798 8049
rect 11850 7997 11862 8049
rect 11914 7997 11926 8049
rect 11978 7997 11990 8049
rect 12042 7997 12054 8049
rect 12106 7997 12118 8049
rect 12170 7997 12182 8049
rect 12234 7997 12246 8049
rect 12298 7997 12310 8049
rect 12362 7997 12374 8049
rect 12426 7997 12438 8049
rect 12490 7997 12502 8049
rect 12554 7997 12566 8049
rect 12618 7997 12630 8049
rect 12682 7997 12694 8049
rect 12746 7997 12758 8049
rect 12810 7997 12868 8049
rect 10048 7965 12868 7997
rect 1117 7959 12868 7965
rect 7684 7763 12868 7770
rect 7684 7647 7698 7763
rect 7814 7647 12868 7763
rect 7684 7640 12868 7647
rect 2977 7532 2983 7584
rect 3035 7532 3047 7584
rect 3099 7532 3111 7584
rect 3163 7532 3175 7584
rect 3227 7532 10320 7584
tri 11575 7476 11600 7501 se
rect 11600 7479 11652 7532
tri 11652 7507 11677 7532 nw
rect 11600 7476 11649 7479
tri 11649 7476 11652 7479 nw
rect 8658 7424 8664 7476
rect 8716 7424 8728 7476
rect 8780 7424 8792 7476
rect 8844 7424 8856 7476
rect 8908 7424 11597 7476
tri 11597 7424 11649 7476 nw
rect 1117 7341 10245 7347
rect 1117 7161 3768 7341
rect 3884 7161 5678 7341
rect 5794 7161 7266 7341
rect 7382 7289 10193 7341
rect 7382 7277 10245 7289
rect 7382 7225 10193 7277
rect 7382 7213 10245 7225
rect 7382 7161 10193 7213
rect 1117 7155 10245 7161
rect 5186 7043 7078 7049
rect 5238 6991 7026 7043
rect 5186 6977 7078 6991
rect 5238 6925 7026 6977
rect 5186 6919 7078 6925
rect 1117 6819 13007 6825
rect 1117 6639 3768 6819
rect 3884 6639 5678 6819
rect 5794 6639 7266 6819
rect 7382 6767 10193 6819
rect 10245 6767 12891 6819
rect 7382 6755 12891 6767
rect 7382 6703 10193 6755
rect 10245 6703 12891 6755
rect 7382 6691 12891 6703
rect 7382 6639 10193 6691
rect 10245 6639 12891 6691
rect 1117 6633 13007 6639
rect 1384 6474 10099 6480
rect 1436 6422 3500 6474
rect 3552 6422 10047 6474
rect 1384 6408 10099 6422
rect 1436 6356 3500 6408
rect 3552 6356 10047 6408
rect 1384 6350 10099 6356
rect 7596 6258 10019 6264
rect 7648 6206 9712 6258
rect 9764 6206 9967 6258
rect 7596 6192 10019 6206
rect 7648 6140 9712 6192
rect 9764 6140 9967 6192
rect 7596 6134 10019 6140
rect 1150 6032 13007 6084
rect 1150 5940 13007 5992
rect 1117 5638 13007 5644
rect 1117 5458 3768 5638
rect 3884 5458 5678 5638
rect 5794 5458 7266 5638
rect 7382 5586 10193 5638
rect 10245 5586 12891 5638
rect 12943 5586 12955 5638
rect 7382 5574 13007 5586
rect 7382 5522 10193 5574
rect 10245 5564 13007 5574
rect 10245 5522 12891 5564
rect 7382 5512 12891 5522
rect 12943 5512 12955 5564
rect 7382 5510 13007 5512
rect 7382 5458 10193 5510
rect 10245 5490 13007 5510
rect 10245 5458 12891 5490
rect 1117 5452 12891 5458
tri 12703 5438 12717 5452 ne
rect 12717 5438 12891 5452
rect 12943 5438 12955 5490
tri 12717 5416 12739 5438 ne
rect 12739 5416 13007 5438
tri 12739 5364 12791 5416 ne
rect 12791 5364 12891 5416
rect 12943 5364 12955 5416
tri 13007 5393 13149 5535 sw
rect 13007 5364 13149 5393
tri 12791 5341 12814 5364 ne
rect 12814 5341 13149 5364
tri 12814 5289 12866 5341 ne
rect 12866 5289 12891 5341
rect 12943 5289 12955 5341
rect 13007 5289 13149 5341
tri 12866 5288 12867 5289 ne
rect 12867 5288 13149 5289
rect 4070 5282 5962 5288
rect 4122 5230 5910 5282
tri 12867 5266 12889 5288 ne
rect 12889 5266 13149 5288
tri 12889 5264 12891 5266 ne
rect 4070 5216 5962 5230
rect 4122 5164 5910 5216
rect 4070 5158 5962 5164
rect 12943 5214 12955 5266
rect 13007 5214 13149 5266
rect 12891 5191 13149 5214
rect 12943 5139 12955 5191
rect 13007 5139 13149 5191
rect 12891 5133 13149 5139
rect 1117 4880 13115 4886
rect 1169 4828 1181 4880
rect 1233 4828 3681 4880
rect 3733 4828 5548 4880
rect 5600 4828 7417 4880
rect 7469 4828 9817 4880
rect 9869 4828 9881 4880
rect 9933 4828 13063 4880
rect 1117 4814 13115 4828
rect 1169 4762 1181 4814
rect 1233 4762 3681 4814
rect 3733 4762 5548 4814
rect 5600 4762 7417 4814
rect 7469 4762 9817 4814
rect 9869 4762 9881 4814
rect 9933 4762 13063 4814
rect 1117 4756 13115 4762
rect 7686 4236 7692 4288
rect 7744 4236 7756 4288
rect 7808 4236 11599 4288
tri 11575 4212 11599 4236 ne
tri 11599 4235 11652 4288 sw
rect 11599 4212 11652 4235
tri 11599 4211 11600 4212 ne
rect 1117 4203 7382 4209
rect 1117 4023 3768 4203
rect 3884 4023 5367 4203
rect 5483 4023 5678 4203
rect 5794 4023 7266 4203
rect 11600 4180 11652 4212
tri 11652 4180 11677 4205 sw
tri 7583 4106 7657 4180 se
rect 7657 4128 10320 4180
tri 7657 4106 7679 4128 nw
tri 7523 4046 7583 4106 se
rect 7583 4046 7597 4106
tri 7597 4046 7657 4106 nw
rect 10047 4046 10163 4052
tri 7509 4032 7523 4046 se
rect 7523 4032 7583 4046
tri 7583 4032 7597 4046 nw
rect 1117 4017 7382 4023
tri 7499 4022 7509 4032 se
rect 7509 4022 7573 4032
tri 7573 4022 7583 4032 nw
rect 9967 4022 10019 4028
tri 7494 4017 7499 4022 se
rect 7499 4017 7521 4022
tri 7447 3970 7494 4017 se
rect 7494 3970 7521 4017
tri 7521 3970 7573 4022 nw
rect 10099 3994 10111 4046
tri 10163 4030 10185 4052 sw
rect 10163 3994 10320 4030
rect 10047 3988 10320 3994
tri 10047 3978 10057 3988 ne
rect 10057 3978 10320 3988
rect 11600 3978 11652 4005
tri 7438 3961 7447 3970 se
rect 7447 3961 7512 3970
tri 7512 3961 7521 3970 nw
rect 3334 3909 3340 3961
rect 3392 3909 3404 3961
rect 3456 3956 7507 3961
tri 7507 3956 7512 3961 nw
rect 9967 3956 10019 3970
rect 3456 3909 7460 3956
tri 7460 3909 7507 3956 nw
tri 10019 3950 10044 3975 sw
tri 11575 3950 11600 3975 se
rect 11600 3950 11649 3978
tri 11649 3950 11677 3978 nw
rect 10019 3904 11597 3950
rect 9967 3898 11597 3904
tri 11597 3898 11649 3950 nw
tri 8023 3376 8123 3476 se
rect 8123 3376 13007 3476
rect 4904 3324 4910 3376
rect 4962 3324 4974 3376
rect 5026 3324 5038 3376
rect 5090 3324 6792 3376
rect 6844 3324 6856 3376
rect 6908 3324 6920 3376
rect 6972 3324 6978 3376
tri 7971 3324 8023 3376 se
rect 8023 3324 13007 3376
tri 7915 3268 7971 3324 se
rect 7971 3268 13007 3324
rect 5209 2666 13007 3268
rect 2342 2066 13007 2072
rect 2342 2060 12891 2066
rect 2342 2008 10193 2060
rect 10245 2014 12891 2060
rect 12943 2014 12955 2066
rect 10245 2008 13007 2014
rect 2342 2001 13007 2008
rect 2342 1996 12891 2001
rect 2342 1944 10193 1996
rect 10245 1949 12891 1996
rect 12943 1949 12955 2001
rect 10245 1944 13007 1949
rect 2342 1936 13007 1944
rect 2342 1932 12891 1936
rect 2342 1880 10193 1932
rect 10245 1884 12891 1932
rect 12943 1884 12955 1936
rect 10245 1880 13007 1884
rect 2342 1870 13007 1880
rect 2342 1868 12891 1870
rect 2342 1816 10193 1868
rect 10245 1818 12891 1868
rect 12943 1818 12955 1870
rect 10245 1816 13007 1818
rect 2342 1804 13007 1816
rect 2342 1752 10193 1804
rect 10245 1752 12891 1804
rect 12943 1752 12955 1804
rect 2342 1746 13007 1752
rect 2342 1588 8809 1623
rect 2342 1536 2354 1588
rect 2406 1536 2420 1588
rect 2472 1536 2486 1588
rect 2538 1536 2552 1588
rect 2604 1536 2618 1588
rect 2670 1536 2684 1588
rect 2736 1536 2749 1588
rect 2801 1536 2814 1588
rect 2866 1536 2879 1588
rect 2931 1536 2944 1588
rect 2996 1536 6794 1588
rect 2342 1524 6794 1536
rect 2342 1472 2354 1524
rect 2406 1472 2420 1524
rect 2472 1472 2486 1524
rect 2538 1472 2552 1524
rect 2604 1472 2618 1524
rect 2670 1472 2684 1524
rect 2736 1472 2749 1524
rect 2801 1472 2814 1524
rect 2866 1472 2879 1524
rect 2931 1472 2944 1524
rect 2996 1472 6794 1524
rect 2342 1460 6794 1472
rect 2342 1408 2354 1460
rect 2406 1408 2420 1460
rect 2472 1408 2486 1460
rect 2538 1408 2552 1460
rect 2604 1408 2618 1460
rect 2670 1408 2684 1460
rect 2736 1408 2749 1460
rect 2801 1408 2814 1460
rect 2866 1408 2879 1460
rect 2931 1408 2944 1460
rect 2996 1408 6794 1460
rect 2342 1396 6794 1408
rect 2342 1344 2354 1396
rect 2406 1344 2420 1396
rect 2472 1344 2486 1396
rect 2538 1344 2552 1396
rect 2604 1344 2618 1396
rect 2670 1344 2684 1396
rect 2736 1344 2749 1396
rect 2801 1344 2814 1396
rect 2866 1344 2879 1396
rect 2931 1344 2944 1396
rect 2996 1344 6794 1396
rect 2342 1332 6794 1344
rect 2342 1280 2354 1332
rect 2406 1280 2420 1332
rect 2472 1280 2486 1332
rect 2538 1280 2552 1332
rect 2604 1280 2618 1332
rect 2670 1280 2684 1332
rect 2736 1280 2749 1332
rect 2801 1280 2814 1332
rect 2866 1280 2879 1332
rect 2931 1280 2944 1332
rect 2996 1280 6794 1332
rect 6974 1280 7266 1588
rect 7382 1536 8151 1588
rect 8203 1536 8217 1588
rect 8269 1536 8283 1588
rect 8335 1536 8349 1588
rect 8401 1536 8415 1588
rect 8467 1536 8481 1588
rect 8533 1536 8546 1588
rect 8598 1536 8611 1588
rect 8663 1536 8676 1588
rect 8728 1536 8741 1588
rect 8793 1536 8809 1588
rect 7382 1524 8809 1536
rect 7382 1472 8151 1524
rect 8203 1472 8217 1524
rect 8269 1472 8283 1524
rect 8335 1472 8349 1524
rect 8401 1472 8415 1524
rect 8467 1472 8481 1524
rect 8533 1472 8546 1524
rect 8598 1472 8611 1524
rect 8663 1472 8676 1524
rect 8728 1472 8741 1524
rect 8793 1472 8809 1524
rect 7382 1460 8809 1472
rect 7382 1408 8151 1460
rect 8203 1408 8217 1460
rect 8269 1408 8283 1460
rect 8335 1408 8349 1460
rect 8401 1408 8415 1460
rect 8467 1408 8481 1460
rect 8533 1408 8546 1460
rect 8598 1408 8611 1460
rect 8663 1408 8676 1460
rect 8728 1408 8741 1460
rect 8793 1408 8809 1460
rect 7382 1396 8809 1408
rect 7382 1344 8151 1396
rect 8203 1344 8217 1396
rect 8269 1344 8283 1396
rect 8335 1344 8349 1396
rect 8401 1344 8415 1396
rect 8467 1344 8481 1396
rect 8533 1344 8546 1396
rect 8598 1344 8611 1396
rect 8663 1344 8676 1396
rect 8728 1344 8741 1396
rect 8793 1344 8809 1396
rect 7382 1332 8809 1344
rect 7382 1280 8151 1332
rect 8203 1280 8217 1332
rect 8269 1280 8283 1332
rect 8335 1280 8349 1332
rect 8401 1280 8415 1332
rect 8467 1280 8481 1332
rect 8533 1280 8546 1332
rect 8598 1280 8611 1332
rect 8663 1280 8676 1332
rect 8728 1280 8741 1332
rect 8793 1280 8809 1332
rect 2342 1247 8809 1280
rect 1384 1185 1985 1191
rect 1436 1133 1933 1185
rect 1384 1121 1985 1133
rect 1436 1069 1933 1121
rect 1384 1063 1985 1069
rect 3073 1185 3552 1191
rect 3125 1133 3500 1185
rect 3073 1121 3552 1133
rect 3125 1069 3500 1121
rect 3073 1063 3552 1069
rect 5188 1185 7568 1191
rect 5240 1133 7020 1185
rect 7072 1133 7452 1185
rect 5188 1121 7452 1133
rect 5240 1069 7020 1121
rect 7072 1069 7452 1121
rect 5188 1063 7568 1069
rect 7596 1185 8075 1191
rect 7648 1133 8023 1185
rect 7596 1121 8075 1133
rect 7648 1069 8023 1121
rect 7596 1063 8075 1069
rect 9163 1185 9764 1191
rect 9215 1133 9712 1185
rect 9163 1121 9764 1133
rect 9215 1069 9712 1121
rect 9163 1063 9764 1069
rect 3334 955 3340 1007
rect 3392 955 3404 1007
rect 3456 996 9294 1007
tri 9294 996 9305 1007 sw
rect 3456 955 9305 996
tri 9272 924 9303 955 ne
rect 9303 924 9305 955
rect 1532 918 1584 924
tri 9303 922 9305 924 ne
tri 9305 922 9379 996 sw
tri 9305 899 9328 922 ne
rect 9328 899 9379 922
tri 3845 873 3871 899 se
rect 3871 873 5369 899
rect 1532 854 1584 866
tri 1584 848 1609 873 sw
tri 3820 848 3845 873 se
rect 3845 848 5369 873
rect 1584 802 3506 848
rect 1532 796 3506 802
rect 3558 796 3570 848
rect 3622 796 3628 848
tri 3768 796 3820 848 se
rect 3820 796 5369 848
tri 3755 783 3768 796 se
rect 3768 783 5369 796
rect 5485 783 5491 899
rect 5669 783 5675 899
rect 5791 783 7277 899
tri 3740 768 3755 783 se
rect 3755 768 3904 783
tri 3904 768 3919 783 nw
tri 7229 768 7244 783 ne
rect 7244 768 7277 783
tri 7277 768 7408 899 sw
tri 9328 848 9379 899 ne
tri 9379 848 9453 922 sw
tri 9379 774 9453 848 ne
tri 9453 774 9527 848 sw
tri 9453 768 9459 774 ne
rect 9459 768 9527 774
rect 2559 716 2565 768
rect 2617 716 3077 768
rect 3129 716 3340 768
rect 2559 704 3340 716
rect 2559 652 2565 704
rect 2617 652 3077 704
rect 3129 652 3340 704
rect 3456 652 3788 768
tri 3788 652 3904 768 nw
tri 7244 735 7277 768 ne
rect 7277 735 7692 768
tri 7277 717 7295 735 ne
rect 7295 717 7692 735
rect 1119 545 1417 597
tri 1394 522 1417 545 ne
tri 1417 522 1492 597 sw
tri 1417 517 1422 522 ne
rect 1422 517 1492 522
rect 1119 508 1365 517
tri 1365 508 1374 517 sw
tri 1422 508 1431 517 ne
rect 1431 508 1492 517
tri 1492 508 1506 522 sw
rect 1827 508 1833 624
rect 1949 572 2309 624
rect 2361 572 2821 624
rect 2873 572 3386 624
rect 1949 560 3386 572
rect 1949 508 2309 560
rect 2361 508 2821 560
rect 2873 508 3264 560
rect 3316 508 3328 560
rect 3380 508 3386 560
rect 5131 537 6374 717
tri 7295 652 7360 717 ne
rect 7360 652 7692 717
rect 7808 716 8019 768
rect 8071 716 8531 768
rect 8583 716 8589 768
rect 7808 704 8589 716
tri 8589 704 8653 768 sw
tri 9459 704 9523 768 ne
rect 9523 704 9527 768
rect 7808 652 8019 704
rect 8071 652 8531 704
rect 8583 666 9356 704
tri 9356 666 9394 704 sw
tri 9523 700 9527 704 ne
tri 9527 700 9601 774 sw
tri 9527 666 9561 700 ne
rect 9561 666 9601 700
rect 8583 652 9394 666
tri 9334 624 9362 652 ne
rect 9362 624 9394 652
rect 7762 585 8275 624
rect 7026 550 7078 556
rect 1119 498 1374 508
tri 1374 498 1384 508 sw
tri 1431 498 1441 508 ne
rect 1441 498 1506 508
tri 1506 498 1516 508 sw
tri 7019 498 7026 505 se
rect 7814 533 7826 585
rect 7878 572 8275 585
rect 8327 572 8787 624
rect 8839 572 9199 624
rect 9251 572 9257 624
tri 9362 592 9394 624 ne
tri 9394 592 9468 666 sw
tri 9561 626 9601 666 ne
tri 9601 626 9675 700 sw
tri 9601 592 9635 626 ne
rect 9635 592 10320 626
rect 7878 560 9257 572
rect 7878 533 8275 560
rect 7762 508 8275 533
rect 8327 508 8787 560
rect 8839 508 9199 560
rect 9251 508 9257 560
tri 9394 518 9468 592 ne
tri 9468 518 9542 592 sw
tri 9635 574 9653 592 ne
rect 9653 574 10320 592
tri 11575 518 11600 543 se
rect 11600 520 11652 579
tri 11652 549 11677 574 nw
rect 11600 518 11650 520
tri 11650 518 11652 520 nw
tri 9468 508 9478 518 ne
rect 9478 508 11598 518
rect 1119 486 1384 498
tri 1384 486 1396 498 sw
tri 1441 486 1453 498 ne
rect 1453 486 1516 498
tri 1516 486 1528 498 sw
tri 7007 486 7019 498 se
rect 7019 486 7078 498
rect 1119 480 1396 486
tri 1396 480 1402 486 sw
tri 1453 480 1459 486 ne
rect 1459 480 1528 486
tri 1528 480 1534 486 sw
tri 7001 480 7007 486 se
rect 7007 480 7026 486
rect 1119 465 1402 480
tri 1342 442 1365 465 ne
rect 1365 442 1402 465
tri 1402 442 1440 480 sw
tri 1459 442 1497 480 ne
rect 1497 442 1618 480
tri 1365 437 1370 442 ne
rect 1370 437 1440 442
rect 1119 428 1313 437
tri 1313 428 1322 437 sw
tri 1370 428 1379 437 ne
rect 1379 428 1440 437
tri 1440 428 1454 442 sw
tri 1497 428 1511 442 ne
rect 1511 428 1618 442
rect 1670 428 1682 480
rect 1734 428 5186 480
rect 5238 428 5250 480
rect 5302 428 5763 480
rect 5815 428 5827 480
rect 5879 434 7026 480
tri 9478 466 9520 508 ne
rect 9520 466 11598 508
tri 11598 466 11650 518 nw
rect 5879 428 7078 434
rect 1119 419 1322 428
tri 1322 419 1331 428 sw
tri 1379 419 1388 428 ne
rect 1388 419 1454 428
rect 1119 388 1331 419
tri 1331 388 1362 419 sw
tri 1388 388 1419 419 ne
rect 1419 388 1454 419
tri 1454 388 1494 428 sw
rect 1119 385 1362 388
tri 1290 362 1313 385 ne
rect 1313 362 1362 385
tri 1362 362 1388 388 sw
tri 1419 362 1445 388 ne
rect 1445 362 13007 388
tri 1313 296 1379 362 ne
rect 1379 353 1388 362
tri 1388 353 1397 362 sw
tri 1445 353 1454 362 ne
rect 1454 353 13007 362
rect 1379 336 1397 353
tri 1397 336 1414 353 sw
tri 1454 336 1471 353 ne
rect 1471 336 13007 353
rect 1379 296 1414 336
tri 1414 296 1454 336 sw
tri 1379 244 1431 296 ne
rect 1431 244 13007 296
rect 1119 -289 5969 31
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_0
timestamp 1704896540
transform 0 1 3175 -1 0 800
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_1
timestamp 1704896540
transform -1 0 7621 0 -1 860
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1704896540
transform 0 -1 7652 -1 0 708
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1704896540
transform 0 1 5712 1 0 2942
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1704896540
transform 0 -1 3540 1 0 599
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1704896540
transform 0 -1 3540 1 0 757
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_4
timestamp 1704896540
transform 1 0 3268 0 -1 553
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_5
timestamp 1704896540
transform 1 0 7774 0 -1 578
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1704896540
transform 0 1 9054 1 0 622
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_1
timestamp 1704896540
transform 0 -1 2094 1 0 622
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_0
timestamp 1704896540
transform -1 0 3118 0 -1 730
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_1
timestamp 1704896540
transform -1 0 2606 0 -1 730
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_2
timestamp 1704896540
transform -1 0 2350 0 -1 708
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_3
timestamp 1704896540
transform -1 0 1828 0 -1 708
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_4
timestamp 1704896540
transform -1 0 1938 0 -1 708
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_5
timestamp 1704896540
transform -1 0 2862 0 -1 708
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_6
timestamp 1704896540
transform -1 0 1572 0 -1 726
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_7
timestamp 1704896540
transform 1 0 8286 0 -1 708
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_8
timestamp 1704896540
transform 1 0 9210 0 -1 708
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_9
timestamp 1704896540
transform 1 0 8798 0 -1 708
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_10
timestamp 1704896540
transform 1 0 8542 0 -1 730
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_11
timestamp 1704896540
transform 1 0 8030 0 -1 730
box 0 0 1 1
use L1M1_CDNS_52468879185326  L1M1_CDNS_52468879185326_0
timestamp 1704896540
transform -1 0 8833 0 1 1770
box -12 -6 694 40
use L1M1_CDNS_52468879185326  L1M1_CDNS_52468879185326_1
timestamp 1704896540
transform -1 0 8833 0 1 914
box -12 -6 694 40
use L1M1_CDNS_52468879185326  L1M1_CDNS_52468879185326_2
timestamp 1704896540
transform 1 0 4153 0 -1 2858
box -12 -6 694 40
use L1M1_CDNS_52468879185326  L1M1_CDNS_52468879185326_3
timestamp 1704896540
transform 1 0 5993 0 -1 2858
box -12 -6 694 40
use L1M1_CDNS_52468879185326  L1M1_CDNS_52468879185326_4
timestamp 1704896540
transform 1 0 2315 0 1 1770
box -12 -6 694 40
use L1M1_CDNS_52468879185326  L1M1_CDNS_52468879185326_5
timestamp 1704896540
transform 1 0 2315 0 1 914
box -12 -6 694 40
use L1M1_CDNS_524688791851014  L1M1_CDNS_524688791851014_0
timestamp 1704896540
transform 0 -1 5123 -1 0 3115
box -12 -6 46 760
use L1M1_CDNS_524688791851014  L1M1_CDNS_524688791851014_1
timestamp 1704896540
transform 0 -1 6963 -1 0 3114
box -12 -6 46 760
use L1M1_CDNS_524688791851015  L1M1_CDNS_524688791851015_0
timestamp 1704896540
transform 0 -1 5123 -1 0 1578
box -12 -6 46 904
use L1M1_CDNS_524688791851015  L1M1_CDNS_524688791851015_1
timestamp 1704896540
transform 0 -1 5123 -1 0 1066
box -12 -6 46 904
use L1M1_CDNS_524688791851015  L1M1_CDNS_524688791851015_2
timestamp 1704896540
transform 0 -1 5123 -1 0 2090
box -12 -6 46 904
use L1M1_CDNS_524688791851015  L1M1_CDNS_524688791851015_3
timestamp 1704896540
transform 0 -1 6963 -1 0 910
box -12 -6 46 904
use L1M1_CDNS_524688791851015  L1M1_CDNS_524688791851015_4
timestamp 1704896540
transform 0 -1 6963 -1 0 2090
box -12 -6 46 904
use L1M1_CDNS_524688791851015  L1M1_CDNS_524688791851015_5
timestamp 1704896540
transform 0 -1 6963 -1 0 1066
box -12 -6 46 904
use L1M1_CDNS_524688791851015  L1M1_CDNS_524688791851015_6
timestamp 1704896540
transform 0 -1 6963 -1 0 1578
box -12 -6 46 904
use L1M1_CDNS_524688791851015  L1M1_CDNS_524688791851015_7
timestamp 1704896540
transform 0 -1 6963 -1 0 800
box -12 -6 46 904
use L1M1_CDNS_524688791851015  L1M1_CDNS_524688791851015_8
timestamp 1704896540
transform 0 -1 6963 -1 0 488
box -12 -6 46 904
use L1M1_CDNS_524688791851015  L1M1_CDNS_524688791851015_9
timestamp 1704896540
transform 0 1 4166 -1 0 488
box -12 -6 46 904
use L1M1_CDNS_524688791851016  L1M1_CDNS_524688791851016_0
timestamp 1704896540
transform 0 -1 4907 -1 0 1322
box -12 -6 46 616
use L1M1_CDNS_524688791851016  L1M1_CDNS_524688791851016_1
timestamp 1704896540
transform 0 -1 4907 -1 0 1834
box -12 -6 46 616
use L1M1_CDNS_524688791851016  L1M1_CDNS_524688791851016_2
timestamp 1704896540
transform 0 -1 4907 -1 0 2346
box -12 -6 46 616
use L1M1_CDNS_524688791851016  L1M1_CDNS_524688791851016_3
timestamp 1704896540
transform 0 -1 5100 -1 0 644
box -12 -6 46 616
use L1M1_CDNS_524688791851016  L1M1_CDNS_524688791851016_4
timestamp 1704896540
transform 0 -1 6747 -1 0 2346
box -12 -6 46 616
use L1M1_CDNS_524688791851016  L1M1_CDNS_524688791851016_5
timestamp 1704896540
transform 0 -1 6747 -1 0 1834
box -12 -6 46 616
use L1M1_CDNS_524688791851016  L1M1_CDNS_524688791851016_6
timestamp 1704896540
transform 0 -1 6747 -1 0 1322
box -12 -6 46 616
use L1M1_CDNS_524688791851018  L1M1_CDNS_524688791851018_0
timestamp 1704896540
transform 0 -1 5123 -1 0 2602
box -12 -6 46 832
use L1M1_CDNS_524688791851018  L1M1_CDNS_524688791851018_1
timestamp 1704896540
transform 0 -1 6963 -1 0 2602
box -12 -6 46 832
use L1M1_CDNS_524688791851064  L1M1_CDNS_524688791851064_0
timestamp 1704896540
transform 0 -1 6963 -1 0 3370
box -12 -6 46 688
use L1M1_CDNS_524688791851064  L1M1_CDNS_524688791851064_1
timestamp 1704896540
transform 0 -1 5136 -1 0 3370
box -12 -6 46 688
use L1M1_CDNS_524688791851064  L1M1_CDNS_524688791851064_2
timestamp 1704896540
transform 0 1 6002 -1 0 644
box -12 -6 46 688
use L1M1_CDNS_524688791851064  L1M1_CDNS_524688791851064_3
timestamp 1704896540
transform 0 1 4166 -1 0 910
box -12 -6 46 688
use L1M1_CDNS_524688791851064  L1M1_CDNS_524688791851064_4
timestamp 1704896540
transform 0 1 4166 -1 0 800
box -12 -6 46 688
use L1M1_CDNS_524688791851579  L1M1_CDNS_524688791851579_0
timestamp 1704896540
transform -1 0 4205 0 1 11997
box -12 -6 478 184
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1704896540
transform 0 -1 3125 -1 0 1191
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_1
timestamp 1704896540
transform 0 -1 3552 -1 0 1191
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_2
timestamp 1704896540
transform 0 -1 9764 -1 0 1191
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_3
timestamp 1704896540
transform 0 -1 9215 -1 0 1191
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_4
timestamp 1704896540
transform 0 1 1933 -1 0 1191
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_5
timestamp 1704896540
transform 0 1 1384 -1 0 1191
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_6
timestamp 1704896540
transform 0 1 7895 -1 0 13079
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_7
timestamp 1704896540
transform 0 1 7596 -1 0 1191
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_8
timestamp 1704896540
transform 0 1 8023 -1 0 1191
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_9
timestamp 1704896540
transform -1 0 5885 0 1 428
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_10
timestamp 1704896540
transform -1 0 5308 0 -1 480
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_11
timestamp 1704896540
transform -1 0 5617 0 -1 12467
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_12
timestamp 1704896540
transform -1 0 1569 0 -1 12467
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_13
timestamp 1704896540
transform 0 1 7026 1 0 428
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_14
timestamp 1704896540
transform 0 -1 3187 1 0 12875
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_15
timestamp 1704896540
transform 0 -1 4527 1 0 12148
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_16
timestamp 1704896540
transform 0 -1 6367 1 0 12148
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_17
timestamp 1704896540
transform 0 -1 3529 1 0 12521
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_18
timestamp 1704896540
transform 0 -1 5499 1 0 12521
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_19
timestamp 1704896540
transform 0 -1 5240 1 0 1063
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_20
timestamp 1704896540
transform 0 -1 7072 1 0 1063
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_21
timestamp 1704896540
transform 0 -1 9658 1 0 12521
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_22
timestamp 1704896540
transform 0 -1 1584 1 0 796
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_23
timestamp 1704896540
transform 1 0 3258 0 -1 560
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_24
timestamp 1704896540
transform 1 0 3500 0 -1 848
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_25
timestamp 1704896540
transform 1 0 3334 0 1 955
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_26
timestamp 1704896540
transform 1 0 3334 0 1 3909
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_27
timestamp 1704896540
transform 1 0 7686 0 1 4236
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_28
timestamp 1704896540
transform 1 0 1612 0 1 428
box 0 0 1 1
use M1M2_CDNS_52468879185197  M1M2_CDNS_52468879185197_0
timestamp 1704896540
transform 0 1 7266 1 0 8285
box 0 0 256 116
use M1M2_CDNS_52468879185197  M1M2_CDNS_52468879185197_1
timestamp 1704896540
transform 0 1 7266 1 0 9363
box 0 0 256 116
use M1M2_CDNS_52468879185197  M1M2_CDNS_52468879185197_2
timestamp 1704896540
transform 0 1 5682 1 0 9363
box 0 0 256 116
use M1M2_CDNS_52468879185197  M1M2_CDNS_52468879185197_3
timestamp 1704896540
transform 0 1 5682 1 0 8285
box 0 0 256 116
use M1M2_CDNS_52468879185197  M1M2_CDNS_52468879185197_4
timestamp 1704896540
transform 0 1 3767 1 0 9363
box 0 0 256 116
use M1M2_CDNS_52468879185197  M1M2_CDNS_52468879185197_5
timestamp 1704896540
transform 0 1 3767 1 0 8285
box 0 0 256 116
use M1M2_CDNS_52468879185197  M1M2_CDNS_52468879185197_6
timestamp 1704896540
transform 1 0 10010 0 1 12004
box 0 0 256 116
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_0
timestamp 1704896540
transform 0 -1 7382 -1 0 4209
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_1
timestamp 1704896540
transform 0 -1 3884 -1 0 4209
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_2
timestamp 1704896540
transform 0 -1 5794 -1 0 4209
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_3
timestamp 1704896540
transform 0 -1 5483 -1 0 4209
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_4
timestamp 1704896540
transform 0 -1 7382 -1 0 6825
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_5
timestamp 1704896540
transform 0 -1 7382 -1 0 5644
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_6
timestamp 1704896540
transform 0 -1 7382 -1 0 7347
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_7
timestamp 1704896540
transform 0 -1 5794 -1 0 5644
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_8
timestamp 1704896540
transform 0 -1 3884 -1 0 5644
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_9
timestamp 1704896540
transform 0 -1 3884 -1 0 6825
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_10
timestamp 1704896540
transform 0 -1 5794 -1 0 6825
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_11
timestamp 1704896540
transform 0 -1 5794 -1 0 7347
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_12
timestamp 1704896540
transform 0 -1 3884 -1 0 7347
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_0
timestamp 1704896540
transform -1 0 1955 0 1 508
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_1
timestamp 1704896540
transform -1 0 5491 0 1 783
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_2
timestamp 1704896540
transform -1 0 3462 0 -1 768
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_3
timestamp 1704896540
transform 0 1 8970 1 0 12148
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_4
timestamp 1704896540
transform 0 1 7452 1 0 1063
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_5
timestamp 1704896540
transform 0 -1 2164 1 0 12148
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_6
timestamp 1704896540
transform 1 0 5669 0 1 783
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_7
timestamp 1704896540
transform 1 0 7686 0 1 652
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_8
timestamp 1704896540
transform 1 0 3761 0 1 12004
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_9
timestamp 1704896540
transform 1 0 2714 0 1 12004
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_10
timestamp 1704896540
transform 1 0 1752 0 1 12004
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_11
timestamp 1704896540
transform 1 0 5472 0 1 12004
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_12
timestamp 1704896540
transform 1 0 7257 0 1 12004
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_13
timestamp 1704896540
transform 1 0 8271 0 1 12004
box 0 0 1 1
use M1M2_CDNS_52468879185201  M1M2_CDNS_52468879185201_0
timestamp 1704896540
transform 0 -1 7683 1 0 13135
box 0 0 320 116
use M1M2_CDNS_52468879185201  M1M2_CDNS_52468879185201_1
timestamp 1704896540
transform 0 -1 3884 1 0 1746
box 0 0 320 116
use M1M2_CDNS_52468879185201  M1M2_CDNS_52468879185201_2
timestamp 1704896540
transform 0 -1 4047 1 0 1247
box 0 0 320 116
use M1M2_CDNS_52468879185201  M1M2_CDNS_52468879185201_3
timestamp 1704896540
transform 0 -1 7382 1 0 1746
box 0 0 320 116
use M1M2_CDNS_52468879185201  M1M2_CDNS_52468879185201_4
timestamp 1704896540
transform 0 -1 5638 1 0 1746
box 0 0 320 116
use M1M2_CDNS_52468879185201  M1M2_CDNS_52468879185201_5
timestamp 1704896540
transform 0 -1 5638 1 0 1286
box 0 0 320 116
use M1M2_CDNS_52468879185201  M1M2_CDNS_52468879185201_6
timestamp 1704896540
transform 0 -1 3886 1 0 1286
box 0 0 320 116
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_0
timestamp 1704896540
transform 0 1 9452 1 0 13135
box 0 0 1 1
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_1
timestamp 1704896540
transform 0 1 9764 1 0 13135
box 0 0 1 1
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_2
timestamp 1704896540
transform 0 -1 10245 1 0 1746
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_0
timestamp 1704896540
transform 0 -1 10245 -1 0 6825
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_1
timestamp 1704896540
transform 0 -1 10245 -1 0 5644
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_2
timestamp 1704896540
transform 0 -1 10245 -1 0 7347
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_3
timestamp 1704896540
transform 1 0 4807 0 1 12951
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_4
timestamp 1704896540
transform 1 0 3969 0 1 12951
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_5
timestamp 1704896540
transform 1 0 6647 0 1 12951
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_6
timestamp 1704896540
transform 1 0 6924 0 1 12951
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_7
timestamp 1704896540
transform 1 0 4904 0 1 3324
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_8
timestamp 1704896540
transform 1 0 6786 0 1 3324
box 0 0 1 1
use M1M2_CDNS_52468879185297  M1M2_CDNS_52468879185297_0
timestamp 1704896540
transform 0 1 7516 1 0 11029
box 0 0 1 1
use M1M2_CDNS_52468879185297  M1M2_CDNS_52468879185297_1
timestamp 1704896540
transform 1 0 2977 0 1 7532
box 0 0 1 1
use M1M2_CDNS_52468879185297  M1M2_CDNS_52468879185297_2
timestamp 1704896540
transform 1 0 8658 0 1 7424
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_0
timestamp 1704896540
transform -1 0 3135 0 1 652
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_1
timestamp 1704896540
transform -1 0 2623 0 1 652
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_2
timestamp 1704896540
transform -1 0 2879 0 1 508
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_3
timestamp 1704896540
transform -1 0 2367 0 1 508
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_4
timestamp 1704896540
transform 0 -1 7878 1 0 527
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_5
timestamp 1704896540
transform 1 0 8781 0 1 508
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_6
timestamp 1704896540
transform 1 0 8269 0 1 508
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_7
timestamp 1704896540
transform 1 0 8525 0 1 652
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_8
timestamp 1704896540
transform 1 0 8013 0 1 652
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_9
timestamp 1704896540
transform 1 0 9193 0 1 508
box 0 0 1 1
use M1M2_CDNS_52468879185967  M1M2_CDNS_52468879185967_0
timestamp 1704896540
transform 1 0 9413 0 1 12004
box 0 0 448 116
use M1M2_CDNS_524688791851077  M1M2_CDNS_524688791851077_0
timestamp 1704896540
transform 0 -1 6975 1 0 1746
box 0 0 320 180
use M1M2_CDNS_524688791851078  M1M2_CDNS_524688791851078_0
timestamp 1704896540
transform -1 0 8771 0 -1 1813
box 0 0 576 52
use M1M2_CDNS_524688791851078  M1M2_CDNS_524688791851078_1
timestamp 1704896540
transform -1 0 2968 0 -1 1813
box 0 0 576 52
use M1M2_CDNS_524688791851081  M1M2_CDNS_524688791851081_0
timestamp 1704896540
transform -1 0 6611 0 1 537
box 0 0 256 180
use M1M2_CDNS_524688791851081  M1M2_CDNS_524688791851081_1
timestamp 1704896540
transform 1 0 4884 0 1 537
box 0 0 256 180
use M1M2_CDNS_524688791851446  M1M2_CDNS_524688791851446_0
timestamp 1704896540
transform -1 0 11204 0 1 12004
box 0 0 704 116
use nfet_CDNS_524688791851024  nfet_CDNS_524688791851024_0
timestamp 1704896540
transform 0 1 5994 -1 0 1533
box -79 -52 535 1052
use nfet_CDNS_524688791851024  nfet_CDNS_524688791851024_1
timestamp 1704896540
transform 0 1 5994 -1 0 2045
box -79 -52 535 1052
use nfet_CDNS_524688791851024  nfet_CDNS_524688791851024_2
timestamp 1704896540
transform 0 1 5994 -1 0 2557
box -79 -52 535 1052
use nfet_CDNS_524688791851025  nfet_CDNS_524688791851025_0
timestamp 1704896540
transform 0 1 4154 -1 0 11201
box -79 -52 179 1052
use nfet_CDNS_524688791851025  nfet_CDNS_524688791851025_1
timestamp 1704896540
transform 0 1 4154 -1 0 4197
box -79 -52 179 1052
use nfet_CDNS_524688791851025  nfet_CDNS_524688791851025_2
timestamp 1704896540
transform 0 1 5994 -1 0 4197
box -79 -52 179 1052
use nfet_CDNS_524688791851025  nfet_CDNS_524688791851025_3
timestamp 1704896540
transform 0 1 5994 -1 0 11201
box -79 -52 179 1052
use nfet_CDNS_524688791851623  nfet_CDNS_524688791851623_0
timestamp 1704896540
transform -1 0 1783 0 1 554
box -79 -26 279 226
use nfet_CDNS_524688791851624  nfet_CDNS_524688791851624_0
timestamp 1704896540
transform 0 1 7680 -1 0 1759
box -79 -26 879 2026
use nfet_CDNS_524688791851624  nfet_CDNS_524688791851624_1
timestamp 1704896540
transform 0 1 1468 1 0 959
box -79 -26 879 2026
use nfet_CDNS_524688791851625  nfet_CDNS_524688791851625_0
timestamp 1704896540
transform 0 -1 5672 1 0 2671
box -79 -26 495 226
use nfet_CDNS_524688791851626  nfet_CDNS_524688791851626_0
timestamp 1704896540
transform 0 1 5994 -1 0 1021
box -79 -52 179 1052
use nfet_CDNS_524688791851626  nfet_CDNS_524688791851626_1
timestamp 1704896540
transform 0 1 4154 1 0 921
box -79 -52 179 1052
use nfet_CDNS_524688791851627  nfet_CDNS_524688791851627_0
timestamp 1704896540
transform 0 1 5994 -1 0 3325
box -79 -52 279 1052
use nfet_CDNS_524688791851627  nfet_CDNS_524688791851627_1
timestamp 1704896540
transform 0 1 4154 -1 0 3325
box -79 -52 279 1052
use nfet_CDNS_524688791851628  nfet_CDNS_524688791851628_0
timestamp 1704896540
transform 0 1 4154 -1 0 1533
box -79 -52 535 1052
use nfet_CDNS_524688791851628  nfet_CDNS_524688791851628_1
timestamp 1704896540
transform 0 1 4154 -1 0 2557
box -79 -52 535 1052
use nfet_CDNS_524688791851628  nfet_CDNS_524688791851628_2
timestamp 1704896540
transform 0 1 4154 -1 0 2045
box -79 -52 535 1052
use nfet_CDNS_524688791851628  nfet_CDNS_524688791851628_3
timestamp 1704896540
transform 0 1 4154 1 0 2613
box -79 -52 535 1052
use nfet_CDNS_524688791851629  nfet_CDNS_524688791851629_0
timestamp 1704896540
transform 0 1 1468 1 0 7412
box -226 -26 1026 2026
use nfet_CDNS_524688791851629  nfet_CDNS_524688791851629_1
timestamp 1704896540
transform 0 1 1468 1 0 2652
box -226 -26 1026 2026
use nfet_CDNS_524688791851629  nfet_CDNS_524688791851629_2
timestamp 1704896540
transform 0 1 1468 1 0 10440
box -226 -26 1026 2026
use nfet_CDNS_524688791851629  nfet_CDNS_524688791851629_3
timestamp 1704896540
transform 0 1 1468 1 0 5680
box -226 -26 1026 2026
use nfet_CDNS_524688791851629  nfet_CDNS_524688791851629_4
timestamp 1704896540
transform 0 -1 9680 1 0 2652
box -226 -26 1026 2026
use nfet_CDNS_524688791851629  nfet_CDNS_524688791851629_5
timestamp 1704896540
transform 0 -1 9680 1 0 7412
box -226 -26 1026 2026
use nfet_CDNS_524688791851629  nfet_CDNS_524688791851629_6
timestamp 1704896540
transform 0 -1 9680 1 0 10440
box -226 -26 1026 2026
use nfet_CDNS_524688791851629  nfet_CDNS_524688791851629_7
timestamp 1704896540
transform 0 -1 9680 1 0 5680
box -226 -26 1026 2026
use nfet_CDNS_524688791851630  nfet_CDNS_524688791851630_0
timestamp 1704896540
transform 0 1 1468 1 0 8498
box -226 -26 1882 2026
use nfet_CDNS_524688791851630  nfet_CDNS_524688791851630_1
timestamp 1704896540
transform 0 1 1468 1 0 3738
box -226 -26 1882 2026
use nfet_CDNS_524688791851630  nfet_CDNS_524688791851630_2
timestamp 1704896540
transform 0 -1 9680 1 0 8498
box -226 -26 1882 2026
use nfet_CDNS_524688791851630  nfet_CDNS_524688791851630_3
timestamp 1704896540
transform 0 -1 9680 1 0 3738
box -226 -26 1882 2026
use nfet_CDNS_524688791851631  nfet_CDNS_524688791851631_0
timestamp 1704896540
transform 0 1 5994 -1 0 5909
box -79 -52 879 1052
use nfet_CDNS_524688791851631  nfet_CDNS_524688791851631_1
timestamp 1704896540
transform 0 1 5994 -1 0 7621
box -79 -52 879 1052
use nfet_CDNS_524688791851631  nfet_CDNS_524688791851631_2
timestamp 1704896540
transform 0 1 5994 -1 0 9333
box -79 -52 879 1052
use nfet_CDNS_524688791851631  nfet_CDNS_524688791851631_3
timestamp 1704896540
transform 0 1 5994 -1 0 11045
box -79 -52 879 1052
use nfet_CDNS_524688791851631  nfet_CDNS_524688791851631_4
timestamp 1704896540
transform 0 1 4154 -1 0 11045
box -79 -52 879 1052
use nfet_CDNS_524688791851631  nfet_CDNS_524688791851631_5
timestamp 1704896540
transform 0 1 4154 -1 0 9333
box -79 -52 879 1052
use nfet_CDNS_524688791851631  nfet_CDNS_524688791851631_6
timestamp 1704896540
transform 0 1 4154 -1 0 7621
box -79 -52 879 1052
use nfet_CDNS_524688791851631  nfet_CDNS_524688791851631_7
timestamp 1704896540
transform 0 1 4154 -1 0 5909
box -79 -52 879 1052
use nfet_CDNS_524688791851631  nfet_CDNS_524688791851631_8
timestamp 1704896540
transform 0 1 5994 1 0 7677
box -79 -52 879 1052
use nfet_CDNS_524688791851631  nfet_CDNS_524688791851631_9
timestamp 1704896540
transform 0 1 5994 1 0 5965
box -79 -52 879 1052
use nfet_CDNS_524688791851631  nfet_CDNS_524688791851631_10
timestamp 1704896540
transform 0 1 5994 1 0 9389
box -79 -52 879 1052
use nfet_CDNS_524688791851631  nfet_CDNS_524688791851631_11
timestamp 1704896540
transform 0 1 5994 1 0 4253
box -79 -52 879 1052
use nfet_CDNS_524688791851631  nfet_CDNS_524688791851631_12
timestamp 1704896540
transform 0 1 4154 1 0 4253
box -79 -52 879 1052
use nfet_CDNS_524688791851631  nfet_CDNS_524688791851631_13
timestamp 1704896540
transform 0 1 4154 1 0 9389
box -79 -52 879 1052
use nfet_CDNS_524688791851631  nfet_CDNS_524688791851631_14
timestamp 1704896540
transform 0 1 4154 1 0 5965
box -79 -52 879 1052
use nfet_CDNS_524688791851631  nfet_CDNS_524688791851631_15
timestamp 1704896540
transform 0 1 4154 1 0 7677
box -79 -52 879 1052
use nfet_CDNS_524688791851632  nfet_CDNS_524688791851632_0
timestamp 1704896540
transform 0 1 5994 1 0 2613
box -79 -52 535 1052
use nfet_CDNS_524688791851633  nfet_CDNS_524688791851633_0
timestamp 1704896540
transform 0 1 4154 -1 0 755
box -79 -26 335 1026
use nfet_CDNS_524688791851633  nfet_CDNS_524688791851633_1
timestamp 1704896540
transform 0 1 5994 -1 0 755
box -79 -26 335 1026
use nfet_CDNS_524688791851634  nfet_CDNS_524688791851634_0
timestamp 1704896540
transform -1 0 8275 0 1 578
box -79 -52 279 202
use nfet_CDNS_524688791851634  nfet_CDNS_524688791851634_1
timestamp 1704896540
transform -1 0 2817 0 1 578
box -79 -52 279 202
use nfet_CDNS_524688791851634  nfet_CDNS_524688791851634_2
timestamp 1704896540
transform -1 0 3329 0 1 578
box -79 -52 279 202
use nfet_CDNS_524688791851634  nfet_CDNS_524688791851634_3
timestamp 1704896540
transform -1 0 8787 0 1 578
box -79 -52 279 202
use nfet_CDNS_524688791851634  nfet_CDNS_524688791851634_4
timestamp 1704896540
transform -1 0 2305 0 1 578
box -79 -52 279 202
use nfet_CDNS_524688791851634  nfet_CDNS_524688791851634_5
timestamp 1704896540
transform 1 0 7819 0 1 578
box -79 -52 279 202
use nfet_CDNS_524688791851634  nfet_CDNS_524688791851634_6
timestamp 1704896540
transform 1 0 8331 0 1 578
box -79 -52 279 202
use nfet_CDNS_524688791851634  nfet_CDNS_524688791851634_7
timestamp 1704896540
transform 1 0 2873 0 1 578
box -79 -52 279 202
use nfet_CDNS_524688791851634  nfet_CDNS_524688791851634_8
timestamp 1704896540
transform 1 0 2361 0 1 578
box -79 -52 279 202
use nfet_CDNS_524688791851634  nfet_CDNS_524688791851634_9
timestamp 1704896540
transform 1 0 8843 0 1 578
box -79 -52 279 202
use nfet_CDNS_524688791851635  nfet_CDNS_524688791851635_0
timestamp 1704896540
transform -1 0 9199 0 1 578
box -79 -52 179 202
use nfet_CDNS_524688791851635  nfet_CDNS_524688791851635_1
timestamp 1704896540
transform -1 0 7763 0 1 578
box -79 -52 179 202
use nfet_CDNS_524688791851635  nfet_CDNS_524688791851635_2
timestamp 1704896540
transform 1 0 3385 0 1 578
box -79 -52 179 202
use nfet_CDNS_524688791851635  nfet_CDNS_524688791851635_3
timestamp 1704896540
transform 1 0 1949 0 1 578
box -79 -52 179 202
use pfet_CDNS_524688791851636  pfet_CDNS_524688791851636_0
timestamp 1704896540
transform -1 0 1602 0 1 12506
box -119 -66 319 666
use pfet_CDNS_524688791851637  pfet_CDNS_524688791851637_0
timestamp 1704896540
transform -1 0 9762 0 -1 13839
box -119 -66 375 1066
use pfet_CDNS_524688791851638  pfet_CDNS_524688791851638_0
timestamp 1704896540
transform 0 1 1839 1 0 12493
box -119 -66 1719 1466
use pfet_CDNS_524688791851639  pfet_CDNS_524688791851639_0
timestamp 1704896540
transform 0 -1 9243 1 0 12493
box -119 -66 1719 1466
use pfet_CDNS_524688791851640  pfet_CDNS_524688791851640_0
timestamp 1704896540
transform -1 0 5603 0 -1 12656
box -119 -66 219 216
use pfet_CDNS_524688791851641  pfet_CDNS_524688791851641_0
timestamp 1704896540
transform 0 -1 4089 -1 0 13779
box -119 -66 319 666
use pfet_CDNS_524688791851641  pfet_CDNS_524688791851641_1
timestamp 1704896540
transform 0 -1 4089 -1 0 13267
box -119 -66 319 666
use pfet_CDNS_524688791851641  pfet_CDNS_524688791851641_2
timestamp 1704896540
transform 0 -1 7605 -1 0 13267
box -119 -66 319 666
use pfet_CDNS_524688791851641  pfet_CDNS_524688791851641_3
timestamp 1704896540
transform 0 -1 7605 -1 0 13779
box -119 -66 319 666
use pfet_CDNS_524688791851641  pfet_CDNS_524688791851641_4
timestamp 1704896540
transform 0 1 4327 -1 0 13361
box -119 -66 319 666
use pfet_CDNS_524688791851641  pfet_CDNS_524688791851641_5
timestamp 1704896540
transform 0 1 4327 -1 0 12849
box -119 -66 319 666
use pfet_CDNS_524688791851641  pfet_CDNS_524688791851641_6
timestamp 1704896540
transform 0 1 4327 -1 0 13873
box -119 -66 319 666
use pfet_CDNS_524688791851641  pfet_CDNS_524688791851641_7
timestamp 1704896540
transform 0 1 6167 -1 0 13873
box -119 -66 319 666
use pfet_CDNS_524688791851641  pfet_CDNS_524688791851641_8
timestamp 1704896540
transform 0 1 6167 -1 0 12849
box -119 -66 319 666
use pfet_CDNS_524688791851641  pfet_CDNS_524688791851641_9
timestamp 1704896540
transform 0 1 6167 -1 0 13361
box -119 -66 319 666
use pfet_CDNS_524688791851641  pfet_CDNS_524688791851641_10
timestamp 1704896540
transform 0 -1 4089 1 0 13323
box -119 -66 319 666
use pfet_CDNS_524688791851641  pfet_CDNS_524688791851641_11
timestamp 1704896540
transform 0 -1 4089 1 0 12811
box -119 -66 319 666
use pfet_CDNS_524688791851641  pfet_CDNS_524688791851641_12
timestamp 1704896540
transform 0 -1 7605 1 0 12811
box -119 -66 319 666
use pfet_CDNS_524688791851641  pfet_CDNS_524688791851641_13
timestamp 1704896540
transform 0 -1 7605 1 0 13323
box -119 -66 319 666
use pfet_CDNS_524688791851642  pfet_CDNS_524688791851642_0
timestamp 1704896540
transform 0 1 4327 1 0 13417
box -119 -66 319 666
use pfet_CDNS_524688791851642  pfet_CDNS_524688791851642_1
timestamp 1704896540
transform 0 1 4327 1 0 12905
box -119 -66 319 666
use pfet_CDNS_524688791851642  pfet_CDNS_524688791851642_2
timestamp 1704896540
transform 0 1 6167 1 0 12905
box -119 -66 319 666
use pfet_CDNS_524688791851642  pfet_CDNS_524688791851642_3
timestamp 1704896540
transform 0 1 6167 1 0 13417
box -119 -66 319 666
use pfet_CDNS_524688791851643  pfet_CDNS_524688791851643_0
timestamp 1704896540
transform 0 1 4327 1 0 12493
box -119 -66 219 666
use pfet_CDNS_524688791851643  pfet_CDNS_524688791851643_1
timestamp 1704896540
transform 0 1 4327 1 0 13929
box -119 -66 219 666
use pfet_CDNS_524688791851643  pfet_CDNS_524688791851643_2
timestamp 1704896540
transform 0 1 6167 1 0 13929
box -119 -66 219 666
use pfet_CDNS_524688791851643  pfet_CDNS_524688791851643_3
timestamp 1704896540
transform 0 1 6167 1 0 12493
box -119 -66 219 666
use pfet_CDNS_524688791851643  pfet_CDNS_524688791851643_4
timestamp 1704896540
transform 0 -1 4089 1 0 13835
box -119 -66 219 666
use pfet_CDNS_524688791851643  pfet_CDNS_524688791851643_5
timestamp 1704896540
transform 0 -1 4089 1 0 12655
box -119 -66 219 666
use pfet_CDNS_524688791851643  pfet_CDNS_524688791851643_6
timestamp 1704896540
transform 0 -1 7605 1 0 12655
box -119 -66 219 666
use pfet_CDNS_524688791851643  pfet_CDNS_524688791851643_7
timestamp 1704896540
transform 0 -1 7605 1 0 13835
box -119 -66 219 666
use pfet_CDNS_524688791851644  pfet_CDNS_524688791851644_0
timestamp 1704896540
transform 1 0 5269 0 1 12839
box -119 -66 687 1066
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_0
timestamp 1704896540
transform 0 1 5486 -1 0 12474
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_1
timestamp 1704896540
transform -1 0 4295 0 1 13929
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_2
timestamp 1704896540
transform -1 0 3457 0 1 13835
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_3
timestamp 1704896540
transform -1 0 6973 0 1 13835
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_4
timestamp 1704896540
transform -1 0 6135 0 1 13929
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_5
timestamp 1704896540
transform -1 0 4295 0 -1 12593
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_6
timestamp 1704896540
transform 1 0 7016 0 -1 1021
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_7
timestamp 1704896540
transform 1 0 5178 0 -1 1021
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_8
timestamp 1704896540
transform 1 0 4959 0 -1 12593
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_9
timestamp 1704896540
transform 1 0 6799 0 -1 12593
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_10
timestamp 1704896540
transform 1 0 5696 0 -1 3064
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_11
timestamp 1704896540
transform 1 0 5178 0 1 1110
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_12
timestamp 1704896540
transform 1 0 5178 0 1 1366
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_13
timestamp 1704896540
transform 1 0 5178 0 1 1878
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_14
timestamp 1704896540
transform 1 0 5178 0 1 1622
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_15
timestamp 1704896540
transform 1 0 5178 0 1 2390
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_16
timestamp 1704896540
transform 1 0 5178 0 1 2134
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_17
timestamp 1704896540
transform 1 0 5178 0 1 2646
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_18
timestamp 1704896540
transform 1 0 7016 0 1 2902
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_19
timestamp 1704896540
transform 1 0 5178 0 1 2902
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_20
timestamp 1704896540
transform 1 0 7016 0 1 2646
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_21
timestamp 1704896540
transform 1 0 7016 0 1 2134
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_22
timestamp 1704896540
transform 1 0 7016 0 1 2390
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_23
timestamp 1704896540
transform 1 0 7016 0 1 1622
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_24
timestamp 1704896540
transform 1 0 7016 0 1 1878
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_25
timestamp 1704896540
transform 1 0 7016 0 1 1366
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_26
timestamp 1704896540
transform 1 0 7016 0 1 1110
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_27
timestamp 1704896540
transform 1 0 4959 0 1 13929
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_28
timestamp 1704896540
transform 1 0 4121 0 1 13835
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_29
timestamp 1704896540
transform 1 0 7637 0 1 13835
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_0
timestamp 1704896540
transform -1 0 7082 0 -1 728
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_1
timestamp 1704896540
transform -1 0 5242 0 -1 728
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_2
timestamp 1704896540
transform 1 0 5178 0 1 3125
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_3
timestamp 1704896540
transform 1 0 7016 0 1 3125
box 0 0 1 1
use sky130_fd_io__sio_opamp_stage_c_c_res  sky130_fd_io__sio_opamp_stage_c_c_res_0
timestamp 1704896540
transform 1 0 10212 0 1 538
box 82 4 1354 3524
use sky130_fd_io__sio_opamp_stage_c_c_res  sky130_fd_io__sio_opamp_stage_c_c_res_1
timestamp 1704896540
transform 1 0 10212 0 1 4092
box 82 4 1354 3524
use sky130_fd_io__sio_opamp_stage_c_c_res  sky130_fd_io__sio_opamp_stage_c_c_res_2
timestamp 1704896540
transform 1 0 11492 0 1 4092
box 82 4 1354 3524
use sky130_fd_io__sio_opamp_stage_c_c_res  sky130_fd_io__sio_opamp_stage_c_c_res_3
timestamp 1704896540
transform 1 0 11492 0 1 538
box 82 4 1354 3524
use sky130_fd_io__tk_em1o_CDNS_52468879185315  sky130_fd_io__tk_em1o_CDNS_52468879185315_0
timestamp 1704896540
transform -1 0 7921 0 1 12951
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185315  sky130_fd_io__tk_em1o_CDNS_52468879185315_1
timestamp 1704896540
transform 1 0 3162 0 1 12951
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185338  sky130_fd_io__tk_em1o_CDNS_52468879185338_0
timestamp 1704896540
transform -1 0 9215 0 1 1063
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185340  sky130_fd_io__tk_em1o_CDNS_52468879185340_0
timestamp 1704896540
transform -1 0 4861 0 1 3930
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185340  sky130_fd_io__tk_em1o_CDNS_52468879185340_1
timestamp 1704896540
transform -1 0 6698 0 1 3930
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185340  sky130_fd_io__tk_em1o_CDNS_52468879185340_2
timestamp 1704896540
transform 1 0 4401 0 1 3930
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185340  sky130_fd_io__tk_em1o_CDNS_52468879185340_3
timestamp 1704896540
transform 1 0 6247 0 1 3930
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_0
timestamp 1704896540
transform 0 1 5973 1 0 2513
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_1
timestamp 1704896540
transform 0 -1 4191 1 0 2512
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_524688791851620  sky130_fd_io__tk_em1o_CDNS_524688791851620_0
timestamp 1704896540
transform 1 0 1932 0 -1 1191
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185314  sky130_fd_io__tk_em1s_CDNS_52468879185314_0
timestamp 1704896540
transform -1 0 3304 0 1 13962
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185314  sky130_fd_io__tk_em1s_CDNS_52468879185314_1
timestamp 1704896540
transform 1 0 7809 0 1 13962
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_524688791851189  sky130_fd_io__tk_em1s_CDNS_524688791851189_0
timestamp 1704896540
transform -1 0 8167 0 1 1063
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_524688791851189  sky130_fd_io__tk_em1s_CDNS_524688791851189_1
timestamp 1704896540
transform 1 0 2981 0 1 1063
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_524688791851621  sky130_fd_io__tk_em1s_CDNS_524688791851621_0
timestamp 1704896540
transform -1 0 4020 0 1 3930
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_524688791851621  sky130_fd_io__tk_em1s_CDNS_524688791851621_1
timestamp 1704896540
transform -1 0 5412 0 1 3930
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_524688791851621  sky130_fd_io__tk_em1s_CDNS_524688791851621_2
timestamp 1704896540
transform -1 0 7273 0 1 3930
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_524688791851621  sky130_fd_io__tk_em1s_CDNS_524688791851621_3
timestamp 1704896540
transform 1 0 5736 0 1 3930
box 0 0 1 1
<< labels >>
flabel comment s 11566 7812 11566 7812 0 FreeSans 1000 0 0 0 condiode
flabel comment s 8702 6760 8702 6760 0 FreeSans 1000 0 0 0 condiode
flabel comment s 8685 11520 8685 11520 0 FreeSans 1000 0 0 0 condiode
flabel comment s 6531 11491 6531 11491 0 FreeSans 1000 0 0 0 condiode
flabel comment s 4609 11481 4609 11481 0 FreeSans 1000 0 0 0 condiode
flabel comment s 2470 1650 2470 1650 0 FreeSans 1000 0 0 0 condiode
flabel comment s 2420 6756 2420 6756 0 FreeSans 1000 0 0 0 condiode
flabel comment s 2317 11520 2317 11520 0 FreeSans 1000 0 0 0 condiode
flabel comment s 13234 12648 13234 12648 3 FreeSans 200 180 0 0 vnb
flabel comment s 5950 -130 5950 -130 3 FreeSans 200 180 0 0 pad
flabel comment s 1142 -130 1142 -130 3 FreeSans 200 0 0 0 pad
flabel comment s 12991 6054 12991 6054 3 FreeSans 200 180 0 0 oe_hs_h
flabel comment s 12991 5964 12991 5964 3 FreeSans 200 180 0 0 od_h
flabel comment s 1236 6054 1236 6054 3 FreeSans 200 0 0 0 oe_hs_h
flabel comment s 1236 5964 1236 5964 3 FreeSans 200 0 0 0 od_h
flabel comment s 12985 3067 12985 3067 3 FreeSans 200 180 0 0 vgnd_io
flabel comment s 11143 14255 11143 14255 3 FreeSans 200 180 0 0 vpwr_ka
flabel comment s 1254 14279 1254 14279 3 FreeSans 200 0 0 0 vpwr_ka
flabel comment s 1132 496 1132 496 3 FreeSans 200 0 0 0 pu_h_n<1>
flabel comment s 3447 688 3447 688 0 FreeSans 1000 0 0 0 500
flabel comment s 4622 1304 4622 1304 0 FreeSans 1000 0 0 0 7
flabel comment s 4622 1809 4622 1809 0 FreeSans 1000 0 0 0 6
flabel comment s 4622 2322 4622 2322 0 FreeSans 1000 0 0 0 5
flabel comment s 4622 2832 4622 2832 0 FreeSans 1000 0 0 0 4
flabel comment s 9164 583 9164 583 0 FreeSans 1000 180 0 0 D
flabel comment s 7701 677 7701 677 0 FreeSans 1000 180 0 0 501
flabel comment s 9164 685 9164 685 0 FreeSans 1000 180 0 0 15
flabel comment s 7927 647 7927 647 0 FreeSans 1000 180 0 0 9
flabel comment s 8192 645 8192 645 0 FreeSans 1000 180 0 0 8
flabel comment s 8462 652 8462 652 0 FreeSans 1000 180 0 0 7
flabel comment s 8709 647 8709 647 0 FreeSans 1000 180 0 0 6
flabel comment s 8974 647 8974 647 0 FreeSans 1000 180 0 0 5
flabel comment s 1984 568 1984 568 0 FreeSans 1000 0 0 0 D
flabel comment s 2174 647 2174 647 0 FreeSans 1000 0 0 0 14
flabel comment s 2439 647 2439 647 0 FreeSans 1000 0 0 0 13
flabel comment s 2686 652 2686 652 0 FreeSans 1000 0 0 0 12
flabel comment s 2956 645 2956 645 0 FreeSans 1000 0 0 0 11
flabel comment s 3221 647 3221 647 0 FreeSans 1000 0 0 0 10
flabel comment s 1132 418 1132 418 3 FreeSans 200 0 0 0 pu_h_n<0>
flabel comment s 6476 12565 6476 12565 0 FreeSans 1000 0 0 0 503 (D)
flabel comment s 6482 14014 6482 14014 0 FreeSans 1000 0 0 0 511
flabel comment s 6476 13552 6476 13552 0 FreeSans 1000 0 0 0 25 (D)
flabel comment s 6443 13009 6443 13009 0 FreeSans 1000 0 0 0 24 (D)
flabel comment s 6497 12737 6497 12737 0 FreeSans 1000 0 0 0 14
flabel comment s 6491 13263 6491 13263 0 FreeSans 1000 0 0 0 13
flabel comment s 6485 13767 6485 13767 0 FreeSans 1000 0 0 0 12
flabel comment s 7290 12703 7290 12703 0 FreeSans 1000 0 0 0 463 (D)
flabel comment s 7290 13913 7290 13913 0 FreeSans 1000 0 0 0 513
flabel comment s 7372 12907 7372 12907 0 FreeSans 1000 0 0 0 08
flabel comment s 7364 13169 7364 13169 0 FreeSans 1000 0 0 0 09
flabel comment s 7378 13417 7378 13417 0 FreeSans 1000 0 0 0 10
flabel comment s 7367 13676 7367 13676 0 FreeSans 1000 0 0 0 11
flabel comment s 1984 685 1984 685 0 FreeSans 1000 0 0 0 16
flabel comment s 3792 13676 3792 13676 0 FreeSans 1000 0 0 0 21
flabel comment s 3803 13417 3803 13417 0 FreeSans 1000 0 0 0 20
flabel comment s 3789 13169 3789 13169 0 FreeSans 1000 0 0 0 19
flabel comment s 3797 12907 3797 12907 0 FreeSans 1000 0 0 0 18
flabel comment s 4614 13767 4614 13767 0 FreeSans 1000 0 0 0 17
flabel comment s 4620 13263 4620 13263 0 FreeSans 1000 0 0 0 16
flabel comment s 4626 12737 4626 12737 0 FreeSans 1000 0 0 0 15
flabel comment s 3715 13913 3715 13913 0 FreeSans 1000 0 0 0 462.1 (D)
flabel comment s 3802 12698 3802 12698 0 FreeSans 1000 0 0 0 462.3 (D)
flabel comment s 4605 12565 4605 12565 0 FreeSans 1000 0 0 0 502 (D)
flabel comment s 4572 13009 4572 13009 0 FreeSans 1000 0 0 0 22 (D)
flabel comment s 4605 13552 4605 13552 0 FreeSans 1000 0 0 0 23 (D)
flabel comment s 4654 13985 4654 13985 0 FreeSans 1000 0 0 0 462.2 (D)
flabel comment s 4584 11166 4584 11166 0 FreeSans 1000 0 0 0 dummy
flabel comment s 6529 11154 6529 11154 0 FreeSans 1000 0 0 0 dummy
flabel comment s 4532 4171 4532 4171 0 FreeSans 1000 0 0 0 dummy
flabel comment s 6517 4158 6517 4158 0 FreeSans 1000 0 0 0 dummy
flabel comment s 6440 4894 6440 4894 0 FreeSans 1600 90 0 0 vsource_0
flabel comment s 7050 4410 7050 4410 0 FreeSans 1600 90 0 0 inp
flabel comment s 5944 4371 5944 4371 0 FreeSans 1600 270 0 0 inn
flabel comment s 12993 281 12993 281 3 FreeSans 200 180 0 0 pu_h_n<0>
flabel comment s 12993 359 12993 359 3 FreeSans 200 180 0 0 pu_h_n<1>
flabel comment s 4638 984 4638 984 0 FreeSans 1000 0 0 0 466 (D)
flabel comment s 4622 3256 4622 3256 0 FreeSans 1000 0 0 0 492 (D)
flabel comment s 4313 4371 4313 4371 0 FreeSans 1600 270 0 0 inn
flabel comment s 5152 4410 5152 4410 0 FreeSans 1600 90 0 0 inp
flabel comment s 4600 4894 4600 4894 0 FreeSans 1600 90 0 0 vsource_1
flabel comment s 6488 3243 6488 3243 0 FreeSans 1000 0 0 0 dummy
flabel comment s 6549 988 6549 988 0 FreeSans 1000 0 0 0 dummy
flabel comment s 9826 10624 9826 10624 3 FreeSans 200 180 0 0 puen_reg_h
flabel comment s 1245 10763 1245 10763 3 FreeSans 200 0 0 0 puen_reg_h
flabel comment s 1235 9152 1235 9152 3 FreeSans 200 0 0 0 slow_h_n
flabel comment s 9826 9152 9826 9152 3 FreeSans 200 180 0 0 slow_h_n
flabel comment s 1227 12855 1227 12855 3 FreeSans 200 0 0 0 drvhi_h
flabel comment s 11158 12851 11158 12851 3 FreeSans 200 180 0 0 drvhi_h
flabel metal1 s 6465 5840 6465 5840 0 FreeSans 1000 90 0 0 vsource_0
flabel metal1 s 4639 5845 4639 5845 0 FreeSans 1000 90 0 0 vsource_1
flabel metal1 s 2097 2442 2097 2442 0 FreeSans 1000 90 0 0 pd_1
flabel metal1 s 9035 2425 9035 2425 0 FreeSans 1000 90 0 0 pd_0
flabel metal1 s 4922 6698 4922 6698 0 FreeSans 1000 90 0 0 pu_1
flabel metal1 s 6808 6692 6808 6692 0 FreeSans 1000 90 0 0 pu_0
flabel metal1 s 1313 7105 1313 7105 0 FreeSans 1000 90 0 0 en_hicc_n
flabel metal1 s 7585 775 7623 856 0 FreeSans 200 0 0 0 vreg_en_h_n
port 2 nsew
flabel metal1 s 7684 1901 7814 2031 0 FreeSans 1000 90 0 0 out
port 3 nsew
flabel metal1 s 1191 12340 1237 12765 0 FreeSans 1000 90 0 0 vpp
port 4 nsew
flabel metal2 s 13182 12356 13266 12486 0 FreeSans 200 0 0 0 ngate
port 5 nsew
flabel metal2 s 13182 12170 13266 12300 0 FreeSans 200 0 0 0 inp
port 6 nsew
flabel metal2 s 1179 11409 1225 11842 0 FreeSans 1000 90 0 0 vpp
port 4 nsew
flabel metal2 s 1117 5452 1179 5644 0 FreeSans 200 0 0 0 vgnd
port 7 nsew
flabel metal2 s 1117 4017 1179 4209 0 FreeSans 200 0 0 0 vgnd
port 7 nsew
flabel metal2 s 2342 1247 2625 1623 0 FreeSans 1000 90 0 0 vgnd
port 7 nsew
flabel metal2 s 1604 13505 1717 13841 0 FreeSans 1000 90 0 0 vcc
port 8 nsew
flabel metal2 s 6130 6940 6192 7019 0 FreeSans 1000 90 0 0 inp
port 6 nsew
flabel metal2 s 4290 5179 4348 5265 0 FreeSans 1000 90 0 0 inn
port 9 nsew
flabel metal2 s 12797 7640 12868 7770 0 FreeSans 200 0 0 0 out
port 3 nsew
flabel metal2 s 1117 9230 1179 9514 0 FreeSans 200 0 0 0 vgnd
port 7 nsew
flabel metal2 s 1117 10056 1179 10249 0 FreeSans 200 0 0 0 vpp
port 4 nsew
flabel metal2 s 1117 8280 1179 8546 0 FreeSans 200 0 0 0 vgnd
port 7 nsew
flabel metal2 s 1119 545 1164 597 0 FreeSans 200 0 0 0 en_hicc
port 10 nsew
flabel metal2 s 1117 4756 1179 4886 0 FreeSans 200 0 0 0 vpp
port 4 nsew
flabel metal2 s 1117 7959 1179 8152 0 FreeSans 200 0 0 0 vpp
port 4 nsew
flabel metal2 s 1117 7155 1179 7347 0 FreeSans 200 0 0 0 vgnd
port 7 nsew
flabel metal2 s 1117 6633 1179 6825 0 FreeSans 200 0 0 0 vgnd
port 7 nsew
flabel metal2 s 5319 1063 5382 1191 0 FreeSans 200 0 0 0 ngate
port 5 nsew
<< properties >>
string GDS_END 97298950
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 96487786
string path 93.775 91.750 139.775 91.750 
<< end >>
