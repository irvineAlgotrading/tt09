magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< pwell >>
rect 15 163 787 1225
<< nmoslvt >>
rect 171 189 201 1199
rect 257 189 287 1199
rect 343 189 373 1199
rect 429 189 459 1199
rect 515 189 545 1199
rect 601 189 631 1199
<< ndiff >>
rect 111 1187 171 1199
rect 111 1153 126 1187
rect 160 1153 171 1187
rect 111 1119 171 1153
rect 111 1085 126 1119
rect 160 1085 171 1119
rect 111 1051 171 1085
rect 111 1017 126 1051
rect 160 1017 171 1051
rect 111 983 171 1017
rect 111 949 126 983
rect 160 949 171 983
rect 111 915 171 949
rect 111 881 126 915
rect 160 881 171 915
rect 111 847 171 881
rect 111 813 126 847
rect 160 813 171 847
rect 111 779 171 813
rect 111 745 126 779
rect 160 745 171 779
rect 111 711 171 745
rect 111 677 126 711
rect 160 677 171 711
rect 111 643 171 677
rect 111 609 126 643
rect 160 609 171 643
rect 111 575 171 609
rect 111 541 126 575
rect 160 541 171 575
rect 111 507 171 541
rect 111 473 126 507
rect 160 473 171 507
rect 111 439 171 473
rect 111 405 126 439
rect 160 405 171 439
rect 111 371 171 405
rect 111 337 126 371
rect 160 337 171 371
rect 111 303 171 337
rect 111 269 126 303
rect 160 269 171 303
rect 111 235 171 269
rect 111 201 126 235
rect 160 201 171 235
rect 111 189 171 201
rect 201 1187 257 1199
rect 201 1153 212 1187
rect 246 1153 257 1187
rect 201 1119 257 1153
rect 201 1085 212 1119
rect 246 1085 257 1119
rect 201 1051 257 1085
rect 201 1017 212 1051
rect 246 1017 257 1051
rect 201 983 257 1017
rect 201 949 212 983
rect 246 949 257 983
rect 201 915 257 949
rect 201 881 212 915
rect 246 881 257 915
rect 201 847 257 881
rect 201 813 212 847
rect 246 813 257 847
rect 201 779 257 813
rect 201 745 212 779
rect 246 745 257 779
rect 201 711 257 745
rect 201 677 212 711
rect 246 677 257 711
rect 201 643 257 677
rect 201 609 212 643
rect 246 609 257 643
rect 201 575 257 609
rect 201 541 212 575
rect 246 541 257 575
rect 201 507 257 541
rect 201 473 212 507
rect 246 473 257 507
rect 201 439 257 473
rect 201 405 212 439
rect 246 405 257 439
rect 201 371 257 405
rect 201 337 212 371
rect 246 337 257 371
rect 201 303 257 337
rect 201 269 212 303
rect 246 269 257 303
rect 201 235 257 269
rect 201 201 212 235
rect 246 201 257 235
rect 201 189 257 201
rect 287 1187 343 1199
rect 287 1153 298 1187
rect 332 1153 343 1187
rect 287 1119 343 1153
rect 287 1085 298 1119
rect 332 1085 343 1119
rect 287 1051 343 1085
rect 287 1017 298 1051
rect 332 1017 343 1051
rect 287 983 343 1017
rect 287 949 298 983
rect 332 949 343 983
rect 287 915 343 949
rect 287 881 298 915
rect 332 881 343 915
rect 287 847 343 881
rect 287 813 298 847
rect 332 813 343 847
rect 287 779 343 813
rect 287 745 298 779
rect 332 745 343 779
rect 287 711 343 745
rect 287 677 298 711
rect 332 677 343 711
rect 287 643 343 677
rect 287 609 298 643
rect 332 609 343 643
rect 287 575 343 609
rect 287 541 298 575
rect 332 541 343 575
rect 287 507 343 541
rect 287 473 298 507
rect 332 473 343 507
rect 287 439 343 473
rect 287 405 298 439
rect 332 405 343 439
rect 287 371 343 405
rect 287 337 298 371
rect 332 337 343 371
rect 287 303 343 337
rect 287 269 298 303
rect 332 269 343 303
rect 287 235 343 269
rect 287 201 298 235
rect 332 201 343 235
rect 287 189 343 201
rect 373 1187 429 1199
rect 373 1153 384 1187
rect 418 1153 429 1187
rect 373 1119 429 1153
rect 373 1085 384 1119
rect 418 1085 429 1119
rect 373 1051 429 1085
rect 373 1017 384 1051
rect 418 1017 429 1051
rect 373 983 429 1017
rect 373 949 384 983
rect 418 949 429 983
rect 373 915 429 949
rect 373 881 384 915
rect 418 881 429 915
rect 373 847 429 881
rect 373 813 384 847
rect 418 813 429 847
rect 373 779 429 813
rect 373 745 384 779
rect 418 745 429 779
rect 373 711 429 745
rect 373 677 384 711
rect 418 677 429 711
rect 373 643 429 677
rect 373 609 384 643
rect 418 609 429 643
rect 373 575 429 609
rect 373 541 384 575
rect 418 541 429 575
rect 373 507 429 541
rect 373 473 384 507
rect 418 473 429 507
rect 373 439 429 473
rect 373 405 384 439
rect 418 405 429 439
rect 373 371 429 405
rect 373 337 384 371
rect 418 337 429 371
rect 373 303 429 337
rect 373 269 384 303
rect 418 269 429 303
rect 373 235 429 269
rect 373 201 384 235
rect 418 201 429 235
rect 373 189 429 201
rect 459 1187 515 1199
rect 459 1153 470 1187
rect 504 1153 515 1187
rect 459 1119 515 1153
rect 459 1085 470 1119
rect 504 1085 515 1119
rect 459 1051 515 1085
rect 459 1017 470 1051
rect 504 1017 515 1051
rect 459 983 515 1017
rect 459 949 470 983
rect 504 949 515 983
rect 459 915 515 949
rect 459 881 470 915
rect 504 881 515 915
rect 459 847 515 881
rect 459 813 470 847
rect 504 813 515 847
rect 459 779 515 813
rect 459 745 470 779
rect 504 745 515 779
rect 459 711 515 745
rect 459 677 470 711
rect 504 677 515 711
rect 459 643 515 677
rect 459 609 470 643
rect 504 609 515 643
rect 459 575 515 609
rect 459 541 470 575
rect 504 541 515 575
rect 459 507 515 541
rect 459 473 470 507
rect 504 473 515 507
rect 459 439 515 473
rect 459 405 470 439
rect 504 405 515 439
rect 459 371 515 405
rect 459 337 470 371
rect 504 337 515 371
rect 459 303 515 337
rect 459 269 470 303
rect 504 269 515 303
rect 459 235 515 269
rect 459 201 470 235
rect 504 201 515 235
rect 459 189 515 201
rect 545 1187 601 1199
rect 545 1153 556 1187
rect 590 1153 601 1187
rect 545 1119 601 1153
rect 545 1085 556 1119
rect 590 1085 601 1119
rect 545 1051 601 1085
rect 545 1017 556 1051
rect 590 1017 601 1051
rect 545 983 601 1017
rect 545 949 556 983
rect 590 949 601 983
rect 545 915 601 949
rect 545 881 556 915
rect 590 881 601 915
rect 545 847 601 881
rect 545 813 556 847
rect 590 813 601 847
rect 545 779 601 813
rect 545 745 556 779
rect 590 745 601 779
rect 545 711 601 745
rect 545 677 556 711
rect 590 677 601 711
rect 545 643 601 677
rect 545 609 556 643
rect 590 609 601 643
rect 545 575 601 609
rect 545 541 556 575
rect 590 541 601 575
rect 545 507 601 541
rect 545 473 556 507
rect 590 473 601 507
rect 545 439 601 473
rect 545 405 556 439
rect 590 405 601 439
rect 545 371 601 405
rect 545 337 556 371
rect 590 337 601 371
rect 545 303 601 337
rect 545 269 556 303
rect 590 269 601 303
rect 545 235 601 269
rect 545 201 556 235
rect 590 201 601 235
rect 545 189 601 201
rect 631 1187 691 1199
rect 631 1153 642 1187
rect 676 1153 691 1187
rect 631 1119 691 1153
rect 631 1085 642 1119
rect 676 1085 691 1119
rect 631 1051 691 1085
rect 631 1017 642 1051
rect 676 1017 691 1051
rect 631 983 691 1017
rect 631 949 642 983
rect 676 949 691 983
rect 631 915 691 949
rect 631 881 642 915
rect 676 881 691 915
rect 631 847 691 881
rect 631 813 642 847
rect 676 813 691 847
rect 631 779 691 813
rect 631 745 642 779
rect 676 745 691 779
rect 631 711 691 745
rect 631 677 642 711
rect 676 677 691 711
rect 631 643 691 677
rect 631 609 642 643
rect 676 609 691 643
rect 631 575 691 609
rect 631 541 642 575
rect 676 541 691 575
rect 631 507 691 541
rect 631 473 642 507
rect 676 473 691 507
rect 631 439 691 473
rect 631 405 642 439
rect 676 405 691 439
rect 631 371 691 405
rect 631 337 642 371
rect 676 337 691 371
rect 631 303 691 337
rect 631 269 642 303
rect 676 269 691 303
rect 631 235 691 269
rect 631 201 642 235
rect 676 201 691 235
rect 631 189 691 201
<< ndiffc >>
rect 126 1153 160 1187
rect 126 1085 160 1119
rect 126 1017 160 1051
rect 126 949 160 983
rect 126 881 160 915
rect 126 813 160 847
rect 126 745 160 779
rect 126 677 160 711
rect 126 609 160 643
rect 126 541 160 575
rect 126 473 160 507
rect 126 405 160 439
rect 126 337 160 371
rect 126 269 160 303
rect 126 201 160 235
rect 212 1153 246 1187
rect 212 1085 246 1119
rect 212 1017 246 1051
rect 212 949 246 983
rect 212 881 246 915
rect 212 813 246 847
rect 212 745 246 779
rect 212 677 246 711
rect 212 609 246 643
rect 212 541 246 575
rect 212 473 246 507
rect 212 405 246 439
rect 212 337 246 371
rect 212 269 246 303
rect 212 201 246 235
rect 298 1153 332 1187
rect 298 1085 332 1119
rect 298 1017 332 1051
rect 298 949 332 983
rect 298 881 332 915
rect 298 813 332 847
rect 298 745 332 779
rect 298 677 332 711
rect 298 609 332 643
rect 298 541 332 575
rect 298 473 332 507
rect 298 405 332 439
rect 298 337 332 371
rect 298 269 332 303
rect 298 201 332 235
rect 384 1153 418 1187
rect 384 1085 418 1119
rect 384 1017 418 1051
rect 384 949 418 983
rect 384 881 418 915
rect 384 813 418 847
rect 384 745 418 779
rect 384 677 418 711
rect 384 609 418 643
rect 384 541 418 575
rect 384 473 418 507
rect 384 405 418 439
rect 384 337 418 371
rect 384 269 418 303
rect 384 201 418 235
rect 470 1153 504 1187
rect 470 1085 504 1119
rect 470 1017 504 1051
rect 470 949 504 983
rect 470 881 504 915
rect 470 813 504 847
rect 470 745 504 779
rect 470 677 504 711
rect 470 609 504 643
rect 470 541 504 575
rect 470 473 504 507
rect 470 405 504 439
rect 470 337 504 371
rect 470 269 504 303
rect 470 201 504 235
rect 556 1153 590 1187
rect 556 1085 590 1119
rect 556 1017 590 1051
rect 556 949 590 983
rect 556 881 590 915
rect 556 813 590 847
rect 556 745 590 779
rect 556 677 590 711
rect 556 609 590 643
rect 556 541 590 575
rect 556 473 590 507
rect 556 405 590 439
rect 556 337 590 371
rect 556 269 590 303
rect 556 201 590 235
rect 642 1153 676 1187
rect 642 1085 676 1119
rect 642 1017 676 1051
rect 642 949 676 983
rect 642 881 676 915
rect 642 813 676 847
rect 642 745 676 779
rect 642 677 676 711
rect 642 609 676 643
rect 642 541 676 575
rect 642 473 676 507
rect 642 405 676 439
rect 642 337 676 371
rect 642 269 676 303
rect 642 201 676 235
<< psubdiff >>
rect 41 1187 111 1199
rect 41 1153 58 1187
rect 92 1153 111 1187
rect 41 1119 111 1153
rect 41 1085 58 1119
rect 92 1085 111 1119
rect 41 1051 111 1085
rect 41 1017 58 1051
rect 92 1017 111 1051
rect 41 983 111 1017
rect 41 949 58 983
rect 92 949 111 983
rect 41 915 111 949
rect 41 881 58 915
rect 92 881 111 915
rect 41 847 111 881
rect 41 813 58 847
rect 92 813 111 847
rect 41 779 111 813
rect 41 745 58 779
rect 92 745 111 779
rect 41 711 111 745
rect 41 677 58 711
rect 92 677 111 711
rect 41 643 111 677
rect 41 609 58 643
rect 92 609 111 643
rect 41 575 111 609
rect 41 541 58 575
rect 92 541 111 575
rect 41 507 111 541
rect 41 473 58 507
rect 92 473 111 507
rect 41 439 111 473
rect 41 405 58 439
rect 92 405 111 439
rect 41 371 111 405
rect 41 337 58 371
rect 92 337 111 371
rect 41 303 111 337
rect 41 269 58 303
rect 92 269 111 303
rect 41 235 111 269
rect 41 201 58 235
rect 92 201 111 235
rect 41 189 111 201
rect 691 1187 761 1199
rect 691 1153 710 1187
rect 744 1153 761 1187
rect 691 1119 761 1153
rect 691 1085 710 1119
rect 744 1085 761 1119
rect 691 1051 761 1085
rect 691 1017 710 1051
rect 744 1017 761 1051
rect 691 983 761 1017
rect 691 949 710 983
rect 744 949 761 983
rect 691 915 761 949
rect 691 881 710 915
rect 744 881 761 915
rect 691 847 761 881
rect 691 813 710 847
rect 744 813 761 847
rect 691 779 761 813
rect 691 745 710 779
rect 744 745 761 779
rect 691 711 761 745
rect 691 677 710 711
rect 744 677 761 711
rect 691 643 761 677
rect 691 609 710 643
rect 744 609 761 643
rect 691 575 761 609
rect 691 541 710 575
rect 744 541 761 575
rect 691 507 761 541
rect 691 473 710 507
rect 744 473 761 507
rect 691 439 761 473
rect 691 405 710 439
rect 744 405 761 439
rect 691 371 761 405
rect 691 337 710 371
rect 744 337 761 371
rect 691 303 761 337
rect 691 269 710 303
rect 744 269 761 303
rect 691 235 761 269
rect 691 201 710 235
rect 744 201 761 235
rect 691 189 761 201
<< psubdiffcont >>
rect 58 1153 92 1187
rect 58 1085 92 1119
rect 58 1017 92 1051
rect 58 949 92 983
rect 58 881 92 915
rect 58 813 92 847
rect 58 745 92 779
rect 58 677 92 711
rect 58 609 92 643
rect 58 541 92 575
rect 58 473 92 507
rect 58 405 92 439
rect 58 337 92 371
rect 58 269 92 303
rect 58 201 92 235
rect 710 1153 744 1187
rect 710 1085 744 1119
rect 710 1017 744 1051
rect 710 949 744 983
rect 710 881 744 915
rect 710 813 744 847
rect 710 745 744 779
rect 710 677 744 711
rect 710 609 744 643
rect 710 541 744 575
rect 710 473 744 507
rect 710 405 744 439
rect 710 337 744 371
rect 710 269 744 303
rect 710 201 744 235
<< poly >>
rect 243 1367 559 1388
rect 243 1333 264 1367
rect 298 1333 344 1367
rect 378 1333 424 1367
rect 458 1333 504 1367
rect 538 1333 559 1367
rect 243 1299 559 1333
rect 120 1275 201 1291
rect 120 1241 136 1275
rect 170 1241 201 1275
rect 243 1265 264 1299
rect 298 1265 344 1299
rect 378 1265 424 1299
rect 458 1265 504 1299
rect 538 1265 559 1299
rect 243 1249 559 1265
rect 601 1275 682 1291
rect 120 1225 201 1241
rect 171 1199 201 1225
rect 257 1199 287 1249
rect 343 1199 373 1249
rect 429 1199 459 1249
rect 515 1199 545 1249
rect 601 1241 632 1275
rect 666 1241 682 1275
rect 601 1225 682 1241
rect 601 1199 631 1225
rect 171 163 201 189
rect 120 147 201 163
rect 120 113 136 147
rect 170 113 201 147
rect 257 139 287 189
rect 343 139 373 189
rect 429 139 459 189
rect 515 139 545 189
rect 601 163 631 189
rect 601 147 682 163
rect 120 97 201 113
rect 243 123 559 139
rect 243 89 264 123
rect 298 89 344 123
rect 378 89 424 123
rect 458 89 504 123
rect 538 89 559 123
rect 601 113 632 147
rect 666 113 682 147
rect 601 97 682 113
rect 243 55 559 89
rect 243 21 264 55
rect 298 21 344 55
rect 378 21 424 55
rect 458 21 504 55
rect 538 21 559 55
rect 243 0 559 21
<< polycont >>
rect 264 1333 298 1367
rect 344 1333 378 1367
rect 424 1333 458 1367
rect 504 1333 538 1367
rect 136 1241 170 1275
rect 264 1265 298 1299
rect 344 1265 378 1299
rect 424 1265 458 1299
rect 504 1265 538 1299
rect 632 1241 666 1275
rect 136 113 170 147
rect 264 89 298 123
rect 344 89 378 123
rect 424 89 458 123
rect 504 89 538 123
rect 632 113 666 147
rect 264 21 298 55
rect 344 21 378 55
rect 424 21 458 55
rect 504 21 538 55
<< locali >>
rect 243 1369 559 1388
rect 243 1335 255 1369
rect 289 1367 337 1369
rect 371 1367 431 1369
rect 465 1367 513 1369
rect 298 1335 337 1367
rect 243 1333 264 1335
rect 298 1333 344 1335
rect 378 1333 424 1367
rect 465 1335 504 1367
rect 547 1335 559 1369
rect 458 1333 504 1335
rect 538 1333 559 1335
rect 243 1299 559 1333
rect 243 1297 264 1299
rect 298 1297 344 1299
rect 120 1275 186 1291
rect 120 1241 136 1275
rect 170 1241 186 1275
rect 243 1263 255 1297
rect 298 1265 337 1297
rect 378 1265 424 1299
rect 458 1297 504 1299
rect 538 1297 559 1299
rect 465 1265 504 1297
rect 289 1263 337 1265
rect 371 1263 431 1265
rect 465 1263 513 1265
rect 547 1263 559 1297
rect 243 1249 559 1263
rect 616 1275 682 1291
rect 120 1225 186 1241
rect 616 1241 632 1275
rect 666 1241 682 1275
rect 616 1225 682 1241
rect 120 1203 160 1225
rect 642 1203 682 1225
rect 41 1187 160 1203
rect 41 1153 58 1187
rect 92 1179 126 1187
rect 94 1153 126 1179
rect 41 1145 60 1153
rect 94 1145 160 1153
rect 41 1119 160 1145
rect 41 1085 58 1119
rect 92 1107 126 1119
rect 94 1085 126 1107
rect 41 1073 60 1085
rect 94 1073 160 1085
rect 41 1051 160 1073
rect 41 1017 58 1051
rect 92 1035 126 1051
rect 94 1017 126 1035
rect 41 1001 60 1017
rect 94 1001 160 1017
rect 41 983 160 1001
rect 41 949 58 983
rect 92 963 126 983
rect 94 949 126 963
rect 41 929 60 949
rect 94 929 160 949
rect 41 915 160 929
rect 41 881 58 915
rect 92 891 126 915
rect 94 881 126 891
rect 41 857 60 881
rect 94 857 160 881
rect 41 847 160 857
rect 41 813 58 847
rect 92 819 126 847
rect 94 813 126 819
rect 41 785 60 813
rect 94 785 160 813
rect 41 779 160 785
rect 41 745 58 779
rect 92 747 126 779
rect 94 745 126 747
rect 41 713 60 745
rect 94 713 160 745
rect 41 711 160 713
rect 41 677 58 711
rect 92 677 126 711
rect 41 675 160 677
rect 41 643 60 675
rect 94 643 160 675
rect 41 609 58 643
rect 94 641 126 643
rect 92 609 126 641
rect 41 603 160 609
rect 41 575 60 603
rect 94 575 160 603
rect 41 541 58 575
rect 94 569 126 575
rect 92 541 126 569
rect 41 531 160 541
rect 41 507 60 531
rect 94 507 160 531
rect 41 473 58 507
rect 94 497 126 507
rect 92 473 126 497
rect 41 459 160 473
rect 41 439 60 459
rect 94 439 160 459
rect 41 405 58 439
rect 94 425 126 439
rect 92 405 126 425
rect 41 387 160 405
rect 41 371 60 387
rect 94 371 160 387
rect 41 337 58 371
rect 94 353 126 371
rect 92 337 126 353
rect 41 315 160 337
rect 41 303 60 315
rect 94 303 160 315
rect 41 269 58 303
rect 94 281 126 303
rect 92 269 126 281
rect 41 243 160 269
rect 41 235 60 243
rect 94 235 160 243
rect 41 201 58 235
rect 94 209 126 235
rect 92 201 126 209
rect 41 185 160 201
rect 212 1187 246 1203
rect 212 1119 246 1145
rect 212 1051 246 1073
rect 212 983 246 1001
rect 212 915 246 929
rect 212 847 246 857
rect 212 779 246 785
rect 212 711 246 713
rect 212 675 246 677
rect 212 603 246 609
rect 212 531 246 541
rect 212 459 246 473
rect 212 387 246 405
rect 212 315 246 337
rect 212 243 246 269
rect 212 185 246 201
rect 298 1187 332 1203
rect 298 1119 332 1145
rect 298 1051 332 1073
rect 298 983 332 1001
rect 298 915 332 929
rect 298 847 332 857
rect 298 779 332 785
rect 298 711 332 713
rect 298 675 332 677
rect 298 603 332 609
rect 298 531 332 541
rect 298 459 332 473
rect 298 387 332 405
rect 298 315 332 337
rect 298 243 332 269
rect 298 185 332 201
rect 384 1187 418 1203
rect 384 1119 418 1145
rect 384 1051 418 1073
rect 384 983 418 1001
rect 384 915 418 929
rect 384 847 418 857
rect 384 779 418 785
rect 384 711 418 713
rect 384 675 418 677
rect 384 603 418 609
rect 384 531 418 541
rect 384 459 418 473
rect 384 387 418 405
rect 384 315 418 337
rect 384 243 418 269
rect 384 185 418 201
rect 470 1187 504 1203
rect 470 1119 504 1145
rect 470 1051 504 1073
rect 470 983 504 1001
rect 470 915 504 929
rect 470 847 504 857
rect 470 779 504 785
rect 470 711 504 713
rect 470 675 504 677
rect 470 603 504 609
rect 470 531 504 541
rect 470 459 504 473
rect 470 387 504 405
rect 470 315 504 337
rect 470 243 504 269
rect 470 185 504 201
rect 556 1187 590 1203
rect 556 1119 590 1145
rect 556 1051 590 1073
rect 556 983 590 1001
rect 556 915 590 929
rect 556 847 590 857
rect 556 779 590 785
rect 556 711 590 713
rect 556 675 590 677
rect 556 603 590 609
rect 556 531 590 541
rect 556 459 590 473
rect 556 387 590 405
rect 556 315 590 337
rect 556 243 590 269
rect 556 185 590 201
rect 642 1187 761 1203
rect 676 1179 710 1187
rect 676 1153 708 1179
rect 744 1153 761 1187
rect 642 1145 708 1153
rect 742 1145 761 1153
rect 642 1119 761 1145
rect 676 1107 710 1119
rect 676 1085 708 1107
rect 744 1085 761 1119
rect 642 1073 708 1085
rect 742 1073 761 1085
rect 642 1051 761 1073
rect 676 1035 710 1051
rect 676 1017 708 1035
rect 744 1017 761 1051
rect 642 1001 708 1017
rect 742 1001 761 1017
rect 642 983 761 1001
rect 676 963 710 983
rect 676 949 708 963
rect 744 949 761 983
rect 642 929 708 949
rect 742 929 761 949
rect 642 915 761 929
rect 676 891 710 915
rect 676 881 708 891
rect 744 881 761 915
rect 642 857 708 881
rect 742 857 761 881
rect 642 847 761 857
rect 676 819 710 847
rect 676 813 708 819
rect 744 813 761 847
rect 642 785 708 813
rect 742 785 761 813
rect 642 779 761 785
rect 676 747 710 779
rect 676 745 708 747
rect 744 745 761 779
rect 642 713 708 745
rect 742 713 761 745
rect 642 711 761 713
rect 676 677 710 711
rect 744 677 761 711
rect 642 675 761 677
rect 642 643 708 675
rect 742 643 761 675
rect 676 641 708 643
rect 676 609 710 641
rect 744 609 761 643
rect 642 603 761 609
rect 642 575 708 603
rect 742 575 761 603
rect 676 569 708 575
rect 676 541 710 569
rect 744 541 761 575
rect 642 531 761 541
rect 642 507 708 531
rect 742 507 761 531
rect 676 497 708 507
rect 676 473 710 497
rect 744 473 761 507
rect 642 459 761 473
rect 642 439 708 459
rect 742 439 761 459
rect 676 425 708 439
rect 676 405 710 425
rect 744 405 761 439
rect 642 387 761 405
rect 642 371 708 387
rect 742 371 761 387
rect 676 353 708 371
rect 676 337 710 353
rect 744 337 761 371
rect 642 315 761 337
rect 642 303 708 315
rect 742 303 761 315
rect 676 281 708 303
rect 676 269 710 281
rect 744 269 761 303
rect 642 243 761 269
rect 642 235 708 243
rect 742 235 761 243
rect 676 209 708 235
rect 676 201 710 209
rect 744 201 761 235
rect 642 185 761 201
rect 120 163 160 185
rect 642 163 682 185
rect 120 147 186 163
rect 120 113 136 147
rect 170 113 186 147
rect 616 147 682 163
rect 120 97 186 113
rect 243 125 559 139
rect 243 91 255 125
rect 289 123 337 125
rect 371 123 431 125
rect 465 123 513 125
rect 298 91 337 123
rect 243 89 264 91
rect 298 89 344 91
rect 378 89 424 123
rect 465 91 504 123
rect 547 91 559 125
rect 616 113 632 147
rect 666 113 682 147
rect 616 97 682 113
rect 458 89 504 91
rect 538 89 559 91
rect 243 55 559 89
rect 243 53 264 55
rect 298 53 344 55
rect 243 19 255 53
rect 298 21 337 53
rect 378 21 424 55
rect 458 53 504 55
rect 538 53 559 55
rect 465 21 504 53
rect 289 19 337 21
rect 371 19 431 21
rect 465 19 513 21
rect 547 19 559 53
rect 243 0 559 19
<< viali >>
rect 255 1367 289 1369
rect 337 1367 371 1369
rect 431 1367 465 1369
rect 513 1367 547 1369
rect 255 1335 264 1367
rect 264 1335 289 1367
rect 337 1335 344 1367
rect 344 1335 371 1367
rect 431 1335 458 1367
rect 458 1335 465 1367
rect 513 1335 538 1367
rect 538 1335 547 1367
rect 255 1265 264 1297
rect 264 1265 289 1297
rect 337 1265 344 1297
rect 344 1265 371 1297
rect 431 1265 458 1297
rect 458 1265 465 1297
rect 513 1265 538 1297
rect 538 1265 547 1297
rect 255 1263 289 1265
rect 337 1263 371 1265
rect 431 1263 465 1265
rect 513 1263 547 1265
rect 60 1153 92 1179
rect 92 1153 94 1179
rect 60 1145 94 1153
rect 60 1085 92 1107
rect 92 1085 94 1107
rect 60 1073 94 1085
rect 60 1017 92 1035
rect 92 1017 94 1035
rect 60 1001 94 1017
rect 60 949 92 963
rect 92 949 94 963
rect 60 929 94 949
rect 60 881 92 891
rect 92 881 94 891
rect 60 857 94 881
rect 60 813 92 819
rect 92 813 94 819
rect 60 785 94 813
rect 60 745 92 747
rect 92 745 94 747
rect 60 713 94 745
rect 60 643 94 675
rect 60 641 92 643
rect 92 641 94 643
rect 60 575 94 603
rect 60 569 92 575
rect 92 569 94 575
rect 60 507 94 531
rect 60 497 92 507
rect 92 497 94 507
rect 60 439 94 459
rect 60 425 92 439
rect 92 425 94 439
rect 60 371 94 387
rect 60 353 92 371
rect 92 353 94 371
rect 60 303 94 315
rect 60 281 92 303
rect 92 281 94 303
rect 60 235 94 243
rect 60 209 92 235
rect 92 209 94 235
rect 212 1153 246 1179
rect 212 1145 246 1153
rect 212 1085 246 1107
rect 212 1073 246 1085
rect 212 1017 246 1035
rect 212 1001 246 1017
rect 212 949 246 963
rect 212 929 246 949
rect 212 881 246 891
rect 212 857 246 881
rect 212 813 246 819
rect 212 785 246 813
rect 212 745 246 747
rect 212 713 246 745
rect 212 643 246 675
rect 212 641 246 643
rect 212 575 246 603
rect 212 569 246 575
rect 212 507 246 531
rect 212 497 246 507
rect 212 439 246 459
rect 212 425 246 439
rect 212 371 246 387
rect 212 353 246 371
rect 212 303 246 315
rect 212 281 246 303
rect 212 235 246 243
rect 212 209 246 235
rect 298 1153 332 1179
rect 298 1145 332 1153
rect 298 1085 332 1107
rect 298 1073 332 1085
rect 298 1017 332 1035
rect 298 1001 332 1017
rect 298 949 332 963
rect 298 929 332 949
rect 298 881 332 891
rect 298 857 332 881
rect 298 813 332 819
rect 298 785 332 813
rect 298 745 332 747
rect 298 713 332 745
rect 298 643 332 675
rect 298 641 332 643
rect 298 575 332 603
rect 298 569 332 575
rect 298 507 332 531
rect 298 497 332 507
rect 298 439 332 459
rect 298 425 332 439
rect 298 371 332 387
rect 298 353 332 371
rect 298 303 332 315
rect 298 281 332 303
rect 298 235 332 243
rect 298 209 332 235
rect 384 1153 418 1179
rect 384 1145 418 1153
rect 384 1085 418 1107
rect 384 1073 418 1085
rect 384 1017 418 1035
rect 384 1001 418 1017
rect 384 949 418 963
rect 384 929 418 949
rect 384 881 418 891
rect 384 857 418 881
rect 384 813 418 819
rect 384 785 418 813
rect 384 745 418 747
rect 384 713 418 745
rect 384 643 418 675
rect 384 641 418 643
rect 384 575 418 603
rect 384 569 418 575
rect 384 507 418 531
rect 384 497 418 507
rect 384 439 418 459
rect 384 425 418 439
rect 384 371 418 387
rect 384 353 418 371
rect 384 303 418 315
rect 384 281 418 303
rect 384 235 418 243
rect 384 209 418 235
rect 470 1153 504 1179
rect 470 1145 504 1153
rect 470 1085 504 1107
rect 470 1073 504 1085
rect 470 1017 504 1035
rect 470 1001 504 1017
rect 470 949 504 963
rect 470 929 504 949
rect 470 881 504 891
rect 470 857 504 881
rect 470 813 504 819
rect 470 785 504 813
rect 470 745 504 747
rect 470 713 504 745
rect 470 643 504 675
rect 470 641 504 643
rect 470 575 504 603
rect 470 569 504 575
rect 470 507 504 531
rect 470 497 504 507
rect 470 439 504 459
rect 470 425 504 439
rect 470 371 504 387
rect 470 353 504 371
rect 470 303 504 315
rect 470 281 504 303
rect 470 235 504 243
rect 470 209 504 235
rect 556 1153 590 1179
rect 556 1145 590 1153
rect 556 1085 590 1107
rect 556 1073 590 1085
rect 556 1017 590 1035
rect 556 1001 590 1017
rect 556 949 590 963
rect 556 929 590 949
rect 556 881 590 891
rect 556 857 590 881
rect 556 813 590 819
rect 556 785 590 813
rect 556 745 590 747
rect 556 713 590 745
rect 556 643 590 675
rect 556 641 590 643
rect 556 575 590 603
rect 556 569 590 575
rect 556 507 590 531
rect 556 497 590 507
rect 556 439 590 459
rect 556 425 590 439
rect 556 371 590 387
rect 556 353 590 371
rect 556 303 590 315
rect 556 281 590 303
rect 556 235 590 243
rect 556 209 590 235
rect 708 1153 710 1179
rect 710 1153 742 1179
rect 708 1145 742 1153
rect 708 1085 710 1107
rect 710 1085 742 1107
rect 708 1073 742 1085
rect 708 1017 710 1035
rect 710 1017 742 1035
rect 708 1001 742 1017
rect 708 949 710 963
rect 710 949 742 963
rect 708 929 742 949
rect 708 881 710 891
rect 710 881 742 891
rect 708 857 742 881
rect 708 813 710 819
rect 710 813 742 819
rect 708 785 742 813
rect 708 745 710 747
rect 710 745 742 747
rect 708 713 742 745
rect 708 643 742 675
rect 708 641 710 643
rect 710 641 742 643
rect 708 575 742 603
rect 708 569 710 575
rect 710 569 742 575
rect 708 507 742 531
rect 708 497 710 507
rect 710 497 742 507
rect 708 439 742 459
rect 708 425 710 439
rect 710 425 742 439
rect 708 371 742 387
rect 708 353 710 371
rect 710 353 742 371
rect 708 303 742 315
rect 708 281 710 303
rect 710 281 742 303
rect 708 235 742 243
rect 708 209 710 235
rect 710 209 742 235
rect 255 123 289 125
rect 337 123 371 125
rect 431 123 465 125
rect 513 123 547 125
rect 255 91 264 123
rect 264 91 289 123
rect 337 91 344 123
rect 344 91 371 123
rect 431 91 458 123
rect 458 91 465 123
rect 513 91 538 123
rect 538 91 547 123
rect 255 21 264 53
rect 264 21 289 53
rect 337 21 344 53
rect 344 21 371 53
rect 431 21 458 53
rect 458 21 465 53
rect 513 21 538 53
rect 538 21 547 53
rect 255 19 289 21
rect 337 19 371 21
rect 431 19 465 21
rect 513 19 547 21
<< metal1 >>
rect 243 1369 559 1388
rect 243 1335 255 1369
rect 289 1335 337 1369
rect 371 1335 431 1369
rect 465 1335 513 1369
rect 547 1335 559 1369
rect 243 1297 559 1335
rect 243 1263 255 1297
rect 289 1263 337 1297
rect 371 1263 431 1297
rect 465 1263 513 1297
rect 547 1263 559 1297
rect 243 1251 559 1263
rect 41 1179 100 1191
rect 41 1145 60 1179
rect 94 1145 100 1179
rect 41 1107 100 1145
rect 41 1073 60 1107
rect 94 1073 100 1107
rect 41 1035 100 1073
rect 41 1001 60 1035
rect 94 1001 100 1035
rect 41 963 100 1001
rect 41 929 60 963
rect 94 929 100 963
rect 41 891 100 929
rect 41 857 60 891
rect 94 857 100 891
rect 41 819 100 857
rect 41 785 60 819
rect 94 785 100 819
rect 41 747 100 785
rect 41 713 60 747
rect 94 713 100 747
rect 41 675 100 713
rect 41 641 60 675
rect 94 641 100 675
rect 41 603 100 641
rect 41 569 60 603
rect 94 569 100 603
rect 41 531 100 569
rect 41 497 60 531
rect 94 497 100 531
rect 41 459 100 497
rect 41 425 60 459
rect 94 425 100 459
rect 41 387 100 425
rect 41 353 60 387
rect 94 353 100 387
rect 41 315 100 353
rect 41 281 60 315
rect 94 281 100 315
rect 41 243 100 281
rect 41 209 60 243
rect 94 209 100 243
rect 41 197 100 209
rect 203 1179 255 1191
rect 203 1145 212 1179
rect 246 1145 255 1179
rect 203 1107 255 1145
rect 203 1073 212 1107
rect 246 1073 255 1107
rect 203 1035 255 1073
rect 203 1001 212 1035
rect 246 1001 255 1035
rect 203 963 255 1001
rect 203 929 212 963
rect 246 929 255 963
rect 203 891 255 929
rect 203 857 212 891
rect 246 857 255 891
rect 203 819 255 857
rect 203 785 212 819
rect 246 785 255 819
rect 203 747 255 785
rect 203 713 212 747
rect 246 713 255 747
rect 203 675 255 713
rect 203 641 212 675
rect 246 641 255 675
rect 203 639 255 641
rect 203 575 212 587
rect 246 575 255 587
rect 203 511 212 523
rect 246 511 255 523
rect 203 447 212 459
rect 246 447 255 459
rect 203 387 255 395
rect 203 383 212 387
rect 246 383 255 387
rect 203 319 255 331
rect 203 255 255 267
rect 203 197 255 203
rect 289 1185 341 1191
rect 289 1121 341 1133
rect 289 1057 341 1069
rect 289 1001 298 1005
rect 332 1001 341 1005
rect 289 993 341 1001
rect 289 929 298 941
rect 332 929 341 941
rect 289 865 298 877
rect 332 865 341 877
rect 289 801 298 813
rect 332 801 341 813
rect 289 747 341 749
rect 289 713 298 747
rect 332 713 341 747
rect 289 675 341 713
rect 289 641 298 675
rect 332 641 341 675
rect 289 603 341 641
rect 289 569 298 603
rect 332 569 341 603
rect 289 531 341 569
rect 289 497 298 531
rect 332 497 341 531
rect 289 459 341 497
rect 289 425 298 459
rect 332 425 341 459
rect 289 387 341 425
rect 289 353 298 387
rect 332 353 341 387
rect 289 315 341 353
rect 289 281 298 315
rect 332 281 341 315
rect 289 243 341 281
rect 289 209 298 243
rect 332 209 341 243
rect 289 197 341 209
rect 375 1179 427 1191
rect 375 1145 384 1179
rect 418 1145 427 1179
rect 375 1107 427 1145
rect 375 1073 384 1107
rect 418 1073 427 1107
rect 375 1035 427 1073
rect 375 1001 384 1035
rect 418 1001 427 1035
rect 375 963 427 1001
rect 375 929 384 963
rect 418 929 427 963
rect 375 891 427 929
rect 375 857 384 891
rect 418 857 427 891
rect 375 819 427 857
rect 375 785 384 819
rect 418 785 427 819
rect 375 747 427 785
rect 375 713 384 747
rect 418 713 427 747
rect 375 675 427 713
rect 375 641 384 675
rect 418 641 427 675
rect 375 639 427 641
rect 375 575 384 587
rect 418 575 427 587
rect 375 511 384 523
rect 418 511 427 523
rect 375 447 384 459
rect 418 447 427 459
rect 375 387 427 395
rect 375 383 384 387
rect 418 383 427 387
rect 375 319 427 331
rect 375 255 427 267
rect 375 197 427 203
rect 461 1185 513 1191
rect 461 1121 513 1133
rect 461 1057 513 1069
rect 461 1001 470 1005
rect 504 1001 513 1005
rect 461 993 513 1001
rect 461 929 470 941
rect 504 929 513 941
rect 461 865 470 877
rect 504 865 513 877
rect 461 801 470 813
rect 504 801 513 813
rect 461 747 513 749
rect 461 713 470 747
rect 504 713 513 747
rect 461 675 513 713
rect 461 641 470 675
rect 504 641 513 675
rect 461 603 513 641
rect 461 569 470 603
rect 504 569 513 603
rect 461 531 513 569
rect 461 497 470 531
rect 504 497 513 531
rect 461 459 513 497
rect 461 425 470 459
rect 504 425 513 459
rect 461 387 513 425
rect 461 353 470 387
rect 504 353 513 387
rect 461 315 513 353
rect 461 281 470 315
rect 504 281 513 315
rect 461 243 513 281
rect 461 209 470 243
rect 504 209 513 243
rect 461 197 513 209
rect 547 1179 599 1191
rect 547 1145 556 1179
rect 590 1145 599 1179
rect 547 1107 599 1145
rect 547 1073 556 1107
rect 590 1073 599 1107
rect 547 1035 599 1073
rect 547 1001 556 1035
rect 590 1001 599 1035
rect 547 963 599 1001
rect 547 929 556 963
rect 590 929 599 963
rect 547 891 599 929
rect 547 857 556 891
rect 590 857 599 891
rect 547 819 599 857
rect 547 785 556 819
rect 590 785 599 819
rect 547 747 599 785
rect 547 713 556 747
rect 590 713 599 747
rect 547 675 599 713
rect 547 641 556 675
rect 590 641 599 675
rect 547 639 599 641
rect 547 575 556 587
rect 590 575 599 587
rect 547 511 556 523
rect 590 511 599 523
rect 547 447 556 459
rect 590 447 599 459
rect 547 387 599 395
rect 547 383 556 387
rect 590 383 599 387
rect 547 319 599 331
rect 547 255 599 267
rect 547 197 599 203
rect 702 1179 761 1191
rect 702 1145 708 1179
rect 742 1145 761 1179
rect 702 1107 761 1145
rect 702 1073 708 1107
rect 742 1073 761 1107
rect 702 1035 761 1073
rect 702 1001 708 1035
rect 742 1001 761 1035
rect 702 963 761 1001
rect 702 929 708 963
rect 742 929 761 963
rect 702 891 761 929
rect 702 857 708 891
rect 742 857 761 891
rect 702 819 761 857
rect 702 785 708 819
rect 742 785 761 819
rect 702 747 761 785
rect 702 713 708 747
rect 742 713 761 747
rect 702 675 761 713
rect 702 641 708 675
rect 742 641 761 675
rect 702 603 761 641
rect 702 569 708 603
rect 742 569 761 603
rect 702 531 761 569
rect 702 497 708 531
rect 742 497 761 531
rect 702 459 761 497
rect 702 425 708 459
rect 742 425 761 459
rect 702 387 761 425
rect 702 353 708 387
rect 742 353 761 387
rect 702 315 761 353
rect 702 281 708 315
rect 742 281 761 315
rect 702 243 761 281
rect 702 209 708 243
rect 742 209 761 243
rect 702 197 761 209
rect 243 125 559 137
rect 243 91 255 125
rect 289 91 337 125
rect 371 91 431 125
rect 465 91 513 125
rect 547 91 559 125
rect 243 53 559 91
rect 243 19 255 53
rect 289 19 337 53
rect 371 19 431 53
rect 465 19 513 53
rect 547 19 559 53
rect 243 0 559 19
<< via1 >>
rect 203 603 255 639
rect 203 587 212 603
rect 212 587 246 603
rect 246 587 255 603
rect 203 569 212 575
rect 212 569 246 575
rect 246 569 255 575
rect 203 531 255 569
rect 203 523 212 531
rect 212 523 246 531
rect 246 523 255 531
rect 203 497 212 511
rect 212 497 246 511
rect 246 497 255 511
rect 203 459 255 497
rect 203 425 212 447
rect 212 425 246 447
rect 246 425 255 447
rect 203 395 255 425
rect 203 353 212 383
rect 212 353 246 383
rect 246 353 255 383
rect 203 331 255 353
rect 203 315 255 319
rect 203 281 212 315
rect 212 281 246 315
rect 246 281 255 315
rect 203 267 255 281
rect 203 243 255 255
rect 203 209 212 243
rect 212 209 246 243
rect 246 209 255 243
rect 203 203 255 209
rect 289 1179 341 1185
rect 289 1145 298 1179
rect 298 1145 332 1179
rect 332 1145 341 1179
rect 289 1133 341 1145
rect 289 1107 341 1121
rect 289 1073 298 1107
rect 298 1073 332 1107
rect 332 1073 341 1107
rect 289 1069 341 1073
rect 289 1035 341 1057
rect 289 1005 298 1035
rect 298 1005 332 1035
rect 332 1005 341 1035
rect 289 963 341 993
rect 289 941 298 963
rect 298 941 332 963
rect 332 941 341 963
rect 289 891 341 929
rect 289 877 298 891
rect 298 877 332 891
rect 332 877 341 891
rect 289 857 298 865
rect 298 857 332 865
rect 332 857 341 865
rect 289 819 341 857
rect 289 813 298 819
rect 298 813 332 819
rect 332 813 341 819
rect 289 785 298 801
rect 298 785 332 801
rect 332 785 341 801
rect 289 749 341 785
rect 375 603 427 639
rect 375 587 384 603
rect 384 587 418 603
rect 418 587 427 603
rect 375 569 384 575
rect 384 569 418 575
rect 418 569 427 575
rect 375 531 427 569
rect 375 523 384 531
rect 384 523 418 531
rect 418 523 427 531
rect 375 497 384 511
rect 384 497 418 511
rect 418 497 427 511
rect 375 459 427 497
rect 375 425 384 447
rect 384 425 418 447
rect 418 425 427 447
rect 375 395 427 425
rect 375 353 384 383
rect 384 353 418 383
rect 418 353 427 383
rect 375 331 427 353
rect 375 315 427 319
rect 375 281 384 315
rect 384 281 418 315
rect 418 281 427 315
rect 375 267 427 281
rect 375 243 427 255
rect 375 209 384 243
rect 384 209 418 243
rect 418 209 427 243
rect 375 203 427 209
rect 461 1179 513 1185
rect 461 1145 470 1179
rect 470 1145 504 1179
rect 504 1145 513 1179
rect 461 1133 513 1145
rect 461 1107 513 1121
rect 461 1073 470 1107
rect 470 1073 504 1107
rect 504 1073 513 1107
rect 461 1069 513 1073
rect 461 1035 513 1057
rect 461 1005 470 1035
rect 470 1005 504 1035
rect 504 1005 513 1035
rect 461 963 513 993
rect 461 941 470 963
rect 470 941 504 963
rect 504 941 513 963
rect 461 891 513 929
rect 461 877 470 891
rect 470 877 504 891
rect 504 877 513 891
rect 461 857 470 865
rect 470 857 504 865
rect 504 857 513 865
rect 461 819 513 857
rect 461 813 470 819
rect 470 813 504 819
rect 504 813 513 819
rect 461 785 470 801
rect 470 785 504 801
rect 504 785 513 801
rect 461 749 513 785
rect 547 603 599 639
rect 547 587 556 603
rect 556 587 590 603
rect 590 587 599 603
rect 547 569 556 575
rect 556 569 590 575
rect 590 569 599 575
rect 547 531 599 569
rect 547 523 556 531
rect 556 523 590 531
rect 590 523 599 531
rect 547 497 556 511
rect 556 497 590 511
rect 590 497 599 511
rect 547 459 599 497
rect 547 425 556 447
rect 556 425 590 447
rect 590 425 599 447
rect 547 395 599 425
rect 547 353 556 383
rect 556 353 590 383
rect 590 353 599 383
rect 547 331 599 353
rect 547 315 599 319
rect 547 281 556 315
rect 556 281 590 315
rect 590 281 599 315
rect 547 267 599 281
rect 547 243 599 255
rect 547 209 556 243
rect 556 209 590 243
rect 590 209 599 243
rect 547 203 599 209
<< metal2 >>
rect 14 1185 788 1191
rect 14 1133 289 1185
rect 341 1133 461 1185
rect 513 1133 788 1185
rect 14 1121 788 1133
rect 14 1069 289 1121
rect 341 1069 461 1121
rect 513 1069 788 1121
rect 14 1057 788 1069
rect 14 1005 289 1057
rect 341 1005 461 1057
rect 513 1005 788 1057
rect 14 993 788 1005
rect 14 941 289 993
rect 341 941 461 993
rect 513 941 788 993
rect 14 929 788 941
rect 14 877 289 929
rect 341 877 461 929
rect 513 877 788 929
rect 14 865 788 877
rect 14 813 289 865
rect 341 813 461 865
rect 513 813 788 865
rect 14 801 788 813
rect 14 749 289 801
rect 341 749 461 801
rect 513 749 788 801
rect 14 719 788 749
rect 14 639 788 669
rect 14 587 203 639
rect 255 587 375 639
rect 427 587 547 639
rect 599 587 788 639
rect 14 575 788 587
rect 14 523 203 575
rect 255 523 375 575
rect 427 523 547 575
rect 599 523 788 575
rect 14 511 788 523
rect 14 459 203 511
rect 255 459 375 511
rect 427 459 547 511
rect 599 459 788 511
rect 14 447 788 459
rect 14 395 203 447
rect 255 395 375 447
rect 427 395 547 447
rect 599 395 788 447
rect 14 383 788 395
rect 14 331 203 383
rect 255 331 375 383
rect 427 331 547 383
rect 599 331 788 383
rect 14 319 788 331
rect 14 267 203 319
rect 255 267 375 319
rect 427 267 547 319
rect 599 267 788 319
rect 14 255 788 267
rect 14 203 203 255
rect 255 203 375 255
rect 427 203 547 255
rect 599 203 788 255
rect 14 197 788 203
<< labels >>
flabel metal1 s 301 42 511 92 0 FreeSans 200 0 0 0 GATE
port 4 nsew
flabel metal1 s 301 1286 511 1336 0 FreeSans 200 0 0 0 GATE
port 4 nsew
flabel metal1 s 41 675 100 705 0 FreeSans 200 90 0 0 SUBSTRATE
port 3 nsew
flabel metal1 s 702 683 761 713 0 FreeSans 200 90 0 0 SUBSTRATE
port 3 nsew
flabel comment s 613 697 613 697 0 FreeSans 180 90 0 0 dummy_poly
flabel comment s 184 703 184 703 0 FreeSans 180 90 0 0 dummy_poly
flabel comment s 315 694 315 694 0 FreeSans 300 0 0 0 D
flabel comment s 229 694 229 694 0 FreeSans 300 0 0 0 S
flabel comment s 487 694 487 694 0 FreeSans 300 0 0 0 S
flabel comment s 401 694 401 694 0 FreeSans 300 0 0 0 S
flabel comment s 315 694 315 694 0 FreeSans 300 0 0 0 S
flabel comment s 229 694 229 694 0 FreeSans 300 0 0 0 S
flabel comment s 573 694 573 694 0 FreeSans 300 0 0 0 S
flabel comment s 487 694 487 694 0 FreeSans 300 0 0 0 D
flabel comment s 401 694 401 694 0 FreeSans 300 0 0 0 S
flabel metal2 s 14 384 35 512 7 FreeSans 300 180 0 0 SOURCE
port 5 nsew
flabel metal2 s 14 908 35 1036 7 FreeSans 300 180 0 0 DRAIN
port 6 nsew
<< properties >>
string GDS_END 6489682
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 6462072
<< end >>
