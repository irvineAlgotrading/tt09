magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -66 1151 102 1251
rect -66 419 3079 1151
rect -66 377 102 419
rect 1883 341 3079 419
rect 3479 409 4339 1219
<< pwell >>
rect -26 1585 5018 1671
rect 449 1353 2439 1585
rect 2748 1353 3006 1585
rect 183 1217 3006 1353
rect 3534 1303 4297 1585
rect 183 43 1175 359
rect 3534 43 4012 325
rect -26 -43 5018 43
<< scnmos >>
rect 3617 1329 3647 1477
rect 3703 1329 3733 1477
rect 3799 1329 3829 1477
rect 3893 1329 3923 1477
rect 4098 1329 4128 1477
rect 4184 1329 4214 1477
rect 3623 151 3653 299
rect 3717 151 3747 299
rect 3813 151 3843 299
rect 3899 151 3929 299
<< scpmoshvt >>
rect 3620 959 3650 1183
rect 3710 959 3740 1183
rect 3800 959 3830 1183
rect 3890 959 3920 1183
rect 4097 959 4127 1183
rect 4187 959 4217 1183
rect 3626 445 3656 669
rect 3716 445 3746 669
rect 3806 445 3836 669
rect 3896 445 3926 669
<< mvnmos >>
rect 262 1243 362 1327
rect 2561 1243 2661 1327
rect 2827 1243 2927 1393
rect 262 133 362 333
rect 418 133 518 333
rect 574 133 674 333
rect 840 133 940 333
rect 996 133 1096 333
<< mvpmos >>
rect 262 485 362 1085
rect 418 485 518 1085
rect 574 485 674 1085
rect 840 485 940 785
rect 996 485 1096 785
rect 1310 571 1410 871
rect 1466 571 1566 871
rect 2092 407 2192 1007
rect 2248 407 2348 1007
rect 2404 407 2504 1007
rect 2560 407 2660 1007
rect 2827 857 2927 1007
<< mvnnmos >>
rect 528 1243 708 1443
rect 764 1243 944 1443
rect 1000 1243 1180 1443
rect 1236 1243 1416 1443
rect 1472 1243 1652 1443
rect 1708 1243 1888 1443
rect 1944 1243 2124 1443
rect 2180 1243 2360 1443
<< ndiff >>
rect 3560 1449 3617 1477
rect 3560 1415 3572 1449
rect 3606 1415 3617 1449
rect 3560 1329 3617 1415
rect 3647 1453 3703 1477
rect 3647 1419 3658 1453
rect 3692 1419 3703 1453
rect 3647 1375 3703 1419
rect 3647 1341 3658 1375
rect 3692 1341 3703 1375
rect 3647 1329 3703 1341
rect 3733 1449 3799 1477
rect 3733 1415 3754 1449
rect 3788 1415 3799 1449
rect 3733 1329 3799 1415
rect 3829 1453 3893 1477
rect 3829 1419 3840 1453
rect 3874 1419 3893 1453
rect 3829 1375 3893 1419
rect 3829 1341 3840 1375
rect 3874 1341 3893 1375
rect 3829 1329 3893 1341
rect 3923 1465 3986 1477
rect 3923 1431 3940 1465
rect 3974 1431 3986 1465
rect 3923 1375 3986 1431
rect 3923 1341 3940 1375
rect 3974 1341 3986 1375
rect 3923 1329 3986 1341
rect 4041 1465 4098 1477
rect 4041 1431 4053 1465
rect 4087 1431 4098 1465
rect 4041 1375 4098 1431
rect 4041 1341 4053 1375
rect 4087 1341 4098 1375
rect 4041 1329 4098 1341
rect 4128 1453 4184 1477
rect 4128 1419 4139 1453
rect 4173 1419 4184 1453
rect 4128 1375 4184 1419
rect 4128 1341 4139 1375
rect 4173 1341 4184 1375
rect 4128 1329 4184 1341
rect 4214 1465 4271 1477
rect 4214 1431 4225 1465
rect 4259 1431 4271 1465
rect 4214 1375 4271 1431
rect 4214 1341 4225 1375
rect 4259 1341 4271 1375
rect 4214 1329 4271 1341
rect 3560 197 3623 299
rect 3560 163 3572 197
rect 3606 163 3623 197
rect 3560 151 3623 163
rect 3653 287 3717 299
rect 3653 253 3672 287
rect 3706 253 3717 287
rect 3653 209 3717 253
rect 3653 175 3672 209
rect 3706 175 3717 209
rect 3653 151 3717 175
rect 3747 213 3813 299
rect 3747 179 3758 213
rect 3792 179 3813 213
rect 3747 151 3813 179
rect 3843 287 3899 299
rect 3843 253 3854 287
rect 3888 253 3899 287
rect 3843 209 3899 253
rect 3843 175 3854 209
rect 3888 175 3899 209
rect 3843 151 3899 175
rect 3929 213 3986 299
rect 3929 179 3940 213
rect 3974 179 3986 213
rect 3929 151 3986 179
<< pdiff >>
rect 3561 1077 3620 1183
rect 3561 1043 3573 1077
rect 3607 1043 3620 1077
rect 3561 1005 3620 1043
rect 3561 971 3573 1005
rect 3607 971 3620 1005
rect 3561 959 3620 971
rect 3650 1145 3710 1183
rect 3650 1111 3663 1145
rect 3697 1111 3710 1145
rect 3650 1075 3710 1111
rect 3650 1041 3663 1075
rect 3697 1041 3710 1075
rect 3650 1005 3710 1041
rect 3650 971 3663 1005
rect 3697 971 3710 1005
rect 3650 959 3710 971
rect 3740 1077 3800 1183
rect 3740 1043 3753 1077
rect 3787 1043 3800 1077
rect 3740 1005 3800 1043
rect 3740 971 3753 1005
rect 3787 971 3800 1005
rect 3740 959 3800 971
rect 3830 1145 3890 1183
rect 3830 1111 3843 1145
rect 3877 1111 3890 1145
rect 3830 1075 3890 1111
rect 3830 1041 3843 1075
rect 3877 1041 3890 1075
rect 3830 1005 3890 1041
rect 3830 971 3843 1005
rect 3877 971 3890 1005
rect 3830 959 3890 971
rect 3920 1145 3979 1183
rect 3920 1111 3933 1145
rect 3967 1111 3979 1145
rect 3920 1075 3979 1111
rect 3920 1041 3933 1075
rect 3967 1041 3979 1075
rect 3920 1005 3979 1041
rect 3920 971 3933 1005
rect 3967 971 3979 1005
rect 3920 959 3979 971
rect 4040 1171 4097 1183
rect 4040 1137 4050 1171
rect 4084 1137 4097 1171
rect 4040 1088 4097 1137
rect 4040 1054 4050 1088
rect 4084 1054 4097 1088
rect 4040 1005 4097 1054
rect 4040 971 4050 1005
rect 4084 971 4097 1005
rect 4040 959 4097 971
rect 4127 1171 4187 1183
rect 4127 1137 4140 1171
rect 4174 1137 4187 1171
rect 4127 1088 4187 1137
rect 4127 1054 4140 1088
rect 4174 1054 4187 1088
rect 4127 1005 4187 1054
rect 4127 971 4140 1005
rect 4174 971 4187 1005
rect 4127 959 4187 971
rect 4217 1145 4274 1183
rect 4217 1111 4230 1145
rect 4264 1111 4274 1145
rect 4217 1075 4274 1111
rect 4217 1041 4230 1075
rect 4264 1041 4274 1075
rect 4217 1005 4274 1041
rect 4217 971 4230 1005
rect 4264 971 4274 1005
rect 4217 959 4274 971
rect 3567 657 3626 669
rect 3567 623 3579 657
rect 3613 623 3626 657
rect 3567 587 3626 623
rect 3567 553 3579 587
rect 3613 553 3626 587
rect 3567 517 3626 553
rect 3567 483 3579 517
rect 3613 483 3626 517
rect 3567 445 3626 483
rect 3656 657 3716 669
rect 3656 623 3669 657
rect 3703 623 3716 657
rect 3656 587 3716 623
rect 3656 553 3669 587
rect 3703 553 3716 587
rect 3656 517 3716 553
rect 3656 483 3669 517
rect 3703 483 3716 517
rect 3656 445 3716 483
rect 3746 657 3806 669
rect 3746 623 3759 657
rect 3793 623 3806 657
rect 3746 585 3806 623
rect 3746 551 3759 585
rect 3793 551 3806 585
rect 3746 445 3806 551
rect 3836 657 3896 669
rect 3836 623 3849 657
rect 3883 623 3896 657
rect 3836 587 3896 623
rect 3836 553 3849 587
rect 3883 553 3896 587
rect 3836 517 3896 553
rect 3836 483 3849 517
rect 3883 483 3896 517
rect 3836 445 3896 483
rect 3926 657 3985 669
rect 3926 623 3939 657
rect 3973 623 3985 657
rect 3926 585 3985 623
rect 3926 551 3939 585
rect 3973 551 3985 585
rect 3926 445 3985 551
<< mvndiff >>
rect 475 1425 528 1443
rect 475 1391 483 1425
rect 517 1391 528 1425
rect 475 1357 528 1391
rect 209 1289 262 1327
rect 209 1255 217 1289
rect 251 1255 262 1289
rect 209 1243 262 1255
rect 362 1289 415 1327
rect 362 1255 373 1289
rect 407 1255 415 1289
rect 362 1243 415 1255
rect 475 1323 483 1357
rect 517 1323 528 1357
rect 475 1289 528 1323
rect 475 1255 483 1289
rect 517 1255 528 1289
rect 475 1243 528 1255
rect 708 1425 764 1443
rect 708 1391 719 1425
rect 753 1391 764 1425
rect 708 1357 764 1391
rect 708 1323 719 1357
rect 753 1323 764 1357
rect 708 1289 764 1323
rect 708 1255 719 1289
rect 753 1255 764 1289
rect 708 1243 764 1255
rect 944 1425 1000 1443
rect 944 1391 955 1425
rect 989 1391 1000 1425
rect 944 1357 1000 1391
rect 944 1323 955 1357
rect 989 1323 1000 1357
rect 944 1289 1000 1323
rect 944 1255 955 1289
rect 989 1255 1000 1289
rect 944 1243 1000 1255
rect 1180 1425 1236 1443
rect 1180 1391 1191 1425
rect 1225 1391 1236 1425
rect 1180 1357 1236 1391
rect 1180 1323 1191 1357
rect 1225 1323 1236 1357
rect 1180 1289 1236 1323
rect 1180 1255 1191 1289
rect 1225 1255 1236 1289
rect 1180 1243 1236 1255
rect 1416 1425 1472 1443
rect 1416 1391 1427 1425
rect 1461 1391 1472 1425
rect 1416 1357 1472 1391
rect 1416 1323 1427 1357
rect 1461 1323 1472 1357
rect 1416 1289 1472 1323
rect 1416 1255 1427 1289
rect 1461 1255 1472 1289
rect 1416 1243 1472 1255
rect 1652 1425 1708 1443
rect 1652 1391 1663 1425
rect 1697 1391 1708 1425
rect 1652 1357 1708 1391
rect 1652 1323 1663 1357
rect 1697 1323 1708 1357
rect 1652 1289 1708 1323
rect 1652 1255 1663 1289
rect 1697 1255 1708 1289
rect 1652 1243 1708 1255
rect 1888 1425 1944 1443
rect 1888 1391 1899 1425
rect 1933 1391 1944 1425
rect 1888 1357 1944 1391
rect 1888 1323 1899 1357
rect 1933 1323 1944 1357
rect 1888 1289 1944 1323
rect 1888 1255 1899 1289
rect 1933 1255 1944 1289
rect 1888 1243 1944 1255
rect 2124 1425 2180 1443
rect 2124 1391 2135 1425
rect 2169 1391 2180 1425
rect 2124 1357 2180 1391
rect 2124 1323 2135 1357
rect 2169 1323 2180 1357
rect 2124 1289 2180 1323
rect 2124 1255 2135 1289
rect 2169 1255 2180 1289
rect 2124 1243 2180 1255
rect 2360 1425 2413 1443
rect 2360 1391 2371 1425
rect 2405 1391 2413 1425
rect 2360 1357 2413 1391
rect 2360 1323 2371 1357
rect 2405 1323 2413 1357
rect 2774 1357 2827 1393
rect 2360 1289 2413 1323
rect 2360 1255 2371 1289
rect 2405 1255 2413 1289
rect 2360 1243 2413 1255
rect 2508 1289 2561 1327
rect 2508 1255 2516 1289
rect 2550 1255 2561 1289
rect 2508 1243 2561 1255
rect 2661 1289 2714 1327
rect 2661 1255 2672 1289
rect 2706 1255 2714 1289
rect 2661 1243 2714 1255
rect 2774 1323 2782 1357
rect 2816 1323 2827 1357
rect 2774 1289 2827 1323
rect 2774 1255 2782 1289
rect 2816 1255 2827 1289
rect 2774 1243 2827 1255
rect 2927 1357 2980 1393
rect 2927 1323 2938 1357
rect 2972 1323 2980 1357
rect 2927 1289 2980 1323
rect 2927 1255 2938 1289
rect 2972 1255 2980 1289
rect 2927 1243 2980 1255
rect 209 315 262 333
rect 209 281 217 315
rect 251 281 262 315
rect 209 247 262 281
rect 209 213 217 247
rect 251 213 262 247
rect 209 179 262 213
rect 209 145 217 179
rect 251 145 262 179
rect 209 133 262 145
rect 362 315 418 333
rect 362 281 373 315
rect 407 281 418 315
rect 362 247 418 281
rect 362 213 373 247
rect 407 213 418 247
rect 362 179 418 213
rect 362 145 373 179
rect 407 145 418 179
rect 362 133 418 145
rect 518 315 574 333
rect 518 281 529 315
rect 563 281 574 315
rect 518 247 574 281
rect 518 213 529 247
rect 563 213 574 247
rect 518 179 574 213
rect 518 145 529 179
rect 563 145 574 179
rect 518 133 574 145
rect 674 315 727 333
rect 674 281 685 315
rect 719 281 727 315
rect 674 247 727 281
rect 674 213 685 247
rect 719 213 727 247
rect 674 179 727 213
rect 674 145 685 179
rect 719 145 727 179
rect 674 133 727 145
rect 787 315 840 333
rect 787 281 795 315
rect 829 281 840 315
rect 787 247 840 281
rect 787 213 795 247
rect 829 213 840 247
rect 787 179 840 213
rect 787 145 795 179
rect 829 145 840 179
rect 787 133 840 145
rect 940 315 996 333
rect 940 281 951 315
rect 985 281 996 315
rect 940 247 996 281
rect 940 213 951 247
rect 985 213 996 247
rect 940 179 996 213
rect 940 145 951 179
rect 985 145 996 179
rect 940 133 996 145
rect 1096 315 1149 333
rect 1096 281 1107 315
rect 1141 281 1149 315
rect 1096 247 1149 281
rect 1096 213 1107 247
rect 1141 213 1149 247
rect 1096 179 1149 213
rect 1096 145 1107 179
rect 1141 145 1149 179
rect 1096 133 1149 145
<< mvpdiff >>
rect 209 1007 262 1085
rect 209 973 217 1007
rect 251 973 262 1007
rect 209 939 262 973
rect 209 905 217 939
rect 251 905 262 939
rect 209 871 262 905
rect 209 837 217 871
rect 251 837 262 871
rect 209 803 262 837
rect 209 769 217 803
rect 251 769 262 803
rect 209 735 262 769
rect 209 701 217 735
rect 251 701 262 735
rect 209 667 262 701
rect 209 633 217 667
rect 251 633 262 667
rect 209 599 262 633
rect 209 565 217 599
rect 251 565 262 599
rect 209 531 262 565
rect 209 497 217 531
rect 251 497 262 531
rect 209 485 262 497
rect 362 1007 418 1085
rect 362 973 373 1007
rect 407 973 418 1007
rect 362 939 418 973
rect 362 905 373 939
rect 407 905 418 939
rect 362 871 418 905
rect 362 837 373 871
rect 407 837 418 871
rect 362 803 418 837
rect 362 769 373 803
rect 407 769 418 803
rect 362 735 418 769
rect 362 701 373 735
rect 407 701 418 735
rect 362 667 418 701
rect 362 633 373 667
rect 407 633 418 667
rect 362 599 418 633
rect 362 565 373 599
rect 407 565 418 599
rect 362 531 418 565
rect 362 497 373 531
rect 407 497 418 531
rect 362 485 418 497
rect 518 1007 574 1085
rect 518 973 529 1007
rect 563 973 574 1007
rect 518 939 574 973
rect 518 905 529 939
rect 563 905 574 939
rect 518 871 574 905
rect 518 837 529 871
rect 563 837 574 871
rect 518 803 574 837
rect 518 769 529 803
rect 563 769 574 803
rect 518 735 574 769
rect 518 701 529 735
rect 563 701 574 735
rect 518 667 574 701
rect 518 633 529 667
rect 563 633 574 667
rect 518 599 574 633
rect 518 565 529 599
rect 563 565 574 599
rect 518 531 574 565
rect 518 497 529 531
rect 563 497 574 531
rect 518 485 574 497
rect 674 1007 727 1085
rect 674 973 685 1007
rect 719 973 727 1007
rect 674 939 727 973
rect 674 905 685 939
rect 719 905 727 939
rect 674 871 727 905
rect 674 837 685 871
rect 719 837 727 871
rect 674 803 727 837
rect 674 769 685 803
rect 719 769 727 803
rect 674 735 727 769
rect 674 701 685 735
rect 719 701 727 735
rect 674 667 727 701
rect 674 633 685 667
rect 719 633 727 667
rect 674 599 727 633
rect 674 565 685 599
rect 719 565 727 599
rect 674 531 727 565
rect 674 497 685 531
rect 719 497 727 531
rect 674 485 727 497
rect 787 735 840 785
rect 787 701 795 735
rect 829 701 840 735
rect 787 667 840 701
rect 787 633 795 667
rect 829 633 840 667
rect 787 599 840 633
rect 787 565 795 599
rect 829 565 840 599
rect 787 531 840 565
rect 787 497 795 531
rect 829 497 840 531
rect 787 485 840 497
rect 940 735 996 785
rect 940 701 951 735
rect 985 701 996 735
rect 940 667 996 701
rect 940 633 951 667
rect 985 633 996 667
rect 940 599 996 633
rect 940 565 951 599
rect 985 565 996 599
rect 940 531 996 565
rect 940 497 951 531
rect 985 497 996 531
rect 940 485 996 497
rect 1096 735 1149 785
rect 1096 701 1107 735
rect 1141 701 1149 735
rect 1096 667 1149 701
rect 1096 633 1107 667
rect 1141 633 1149 667
rect 1096 599 1149 633
rect 1096 565 1107 599
rect 1141 565 1149 599
rect 1096 531 1149 565
rect 1096 497 1107 531
rect 1141 497 1149 531
rect 1096 485 1149 497
rect 1257 821 1310 871
rect 1257 787 1265 821
rect 1299 787 1310 821
rect 1257 753 1310 787
rect 1257 719 1265 753
rect 1299 719 1310 753
rect 1257 685 1310 719
rect 1257 651 1265 685
rect 1299 651 1310 685
rect 1257 617 1310 651
rect 1257 583 1265 617
rect 1299 583 1310 617
rect 1257 571 1310 583
rect 1410 821 1466 871
rect 1410 787 1421 821
rect 1455 787 1466 821
rect 1410 753 1466 787
rect 1410 719 1421 753
rect 1455 719 1466 753
rect 1410 685 1466 719
rect 1410 651 1421 685
rect 1455 651 1466 685
rect 1410 617 1466 651
rect 1410 583 1421 617
rect 1455 583 1466 617
rect 1410 571 1466 583
rect 1566 821 1619 871
rect 1566 787 1577 821
rect 1611 787 1619 821
rect 1566 753 1619 787
rect 1566 719 1577 753
rect 1611 719 1619 753
rect 1566 685 1619 719
rect 1566 651 1577 685
rect 1611 651 1619 685
rect 1566 617 1619 651
rect 1566 583 1577 617
rect 1611 583 1619 617
rect 1566 571 1619 583
rect 2039 929 2092 1007
rect 2039 895 2047 929
rect 2081 895 2092 929
rect 2039 861 2092 895
rect 2039 827 2047 861
rect 2081 827 2092 861
rect 2039 793 2092 827
rect 2039 759 2047 793
rect 2081 759 2092 793
rect 2039 725 2092 759
rect 2039 691 2047 725
rect 2081 691 2092 725
rect 2039 657 2092 691
rect 2039 623 2047 657
rect 2081 623 2092 657
rect 2039 589 2092 623
rect 2039 555 2047 589
rect 2081 555 2092 589
rect 2039 521 2092 555
rect 2039 487 2047 521
rect 2081 487 2092 521
rect 2039 453 2092 487
rect 2039 419 2047 453
rect 2081 419 2092 453
rect 2039 407 2092 419
rect 2192 929 2248 1007
rect 2192 895 2203 929
rect 2237 895 2248 929
rect 2192 861 2248 895
rect 2192 827 2203 861
rect 2237 827 2248 861
rect 2192 793 2248 827
rect 2192 759 2203 793
rect 2237 759 2248 793
rect 2192 725 2248 759
rect 2192 691 2203 725
rect 2237 691 2248 725
rect 2192 657 2248 691
rect 2192 623 2203 657
rect 2237 623 2248 657
rect 2192 589 2248 623
rect 2192 555 2203 589
rect 2237 555 2248 589
rect 2192 521 2248 555
rect 2192 487 2203 521
rect 2237 487 2248 521
rect 2192 453 2248 487
rect 2192 419 2203 453
rect 2237 419 2248 453
rect 2192 407 2248 419
rect 2348 929 2404 1007
rect 2348 895 2359 929
rect 2393 895 2404 929
rect 2348 861 2404 895
rect 2348 827 2359 861
rect 2393 827 2404 861
rect 2348 793 2404 827
rect 2348 759 2359 793
rect 2393 759 2404 793
rect 2348 725 2404 759
rect 2348 691 2359 725
rect 2393 691 2404 725
rect 2348 657 2404 691
rect 2348 623 2359 657
rect 2393 623 2404 657
rect 2348 589 2404 623
rect 2348 555 2359 589
rect 2393 555 2404 589
rect 2348 521 2404 555
rect 2348 487 2359 521
rect 2393 487 2404 521
rect 2348 453 2404 487
rect 2348 419 2359 453
rect 2393 419 2404 453
rect 2348 407 2404 419
rect 2504 929 2560 1007
rect 2504 895 2515 929
rect 2549 895 2560 929
rect 2504 861 2560 895
rect 2504 827 2515 861
rect 2549 827 2560 861
rect 2504 793 2560 827
rect 2504 759 2515 793
rect 2549 759 2560 793
rect 2504 725 2560 759
rect 2504 691 2515 725
rect 2549 691 2560 725
rect 2504 657 2560 691
rect 2504 623 2515 657
rect 2549 623 2560 657
rect 2504 589 2560 623
rect 2504 555 2515 589
rect 2549 555 2560 589
rect 2504 521 2560 555
rect 2504 487 2515 521
rect 2549 487 2560 521
rect 2504 453 2560 487
rect 2504 419 2515 453
rect 2549 419 2560 453
rect 2504 407 2560 419
rect 2660 929 2713 1007
rect 2660 895 2671 929
rect 2705 895 2713 929
rect 2660 861 2713 895
rect 2660 827 2671 861
rect 2705 827 2713 861
rect 2774 971 2827 1007
rect 2774 937 2782 971
rect 2816 937 2827 971
rect 2774 903 2827 937
rect 2774 869 2782 903
rect 2816 869 2827 903
rect 2774 857 2827 869
rect 2927 971 2980 1007
rect 2927 937 2938 971
rect 2972 937 2980 971
rect 2927 903 2980 937
rect 2927 869 2938 903
rect 2972 869 2980 903
rect 2927 857 2980 869
rect 2660 793 2713 827
rect 2660 759 2671 793
rect 2705 759 2713 793
rect 2660 725 2713 759
rect 2660 691 2671 725
rect 2705 691 2713 725
rect 2660 657 2713 691
rect 2660 623 2671 657
rect 2705 623 2713 657
rect 2660 589 2713 623
rect 2660 555 2671 589
rect 2705 555 2713 589
rect 2660 521 2713 555
rect 2660 487 2671 521
rect 2705 487 2713 521
rect 2660 453 2713 487
rect 2660 419 2671 453
rect 2705 419 2713 453
rect 2660 407 2713 419
<< ndiffc >>
rect 3572 1415 3606 1449
rect 3658 1419 3692 1453
rect 3658 1341 3692 1375
rect 3754 1415 3788 1449
rect 3840 1419 3874 1453
rect 3840 1341 3874 1375
rect 3940 1431 3974 1465
rect 3940 1341 3974 1375
rect 4053 1431 4087 1465
rect 4053 1341 4087 1375
rect 4139 1419 4173 1453
rect 4139 1341 4173 1375
rect 4225 1431 4259 1465
rect 4225 1341 4259 1375
rect 3572 163 3606 197
rect 3672 253 3706 287
rect 3672 175 3706 209
rect 3758 179 3792 213
rect 3854 253 3888 287
rect 3854 175 3888 209
rect 3940 179 3974 213
<< pdiffc >>
rect 3573 1043 3607 1077
rect 3573 971 3607 1005
rect 3663 1111 3697 1145
rect 3663 1041 3697 1075
rect 3663 971 3697 1005
rect 3753 1043 3787 1077
rect 3753 971 3787 1005
rect 3843 1111 3877 1145
rect 3843 1041 3877 1075
rect 3843 971 3877 1005
rect 3933 1111 3967 1145
rect 3933 1041 3967 1075
rect 3933 971 3967 1005
rect 4050 1137 4084 1171
rect 4050 1054 4084 1088
rect 4050 971 4084 1005
rect 4140 1137 4174 1171
rect 4140 1054 4174 1088
rect 4140 971 4174 1005
rect 4230 1111 4264 1145
rect 4230 1041 4264 1075
rect 4230 971 4264 1005
rect 3579 623 3613 657
rect 3579 553 3613 587
rect 3579 483 3613 517
rect 3669 623 3703 657
rect 3669 553 3703 587
rect 3669 483 3703 517
rect 3759 623 3793 657
rect 3759 551 3793 585
rect 3849 623 3883 657
rect 3849 553 3883 587
rect 3849 483 3883 517
rect 3939 623 3973 657
rect 3939 551 3973 585
<< mvndiffc >>
rect 483 1391 517 1425
rect 217 1255 251 1289
rect 373 1255 407 1289
rect 483 1323 517 1357
rect 483 1255 517 1289
rect 719 1391 753 1425
rect 719 1323 753 1357
rect 719 1255 753 1289
rect 955 1391 989 1425
rect 955 1323 989 1357
rect 955 1255 989 1289
rect 1191 1391 1225 1425
rect 1191 1323 1225 1357
rect 1191 1255 1225 1289
rect 1427 1391 1461 1425
rect 1427 1323 1461 1357
rect 1427 1255 1461 1289
rect 1663 1391 1697 1425
rect 1663 1323 1697 1357
rect 1663 1255 1697 1289
rect 1899 1391 1933 1425
rect 1899 1323 1933 1357
rect 1899 1255 1933 1289
rect 2135 1391 2169 1425
rect 2135 1323 2169 1357
rect 2135 1255 2169 1289
rect 2371 1391 2405 1425
rect 2371 1323 2405 1357
rect 2371 1255 2405 1289
rect 2516 1255 2550 1289
rect 2672 1255 2706 1289
rect 2782 1323 2816 1357
rect 2782 1255 2816 1289
rect 2938 1323 2972 1357
rect 2938 1255 2972 1289
rect 217 281 251 315
rect 217 213 251 247
rect 217 145 251 179
rect 373 281 407 315
rect 373 213 407 247
rect 373 145 407 179
rect 529 281 563 315
rect 529 213 563 247
rect 529 145 563 179
rect 685 281 719 315
rect 685 213 719 247
rect 685 145 719 179
rect 795 281 829 315
rect 795 213 829 247
rect 795 145 829 179
rect 951 281 985 315
rect 951 213 985 247
rect 951 145 985 179
rect 1107 281 1141 315
rect 1107 213 1141 247
rect 1107 145 1141 179
<< mvpdiffc >>
rect 217 973 251 1007
rect 217 905 251 939
rect 217 837 251 871
rect 217 769 251 803
rect 217 701 251 735
rect 217 633 251 667
rect 217 565 251 599
rect 217 497 251 531
rect 373 973 407 1007
rect 373 905 407 939
rect 373 837 407 871
rect 373 769 407 803
rect 373 701 407 735
rect 373 633 407 667
rect 373 565 407 599
rect 373 497 407 531
rect 529 973 563 1007
rect 529 905 563 939
rect 529 837 563 871
rect 529 769 563 803
rect 529 701 563 735
rect 529 633 563 667
rect 529 565 563 599
rect 529 497 563 531
rect 685 973 719 1007
rect 685 905 719 939
rect 685 837 719 871
rect 685 769 719 803
rect 685 701 719 735
rect 685 633 719 667
rect 685 565 719 599
rect 685 497 719 531
rect 795 701 829 735
rect 795 633 829 667
rect 795 565 829 599
rect 795 497 829 531
rect 951 701 985 735
rect 951 633 985 667
rect 951 565 985 599
rect 951 497 985 531
rect 1107 701 1141 735
rect 1107 633 1141 667
rect 1107 565 1141 599
rect 1107 497 1141 531
rect 1265 787 1299 821
rect 1265 719 1299 753
rect 1265 651 1299 685
rect 1265 583 1299 617
rect 1421 787 1455 821
rect 1421 719 1455 753
rect 1421 651 1455 685
rect 1421 583 1455 617
rect 1577 787 1611 821
rect 1577 719 1611 753
rect 1577 651 1611 685
rect 1577 583 1611 617
rect 2047 895 2081 929
rect 2047 827 2081 861
rect 2047 759 2081 793
rect 2047 691 2081 725
rect 2047 623 2081 657
rect 2047 555 2081 589
rect 2047 487 2081 521
rect 2047 419 2081 453
rect 2203 895 2237 929
rect 2203 827 2237 861
rect 2203 759 2237 793
rect 2203 691 2237 725
rect 2203 623 2237 657
rect 2203 555 2237 589
rect 2203 487 2237 521
rect 2203 419 2237 453
rect 2359 895 2393 929
rect 2359 827 2393 861
rect 2359 759 2393 793
rect 2359 691 2393 725
rect 2359 623 2393 657
rect 2359 555 2393 589
rect 2359 487 2393 521
rect 2359 419 2393 453
rect 2515 895 2549 929
rect 2515 827 2549 861
rect 2515 759 2549 793
rect 2515 691 2549 725
rect 2515 623 2549 657
rect 2515 555 2549 589
rect 2515 487 2549 521
rect 2515 419 2549 453
rect 2671 895 2705 929
rect 2671 827 2705 861
rect 2782 937 2816 971
rect 2782 869 2816 903
rect 2938 937 2972 971
rect 2938 869 2972 903
rect 2671 759 2705 793
rect 2671 691 2705 725
rect 2671 623 2705 657
rect 2671 555 2705 589
rect 2671 487 2705 521
rect 2671 419 2705 453
<< nsubdiff >>
rect 3559 797 3589 831
rect 3623 797 3661 831
rect 3695 797 3726 831
<< mvpsubdiff >>
rect 0 1611 31 1645
rect 65 1611 127 1645
rect 161 1611 223 1645
rect 257 1611 319 1645
rect 353 1611 415 1645
rect 449 1611 511 1645
rect 545 1611 607 1645
rect 641 1611 703 1645
rect 737 1611 799 1645
rect 833 1611 895 1645
rect 929 1611 991 1645
rect 1025 1611 1087 1645
rect 1121 1611 1183 1645
rect 1217 1611 1279 1645
rect 1313 1611 1375 1645
rect 1409 1611 1471 1645
rect 1505 1611 1567 1645
rect 1601 1611 1663 1645
rect 1697 1611 1759 1645
rect 1793 1611 1855 1645
rect 1889 1611 1951 1645
rect 1985 1611 2047 1645
rect 2081 1611 2143 1645
rect 2177 1611 2239 1645
rect 2273 1611 2335 1645
rect 2369 1611 2431 1645
rect 2465 1611 2527 1645
rect 2561 1611 2623 1645
rect 2657 1611 2719 1645
rect 2753 1611 2815 1645
rect 2849 1611 2911 1645
rect 2945 1611 3007 1645
rect 3041 1611 3103 1645
rect 3137 1611 3199 1645
rect 3233 1611 3295 1645
rect 3329 1611 3391 1645
rect 3425 1611 3487 1645
rect 3521 1611 3583 1645
rect 3617 1611 3679 1645
rect 3713 1611 3775 1645
rect 3809 1611 3871 1645
rect 3905 1611 3967 1645
rect 4001 1611 4063 1645
rect 4097 1611 4159 1645
rect 4193 1611 4255 1645
rect 4289 1611 4351 1645
rect 4385 1611 4447 1645
rect 4481 1611 4543 1645
rect 4577 1611 4639 1645
rect 4673 1611 4735 1645
rect 4769 1611 4831 1645
rect 4865 1611 4927 1645
rect 4961 1611 4992 1645
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3679 17
rect 3713 -17 3775 17
rect 3809 -17 3871 17
rect 3905 -17 3967 17
rect 4001 -17 4063 17
rect 4097 -17 4159 17
rect 4193 -17 4255 17
rect 4289 -17 4351 17
rect 4385 -17 4447 17
rect 4481 -17 4543 17
rect 4577 -17 4639 17
rect 4673 -17 4735 17
rect 4769 -17 4831 17
rect 4865 -17 4927 17
rect 4961 -17 4992 17
<< mvnsubdiff >>
rect 72 992 106 1036
rect 72 831 106 958
rect 0 797 31 831
rect 65 797 137 831
rect 1827 797 1853 831
rect 1887 797 1925 831
rect 1959 797 1985 831
<< nsubdiffcont >>
rect 3589 797 3623 831
rect 3661 797 3695 831
<< mvpsubdiffcont >>
rect 31 1611 65 1645
rect 127 1611 161 1645
rect 223 1611 257 1645
rect 319 1611 353 1645
rect 415 1611 449 1645
rect 511 1611 545 1645
rect 607 1611 641 1645
rect 703 1611 737 1645
rect 799 1611 833 1645
rect 895 1611 929 1645
rect 991 1611 1025 1645
rect 1087 1611 1121 1645
rect 1183 1611 1217 1645
rect 1279 1611 1313 1645
rect 1375 1611 1409 1645
rect 1471 1611 1505 1645
rect 1567 1611 1601 1645
rect 1663 1611 1697 1645
rect 1759 1611 1793 1645
rect 1855 1611 1889 1645
rect 1951 1611 1985 1645
rect 2047 1611 2081 1645
rect 2143 1611 2177 1645
rect 2239 1611 2273 1645
rect 2335 1611 2369 1645
rect 2431 1611 2465 1645
rect 2527 1611 2561 1645
rect 2623 1611 2657 1645
rect 2719 1611 2753 1645
rect 2815 1611 2849 1645
rect 2911 1611 2945 1645
rect 3007 1611 3041 1645
rect 3103 1611 3137 1645
rect 3199 1611 3233 1645
rect 3295 1611 3329 1645
rect 3391 1611 3425 1645
rect 3487 1611 3521 1645
rect 3583 1611 3617 1645
rect 3679 1611 3713 1645
rect 3775 1611 3809 1645
rect 3871 1611 3905 1645
rect 3967 1611 4001 1645
rect 4063 1611 4097 1645
rect 4159 1611 4193 1645
rect 4255 1611 4289 1645
rect 4351 1611 4385 1645
rect 4447 1611 4481 1645
rect 4543 1611 4577 1645
rect 4639 1611 4673 1645
rect 4735 1611 4769 1645
rect 4831 1611 4865 1645
rect 4927 1611 4961 1645
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
rect 3391 -17 3425 17
rect 3487 -17 3521 17
rect 3583 -17 3617 17
rect 3679 -17 3713 17
rect 3775 -17 3809 17
rect 3871 -17 3905 17
rect 3967 -17 4001 17
rect 4063 -17 4097 17
rect 4159 -17 4193 17
rect 4255 -17 4289 17
rect 4351 -17 4385 17
rect 4447 -17 4481 17
rect 4543 -17 4577 17
rect 4639 -17 4673 17
rect 4735 -17 4769 17
rect 4831 -17 4865 17
rect 4927 -17 4961 17
<< mvnsubdiffcont >>
rect 72 958 106 992
rect 31 797 65 831
rect 1853 797 1887 831
rect 1925 797 1959 831
<< poly >>
rect 3617 1477 3647 1503
rect 3703 1477 3733 1503
rect 3799 1477 3829 1503
rect 3893 1477 3923 1503
rect 4098 1477 4128 1503
rect 4184 1477 4214 1503
rect 528 1443 708 1475
rect 764 1443 944 1475
rect 1000 1443 1180 1475
rect 1236 1443 1416 1475
rect 1472 1443 1652 1475
rect 1708 1443 1888 1475
rect 1944 1443 2124 1475
rect 2180 1443 2360 1475
rect 224 1420 362 1436
rect 224 1386 240 1420
rect 274 1386 308 1420
rect 342 1386 362 1420
rect 224 1370 362 1386
rect 262 1327 362 1370
rect 2827 1393 2927 1419
rect 2561 1327 2661 1353
rect 3617 1281 3647 1329
rect 3703 1281 3733 1329
rect 3799 1281 3829 1329
rect 3893 1281 3923 1329
rect 4098 1291 4128 1329
rect 4184 1291 4214 1329
rect 3617 1265 3923 1281
rect 262 1217 362 1243
rect 528 1211 708 1243
rect 764 1211 944 1243
rect 1000 1211 1180 1243
rect 1236 1211 1416 1243
rect 528 1171 1416 1211
rect 1472 1211 1652 1243
rect 1708 1211 1888 1243
rect 1944 1211 2124 1243
rect 2180 1211 2360 1243
rect 1472 1171 2360 1211
rect 1376 1129 1416 1171
rect 262 1085 362 1111
rect 418 1085 518 1111
rect 574 1085 674 1111
rect 1376 1089 1693 1129
rect 1183 1031 1611 1047
rect 1183 997 1489 1031
rect 1523 997 1557 1031
rect 1591 997 1611 1031
rect 1183 981 1611 997
rect 840 785 940 811
rect 996 785 1096 811
rect 262 426 362 485
rect 418 426 518 485
rect 574 439 674 485
rect 574 426 736 439
rect 262 423 736 426
rect 262 389 618 423
rect 652 389 686 423
rect 720 389 736 423
rect 262 386 736 389
rect 262 333 362 386
rect 418 333 518 386
rect 574 373 736 386
rect 840 422 940 485
rect 996 422 1096 485
rect 1183 422 1223 981
rect 1310 871 1410 981
rect 1466 871 1566 897
rect 1310 545 1410 571
rect 1466 503 1566 571
rect 1265 487 1566 503
rect 1265 453 1281 487
rect 1315 453 1349 487
rect 1383 453 1566 487
rect 1265 437 1566 453
rect 840 382 1223 422
rect 574 333 674 373
rect 840 333 940 382
rect 996 333 1096 382
rect 1653 225 1693 1089
rect 1753 307 1793 1171
rect 2561 1151 2661 1243
rect 2827 1175 2927 1243
rect 3617 1231 3669 1265
rect 3703 1231 3737 1265
rect 3771 1231 3805 1265
rect 3839 1231 3873 1265
rect 3907 1231 3923 1265
rect 3617 1215 3923 1231
rect 3617 1198 3653 1215
rect 3707 1198 3743 1215
rect 3797 1198 3833 1215
rect 3887 1198 3923 1215
rect 4094 1275 4280 1291
rect 4094 1261 4230 1275
rect 4094 1198 4130 1261
rect 4184 1241 4230 1261
rect 4264 1241 4280 1275
rect 4184 1225 4280 1241
rect 4184 1198 4220 1225
rect 3620 1183 3650 1198
rect 3710 1183 3740 1198
rect 3800 1183 3830 1198
rect 3890 1183 3920 1198
rect 4097 1183 4127 1198
rect 4187 1183 4217 1198
rect 2827 1159 2997 1175
rect 2561 1135 2752 1151
rect 2561 1129 2634 1135
rect 2092 1101 2634 1129
rect 2668 1101 2702 1135
rect 2736 1101 2752 1135
rect 2092 1085 2752 1101
rect 2827 1125 2879 1159
rect 2913 1125 2947 1159
rect 2981 1125 2997 1159
rect 2827 1109 2997 1125
rect 2092 1007 2192 1085
rect 2248 1007 2348 1085
rect 2404 1007 2504 1085
rect 2560 1007 2660 1085
rect 2827 1007 2927 1109
rect 3620 933 3650 959
rect 3710 933 3740 959
rect 3800 933 3830 959
rect 3890 933 3920 959
rect 4097 933 4127 959
rect 4187 933 4217 959
rect 2827 831 2927 857
rect 3626 669 3656 695
rect 3716 669 3746 695
rect 3806 669 3836 695
rect 3896 669 3926 695
rect 2793 441 2859 457
rect 2793 407 2809 441
rect 2843 407 2859 441
rect 3626 430 3656 445
rect 3716 430 3746 445
rect 3806 430 3836 445
rect 3896 430 3926 445
rect 3623 413 3659 430
rect 3713 413 3749 430
rect 3803 413 3839 430
rect 3893 413 3929 430
rect 2092 381 2192 407
rect 2248 381 2348 407
rect 2404 381 2504 407
rect 2560 381 2660 407
rect 2793 373 2859 407
rect 2793 339 2809 373
rect 2843 339 2859 373
rect 2793 307 2859 339
rect 1753 267 2859 307
rect 3493 397 3929 413
rect 3493 363 3639 397
rect 3673 363 3707 397
rect 3741 363 3775 397
rect 3809 363 3843 397
rect 3877 363 3929 397
rect 3493 347 3929 363
rect 3493 225 3533 347
rect 3623 299 3653 347
rect 3717 299 3747 347
rect 3813 299 3843 347
rect 3899 299 3929 347
rect 1653 184 3533 225
rect 262 107 362 133
rect 418 107 518 133
rect 574 107 674 133
rect 840 107 940 133
rect 996 107 1096 133
rect 3623 125 3653 151
rect 3717 125 3747 151
rect 3813 125 3843 151
rect 3899 125 3929 151
<< polycont >>
rect 240 1386 274 1420
rect 308 1386 342 1420
rect 1489 997 1523 1031
rect 1557 997 1591 1031
rect 618 389 652 423
rect 686 389 720 423
rect 1281 453 1315 487
rect 1349 453 1383 487
rect 3669 1231 3703 1265
rect 3737 1231 3771 1265
rect 3805 1231 3839 1265
rect 3873 1231 3907 1265
rect 4230 1241 4264 1275
rect 2634 1101 2668 1135
rect 2702 1101 2736 1135
rect 2879 1125 2913 1159
rect 2947 1125 2981 1159
rect 2809 407 2843 441
rect 2809 339 2843 373
rect 3639 363 3673 397
rect 3707 363 3741 397
rect 3775 363 3809 397
rect 3843 363 3877 397
<< locali >>
rect 0 1611 31 1645
rect 65 1611 127 1645
rect 161 1611 223 1645
rect 257 1611 319 1645
rect 353 1611 415 1645
rect 449 1611 511 1645
rect 545 1611 607 1645
rect 641 1611 703 1645
rect 737 1611 799 1645
rect 833 1611 895 1645
rect 929 1611 991 1645
rect 1025 1611 1087 1645
rect 1121 1611 1183 1645
rect 1217 1611 1279 1645
rect 1313 1611 1375 1645
rect 1409 1611 1471 1645
rect 1505 1611 1567 1645
rect 1601 1611 1663 1645
rect 1697 1611 1759 1645
rect 1793 1611 1855 1645
rect 1889 1611 1951 1645
rect 1985 1611 2047 1645
rect 2081 1611 2143 1645
rect 2177 1611 2239 1645
rect 2273 1611 2335 1645
rect 2369 1611 2431 1645
rect 2465 1611 2527 1645
rect 2561 1611 2623 1645
rect 2657 1611 2719 1645
rect 2753 1611 2815 1645
rect 2849 1611 2911 1645
rect 2945 1611 3007 1645
rect 3041 1611 3103 1645
rect 3137 1611 3199 1645
rect 3233 1611 3295 1645
rect 3329 1611 3391 1645
rect 3425 1611 3487 1645
rect 3521 1611 3583 1645
rect 3617 1611 3679 1645
rect 3713 1611 3775 1645
rect 3809 1611 3871 1645
rect 3905 1611 3967 1645
rect 4001 1611 4063 1645
rect 4097 1611 4159 1645
rect 4193 1611 4255 1645
rect 4289 1611 4351 1645
rect 4385 1611 4447 1645
rect 4481 1611 4543 1645
rect 4577 1611 4639 1645
rect 4673 1611 4735 1645
rect 4769 1611 4831 1645
rect 4865 1611 4927 1645
rect 4961 1611 4992 1645
rect 212 1554 2977 1560
rect 212 1520 223 1554
rect 257 1520 319 1554
rect 353 1520 415 1554
rect 449 1520 511 1554
rect 545 1520 607 1554
rect 641 1520 703 1554
rect 737 1520 799 1554
rect 833 1520 895 1554
rect 929 1520 991 1554
rect 1025 1520 1087 1554
rect 1121 1520 1183 1554
rect 1217 1520 1279 1554
rect 1313 1520 1375 1554
rect 1409 1520 1471 1554
rect 1505 1520 1567 1554
rect 1601 1520 1663 1554
rect 1697 1520 1759 1554
rect 1793 1520 1855 1554
rect 1889 1520 1951 1554
rect 1985 1520 2047 1554
rect 2081 1520 2143 1554
rect 2177 1520 2239 1554
rect 2273 1520 2335 1554
rect 2369 1520 2431 1554
rect 2465 1520 2527 1554
rect 2561 1520 2623 1554
rect 2657 1520 2718 1554
rect 2752 1520 2815 1554
rect 2849 1520 2911 1554
rect 2945 1520 2977 1554
rect 212 1514 2977 1520
rect 212 1436 256 1514
rect 472 1441 516 1514
rect 212 1420 362 1436
rect 212 1386 240 1420
rect 274 1386 308 1420
rect 342 1386 362 1420
rect 212 1370 362 1386
rect 472 1425 517 1441
rect 472 1391 483 1425
rect 212 1289 256 1370
rect 472 1357 517 1391
rect 472 1323 483 1357
rect 212 1255 217 1289
rect 251 1255 256 1289
rect 212 1239 256 1255
rect 368 1289 412 1305
rect 368 1255 373 1289
rect 407 1255 412 1289
rect 368 1195 412 1255
rect 472 1289 517 1323
rect 472 1255 483 1289
rect 472 1239 517 1255
rect 714 1425 758 1441
rect 714 1391 719 1425
rect 753 1391 758 1425
rect 714 1357 758 1391
rect 714 1323 719 1357
rect 753 1323 758 1357
rect 714 1289 758 1323
rect 714 1255 719 1289
rect 753 1255 758 1289
rect 714 1195 758 1255
rect 950 1425 994 1514
rect 950 1391 955 1425
rect 989 1391 994 1425
rect 950 1357 994 1391
rect 950 1323 955 1357
rect 989 1323 994 1357
rect 950 1289 994 1323
rect 950 1255 955 1289
rect 989 1255 994 1289
rect 950 1239 994 1255
rect 1186 1425 1230 1441
rect 1186 1391 1191 1425
rect 1225 1391 1230 1425
rect 1186 1357 1230 1391
rect 1186 1323 1191 1357
rect 1225 1323 1230 1357
rect 1186 1289 1230 1323
rect 1186 1255 1191 1289
rect 1225 1255 1230 1289
rect 1186 1195 1230 1255
rect 1422 1425 1466 1514
rect 1422 1391 1427 1425
rect 1461 1391 1466 1425
rect 1422 1357 1466 1391
rect 1422 1323 1427 1357
rect 1461 1323 1466 1357
rect 1422 1289 1466 1323
rect 1422 1255 1427 1289
rect 1461 1255 1466 1289
rect 1422 1239 1466 1255
rect 1658 1425 1702 1441
rect 1658 1391 1663 1425
rect 1697 1391 1702 1425
rect 1658 1357 1702 1391
rect 1658 1323 1663 1357
rect 1697 1323 1702 1357
rect 1658 1289 1702 1323
rect 1658 1255 1663 1289
rect 1697 1255 1702 1289
rect 1658 1195 1702 1255
rect 1894 1425 1938 1514
rect 1894 1391 1899 1425
rect 1933 1391 1938 1425
rect 1894 1357 1938 1391
rect 1894 1323 1899 1357
rect 1933 1323 1938 1357
rect 1894 1289 1938 1323
rect 1894 1255 1899 1289
rect 1933 1255 1938 1289
rect 1894 1239 1938 1255
rect 2130 1425 2174 1441
rect 2130 1391 2135 1425
rect 2169 1391 2174 1425
rect 2130 1357 2174 1391
rect 2130 1323 2135 1357
rect 2169 1323 2174 1357
rect 2130 1289 2174 1323
rect 2130 1255 2135 1289
rect 2169 1255 2174 1289
rect 2130 1195 2174 1255
rect 2366 1425 2410 1514
rect 2366 1391 2371 1425
rect 2405 1391 2410 1425
rect 2366 1357 2410 1391
rect 2366 1323 2371 1357
rect 2405 1323 2410 1357
rect 2366 1289 2410 1323
rect 2366 1255 2371 1289
rect 2405 1255 2410 1289
rect 2366 1239 2410 1255
rect 2511 1289 2555 1305
rect 2511 1255 2516 1289
rect 2550 1255 2555 1289
rect 2511 1195 2555 1255
rect 2667 1289 2711 1514
rect 2667 1255 2672 1289
rect 2706 1255 2711 1289
rect 2667 1239 2711 1255
rect 2777 1357 2821 1373
rect 2777 1323 2782 1357
rect 2816 1323 2821 1357
rect 2777 1289 2821 1323
rect 2777 1255 2782 1289
rect 2816 1255 2821 1289
rect 368 1151 1304 1195
rect 72 992 106 1036
rect 72 831 106 958
rect 212 1007 256 1023
rect 212 973 217 1007
rect 251 973 256 1007
rect 212 939 256 973
rect 212 905 217 939
rect 251 905 256 939
rect 367 1007 413 1023
rect 367 973 373 1007
rect 407 973 413 1007
rect 367 939 413 973
rect 367 925 373 939
rect 212 871 256 905
rect 331 919 373 925
rect 331 885 337 919
rect 371 905 373 919
rect 407 925 413 939
rect 524 1007 568 1023
rect 524 973 529 1007
rect 563 973 568 1007
rect 524 939 568 973
rect 407 919 449 925
rect 407 905 409 919
rect 371 885 409 905
rect 443 885 449 919
rect 331 879 449 885
rect 524 905 529 939
rect 563 905 568 939
rect 679 1007 725 1023
rect 679 973 685 1007
rect 719 973 725 1007
rect 679 939 725 973
rect 679 925 685 939
rect 212 837 217 871
rect 251 837 256 871
rect 0 797 31 831
rect 65 797 103 831
rect 212 803 256 837
rect 212 769 217 803
rect 251 769 256 803
rect 212 735 256 769
rect 212 701 217 735
rect 251 701 256 735
rect 212 667 256 701
rect 212 633 217 667
rect 251 633 256 667
rect 212 599 256 633
rect 212 565 217 599
rect 251 565 256 599
rect 212 531 256 565
rect 212 497 217 531
rect 251 497 256 531
rect 212 428 256 497
rect 367 871 413 879
rect 367 837 373 871
rect 407 837 413 871
rect 367 803 413 837
rect 367 769 373 803
rect 407 769 413 803
rect 367 735 413 769
rect 367 701 373 735
rect 407 701 413 735
rect 367 667 413 701
rect 367 633 373 667
rect 407 633 413 667
rect 367 599 413 633
rect 367 565 373 599
rect 407 565 413 599
rect 367 531 413 565
rect 367 497 373 531
rect 407 497 413 531
rect 367 481 413 497
rect 524 871 568 905
rect 643 919 685 925
rect 643 885 649 919
rect 683 905 685 919
rect 719 925 725 939
rect 719 919 761 925
rect 719 905 721 919
rect 683 885 721 905
rect 755 885 761 919
rect 643 879 761 885
rect 524 837 529 871
rect 563 837 568 871
rect 524 803 568 837
rect 524 769 529 803
rect 563 769 568 803
rect 524 735 568 769
rect 524 701 529 735
rect 563 701 568 735
rect 524 667 568 701
rect 524 633 529 667
rect 563 633 568 667
rect 524 599 568 633
rect 524 565 529 599
rect 563 565 568 599
rect 524 531 568 565
rect 524 497 529 531
rect 563 497 568 531
rect 524 428 568 497
rect 679 871 725 879
rect 679 837 685 871
rect 719 837 725 871
rect 679 803 725 837
rect 679 769 685 803
rect 719 769 725 803
rect 679 735 725 769
rect 1260 821 1304 1151
rect 1572 1151 2555 1195
rect 2777 1151 2821 1255
rect 2933 1357 2977 1514
rect 3556 1543 4275 1549
rect 3556 1509 3564 1543
rect 3598 1509 3660 1543
rect 3694 1509 3756 1543
rect 3790 1509 3852 1543
rect 3886 1509 3948 1543
rect 3982 1509 4044 1543
rect 4078 1509 4140 1543
rect 4174 1509 4236 1543
rect 4270 1509 4275 1543
rect 3556 1503 4275 1509
rect 3556 1449 3622 1503
rect 3556 1415 3572 1449
rect 3606 1415 3622 1449
rect 3556 1383 3622 1415
rect 3658 1453 3692 1469
rect 2933 1323 2938 1357
rect 2972 1323 2977 1357
rect 3658 1375 3692 1419
rect 3738 1449 3804 1503
rect 3738 1415 3754 1449
rect 3788 1415 3804 1449
rect 3738 1383 3804 1415
rect 3840 1453 3890 1469
rect 3874 1419 3890 1453
rect 2933 1289 2977 1323
rect 2933 1255 2938 1289
rect 2972 1255 2977 1289
rect 2933 1239 2977 1255
rect 3558 1341 3658 1349
rect 3840 1375 3890 1419
rect 3692 1341 3840 1349
rect 3874 1341 3890 1375
rect 3558 1315 3890 1341
rect 3924 1465 3990 1503
rect 3924 1431 3940 1465
rect 3974 1431 3990 1465
rect 3924 1375 3990 1431
rect 3924 1341 3940 1375
rect 3974 1341 3990 1375
rect 3924 1325 3990 1341
rect 4037 1465 4087 1503
rect 4037 1431 4053 1465
rect 4037 1375 4087 1431
rect 4037 1341 4053 1375
rect 4037 1325 4087 1341
rect 4123 1453 4189 1469
rect 4123 1419 4139 1453
rect 4173 1419 4189 1453
rect 4123 1375 4189 1419
rect 4123 1341 4139 1375
rect 4173 1341 4189 1375
rect 4123 1325 4189 1341
rect 4225 1465 4275 1503
rect 4259 1431 4275 1465
rect 4225 1375 4275 1431
rect 4259 1341 4275 1375
rect 4225 1325 4275 1341
rect 1572 1047 1616 1151
rect 2618 1135 2821 1151
rect 2618 1101 2634 1135
rect 2668 1101 2702 1135
rect 2736 1101 2821 1135
rect 2863 1159 2997 1175
rect 3558 1171 3604 1315
rect 4123 1281 4180 1325
rect 3653 1265 4180 1281
rect 3653 1231 3669 1265
rect 3703 1231 3737 1265
rect 3771 1231 3805 1265
rect 3839 1231 3873 1265
rect 3907 1237 4180 1265
rect 3907 1231 3988 1237
rect 3653 1195 3988 1231
rect 2863 1125 2879 1159
rect 2913 1125 2947 1159
rect 2981 1125 2997 1159
rect 2863 1109 2997 1125
rect 3432 1161 3604 1171
rect 4034 1171 4084 1187
rect 4034 1161 4050 1171
rect 3432 1145 3893 1161
rect 3432 1127 3663 1145
rect 2618 1085 2821 1101
rect 1469 1031 1616 1047
rect 1469 997 1489 1031
rect 1523 997 1557 1031
rect 1591 997 1616 1031
rect 1469 981 1616 997
rect 1260 787 1265 821
rect 1299 787 1304 821
rect 1260 753 1304 787
rect 679 701 685 735
rect 719 701 725 735
rect 679 667 725 701
rect 679 633 685 667
rect 719 633 725 667
rect 679 599 725 633
rect 679 565 685 599
rect 719 565 725 599
rect 679 531 725 565
rect 679 497 685 531
rect 719 497 725 531
rect 679 481 725 497
rect 790 735 834 751
rect 790 701 795 735
rect 829 701 834 735
rect 790 667 834 701
rect 790 633 795 667
rect 829 633 834 667
rect 790 599 834 633
rect 790 565 795 599
rect 829 565 834 599
rect 790 531 834 565
rect 790 497 795 531
rect 829 497 834 531
rect 790 439 834 497
rect 945 743 1062 751
rect 945 709 950 743
rect 984 735 1022 743
rect 985 709 1022 735
rect 1056 709 1062 743
rect 945 701 951 709
rect 985 703 1062 709
rect 1102 735 1146 751
rect 985 701 991 703
rect 945 667 991 701
rect 945 633 951 667
rect 985 633 991 667
rect 945 599 991 633
rect 945 565 951 599
rect 985 565 991 599
rect 945 531 991 565
rect 945 497 951 531
rect 985 497 991 531
rect 945 481 991 497
rect 1102 701 1107 735
rect 1141 701 1146 735
rect 1102 667 1146 701
rect 1102 633 1107 667
rect 1141 633 1146 667
rect 1102 599 1146 633
rect 1102 565 1107 599
rect 1141 565 1146 599
rect 1102 531 1146 565
rect 1102 497 1107 531
rect 1141 497 1146 531
rect 212 384 568 428
rect 212 315 256 384
rect 212 281 217 315
rect 251 281 256 315
rect 212 247 256 281
rect 212 213 217 247
rect 251 213 256 247
rect 212 179 256 213
rect 212 145 217 179
rect 251 145 256 179
rect 212 129 256 145
rect 367 315 413 331
rect 367 281 373 315
rect 407 281 413 315
rect 367 247 413 281
rect 367 213 373 247
rect 407 213 413 247
rect 367 179 413 213
rect 367 145 373 179
rect 407 145 413 179
rect 367 97 413 145
rect 524 315 568 384
rect 602 428 834 439
rect 1102 428 1146 497
rect 1260 719 1265 753
rect 1299 719 1304 753
rect 1260 685 1304 719
rect 1260 651 1265 685
rect 1299 651 1304 685
rect 1260 617 1304 651
rect 1260 583 1265 617
rect 1299 583 1304 617
rect 1260 503 1304 583
rect 1415 821 1461 869
rect 1415 787 1421 821
rect 1455 787 1461 821
rect 1415 753 1461 787
rect 1415 719 1421 753
rect 1455 719 1461 753
rect 1415 685 1461 719
rect 1415 651 1421 685
rect 1455 651 1461 685
rect 1415 617 1461 651
rect 1415 583 1421 617
rect 1455 613 1461 617
rect 1572 821 1616 981
rect 2042 1007 2710 1051
rect 2042 929 2086 1007
rect 2042 895 2047 929
rect 2081 895 2086 929
rect 2042 861 2086 895
rect 1572 787 1577 821
rect 1611 787 1616 821
rect 1827 797 1853 831
rect 1887 797 1925 831
rect 1959 797 1985 831
rect 2042 827 2047 861
rect 2081 827 2086 861
rect 1572 753 1616 787
rect 1572 719 1577 753
rect 1611 719 1616 753
rect 2042 793 2086 827
rect 2042 759 2047 793
rect 2081 759 2086 793
rect 2042 749 2086 759
rect 2198 929 2242 945
rect 2198 895 2203 929
rect 2237 895 2242 929
rect 2198 861 2242 895
rect 2198 827 2203 861
rect 2237 827 2242 861
rect 2198 793 2242 827
rect 2198 759 2203 793
rect 2237 759 2242 793
rect 1572 685 1616 719
rect 2005 743 2123 749
rect 2005 709 2011 743
rect 2045 725 2083 743
rect 2045 709 2047 725
rect 2005 703 2047 709
rect 1572 651 1577 685
rect 1611 651 1616 685
rect 1572 617 1616 651
rect 1455 583 1487 613
rect 1415 567 1487 583
rect 1572 583 1577 617
rect 1611 583 1616 617
rect 1572 567 1616 583
rect 2042 691 2047 703
rect 2081 709 2083 725
rect 2117 709 2123 743
rect 2081 703 2123 709
rect 2198 725 2242 759
rect 2354 929 2398 1007
rect 2354 895 2359 929
rect 2393 895 2398 929
rect 2354 861 2398 895
rect 2354 827 2359 861
rect 2393 827 2398 861
rect 2354 793 2398 827
rect 2354 759 2359 793
rect 2393 759 2398 793
rect 2354 749 2398 759
rect 2510 929 2554 945
rect 2510 895 2515 929
rect 2549 895 2554 929
rect 2510 861 2554 895
rect 2510 827 2515 861
rect 2549 827 2554 861
rect 2510 793 2554 827
rect 2510 759 2515 793
rect 2549 759 2554 793
rect 2081 691 2086 703
rect 2042 657 2086 691
rect 2042 623 2047 657
rect 2081 623 2086 657
rect 2042 589 2086 623
rect 1441 531 1487 567
rect 2042 555 2047 589
rect 2081 555 2086 589
rect 1260 487 1399 503
rect 1260 453 1281 487
rect 1315 453 1349 487
rect 1383 453 1399 487
rect 1441 485 1561 531
rect 1260 437 1399 453
rect 602 423 1146 428
rect 602 389 618 423
rect 652 389 686 423
rect 720 389 1146 423
rect 602 384 1146 389
rect 602 373 834 384
rect 524 281 529 315
rect 563 281 568 315
rect 524 247 568 281
rect 524 213 529 247
rect 563 213 568 247
rect 524 179 568 213
rect 524 145 529 179
rect 563 145 568 179
rect 524 129 568 145
rect 679 315 725 331
rect 679 281 685 315
rect 719 281 725 315
rect 679 247 725 281
rect 679 213 685 247
rect 719 213 725 247
rect 679 179 725 213
rect 679 145 685 179
rect 719 145 725 179
rect 679 97 725 145
rect 790 315 834 373
rect 790 281 795 315
rect 829 281 834 315
rect 790 247 834 281
rect 790 213 795 247
rect 829 213 834 247
rect 790 179 834 213
rect 790 145 795 179
rect 829 145 834 179
rect 790 129 834 145
rect 945 315 991 331
rect 945 281 951 315
rect 985 281 991 315
rect 945 247 991 281
rect 945 213 951 247
rect 985 213 991 247
rect 945 179 991 213
rect 945 145 951 179
rect 985 145 991 179
rect 945 97 991 145
rect 1102 315 1146 384
rect 1515 361 1561 485
rect 2042 521 2086 555
rect 2042 487 2047 521
rect 2081 487 2086 521
rect 2042 453 2086 487
rect 2042 419 2047 453
rect 2081 419 2086 453
rect 2042 403 2086 419
rect 2198 691 2203 725
rect 2237 691 2242 725
rect 2317 743 2435 749
rect 2317 709 2323 743
rect 2357 725 2395 743
rect 2357 709 2359 725
rect 2317 703 2359 709
rect 2198 657 2242 691
rect 2198 623 2203 657
rect 2237 623 2242 657
rect 2198 589 2242 623
rect 2198 555 2203 589
rect 2237 555 2242 589
rect 2198 521 2242 555
rect 2198 487 2203 521
rect 2237 487 2242 521
rect 2198 453 2242 487
rect 2198 419 2203 453
rect 2237 419 2242 453
rect 2198 361 2242 419
rect 2354 691 2359 703
rect 2393 709 2395 725
rect 2429 709 2435 743
rect 2393 703 2435 709
rect 2510 725 2554 759
rect 2666 929 2710 1007
rect 2666 895 2671 929
rect 2705 895 2710 929
rect 2666 861 2710 895
rect 2666 827 2671 861
rect 2705 827 2710 861
rect 2777 971 2821 1085
rect 2777 937 2782 971
rect 2816 937 2821 971
rect 2777 903 2821 937
rect 2931 971 2977 1011
rect 2931 937 2938 971
rect 2972 937 2977 971
rect 2931 925 2977 937
rect 2777 869 2782 903
rect 2816 869 2821 903
rect 2859 919 2977 925
rect 2859 885 2865 919
rect 2899 885 2937 919
rect 2971 903 2977 919
rect 2859 879 2938 885
rect 2777 853 2821 869
rect 2931 869 2938 879
rect 2972 869 2977 903
rect 2931 853 2977 869
rect 2666 793 2710 827
rect 2666 759 2671 793
rect 2705 759 2710 793
rect 2666 749 2710 759
rect 2393 691 2398 703
rect 2354 657 2398 691
rect 2354 623 2359 657
rect 2393 623 2398 657
rect 2354 589 2398 623
rect 2354 555 2359 589
rect 2393 555 2398 589
rect 2354 521 2398 555
rect 2354 487 2359 521
rect 2393 487 2398 521
rect 2354 453 2398 487
rect 2354 419 2359 453
rect 2393 419 2398 453
rect 2354 403 2398 419
rect 2510 691 2515 725
rect 2549 691 2554 725
rect 2629 743 2747 749
rect 2629 709 2635 743
rect 2669 725 2707 743
rect 2669 709 2671 725
rect 2629 703 2671 709
rect 2510 657 2554 691
rect 2510 623 2515 657
rect 2549 623 2554 657
rect 2510 589 2554 623
rect 2510 555 2515 589
rect 2549 555 2554 589
rect 2510 521 2554 555
rect 2510 487 2515 521
rect 2549 487 2554 521
rect 2510 453 2554 487
rect 2510 419 2515 453
rect 2549 419 2554 453
rect 2510 361 2554 419
rect 2666 691 2671 703
rect 2705 709 2707 725
rect 2741 709 2747 743
rect 2705 703 2747 709
rect 2705 691 2710 703
rect 2666 657 2710 691
rect 2666 623 2671 657
rect 2705 623 2710 657
rect 2666 589 2710 623
rect 2666 555 2671 589
rect 2705 555 2710 589
rect 2666 521 2710 555
rect 2666 487 2671 521
rect 2705 487 2710 521
rect 2666 453 2710 487
rect 2666 419 2671 453
rect 2705 419 2710 453
rect 2666 403 2710 419
rect 2793 441 2859 457
rect 2793 407 2809 441
rect 2843 407 2859 441
rect 1515 317 2554 361
rect 2793 373 2859 407
rect 2793 339 2809 373
rect 2843 339 2859 373
rect 3432 433 3476 1127
rect 3647 1111 3663 1127
rect 3697 1127 3843 1145
rect 3697 1111 3713 1127
rect 3557 1077 3607 1093
rect 3557 1043 3573 1077
rect 3557 1005 3607 1043
rect 3557 971 3573 1005
rect 3557 921 3607 971
rect 3647 1075 3713 1111
rect 3827 1111 3843 1127
rect 3877 1111 3893 1145
rect 3647 1041 3663 1075
rect 3697 1041 3713 1075
rect 3647 1005 3713 1041
rect 3647 971 3663 1005
rect 3697 971 3713 1005
rect 3647 955 3713 971
rect 3753 1077 3787 1093
rect 3753 1005 3787 1043
rect 3753 921 3787 971
rect 3827 1075 3893 1111
rect 3827 1041 3843 1075
rect 3877 1041 3893 1075
rect 3827 1005 3893 1041
rect 3827 971 3843 1005
rect 3877 971 3893 1005
rect 3827 955 3893 971
rect 3933 1145 4050 1161
rect 3967 1137 4050 1145
rect 3967 1111 4084 1137
rect 3933 1088 4084 1111
rect 3933 1075 4050 1088
rect 3967 1054 4050 1075
rect 3967 1041 4084 1054
rect 3933 1005 4084 1041
rect 3967 971 4050 1005
rect 3933 921 4084 971
rect 4123 1171 4180 1237
rect 4214 1275 4280 1291
rect 4214 1241 4230 1275
rect 4264 1241 4280 1275
rect 4214 1195 4280 1241
rect 4123 1137 4140 1171
rect 4174 1137 4180 1171
rect 4123 1088 4180 1137
rect 4123 1054 4140 1088
rect 4174 1054 4180 1088
rect 4123 1005 4180 1054
rect 4123 971 4140 1005
rect 4174 971 4180 1005
rect 4123 955 4180 971
rect 4214 1145 4280 1161
rect 4214 1111 4230 1145
rect 4264 1111 4280 1145
rect 4214 1075 4280 1111
rect 4214 1041 4230 1075
rect 4264 1041 4280 1075
rect 4214 1005 4280 1041
rect 4214 971 4230 1005
rect 4264 971 4280 1005
rect 4214 921 4280 971
rect 3557 887 4280 921
rect 3933 847 4084 887
rect 3559 831 4084 847
rect 3559 797 3589 831
rect 3623 797 3661 831
rect 3695 797 4084 831
rect 3559 781 4084 797
rect 3933 741 4084 781
rect 3563 707 4084 741
rect 3563 657 3613 707
rect 3563 623 3579 657
rect 3563 587 3613 623
rect 3563 553 3579 587
rect 3563 517 3613 553
rect 3563 483 3579 517
rect 3563 467 3613 483
rect 3653 657 3719 673
rect 3653 623 3669 657
rect 3703 623 3719 657
rect 3653 587 3719 623
rect 3653 553 3669 587
rect 3703 553 3719 587
rect 3653 517 3719 553
rect 3759 657 3793 707
rect 3759 585 3793 623
rect 3759 535 3793 551
rect 3833 657 3899 673
rect 3833 623 3849 657
rect 3883 623 3899 657
rect 3833 587 3899 623
rect 3833 553 3849 587
rect 3883 553 3899 587
rect 3653 483 3669 517
rect 3703 501 3719 517
rect 3833 517 3899 553
rect 3939 657 4084 707
rect 3973 648 4084 657
rect 3939 614 3960 623
rect 3994 614 4032 648
rect 4066 614 4084 648
rect 3939 604 4084 614
rect 3939 585 3989 604
rect 3973 551 3989 585
rect 3939 535 3989 551
rect 3833 501 3849 517
rect 3703 483 3849 501
rect 3883 501 3899 517
rect 3883 483 3988 501
rect 3653 467 3988 483
rect 3432 397 3893 433
rect 3432 363 3639 397
rect 3673 363 3707 397
rect 3741 363 3775 397
rect 3809 363 3843 397
rect 3877 363 3893 397
rect 3432 347 3893 363
rect 1102 281 1107 315
rect 1141 281 1146 315
rect 1102 247 1146 281
rect 2793 313 2859 339
rect 3942 313 3988 467
rect 2793 287 3988 313
rect 2793 269 3672 287
rect 1102 213 1107 247
rect 1141 213 1146 247
rect 3656 253 3672 269
rect 3706 279 3854 287
rect 1102 179 1146 213
rect 1102 145 1107 179
rect 1141 145 1146 179
rect 1102 129 1146 145
rect 3556 197 3622 235
rect 3556 163 3572 197
rect 3606 163 3622 197
rect 3556 125 3622 163
rect 3656 209 3706 253
rect 3888 279 3988 287
rect 3656 175 3672 209
rect 3656 159 3706 175
rect 3742 213 3808 245
rect 3742 179 3758 213
rect 3792 179 3808 213
rect 3742 125 3808 179
rect 3854 209 3888 253
rect 3854 159 3888 175
rect 3924 213 3990 245
rect 3924 179 3940 213
rect 3974 179 3990 213
rect 3924 125 3990 179
rect 3556 119 3990 125
rect 367 91 485 97
rect 367 57 373 91
rect 407 57 445 91
rect 479 57 485 91
rect 367 51 485 57
rect 607 91 725 97
rect 607 57 613 91
rect 647 57 685 91
rect 719 57 725 91
rect 607 51 725 57
rect 909 91 1027 97
rect 909 57 915 91
rect 949 57 987 91
rect 1021 57 1027 91
rect 3556 85 3564 119
rect 3598 85 3660 119
rect 3694 85 3756 119
rect 3790 85 3852 119
rect 3886 85 3948 119
rect 3982 85 3990 119
rect 3556 79 3990 85
rect 909 51 1027 57
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3679 17
rect 3713 -17 3775 17
rect 3809 -17 3871 17
rect 3905 -17 3967 17
rect 4001 -17 4063 17
rect 4097 -17 4159 17
rect 4193 -17 4255 17
rect 4289 -17 4351 17
rect 4385 -17 4447 17
rect 4481 -17 4543 17
rect 4577 -17 4639 17
rect 4673 -17 4735 17
rect 4769 -17 4831 17
rect 4865 -17 4927 17
rect 4961 -17 4992 17
<< viali >>
rect 31 1611 65 1645
rect 127 1611 161 1645
rect 223 1611 257 1645
rect 319 1611 353 1645
rect 415 1611 449 1645
rect 511 1611 545 1645
rect 607 1611 641 1645
rect 703 1611 737 1645
rect 799 1611 833 1645
rect 895 1611 929 1645
rect 991 1611 1025 1645
rect 1087 1611 1121 1645
rect 1183 1611 1217 1645
rect 1279 1611 1313 1645
rect 1375 1611 1409 1645
rect 1471 1611 1505 1645
rect 1567 1611 1601 1645
rect 1663 1611 1697 1645
rect 1759 1611 1793 1645
rect 1855 1611 1889 1645
rect 1951 1611 1985 1645
rect 2047 1611 2081 1645
rect 2143 1611 2177 1645
rect 2239 1611 2273 1645
rect 2335 1611 2369 1645
rect 2431 1611 2465 1645
rect 2527 1611 2561 1645
rect 2623 1611 2657 1645
rect 2719 1611 2753 1645
rect 2815 1611 2849 1645
rect 2911 1611 2945 1645
rect 3007 1611 3041 1645
rect 3103 1611 3137 1645
rect 3199 1611 3233 1645
rect 3295 1611 3329 1645
rect 3391 1611 3425 1645
rect 3487 1611 3521 1645
rect 3583 1611 3617 1645
rect 3679 1611 3713 1645
rect 3775 1611 3809 1645
rect 3871 1611 3905 1645
rect 3967 1611 4001 1645
rect 4063 1611 4097 1645
rect 4159 1611 4193 1645
rect 4255 1611 4289 1645
rect 4351 1611 4385 1645
rect 4447 1611 4481 1645
rect 4543 1611 4577 1645
rect 4639 1611 4673 1645
rect 4735 1611 4769 1645
rect 4831 1611 4865 1645
rect 4927 1611 4961 1645
rect 223 1520 257 1554
rect 319 1520 353 1554
rect 415 1520 449 1554
rect 511 1520 545 1554
rect 607 1520 641 1554
rect 703 1520 737 1554
rect 799 1520 833 1554
rect 895 1520 929 1554
rect 991 1520 1025 1554
rect 1087 1520 1121 1554
rect 1183 1520 1217 1554
rect 1279 1520 1313 1554
rect 1375 1520 1409 1554
rect 1471 1520 1505 1554
rect 1567 1520 1601 1554
rect 1663 1520 1697 1554
rect 1759 1520 1793 1554
rect 1855 1520 1889 1554
rect 1951 1520 1985 1554
rect 2047 1520 2081 1554
rect 2143 1520 2177 1554
rect 2239 1520 2273 1554
rect 2335 1520 2369 1554
rect 2431 1520 2465 1554
rect 2527 1520 2561 1554
rect 2623 1520 2657 1554
rect 2718 1520 2752 1554
rect 2815 1520 2849 1554
rect 2911 1520 2945 1554
rect 337 885 371 919
rect 409 885 443 919
rect 31 797 65 831
rect 103 797 137 831
rect 649 885 683 919
rect 721 885 755 919
rect 3564 1509 3598 1543
rect 3660 1509 3694 1543
rect 3756 1509 3790 1543
rect 3852 1509 3886 1543
rect 3948 1509 3982 1543
rect 4044 1509 4078 1543
rect 4140 1509 4174 1543
rect 4236 1509 4270 1543
rect 950 735 984 743
rect 950 709 951 735
rect 951 709 984 735
rect 1022 709 1056 743
rect 1853 797 1887 831
rect 1925 797 1959 831
rect 2011 709 2045 743
rect 2083 709 2117 743
rect 2323 709 2357 743
rect 2395 709 2429 743
rect 2865 885 2899 919
rect 2937 903 2971 919
rect 2937 885 2938 903
rect 2938 885 2971 903
rect 2635 709 2669 743
rect 2707 709 2741 743
rect 3960 623 3973 648
rect 3973 623 3994 648
rect 3960 614 3994 623
rect 4032 614 4066 648
rect 373 57 407 91
rect 445 57 479 91
rect 613 57 647 91
rect 685 57 719 91
rect 915 57 949 91
rect 987 57 1021 91
rect 3564 85 3598 119
rect 3660 85 3694 119
rect 3756 85 3790 119
rect 3852 85 3886 119
rect 3948 85 3982 119
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
rect 1663 -17 1697 17
rect 1759 -17 1793 17
rect 1855 -17 1889 17
rect 1951 -17 1985 17
rect 2047 -17 2081 17
rect 2143 -17 2177 17
rect 2239 -17 2273 17
rect 2335 -17 2369 17
rect 2431 -17 2465 17
rect 2527 -17 2561 17
rect 2623 -17 2657 17
rect 2719 -17 2753 17
rect 2815 -17 2849 17
rect 2911 -17 2945 17
rect 3007 -17 3041 17
rect 3103 -17 3137 17
rect 3199 -17 3233 17
rect 3295 -17 3329 17
rect 3391 -17 3425 17
rect 3487 -17 3521 17
rect 3583 -17 3617 17
rect 3679 -17 3713 17
rect 3775 -17 3809 17
rect 3871 -17 3905 17
rect 3967 -17 4001 17
rect 4063 -17 4097 17
rect 4159 -17 4193 17
rect 4255 -17 4289 17
rect 4351 -17 4385 17
rect 4447 -17 4481 17
rect 4543 -17 4577 17
rect 4639 -17 4673 17
rect 4735 -17 4769 17
rect 4831 -17 4865 17
rect 4927 -17 4961 17
<< metal1 >>
rect 0 1645 4992 1651
rect 0 1611 31 1645
rect 65 1611 127 1645
rect 161 1611 223 1645
rect 257 1611 319 1645
rect 353 1611 415 1645
rect 449 1611 511 1645
rect 545 1611 607 1645
rect 641 1611 703 1645
rect 737 1611 799 1645
rect 833 1611 895 1645
rect 929 1611 991 1645
rect 1025 1611 1087 1645
rect 1121 1611 1183 1645
rect 1217 1611 1279 1645
rect 1313 1611 1375 1645
rect 1409 1611 1471 1645
rect 1505 1611 1567 1645
rect 1601 1611 1663 1645
rect 1697 1611 1759 1645
rect 1793 1611 1855 1645
rect 1889 1611 1951 1645
rect 1985 1611 2047 1645
rect 2081 1611 2143 1645
rect 2177 1611 2239 1645
rect 2273 1611 2335 1645
rect 2369 1611 2431 1645
rect 2465 1611 2527 1645
rect 2561 1611 2623 1645
rect 2657 1611 2719 1645
rect 2753 1611 2815 1645
rect 2849 1611 2911 1645
rect 2945 1611 3007 1645
rect 3041 1611 3103 1645
rect 3137 1611 3199 1645
rect 3233 1611 3295 1645
rect 3329 1611 3391 1645
rect 3425 1611 3487 1645
rect 3521 1611 3583 1645
rect 3617 1611 3679 1645
rect 3713 1611 3775 1645
rect 3809 1611 3871 1645
rect 3905 1611 3967 1645
rect 4001 1611 4063 1645
rect 4097 1611 4159 1645
rect 4193 1611 4255 1645
rect 4289 1611 4351 1645
rect 4385 1611 4447 1645
rect 4481 1611 4543 1645
rect 4577 1611 4639 1645
rect 4673 1611 4735 1645
rect 4769 1611 4831 1645
rect 4865 1611 4927 1645
rect 4961 1611 4992 1645
rect 0 1605 4992 1611
rect 0 1554 4992 1577
rect 0 1520 223 1554
rect 257 1520 319 1554
rect 353 1520 415 1554
rect 449 1520 511 1554
rect 545 1520 607 1554
rect 641 1520 703 1554
rect 737 1520 799 1554
rect 833 1520 895 1554
rect 929 1520 991 1554
rect 1025 1520 1087 1554
rect 1121 1520 1183 1554
rect 1217 1520 1279 1554
rect 1313 1520 1375 1554
rect 1409 1520 1471 1554
rect 1505 1520 1567 1554
rect 1601 1520 1663 1554
rect 1697 1520 1759 1554
rect 1793 1520 1855 1554
rect 1889 1520 1951 1554
rect 1985 1520 2047 1554
rect 2081 1520 2143 1554
rect 2177 1520 2239 1554
rect 2273 1520 2335 1554
rect 2369 1520 2431 1554
rect 2465 1520 2527 1554
rect 2561 1520 2623 1554
rect 2657 1520 2718 1554
rect 2752 1520 2815 1554
rect 2849 1520 2911 1554
rect 2945 1543 4992 1554
rect 2945 1520 3564 1543
rect 0 1509 3564 1520
rect 3598 1509 3660 1543
rect 3694 1509 3756 1543
rect 3790 1509 3852 1543
rect 3886 1509 3948 1543
rect 3982 1509 4044 1543
rect 4078 1509 4140 1543
rect 4174 1509 4236 1543
rect 4270 1509 4992 1543
rect 0 1503 4992 1509
rect 0 919 4992 939
rect 0 885 337 919
rect 371 885 409 919
rect 443 885 649 919
rect 683 885 721 919
rect 755 885 2865 919
rect 2899 885 2937 919
rect 2971 885 4992 919
rect 0 865 4992 885
rect 0 831 4992 837
rect 0 797 31 831
rect 65 797 103 831
rect 137 797 1853 831
rect 1887 797 1925 831
rect 1959 797 4992 831
rect 0 791 4992 797
rect 0 743 4992 763
rect 0 709 950 743
rect 984 709 1022 743
rect 1056 709 2011 743
rect 2045 709 2083 743
rect 2117 709 2323 743
rect 2357 709 2395 743
rect 2429 709 2635 743
rect 2669 709 2707 743
rect 2741 709 4992 743
rect 0 689 4992 709
rect 14 648 4978 661
rect 14 614 3960 648
rect 3994 614 4032 648
rect 4066 614 4978 648
rect 14 604 4978 614
rect 0 119 4992 125
rect 0 91 3564 119
rect 0 57 373 91
rect 407 57 445 91
rect 479 57 613 91
rect 647 57 685 91
rect 719 57 915 91
rect 949 57 987 91
rect 1021 85 3564 91
rect 3598 85 3660 119
rect 3694 85 3756 119
rect 3790 85 3852 119
rect 3886 85 3948 119
rect 3982 85 4992 119
rect 1021 57 4992 85
rect 0 51 4992 57
rect 0 17 4992 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1663 17
rect 1697 -17 1759 17
rect 1793 -17 1855 17
rect 1889 -17 1951 17
rect 1985 -17 2047 17
rect 2081 -17 2143 17
rect 2177 -17 2239 17
rect 2273 -17 2335 17
rect 2369 -17 2431 17
rect 2465 -17 2527 17
rect 2561 -17 2623 17
rect 2657 -17 2719 17
rect 2753 -17 2815 17
rect 2849 -17 2911 17
rect 2945 -17 3007 17
rect 3041 -17 3103 17
rect 3137 -17 3199 17
rect 3233 -17 3295 17
rect 3329 -17 3391 17
rect 3425 -17 3487 17
rect 3521 -17 3583 17
rect 3617 -17 3679 17
rect 3713 -17 3775 17
rect 3809 -17 3871 17
rect 3905 -17 3967 17
rect 4001 -17 4063 17
rect 4097 -17 4159 17
rect 4193 -17 4255 17
rect 4289 -17 4351 17
rect 4385 -17 4447 17
rect 4481 -17 4543 17
rect 4577 -17 4639 17
rect 4673 -17 4735 17
rect 4769 -17 4831 17
rect 4865 -17 4927 17
rect 4961 -17 4992 17
rect 0 -23 4992 -17
<< labels >>
flabel locali s 2913 1125 2947 1159 0 FreeSans 400 0 0 0 SLEEP_B
port 2 nsew signal input
flabel locali s 4230 1241 4264 1275 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 217 396 251 430 0 FreeSans 400 90 0 0 X
port 8 nsew signal output
flabel metal1 s 0 1605 4992 1628 0 FreeSans 340 0 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 0 0 4992 23 0 FreeSans 340 0 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 0 51 4992 125 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel metal1 s 0 1503 4992 1577 0 FreeSans 340 0 0 0 VGND
port 4 nsew ground bidirectional
flabel metal1 s 0 791 4992 837 0 FreeSans 520 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 0 865 4992 939 0 FreeSans 520 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 0 689 4992 763 0 FreeSans 520 0 0 0 VPWR
port 7 nsew power bidirectional
flabel metal1 s 14 604 4978 661 0 FreeSans 520 0 0 0 LVPWR
port 3 nsew power bidirectional
flabel comment s 812 616 812 616 0 FreeSans 300 180 0 0 D
flabel comment s 968 616 968 616 0 FreeSans 300 180 0 0 S
flabel comment s 1124 616 1124 616 0 FreeSans 300 180 0 0 D
flabel comment s 500 1340 500 1340 0 FreeSans 300 0 0 0 S
flabel comment s 854 1340 854 1340 0 FreeSans 200 0 0 0 I16
flabel comment s 736 1340 736 1340 0 FreeSans 300 0 0 0 D
flabel comment s 890 616 890 616 0 FreeSans 200 0 0 0 I46
flabel comment s 2132 504 2132 504 0 FreeSans 200 0 0 0 I23
flabel comment s 1046 616 1046 616 0 FreeSans 200 0 0 0 I46
flabel comment s 890 230 890 230 0 FreeSans 200 0 0 0 I45
flabel comment s 2444 504 2444 504 0 FreeSans 200 0 0 0 I23
rlabel comment s 4301 1551 4301 1551 4 inv_2
rlabel comment s 4013 1551 4013 1551 4 inv_4
flabel comment s 1326 1340 1326 1340 0 FreeSans 200 0 0 0 I16
rlabel comment s 3533 77 3533 77 4 inv_4
flabel comment s 2710 288 2710 288 0 FreeSans 400 0 0 0 t4
flabel comment s 1090 1340 1090 1340 0 FreeSans 200 0 0 0 I16
flabel comment s 312 752 312 752 0 FreeSans 200 0 0 0 I48
flabel comment s 2270 1340 2270 1340 0 FreeSans 200 0 0 0 I15
flabel comment s 2034 1340 2034 1340 0 FreeSans 200 0 0 0 I15
flabel comment s 2288 504 2288 504 0 FreeSans 200 0 0 0 I23
flabel comment s 1798 1340 1798 1340 0 FreeSans 200 0 0 0 I15
flabel comment s 468 752 468 752 0 FreeSans 200 0 0 0 I48
flabel comment s 624 230 624 230 0 FreeSans 200 0 0 0 I47
flabel comment s 468 230 468 230 0 FreeSans 200 0 0 0 I47
flabel comment s 1562 1340 1562 1340 0 FreeSans 200 0 0 0 I15
flabel comment s 1516 702 1516 702 0 FreeSans 200 0 0 0 M3
flabel comment s 2647 1272 2647 1272 0 FreeSans 200 0 0 0 M9
flabel comment s 1444 1340 1444 1340 0 FreeSans 300 0 0 0 S
flabel comment s 1360 702 1360 702 0 FreeSans 200 0 0 0 M4
flabel comment s 2600 504 2600 504 0 FreeSans 200 0 0 0 I23
flabel comment s 1046 230 1046 230 0 FreeSans 200 0 0 0 I45
flabel comment s 312 230 312 230 0 FreeSans 200 0 0 0 I47
flabel comment s 624 752 624 752 0 FreeSans 200 0 0 0 I48
flabel comment s 618 1340 618 1340 0 FreeSans 200 0 0 0 I16
flabel comment s 1124 230 1124 230 0 FreeSans 300 180 0 0 D
flabel comment s 968 230 968 230 0 FreeSans 300 180 0 0 S
flabel comment s 812 230 812 230 0 FreeSans 300 180 0 0 D
flabel comment s 702 230 702 230 0 FreeSans 300 180 0 0 S
flabel comment s 546 230 546 230 0 FreeSans 300 180 0 0 D
flabel comment s 390 230 390 230 0 FreeSans 300 180 0 0 S
flabel comment s 234 230 234 230 0 FreeSans 300 180 0 0 D
flabel comment s 312 1272 312 1272 0 FreeSans 200 0 0 0 I44
flabel comment s 1438 702 1438 702 0 FreeSans 300 180 0 0 S
flabel comment s 1282 702 1282 702 0 FreeSans 300 180 0 0 D
flabel comment s 2064 674 2064 674 0 FreeSans 300 0 0 0 S
flabel comment s 2220 674 2220 674 0 FreeSans 300 0 0 0 D
flabel comment s 2376 674 2376 674 0 FreeSans 300 0 0 0 S
flabel comment s 2532 674 2532 674 0 FreeSans 300 0 0 0 D
flabel comment s 2688 674 2688 674 0 FreeSans 300 0 0 0 S
flabel comment s 1438 702 1438 702 0 FreeSans 300 0 0 0 S
flabel comment s 1594 702 1594 702 0 FreeSans 300 0 0 0 D
flabel comment s 702 752 702 752 0 FreeSans 300 180 0 0 S
flabel comment s 546 752 546 752 0 FreeSans 300 180 0 0 D
flabel comment s 390 752 390 752 0 FreeSans 300 180 0 0 S
flabel comment s 234 752 234 752 0 FreeSans 300 180 0 0 D
flabel comment s 2955 920 2955 920 0 FreeSans 300 180 0 0 S
flabel comment s 2799 920 2799 920 0 FreeSans 300 180 0 0 D
flabel comment s 234 1272 234 1272 0 FreeSans 300 0 0 0 S
flabel comment s 390 1272 390 1272 0 FreeSans 300 0 0 0 D
flabel comment s 2689 1272 2689 1272 0 FreeSans 300 180 0 0 S
flabel comment s 2533 1272 2533 1272 0 FreeSans 300 180 0 0 D
flabel comment s 2955 1306 2955 1306 0 FreeSans 300 180 0 0 S
flabel comment s 2799 1306 2799 1306 0 FreeSans 300 180 0 0 D
flabel comment s 972 1340 972 1340 0 FreeSans 300 0 0 0 S
flabel comment s 1208 1340 1208 1340 0 FreeSans 300 0 0 0 D
flabel comment s 1282 1173 1282 1173 0 FreeSans 400 0 0 0 t2
flabel comment s 1594 1173 1594 1173 0 FreeSans 400 0 0 0 t1
flabel comment s 2710 190 2710 190 0 FreeSans 400 0 0 0 t3
flabel comment s 1444 1340 1444 1340 0 FreeSans 300 0 0 0 S
flabel comment s 1680 1340 1680 1340 0 FreeSans 300 0 0 0 D
flabel comment s 1916 1340 1916 1340 0 FreeSans 300 0 0 0 S
flabel comment s 2152 1340 2152 1340 0 FreeSans 300 0 0 0 D
flabel comment s 2388 1340 2388 1340 0 FreeSans 300 0 0 0 S
flabel comment s 2877 920 2877 920 0 FreeSans 200 0 0 0 I36
flabel comment s 2877 1306 2877 1306 0 FreeSans 200 0 0 0 I35
rlabel viali s 4032 614 4066 648 1 LVPWR
port 3 nsew power bidirectional
rlabel viali s 3960 614 3994 648 1 LVPWR
port 3 nsew power bidirectional
rlabel metal1 s 14 604 4978 661 1 LVPWR
port 3 nsew power bidirectional
rlabel locali s 367 97 413 331 1 VGND
port 4 nsew ground bidirectional
rlabel locali s 367 51 485 97 1 VGND
port 4 nsew ground bidirectional
rlabel locali s 3924 125 3990 245 1 VGND
port 4 nsew ground bidirectional
rlabel locali s 3742 125 3808 245 1 VGND
port 4 nsew ground bidirectional
rlabel locali s 3556 125 3622 235 1 VGND
port 4 nsew ground bidirectional
rlabel locali s 3556 79 3990 125 1 VGND
port 4 nsew ground bidirectional
rlabel locali s 4225 1325 4275 1503 1 VGND
port 4 nsew ground bidirectional
rlabel locali s 4037 1325 4087 1503 1 VGND
port 4 nsew ground bidirectional
rlabel locali s 3924 1325 3990 1503 1 VGND
port 4 nsew ground bidirectional
rlabel locali s 3738 1383 3804 1503 1 VGND
port 4 nsew ground bidirectional
rlabel locali s 3556 1503 4275 1549 1 VGND
port 4 nsew ground bidirectional
rlabel locali s 3556 1383 3622 1503 1 VGND
port 4 nsew ground bidirectional
rlabel locali s 679 97 725 331 1 VGND
port 4 nsew ground bidirectional
rlabel locali s 607 51 725 97 1 VGND
port 4 nsew ground bidirectional
rlabel locali s 945 97 991 331 1 VGND
port 4 nsew ground bidirectional
rlabel locali s 909 51 1027 97 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 4236 1509 4270 1543 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 4140 1509 4174 1543 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 4044 1509 4078 1543 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 3948 1509 3982 1543 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 3948 85 3982 119 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 3852 1509 3886 1543 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 3852 85 3886 119 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 3756 1509 3790 1543 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 3756 85 3790 119 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 3660 1509 3694 1543 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 3660 85 3694 119 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 3564 1509 3598 1543 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 3564 85 3598 119 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 2911 1520 2945 1554 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 2815 1520 2849 1554 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 2718 1520 2752 1554 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 2623 1520 2657 1554 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 2527 1520 2561 1554 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 2431 1520 2465 1554 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 2335 1520 2369 1554 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 2239 1520 2273 1554 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 2143 1520 2177 1554 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 2047 1520 2081 1554 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 1951 1520 1985 1554 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 1855 1520 1889 1554 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 1759 1520 1793 1554 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 1663 1520 1697 1554 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 1567 1520 1601 1554 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 1471 1520 1505 1554 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 1375 1520 1409 1554 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 1279 1520 1313 1554 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 1183 1520 1217 1554 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 1087 1520 1121 1554 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 991 1520 1025 1554 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 987 57 1021 91 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 915 57 949 91 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 895 1520 929 1554 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 799 1520 833 1554 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 703 1520 737 1554 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 685 57 719 91 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 613 57 647 91 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 607 1520 641 1554 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 511 1520 545 1554 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 445 57 479 91 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 415 1520 449 1554 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 373 57 407 91 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 319 1520 353 1554 1 VGND
port 4 nsew ground bidirectional
rlabel viali s 223 1520 257 1554 1 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 51 4992 125 1 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 1503 4992 1577 1 VGND
port 4 nsew ground bidirectional
rlabel locali s 0 1611 4992 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 4927 1611 4961 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 4927 -17 4961 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 4831 1611 4865 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 4831 -17 4865 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 4735 1611 4769 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 4735 -17 4769 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 4639 1611 4673 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 4639 -17 4673 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 4543 1611 4577 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 4543 -17 4577 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 4447 1611 4481 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 4447 -17 4481 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 4351 1611 4385 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 4351 -17 4385 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 4255 1611 4289 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 4255 -17 4289 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 4159 1611 4193 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 4159 -17 4193 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 4063 1611 4097 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 4063 -17 4097 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 3967 1611 4001 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 3967 -17 4001 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 3871 1611 3905 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 3871 -17 3905 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 3775 1611 3809 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 3775 -17 3809 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 3679 1611 3713 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 3679 -17 3713 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 3583 1611 3617 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 3583 -17 3617 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 3487 1611 3521 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 3487 -17 3521 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 3391 1611 3425 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 3391 -17 3425 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 3295 1611 3329 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 3295 -17 3329 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 3199 1611 3233 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 3199 -17 3233 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 3103 1611 3137 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 3103 -17 3137 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 3007 1611 3041 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 3007 -17 3041 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 2911 1611 2945 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 2911 -17 2945 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 2815 1611 2849 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 2815 -17 2849 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 2719 1611 2753 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 2719 -17 2753 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 2623 1611 2657 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 2623 -17 2657 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 2527 1611 2561 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 2527 -17 2561 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 2431 1611 2465 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 2431 -17 2465 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 2335 1611 2369 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 2335 -17 2369 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 2239 1611 2273 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 2239 -17 2273 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 2143 1611 2177 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 2143 -17 2177 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 2047 1611 2081 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 2047 -17 2081 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 1951 1611 1985 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 1951 -17 1985 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 1855 1611 1889 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 1855 -17 1889 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 1759 1611 1793 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 1759 -17 1793 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 1663 1611 1697 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 1663 -17 1697 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 1567 1611 1601 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 1567 -17 1601 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 1471 1611 1505 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 1471 -17 1505 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 1375 1611 1409 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 1375 -17 1409 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 1279 1611 1313 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 1279 -17 1313 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 1183 1611 1217 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 1183 -17 1217 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 1087 1611 1121 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 1087 -17 1121 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 991 1611 1025 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 991 -17 1025 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 895 1611 929 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 895 -17 929 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 799 1611 833 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 799 -17 833 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 703 1611 737 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 703 -17 737 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 607 1611 641 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 607 -17 641 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 511 1611 545 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 511 -17 545 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 415 1611 449 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 415 -17 449 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 319 1611 353 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 319 -17 353 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 223 1611 257 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 223 -17 257 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 127 1611 161 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 127 -17 161 17 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 31 1611 65 1645 1 VNB
port 5 nsew ground bidirectional
rlabel viali s 31 -17 65 17 1 VNB
port 5 nsew ground bidirectional
rlabel metal1 s 0 -23 4992 23 1 VNB
port 5 nsew ground bidirectional
rlabel metal1 s 0 1605 4992 1651 1 VNB
port 5 nsew ground bidirectional
rlabel locali s 1827 797 1985 831 1 VPB
port 6 nsew power bidirectional
rlabel viali s 1925 797 1959 831 1 VPB
port 6 nsew power bidirectional
rlabel viali s 1853 797 1887 831 1 VPB
port 6 nsew power bidirectional
rlabel viali s 103 797 137 831 1 VPB
port 6 nsew power bidirectional
rlabel viali s 31 797 65 831 1 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 791 4992 837 1 VPB
port 6 nsew power bidirectional
rlabel locali s 2666 749 2710 1007 1 VPWR
port 7 nsew power bidirectional
rlabel locali s 2666 403 2710 703 1 VPWR
port 7 nsew power bidirectional
rlabel locali s 2629 703 2747 749 1 VPWR
port 7 nsew power bidirectional
rlabel locali s 2354 749 2398 1007 1 VPWR
port 7 nsew power bidirectional
rlabel locali s 2354 403 2398 703 1 VPWR
port 7 nsew power bidirectional
rlabel locali s 2317 703 2435 749 1 VPWR
port 7 nsew power bidirectional
rlabel locali s 2042 1007 2710 1051 1 VPWR
port 7 nsew power bidirectional
rlabel locali s 2042 749 2086 1007 1 VPWR
port 7 nsew power bidirectional
rlabel locali s 2042 403 2086 703 1 VPWR
port 7 nsew power bidirectional
rlabel locali s 2005 703 2123 749 1 VPWR
port 7 nsew power bidirectional
rlabel locali s 2931 925 2977 1011 1 VPWR
port 7 nsew power bidirectional
rlabel locali s 2931 853 2977 879 1 VPWR
port 7 nsew power bidirectional
rlabel locali s 2859 879 2977 925 1 VPWR
port 7 nsew power bidirectional
rlabel locali s 679 925 725 1023 1 VPWR
port 7 nsew power bidirectional
rlabel locali s 679 481 725 879 1 VPWR
port 7 nsew power bidirectional
rlabel locali s 643 879 761 925 1 VPWR
port 7 nsew power bidirectional
rlabel locali s 945 703 1062 751 1 VPWR
port 7 nsew power bidirectional
rlabel locali s 945 481 991 703 1 VPWR
port 7 nsew power bidirectional
rlabel viali s 2937 885 2971 919 1 VPWR
port 7 nsew power bidirectional
rlabel viali s 2865 885 2899 919 1 VPWR
port 7 nsew power bidirectional
rlabel viali s 2707 709 2741 743 1 VPWR
port 7 nsew power bidirectional
rlabel viali s 2635 709 2669 743 1 VPWR
port 7 nsew power bidirectional
rlabel viali s 2395 709 2429 743 1 VPWR
port 7 nsew power bidirectional
rlabel viali s 2323 709 2357 743 1 VPWR
port 7 nsew power bidirectional
rlabel viali s 2083 709 2117 743 1 VPWR
port 7 nsew power bidirectional
rlabel viali s 2011 709 2045 743 1 VPWR
port 7 nsew power bidirectional
rlabel viali s 1022 709 1056 743 1 VPWR
port 7 nsew power bidirectional
rlabel viali s 950 709 984 743 1 VPWR
port 7 nsew power bidirectional
rlabel viali s 721 885 755 919 1 VPWR
port 7 nsew power bidirectional
rlabel viali s 649 885 683 919 1 VPWR
port 7 nsew power bidirectional
rlabel viali s 409 885 443 919 1 VPWR
port 7 nsew power bidirectional
rlabel viali s 337 885 371 919 1 VPWR
port 7 nsew power bidirectional
rlabel metal1 s 0 689 4992 763 1 VPWR
port 7 nsew power bidirectional
rlabel metal1 s 0 865 4992 939 1 VPWR
port 7 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 4992 1628
string GDS_END 531566
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 478572
string LEFclass CORE
string LEFsite unithvdbl
string LEFsymmetry X Y
<< end >>
