magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< pwell >>
rect -26 -26 79 1426
<< ndiff >>
rect 0 1338 53 1400
rect 0 1304 11 1338
rect 45 1304 53 1338
rect 0 1270 53 1304
rect 0 1236 11 1270
rect 45 1236 53 1270
rect 0 1202 53 1236
rect 0 1168 11 1202
rect 45 1168 53 1202
rect 0 1134 53 1168
rect 0 1100 11 1134
rect 45 1100 53 1134
rect 0 1066 53 1100
rect 0 1032 11 1066
rect 45 1032 53 1066
rect 0 998 53 1032
rect 0 964 11 998
rect 45 964 53 998
rect 0 930 53 964
rect 0 896 11 930
rect 45 896 53 930
rect 0 862 53 896
rect 0 828 11 862
rect 45 828 53 862
rect 0 794 53 828
rect 0 760 11 794
rect 45 760 53 794
rect 0 726 53 760
rect 0 692 11 726
rect 45 692 53 726
rect 0 658 53 692
rect 0 624 11 658
rect 45 624 53 658
rect 0 590 53 624
rect 0 556 11 590
rect 45 556 53 590
rect 0 522 53 556
rect 0 488 11 522
rect 45 488 53 522
rect 0 454 53 488
rect 0 420 11 454
rect 45 420 53 454
rect 0 386 53 420
rect 0 352 11 386
rect 45 352 53 386
rect 0 318 53 352
rect 0 284 11 318
rect 45 284 53 318
rect 0 250 53 284
rect 0 216 11 250
rect 45 216 53 250
rect 0 182 53 216
rect 0 148 11 182
rect 45 148 53 182
rect 0 114 53 148
rect 0 80 11 114
rect 45 80 53 114
rect 0 46 53 80
rect 0 12 11 46
rect 45 12 53 46
rect 0 0 53 12
<< ndiffc >>
rect 11 1304 45 1338
rect 11 1236 45 1270
rect 11 1168 45 1202
rect 11 1100 45 1134
rect 11 1032 45 1066
rect 11 964 45 998
rect 11 896 45 930
rect 11 828 45 862
rect 11 760 45 794
rect 11 692 45 726
rect 11 624 45 658
rect 11 556 45 590
rect 11 488 45 522
rect 11 420 45 454
rect 11 352 45 386
rect 11 284 45 318
rect 11 216 45 250
rect 11 148 45 182
rect 11 80 45 114
rect 11 12 45 46
<< locali >>
rect 11 1338 45 1354
rect 11 1270 45 1304
rect 11 1202 45 1236
rect 11 1134 45 1168
rect 11 1066 45 1100
rect 11 998 45 1032
rect 11 930 45 964
rect 11 862 45 896
rect 11 794 45 828
rect 11 726 45 760
rect 11 658 45 692
rect 11 590 45 624
rect 11 522 45 556
rect 11 454 45 488
rect 11 386 45 420
rect 11 318 45 352
rect 11 250 45 284
rect 11 182 45 216
rect 11 114 45 148
rect 11 46 45 80
rect 11 -4 45 12
<< properties >>
string GDS_END 34504456
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 34502980
<< end >>
