magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< dnwell >>
rect -7428 -1830 -381 253
rect -2055 -4494 -1489 -1830
<< nwell >>
rect -6263 1543 554 2461
rect -7015 -1836 -1569 -1015
rect -7015 -2018 -1377 -1836
<< pwell >>
rect -6186 -495 -372 -393
<< psubdiff >>
rect -6160 -427 -398 -419
rect -6160 -461 -6136 -427
rect -6102 -461 -6068 -427
rect -6034 -461 -6000 -427
rect -5966 -461 -5932 -427
rect -5898 -461 -5864 -427
rect -5830 -461 -5796 -427
rect -5762 -461 -5728 -427
rect -5694 -461 -5660 -427
rect -5626 -461 -5592 -427
rect -5558 -461 -5524 -427
rect -5490 -461 -5456 -427
rect -5422 -461 -5388 -427
rect -5354 -461 -5320 -427
rect -5286 -461 -5252 -427
rect -5218 -461 -5184 -427
rect -5150 -461 -5116 -427
rect -5082 -461 -5048 -427
rect -5014 -461 -4980 -427
rect -4946 -461 -4912 -427
rect -4878 -461 -4844 -427
rect -4810 -461 -4776 -427
rect -4742 -461 -4708 -427
rect -4674 -461 -4640 -427
rect -4606 -461 -4572 -427
rect -4538 -461 -4504 -427
rect -4470 -461 -4436 -427
rect -4402 -461 -4368 -427
rect -4334 -461 -4300 -427
rect -4266 -461 -4232 -427
rect -4198 -461 -4164 -427
rect -4130 -461 -4096 -427
rect -4062 -461 -4028 -427
rect -3994 -461 -3960 -427
rect -3926 -461 -3892 -427
rect -3858 -461 -3824 -427
rect -3790 -461 -3756 -427
rect -3722 -461 -3688 -427
rect -3654 -461 -3620 -427
rect -3586 -461 -3552 -427
rect -3518 -461 -3484 -427
rect -3450 -461 -3416 -427
rect -3382 -461 -3348 -427
rect -3314 -461 -3280 -427
rect -3246 -461 -3212 -427
rect -3178 -461 -3144 -427
rect -3110 -461 -3076 -427
rect -3042 -461 -3008 -427
rect -2974 -461 -2940 -427
rect -2906 -461 -2872 -427
rect -2838 -461 -2804 -427
rect -2770 -461 -2736 -427
rect -2702 -461 -2668 -427
rect -2634 -461 -2600 -427
rect -2566 -461 -2532 -427
rect -2498 -461 -2464 -427
rect -2430 -461 -2396 -427
rect -2362 -461 -2328 -427
rect -2294 -461 -2260 -427
rect -2226 -461 -2192 -427
rect -2158 -461 -2124 -427
rect -2090 -461 -2056 -427
rect -2022 -461 -1988 -427
rect -1954 -461 -1920 -427
rect -1886 -461 -1852 -427
rect -1818 -461 -1784 -427
rect -1750 -461 -1716 -427
rect -1682 -461 -1648 -427
rect -1614 -461 -1580 -427
rect -1546 -461 -1512 -427
rect -1478 -461 -1444 -427
rect -1410 -461 -1376 -427
rect -1342 -461 -1308 -427
rect -1274 -461 -1240 -427
rect -1206 -461 -1172 -427
rect -1138 -461 -1104 -427
rect -1070 -461 -1036 -427
rect -1002 -461 -968 -427
rect -934 -461 -900 -427
rect -866 -461 -832 -427
rect -798 -461 -764 -427
rect -730 -461 -696 -427
rect -662 -461 -628 -427
rect -594 -461 -560 -427
rect -526 -461 -492 -427
rect -458 -461 -398 -427
rect -6160 -469 -398 -461
<< nsubdiff >>
rect -6949 -1910 -1443 -1902
rect -6949 -1944 -6925 -1910
rect -6891 -1944 -6857 -1910
rect -6823 -1944 -6789 -1910
rect -6755 -1944 -6721 -1910
rect -6687 -1944 -6653 -1910
rect -6619 -1944 -6585 -1910
rect -6551 -1944 -6517 -1910
rect -6483 -1944 -6449 -1910
rect -6415 -1944 -6381 -1910
rect -6347 -1944 -6313 -1910
rect -6279 -1944 -6245 -1910
rect -6211 -1944 -6177 -1910
rect -6143 -1944 -6109 -1910
rect -6075 -1944 -6041 -1910
rect -6007 -1944 -5973 -1910
rect -5939 -1944 -5905 -1910
rect -5871 -1944 -5837 -1910
rect -5803 -1944 -5769 -1910
rect -5735 -1944 -5701 -1910
rect -5667 -1944 -5633 -1910
rect -5599 -1944 -5565 -1910
rect -5531 -1944 -5497 -1910
rect -5463 -1944 -5429 -1910
rect -5395 -1944 -5361 -1910
rect -5327 -1944 -5293 -1910
rect -5259 -1944 -5225 -1910
rect -5191 -1944 -5157 -1910
rect -5123 -1944 -5089 -1910
rect -5055 -1944 -5021 -1910
rect -4987 -1944 -4953 -1910
rect -4919 -1944 -4885 -1910
rect -4851 -1944 -4817 -1910
rect -4783 -1944 -4749 -1910
rect -4715 -1944 -4681 -1910
rect -4647 -1944 -4613 -1910
rect -4579 -1944 -4545 -1910
rect -4511 -1944 -4477 -1910
rect -4443 -1944 -4409 -1910
rect -4375 -1944 -4341 -1910
rect -4307 -1944 -4273 -1910
rect -4239 -1944 -4205 -1910
rect -4171 -1944 -4137 -1910
rect -4103 -1944 -4069 -1910
rect -4035 -1944 -4001 -1910
rect -3967 -1944 -3933 -1910
rect -3899 -1944 -3865 -1910
rect -3831 -1944 -3797 -1910
rect -3763 -1944 -3729 -1910
rect -3695 -1944 -3661 -1910
rect -3627 -1944 -3593 -1910
rect -3559 -1944 -3525 -1910
rect -3491 -1944 -3457 -1910
rect -3423 -1944 -3389 -1910
rect -3355 -1944 -3321 -1910
rect -3287 -1944 -3253 -1910
rect -3219 -1944 -3185 -1910
rect -3151 -1944 -3117 -1910
rect -3083 -1944 -3049 -1910
rect -3015 -1944 -2981 -1910
rect -2947 -1944 -2913 -1910
rect -2879 -1944 -2845 -1910
rect -2811 -1944 -2777 -1910
rect -2743 -1944 -2709 -1910
rect -2675 -1944 -2641 -1910
rect -2607 -1944 -2573 -1910
rect -2539 -1944 -2505 -1910
rect -2471 -1944 -2437 -1910
rect -2403 -1944 -2369 -1910
rect -2335 -1944 -2301 -1910
rect -2267 -1944 -2233 -1910
rect -2199 -1944 -2165 -1910
rect -2131 -1944 -2097 -1910
rect -2063 -1944 -2029 -1910
rect -1995 -1944 -1961 -1910
rect -1927 -1944 -1893 -1910
rect -1859 -1944 -1825 -1910
rect -1791 -1944 -1757 -1910
rect -1723 -1944 -1689 -1910
rect -1655 -1944 -1621 -1910
rect -1587 -1944 -1553 -1910
rect -1519 -1944 -1443 -1910
rect -6949 -1952 -1443 -1944
<< mvnsubdiff >>
rect -6197 2387 488 2395
rect -6197 2353 -6173 2387
rect -6139 2353 -6105 2387
rect -6071 2353 -6037 2387
rect -6003 2353 -5969 2387
rect -5935 2353 -5901 2387
rect -5867 2353 -5833 2387
rect -5799 2353 -5765 2387
rect -5731 2353 -5697 2387
rect -5663 2353 -5629 2387
rect -5595 2353 -5561 2387
rect -5527 2353 -5493 2387
rect -5459 2353 -5425 2387
rect -5391 2353 -5357 2387
rect -5323 2353 -5289 2387
rect -5255 2353 -5221 2387
rect -5187 2353 -5153 2387
rect -5119 2353 -5085 2387
rect -5051 2353 -5017 2387
rect -4983 2353 -4949 2387
rect -4915 2353 -4881 2387
rect -4847 2353 -4813 2387
rect -4779 2353 -4745 2387
rect -4711 2353 -4677 2387
rect -4643 2353 -4609 2387
rect -4575 2353 -4541 2387
rect -4507 2353 -4473 2387
rect -4439 2353 -4405 2387
rect -4371 2353 -4337 2387
rect -4303 2353 -4269 2387
rect -4235 2353 -4201 2387
rect -4167 2353 -4133 2387
rect -4099 2353 -4065 2387
rect -4031 2353 -3997 2387
rect -3963 2353 -3929 2387
rect -3895 2353 -3861 2387
rect -3827 2353 -3793 2387
rect -3759 2353 -3725 2387
rect -3691 2353 -3657 2387
rect -3623 2353 -3589 2387
rect -3555 2353 -3521 2387
rect -3487 2353 -3453 2387
rect -3419 2353 -3385 2387
rect -3351 2353 -3317 2387
rect -3283 2353 -3249 2387
rect -3215 2353 -3181 2387
rect -3147 2353 -3113 2387
rect -3079 2353 -3045 2387
rect -3011 2353 -2977 2387
rect -2943 2353 -2909 2387
rect -2875 2353 -2841 2387
rect -2807 2353 -2773 2387
rect -2739 2353 -2705 2387
rect -2671 2353 -2637 2387
rect -2603 2353 -2569 2387
rect -2535 2353 -2501 2387
rect -2467 2353 -2433 2387
rect -2399 2353 -2365 2387
rect -2331 2353 -2297 2387
rect -2263 2353 -2229 2387
rect -2195 2353 -2161 2387
rect -2127 2353 -2093 2387
rect -2059 2353 -2025 2387
rect -1991 2353 -1957 2387
rect -1923 2353 -1889 2387
rect -1855 2353 -1821 2387
rect -1787 2353 -1753 2387
rect -1719 2353 -1685 2387
rect -1651 2353 -1617 2387
rect -1583 2353 -1549 2387
rect -1515 2353 -1481 2387
rect -1447 2353 -1413 2387
rect -1379 2353 -1345 2387
rect -1311 2353 -1277 2387
rect -1243 2353 -1209 2387
rect -1175 2353 -1141 2387
rect -1107 2353 -1073 2387
rect -1039 2353 -1005 2387
rect -971 2353 -937 2387
rect -903 2353 -869 2387
rect -835 2353 -801 2387
rect -767 2353 -733 2387
rect -699 2353 -665 2387
rect -631 2353 -597 2387
rect -563 2353 -529 2387
rect -495 2353 -461 2387
rect -427 2353 -393 2387
rect -359 2353 -325 2387
rect -291 2353 -257 2387
rect -223 2353 -189 2387
rect -155 2353 -121 2387
rect -87 2353 -53 2387
rect -19 2353 15 2387
rect 49 2353 83 2387
rect 117 2353 151 2387
rect 185 2353 219 2387
rect 253 2353 287 2387
rect 321 2353 355 2387
rect 389 2353 423 2387
rect 457 2353 488 2387
rect -6197 2345 488 2353
<< psubdiffcont >>
rect -6136 -461 -6102 -427
rect -6068 -461 -6034 -427
rect -6000 -461 -5966 -427
rect -5932 -461 -5898 -427
rect -5864 -461 -5830 -427
rect -5796 -461 -5762 -427
rect -5728 -461 -5694 -427
rect -5660 -461 -5626 -427
rect -5592 -461 -5558 -427
rect -5524 -461 -5490 -427
rect -5456 -461 -5422 -427
rect -5388 -461 -5354 -427
rect -5320 -461 -5286 -427
rect -5252 -461 -5218 -427
rect -5184 -461 -5150 -427
rect -5116 -461 -5082 -427
rect -5048 -461 -5014 -427
rect -4980 -461 -4946 -427
rect -4912 -461 -4878 -427
rect -4844 -461 -4810 -427
rect -4776 -461 -4742 -427
rect -4708 -461 -4674 -427
rect -4640 -461 -4606 -427
rect -4572 -461 -4538 -427
rect -4504 -461 -4470 -427
rect -4436 -461 -4402 -427
rect -4368 -461 -4334 -427
rect -4300 -461 -4266 -427
rect -4232 -461 -4198 -427
rect -4164 -461 -4130 -427
rect -4096 -461 -4062 -427
rect -4028 -461 -3994 -427
rect -3960 -461 -3926 -427
rect -3892 -461 -3858 -427
rect -3824 -461 -3790 -427
rect -3756 -461 -3722 -427
rect -3688 -461 -3654 -427
rect -3620 -461 -3586 -427
rect -3552 -461 -3518 -427
rect -3484 -461 -3450 -427
rect -3416 -461 -3382 -427
rect -3348 -461 -3314 -427
rect -3280 -461 -3246 -427
rect -3212 -461 -3178 -427
rect -3144 -461 -3110 -427
rect -3076 -461 -3042 -427
rect -3008 -461 -2974 -427
rect -2940 -461 -2906 -427
rect -2872 -461 -2838 -427
rect -2804 -461 -2770 -427
rect -2736 -461 -2702 -427
rect -2668 -461 -2634 -427
rect -2600 -461 -2566 -427
rect -2532 -461 -2498 -427
rect -2464 -461 -2430 -427
rect -2396 -461 -2362 -427
rect -2328 -461 -2294 -427
rect -2260 -461 -2226 -427
rect -2192 -461 -2158 -427
rect -2124 -461 -2090 -427
rect -2056 -461 -2022 -427
rect -1988 -461 -1954 -427
rect -1920 -461 -1886 -427
rect -1852 -461 -1818 -427
rect -1784 -461 -1750 -427
rect -1716 -461 -1682 -427
rect -1648 -461 -1614 -427
rect -1580 -461 -1546 -427
rect -1512 -461 -1478 -427
rect -1444 -461 -1410 -427
rect -1376 -461 -1342 -427
rect -1308 -461 -1274 -427
rect -1240 -461 -1206 -427
rect -1172 -461 -1138 -427
rect -1104 -461 -1070 -427
rect -1036 -461 -1002 -427
rect -968 -461 -934 -427
rect -900 -461 -866 -427
rect -832 -461 -798 -427
rect -764 -461 -730 -427
rect -696 -461 -662 -427
rect -628 -461 -594 -427
rect -560 -461 -526 -427
rect -492 -461 -458 -427
<< nsubdiffcont >>
rect -6925 -1944 -6891 -1910
rect -6857 -1944 -6823 -1910
rect -6789 -1944 -6755 -1910
rect -6721 -1944 -6687 -1910
rect -6653 -1944 -6619 -1910
rect -6585 -1944 -6551 -1910
rect -6517 -1944 -6483 -1910
rect -6449 -1944 -6415 -1910
rect -6381 -1944 -6347 -1910
rect -6313 -1944 -6279 -1910
rect -6245 -1944 -6211 -1910
rect -6177 -1944 -6143 -1910
rect -6109 -1944 -6075 -1910
rect -6041 -1944 -6007 -1910
rect -5973 -1944 -5939 -1910
rect -5905 -1944 -5871 -1910
rect -5837 -1944 -5803 -1910
rect -5769 -1944 -5735 -1910
rect -5701 -1944 -5667 -1910
rect -5633 -1944 -5599 -1910
rect -5565 -1944 -5531 -1910
rect -5497 -1944 -5463 -1910
rect -5429 -1944 -5395 -1910
rect -5361 -1944 -5327 -1910
rect -5293 -1944 -5259 -1910
rect -5225 -1944 -5191 -1910
rect -5157 -1944 -5123 -1910
rect -5089 -1944 -5055 -1910
rect -5021 -1944 -4987 -1910
rect -4953 -1944 -4919 -1910
rect -4885 -1944 -4851 -1910
rect -4817 -1944 -4783 -1910
rect -4749 -1944 -4715 -1910
rect -4681 -1944 -4647 -1910
rect -4613 -1944 -4579 -1910
rect -4545 -1944 -4511 -1910
rect -4477 -1944 -4443 -1910
rect -4409 -1944 -4375 -1910
rect -4341 -1944 -4307 -1910
rect -4273 -1944 -4239 -1910
rect -4205 -1944 -4171 -1910
rect -4137 -1944 -4103 -1910
rect -4069 -1944 -4035 -1910
rect -4001 -1944 -3967 -1910
rect -3933 -1944 -3899 -1910
rect -3865 -1944 -3831 -1910
rect -3797 -1944 -3763 -1910
rect -3729 -1944 -3695 -1910
rect -3661 -1944 -3627 -1910
rect -3593 -1944 -3559 -1910
rect -3525 -1944 -3491 -1910
rect -3457 -1944 -3423 -1910
rect -3389 -1944 -3355 -1910
rect -3321 -1944 -3287 -1910
rect -3253 -1944 -3219 -1910
rect -3185 -1944 -3151 -1910
rect -3117 -1944 -3083 -1910
rect -3049 -1944 -3015 -1910
rect -2981 -1944 -2947 -1910
rect -2913 -1944 -2879 -1910
rect -2845 -1944 -2811 -1910
rect -2777 -1944 -2743 -1910
rect -2709 -1944 -2675 -1910
rect -2641 -1944 -2607 -1910
rect -2573 -1944 -2539 -1910
rect -2505 -1944 -2471 -1910
rect -2437 -1944 -2403 -1910
rect -2369 -1944 -2335 -1910
rect -2301 -1944 -2267 -1910
rect -2233 -1944 -2199 -1910
rect -2165 -1944 -2131 -1910
rect -2097 -1944 -2063 -1910
rect -2029 -1944 -1995 -1910
rect -1961 -1944 -1927 -1910
rect -1893 -1944 -1859 -1910
rect -1825 -1944 -1791 -1910
rect -1757 -1944 -1723 -1910
rect -1689 -1944 -1655 -1910
rect -1621 -1944 -1587 -1910
rect -1553 -1944 -1519 -1910
<< mvnsubdiffcont >>
rect -6173 2353 -6139 2387
rect -6105 2353 -6071 2387
rect -6037 2353 -6003 2387
rect -5969 2353 -5935 2387
rect -5901 2353 -5867 2387
rect -5833 2353 -5799 2387
rect -5765 2353 -5731 2387
rect -5697 2353 -5663 2387
rect -5629 2353 -5595 2387
rect -5561 2353 -5527 2387
rect -5493 2353 -5459 2387
rect -5425 2353 -5391 2387
rect -5357 2353 -5323 2387
rect -5289 2353 -5255 2387
rect -5221 2353 -5187 2387
rect -5153 2353 -5119 2387
rect -5085 2353 -5051 2387
rect -5017 2353 -4983 2387
rect -4949 2353 -4915 2387
rect -4881 2353 -4847 2387
rect -4813 2353 -4779 2387
rect -4745 2353 -4711 2387
rect -4677 2353 -4643 2387
rect -4609 2353 -4575 2387
rect -4541 2353 -4507 2387
rect -4473 2353 -4439 2387
rect -4405 2353 -4371 2387
rect -4337 2353 -4303 2387
rect -4269 2353 -4235 2387
rect -4201 2353 -4167 2387
rect -4133 2353 -4099 2387
rect -4065 2353 -4031 2387
rect -3997 2353 -3963 2387
rect -3929 2353 -3895 2387
rect -3861 2353 -3827 2387
rect -3793 2353 -3759 2387
rect -3725 2353 -3691 2387
rect -3657 2353 -3623 2387
rect -3589 2353 -3555 2387
rect -3521 2353 -3487 2387
rect -3453 2353 -3419 2387
rect -3385 2353 -3351 2387
rect -3317 2353 -3283 2387
rect -3249 2353 -3215 2387
rect -3181 2353 -3147 2387
rect -3113 2353 -3079 2387
rect -3045 2353 -3011 2387
rect -2977 2353 -2943 2387
rect -2909 2353 -2875 2387
rect -2841 2353 -2807 2387
rect -2773 2353 -2739 2387
rect -2705 2353 -2671 2387
rect -2637 2353 -2603 2387
rect -2569 2353 -2535 2387
rect -2501 2353 -2467 2387
rect -2433 2353 -2399 2387
rect -2365 2353 -2331 2387
rect -2297 2353 -2263 2387
rect -2229 2353 -2195 2387
rect -2161 2353 -2127 2387
rect -2093 2353 -2059 2387
rect -2025 2353 -1991 2387
rect -1957 2353 -1923 2387
rect -1889 2353 -1855 2387
rect -1821 2353 -1787 2387
rect -1753 2353 -1719 2387
rect -1685 2353 -1651 2387
rect -1617 2353 -1583 2387
rect -1549 2353 -1515 2387
rect -1481 2353 -1447 2387
rect -1413 2353 -1379 2387
rect -1345 2353 -1311 2387
rect -1277 2353 -1243 2387
rect -1209 2353 -1175 2387
rect -1141 2353 -1107 2387
rect -1073 2353 -1039 2387
rect -1005 2353 -971 2387
rect -937 2353 -903 2387
rect -869 2353 -835 2387
rect -801 2353 -767 2387
rect -733 2353 -699 2387
rect -665 2353 -631 2387
rect -597 2353 -563 2387
rect -529 2353 -495 2387
rect -461 2353 -427 2387
rect -393 2353 -359 2387
rect -325 2353 -291 2387
rect -257 2353 -223 2387
rect -189 2353 -155 2387
rect -121 2353 -87 2387
rect -53 2353 -19 2387
rect 15 2353 49 2387
rect 83 2353 117 2387
rect 151 2353 185 2387
rect 219 2353 253 2387
rect 287 2353 321 2387
rect 355 2353 389 2387
rect 423 2353 457 2387
<< poly >>
rect -6135 2291 -6001 2307
rect -6135 2257 -6119 2291
rect -6085 2257 -6051 2291
rect -6017 2257 -6001 2291
rect -6135 2241 -6001 2257
rect -5835 2291 -5701 2307
rect -5835 2257 -5819 2291
rect -5785 2257 -5751 2291
rect -5717 2257 -5701 2291
rect -5835 2241 -5701 2257
rect -5535 2291 -5401 2307
rect -5535 2257 -5519 2291
rect -5485 2257 -5451 2291
rect -5417 2257 -5401 2291
rect -6128 2235 -6008 2241
rect -5828 2235 -5708 2241
rect -5535 2235 -5401 2257
rect -5359 2291 -5225 2307
rect -5359 2257 -5343 2291
rect -5309 2257 -5275 2291
rect -5241 2257 -5225 2291
rect -5359 2235 -5225 2257
rect -5059 2291 -4925 2307
rect -5059 2257 -5043 2291
rect -5009 2257 -4975 2291
rect -4941 2257 -4925 2291
rect -5059 2241 -4925 2257
rect -4759 2291 -4625 2307
rect -4759 2257 -4743 2291
rect -4709 2257 -4675 2291
rect -4641 2257 -4625 2291
rect -5052 2235 -4932 2241
rect -4759 2235 -4625 2257
rect -4583 2291 -4449 2307
rect -4583 2257 -4567 2291
rect -4533 2257 -4499 2291
rect -4465 2257 -4449 2291
rect -4583 2235 -4449 2257
rect -4283 2291 -4149 2307
rect -4283 2257 -4267 2291
rect -4233 2257 -4199 2291
rect -4165 2257 -4149 2291
rect -4283 2241 -4149 2257
rect -3683 2291 -3549 2307
rect -3683 2257 -3667 2291
rect -3633 2257 -3599 2291
rect -3565 2257 -3549 2291
rect -4276 2235 -4156 2241
rect -3683 2235 -3549 2257
rect -3507 2291 -3373 2307
rect -3507 2257 -3491 2291
rect -3457 2257 -3423 2291
rect -3389 2257 -3373 2291
rect -3507 2235 -3373 2257
rect -3207 2291 -3073 2307
rect -3207 2257 -3191 2291
rect -3157 2257 -3123 2291
rect -3089 2257 -3073 2291
rect -3207 2241 -3073 2257
rect -2907 2291 -2773 2307
rect -2907 2257 -2891 2291
rect -2857 2257 -2823 2291
rect -2789 2257 -2773 2291
rect -3200 2235 -3080 2241
rect -2907 2235 -2773 2257
rect -2731 2291 -2597 2307
rect -2731 2257 -2715 2291
rect -2681 2257 -2647 2291
rect -2613 2257 -2597 2291
rect -2731 2235 -2597 2257
rect -2431 2291 -2297 2307
rect -2431 2257 -2415 2291
rect -2381 2257 -2347 2291
rect -2313 2257 -2297 2291
rect -2431 2241 -2297 2257
rect -1830 2291 -1696 2307
rect -1830 2257 -1814 2291
rect -1780 2257 -1746 2291
rect -1712 2257 -1696 2291
rect -2424 2235 -2304 2241
rect -1830 2235 -1696 2257
rect -1654 2291 -1520 2307
rect -1654 2257 -1638 2291
rect -1604 2257 -1570 2291
rect -1536 2257 -1520 2291
rect -1654 2235 -1520 2257
rect -1354 2291 -1220 2307
rect -1354 2257 -1338 2291
rect -1304 2257 -1270 2291
rect -1236 2257 -1220 2291
rect -1354 2241 -1220 2257
rect -1054 2291 -920 2307
rect -1054 2257 -1038 2291
rect -1004 2257 -970 2291
rect -936 2257 -920 2291
rect -1347 2235 -1227 2241
rect -1054 2235 -920 2257
rect -878 2291 -744 2307
rect -878 2257 -862 2291
rect -828 2257 -794 2291
rect -760 2257 -744 2291
rect -878 2235 -744 2257
rect -578 2291 -444 2307
rect -578 2257 -562 2291
rect -528 2257 -494 2291
rect -460 2257 -444 2291
rect -578 2241 -444 2257
rect -571 2235 -451 2241
rect -213 1561 435 1577
rect -213 1527 -197 1561
rect -163 1527 -124 1561
rect -90 1527 -51 1561
rect -17 1527 22 1561
rect 56 1527 95 1561
rect 129 1527 168 1561
rect 202 1527 241 1561
rect 275 1527 313 1561
rect 347 1527 385 1561
rect 419 1527 435 1561
rect -213 1511 435 1527
rect -6128 -284 -6008 -278
rect -5828 -284 -5708 -278
rect -6135 -300 -6001 -284
rect -6135 -334 -6119 -300
rect -6085 -334 -6051 -300
rect -6017 -334 -6001 -300
rect -6135 -350 -6001 -334
rect -5835 -300 -5701 -284
rect -5835 -334 -5819 -300
rect -5785 -334 -5751 -300
rect -5717 -334 -5701 -300
rect -5835 -350 -5701 -334
rect -5535 -300 -5401 -278
rect -5535 -334 -5519 -300
rect -5485 -334 -5451 -300
rect -5417 -334 -5401 -300
rect -5535 -350 -5401 -334
rect -5359 -300 -5225 -278
rect -5052 -284 -4932 -278
rect -5359 -334 -5343 -300
rect -5309 -334 -5275 -300
rect -5241 -334 -5225 -300
rect -5359 -350 -5225 -334
rect -5059 -300 -4925 -284
rect -5059 -334 -5043 -300
rect -5009 -334 -4975 -300
rect -4941 -334 -4925 -300
rect -5059 -350 -4925 -334
rect -4759 -300 -4625 -278
rect -4759 -334 -4743 -300
rect -4709 -334 -4675 -300
rect -4641 -334 -4625 -300
rect -4759 -350 -4625 -334
rect -4583 -300 -4449 -278
rect -4276 -284 -4156 -278
rect -4583 -334 -4567 -300
rect -4533 -334 -4499 -300
rect -4465 -334 -4449 -300
rect -4583 -350 -4449 -334
rect -4283 -300 -4149 -284
rect -4283 -334 -4267 -300
rect -4233 -334 -4199 -300
rect -4165 -334 -4149 -300
rect -4283 -350 -4149 -334
rect -3683 -300 -3549 -278
rect -3683 -334 -3667 -300
rect -3633 -334 -3599 -300
rect -3565 -334 -3549 -300
rect -3683 -350 -3549 -334
rect -3507 -300 -3373 -278
rect -3200 -284 -3080 -278
rect -3507 -334 -3491 -300
rect -3457 -334 -3423 -300
rect -3389 -334 -3373 -300
rect -3507 -350 -3373 -334
rect -3207 -300 -3073 -284
rect -3207 -334 -3191 -300
rect -3157 -334 -3123 -300
rect -3089 -334 -3073 -300
rect -3207 -350 -3073 -334
rect -2907 -300 -2773 -278
rect -2907 -334 -2891 -300
rect -2857 -334 -2823 -300
rect -2789 -334 -2773 -300
rect -2907 -350 -2773 -334
rect -2731 -300 -2597 -278
rect -2424 -284 -2304 -278
rect -2731 -334 -2715 -300
rect -2681 -334 -2647 -300
rect -2613 -334 -2597 -300
rect -2731 -350 -2597 -334
rect -2431 -300 -2297 -284
rect -2431 -334 -2415 -300
rect -2381 -334 -2347 -300
rect -2313 -334 -2297 -300
rect -2431 -350 -2297 -334
rect -1830 -300 -1696 -278
rect -1830 -334 -1814 -300
rect -1780 -334 -1746 -300
rect -1712 -334 -1696 -300
rect -1830 -350 -1696 -334
rect -1654 -300 -1520 -278
rect -1347 -284 -1227 -278
rect -1654 -334 -1638 -300
rect -1604 -334 -1570 -300
rect -1536 -334 -1520 -300
rect -1654 -350 -1520 -334
rect -1354 -300 -1220 -284
rect -1354 -334 -1338 -300
rect -1304 -334 -1270 -300
rect -1236 -334 -1220 -300
rect -1354 -350 -1220 -334
rect -1054 -300 -920 -278
rect -1054 -334 -1038 -300
rect -1004 -334 -970 -300
rect -936 -334 -920 -300
rect -1054 -350 -920 -334
rect -878 -300 -744 -278
rect -571 -284 -451 -278
rect -878 -334 -862 -300
rect -828 -334 -794 -300
rect -760 -334 -744 -300
rect -878 -350 -744 -334
rect -578 -300 -444 -284
rect -578 -334 -562 -300
rect -528 -334 -494 -300
rect -460 -334 -444 -300
rect -578 -350 -444 -334
rect -231 -290 -97 -274
rect -231 -324 -215 -290
rect -181 -324 -147 -290
rect -113 -324 -97 -290
rect -231 -340 -97 -324
rect -6017 -537 -5883 -521
rect -6017 -571 -6001 -537
rect -5967 -571 -5933 -537
rect -5899 -571 -5883 -537
rect -6017 -587 -5883 -571
rect -5717 -537 -5583 -521
rect -5717 -571 -5701 -537
rect -5667 -571 -5633 -537
rect -5599 -571 -5583 -537
rect -5717 -587 -5583 -571
rect -5417 -537 -5283 -521
rect -5417 -571 -5401 -537
rect -5367 -571 -5333 -537
rect -5299 -571 -5283 -537
rect -6010 -593 -5890 -587
rect -5710 -593 -5590 -587
rect -5417 -593 -5283 -571
rect -5241 -537 -5107 -521
rect -5241 -571 -5225 -537
rect -5191 -571 -5157 -537
rect -5123 -571 -5107 -537
rect -5241 -593 -5107 -571
rect -4941 -537 -4807 -521
rect -4941 -571 -4925 -537
rect -4891 -571 -4857 -537
rect -4823 -571 -4807 -537
rect -4941 -593 -4807 -571
rect -4765 -537 -4631 -521
rect -4765 -571 -4749 -537
rect -4715 -571 -4681 -537
rect -4647 -571 -4631 -537
rect -4765 -593 -4631 -571
rect -4465 -537 -4331 -521
rect -4465 -571 -4449 -537
rect -4415 -571 -4381 -537
rect -4347 -571 -4331 -537
rect -4465 -587 -4331 -571
rect -4165 -537 -4031 -521
rect -4165 -571 -4149 -537
rect -4115 -571 -4081 -537
rect -4047 -571 -4031 -537
rect -4458 -593 -4338 -587
rect -4165 -593 -4031 -571
rect -3989 -537 -3855 -521
rect -3989 -571 -3973 -537
rect -3939 -571 -3905 -537
rect -3871 -571 -3855 -537
rect -3989 -593 -3855 -571
rect -3689 -537 -3555 -521
rect -3689 -571 -3673 -537
rect -3639 -571 -3605 -537
rect -3571 -571 -3555 -537
rect -3689 -593 -3555 -571
rect -3513 -537 -3379 -521
rect -3513 -571 -3497 -537
rect -3463 -571 -3429 -537
rect -3395 -571 -3379 -537
rect -3513 -593 -3379 -571
rect -3213 -537 -3079 -521
rect -3213 -571 -3197 -537
rect -3163 -571 -3129 -537
rect -3095 -571 -3079 -537
rect -3213 -587 -3079 -571
rect -2913 -537 -2779 -521
rect -2913 -571 -2897 -537
rect -2863 -571 -2829 -537
rect -2795 -571 -2779 -537
rect -3206 -593 -3086 -587
rect -2913 -593 -2779 -571
rect -2737 -537 -2603 -521
rect -2737 -571 -2721 -537
rect -2687 -571 -2653 -537
rect -2619 -571 -2603 -537
rect -2737 -593 -2603 -571
rect -2437 -537 -2303 -521
rect -2437 -571 -2421 -537
rect -2387 -571 -2353 -537
rect -2319 -571 -2303 -537
rect -2437 -593 -2303 -571
rect -2261 -537 -2127 -521
rect -2261 -571 -2245 -537
rect -2211 -571 -2177 -537
rect -2143 -571 -2127 -537
rect -2261 -593 -2127 -571
rect -1961 -537 -1827 -521
rect -1961 -571 -1945 -537
rect -1911 -571 -1877 -537
rect -1843 -571 -1827 -537
rect -1961 -587 -1827 -571
rect -1954 -593 -1834 -587
rect -6633 -867 -6499 -851
rect -6633 -901 -6617 -867
rect -6583 -901 -6549 -867
rect -6515 -901 -6499 -867
rect -6633 -917 -6499 -901
rect -6896 -1089 -6248 -1073
rect -6896 -1123 -6880 -1089
rect -6846 -1123 -6807 -1089
rect -6773 -1123 -6734 -1089
rect -6700 -1123 -6661 -1089
rect -6627 -1123 -6588 -1089
rect -6554 -1123 -6515 -1089
rect -6481 -1123 -6442 -1089
rect -6408 -1123 -6370 -1089
rect -6336 -1123 -6298 -1089
rect -6264 -1123 -6248 -1089
rect -6896 -1139 -6248 -1123
rect -5986 -1145 -5890 -845
rect -5686 -1145 -5590 -845
rect -5386 -1145 -5290 -819
rect -5234 -1145 -5138 -819
rect -4910 -1145 -4814 -819
rect -4758 -1145 -4662 -819
rect -4434 -1145 -4338 -845
rect -4134 -1145 -4038 -819
rect -3982 -1145 -3886 -819
rect -3658 -1145 -3562 -819
rect -3506 -1145 -3410 -819
rect -3182 -1145 -3086 -845
rect -2882 -1145 -2786 -819
rect -2730 -1145 -2634 -819
rect -2406 -1145 -2310 -819
rect -2254 -1145 -2158 -819
rect -1930 -1145 -1834 -845
rect -6010 -1803 -5890 -1797
rect -5710 -1803 -5590 -1797
rect -6017 -1819 -5883 -1803
rect -6017 -1853 -6001 -1819
rect -5967 -1853 -5933 -1819
rect -5899 -1853 -5883 -1819
rect -6017 -1869 -5883 -1853
rect -5717 -1819 -5583 -1803
rect -5717 -1853 -5701 -1819
rect -5667 -1853 -5633 -1819
rect -5599 -1853 -5583 -1819
rect -5717 -1869 -5583 -1853
rect -5417 -1819 -5283 -1797
rect -5417 -1853 -5401 -1819
rect -5367 -1853 -5333 -1819
rect -5299 -1853 -5283 -1819
rect -5417 -1869 -5283 -1853
rect -5241 -1819 -5107 -1797
rect -5241 -1853 -5225 -1819
rect -5191 -1853 -5157 -1819
rect -5123 -1853 -5107 -1819
rect -5241 -1869 -5107 -1853
rect -4941 -1819 -4807 -1797
rect -4941 -1853 -4925 -1819
rect -4891 -1853 -4857 -1819
rect -4823 -1853 -4807 -1819
rect -4941 -1869 -4807 -1853
rect -4765 -1819 -4631 -1797
rect -4458 -1803 -4338 -1797
rect -4765 -1853 -4749 -1819
rect -4715 -1853 -4681 -1819
rect -4647 -1853 -4631 -1819
rect -4765 -1869 -4631 -1853
rect -4465 -1819 -4331 -1803
rect -4465 -1853 -4449 -1819
rect -4415 -1853 -4381 -1819
rect -4347 -1853 -4331 -1819
rect -4465 -1869 -4331 -1853
rect -4165 -1819 -4031 -1797
rect -4165 -1853 -4149 -1819
rect -4115 -1853 -4081 -1819
rect -4047 -1853 -4031 -1819
rect -4165 -1869 -4031 -1853
rect -3989 -1819 -3855 -1797
rect -3989 -1853 -3973 -1819
rect -3939 -1853 -3905 -1819
rect -3871 -1853 -3855 -1819
rect -3989 -1869 -3855 -1853
rect -3689 -1819 -3555 -1797
rect -3689 -1853 -3673 -1819
rect -3639 -1853 -3605 -1819
rect -3571 -1853 -3555 -1819
rect -3689 -1869 -3555 -1853
rect -3513 -1819 -3379 -1797
rect -3206 -1803 -3086 -1797
rect -3513 -1853 -3497 -1819
rect -3463 -1853 -3429 -1819
rect -3395 -1853 -3379 -1819
rect -3513 -1869 -3379 -1853
rect -3213 -1819 -3079 -1803
rect -3213 -1853 -3197 -1819
rect -3163 -1853 -3129 -1819
rect -3095 -1853 -3079 -1819
rect -3213 -1869 -3079 -1853
rect -2913 -1819 -2779 -1797
rect -2913 -1853 -2897 -1819
rect -2863 -1853 -2829 -1819
rect -2795 -1853 -2779 -1819
rect -2913 -1869 -2779 -1853
rect -2737 -1819 -2603 -1797
rect -2737 -1853 -2721 -1819
rect -2687 -1853 -2653 -1819
rect -2619 -1853 -2603 -1819
rect -2737 -1869 -2603 -1853
rect -2437 -1819 -2303 -1797
rect -2437 -1853 -2421 -1819
rect -2387 -1853 -2353 -1819
rect -2319 -1853 -2303 -1819
rect -2437 -1869 -2303 -1853
rect -2261 -1819 -2127 -1797
rect -1954 -1803 -1834 -1797
rect -2261 -1853 -2245 -1819
rect -2211 -1853 -2177 -1819
rect -2143 -1853 -2127 -1819
rect -2261 -1869 -2127 -1853
rect -1961 -1819 -1827 -1803
rect -1961 -1853 -1945 -1819
rect -1911 -1853 -1877 -1819
rect -1843 -1853 -1827 -1819
rect -1961 -1869 -1827 -1853
<< polycont >>
rect -6119 2257 -6085 2291
rect -6051 2257 -6017 2291
rect -5819 2257 -5785 2291
rect -5751 2257 -5717 2291
rect -5519 2257 -5485 2291
rect -5451 2257 -5417 2291
rect -5343 2257 -5309 2291
rect -5275 2257 -5241 2291
rect -5043 2257 -5009 2291
rect -4975 2257 -4941 2291
rect -4743 2257 -4709 2291
rect -4675 2257 -4641 2291
rect -4567 2257 -4533 2291
rect -4499 2257 -4465 2291
rect -4267 2257 -4233 2291
rect -4199 2257 -4165 2291
rect -3667 2257 -3633 2291
rect -3599 2257 -3565 2291
rect -3491 2257 -3457 2291
rect -3423 2257 -3389 2291
rect -3191 2257 -3157 2291
rect -3123 2257 -3089 2291
rect -2891 2257 -2857 2291
rect -2823 2257 -2789 2291
rect -2715 2257 -2681 2291
rect -2647 2257 -2613 2291
rect -2415 2257 -2381 2291
rect -2347 2257 -2313 2291
rect -1814 2257 -1780 2291
rect -1746 2257 -1712 2291
rect -1638 2257 -1604 2291
rect -1570 2257 -1536 2291
rect -1338 2257 -1304 2291
rect -1270 2257 -1236 2291
rect -1038 2257 -1004 2291
rect -970 2257 -936 2291
rect -862 2257 -828 2291
rect -794 2257 -760 2291
rect -562 2257 -528 2291
rect -494 2257 -460 2291
rect -197 1527 -163 1561
rect -124 1527 -90 1561
rect -51 1527 -17 1561
rect 22 1527 56 1561
rect 95 1527 129 1561
rect 168 1527 202 1561
rect 241 1527 275 1561
rect 313 1527 347 1561
rect 385 1527 419 1561
rect -6119 -334 -6085 -300
rect -6051 -334 -6017 -300
rect -5819 -334 -5785 -300
rect -5751 -334 -5717 -300
rect -5519 -334 -5485 -300
rect -5451 -334 -5417 -300
rect -5343 -334 -5309 -300
rect -5275 -334 -5241 -300
rect -5043 -334 -5009 -300
rect -4975 -334 -4941 -300
rect -4743 -334 -4709 -300
rect -4675 -334 -4641 -300
rect -4567 -334 -4533 -300
rect -4499 -334 -4465 -300
rect -4267 -334 -4233 -300
rect -4199 -334 -4165 -300
rect -3667 -334 -3633 -300
rect -3599 -334 -3565 -300
rect -3491 -334 -3457 -300
rect -3423 -334 -3389 -300
rect -3191 -334 -3157 -300
rect -3123 -334 -3089 -300
rect -2891 -334 -2857 -300
rect -2823 -334 -2789 -300
rect -2715 -334 -2681 -300
rect -2647 -334 -2613 -300
rect -2415 -334 -2381 -300
rect -2347 -334 -2313 -300
rect -1814 -334 -1780 -300
rect -1746 -334 -1712 -300
rect -1638 -334 -1604 -300
rect -1570 -334 -1536 -300
rect -1338 -334 -1304 -300
rect -1270 -334 -1236 -300
rect -1038 -334 -1004 -300
rect -970 -334 -936 -300
rect -862 -334 -828 -300
rect -794 -334 -760 -300
rect -562 -334 -528 -300
rect -494 -334 -460 -300
rect -215 -324 -181 -290
rect -147 -324 -113 -290
rect -6001 -571 -5967 -537
rect -5933 -571 -5899 -537
rect -5701 -571 -5667 -537
rect -5633 -571 -5599 -537
rect -5401 -571 -5367 -537
rect -5333 -571 -5299 -537
rect -5225 -571 -5191 -537
rect -5157 -571 -5123 -537
rect -4925 -571 -4891 -537
rect -4857 -571 -4823 -537
rect -4749 -571 -4715 -537
rect -4681 -571 -4647 -537
rect -4449 -571 -4415 -537
rect -4381 -571 -4347 -537
rect -4149 -571 -4115 -537
rect -4081 -571 -4047 -537
rect -3973 -571 -3939 -537
rect -3905 -571 -3871 -537
rect -3673 -571 -3639 -537
rect -3605 -571 -3571 -537
rect -3497 -571 -3463 -537
rect -3429 -571 -3395 -537
rect -3197 -571 -3163 -537
rect -3129 -571 -3095 -537
rect -2897 -571 -2863 -537
rect -2829 -571 -2795 -537
rect -2721 -571 -2687 -537
rect -2653 -571 -2619 -537
rect -2421 -571 -2387 -537
rect -2353 -571 -2319 -537
rect -2245 -571 -2211 -537
rect -2177 -571 -2143 -537
rect -1945 -571 -1911 -537
rect -1877 -571 -1843 -537
rect -6617 -901 -6583 -867
rect -6549 -901 -6515 -867
rect -6880 -1123 -6846 -1089
rect -6807 -1123 -6773 -1089
rect -6734 -1123 -6700 -1089
rect -6661 -1123 -6627 -1089
rect -6588 -1123 -6554 -1089
rect -6515 -1123 -6481 -1089
rect -6442 -1123 -6408 -1089
rect -6370 -1123 -6336 -1089
rect -6298 -1123 -6264 -1089
rect -6001 -1853 -5967 -1819
rect -5933 -1853 -5899 -1819
rect -5701 -1853 -5667 -1819
rect -5633 -1853 -5599 -1819
rect -5401 -1853 -5367 -1819
rect -5333 -1853 -5299 -1819
rect -5225 -1853 -5191 -1819
rect -5157 -1853 -5123 -1819
rect -4925 -1853 -4891 -1819
rect -4857 -1853 -4823 -1819
rect -4749 -1853 -4715 -1819
rect -4681 -1853 -4647 -1819
rect -4449 -1853 -4415 -1819
rect -4381 -1853 -4347 -1819
rect -4149 -1853 -4115 -1819
rect -4081 -1853 -4047 -1819
rect -3973 -1853 -3939 -1819
rect -3905 -1853 -3871 -1819
rect -3673 -1853 -3639 -1819
rect -3605 -1853 -3571 -1819
rect -3497 -1853 -3463 -1819
rect -3429 -1853 -3395 -1819
rect -3197 -1853 -3163 -1819
rect -3129 -1853 -3095 -1819
rect -2897 -1853 -2863 -1819
rect -2829 -1853 -2795 -1819
rect -2721 -1853 -2687 -1819
rect -2653 -1853 -2619 -1819
rect -2421 -1853 -2387 -1819
rect -2353 -1853 -2319 -1819
rect -2245 -1853 -2211 -1819
rect -2177 -1853 -2143 -1819
rect -1945 -1853 -1911 -1819
rect -1877 -1853 -1843 -1819
<< locali >>
rect -6197 2387 488 2395
rect -6139 2353 -6124 2387
rect -6071 2353 -6051 2387
rect -6003 2353 -5978 2387
rect -5935 2353 -5905 2387
rect -5867 2353 -5833 2387
rect -5798 2353 -5765 2387
rect -5725 2353 -5697 2387
rect -5652 2353 -5629 2387
rect -5579 2353 -5561 2387
rect -5506 2353 -5493 2387
rect -5433 2353 -5425 2387
rect -5360 2353 -5357 2387
rect -5323 2353 -5321 2387
rect -5255 2353 -5248 2387
rect -5187 2353 -5175 2387
rect -5119 2353 -5102 2387
rect -5051 2353 -5030 2387
rect -4983 2353 -4958 2387
rect -4915 2353 -4886 2387
rect -4847 2353 -4814 2387
rect -4779 2353 -4745 2387
rect -4708 2353 -4677 2387
rect -4636 2353 -4609 2387
rect -4564 2353 -4541 2387
rect -4492 2353 -4473 2387
rect -4420 2353 -4405 2387
rect -4348 2353 -4337 2387
rect -4276 2353 -4269 2387
rect -4204 2353 -4201 2387
rect -4167 2353 -4166 2387
rect -4099 2353 -4094 2387
rect -4031 2353 -4022 2387
rect -3963 2353 -3950 2387
rect -3895 2353 -3878 2387
rect -3827 2353 -3806 2387
rect -3759 2353 -3734 2387
rect -3691 2353 -3662 2387
rect -3623 2353 -3590 2387
rect -3555 2353 -3521 2387
rect -3484 2353 -3453 2387
rect -3412 2353 -3385 2387
rect -3340 2353 -3317 2387
rect -3268 2353 -3249 2387
rect -3196 2353 -3181 2387
rect -3124 2353 -3113 2387
rect -3052 2353 -3045 2387
rect -2980 2353 -2977 2387
rect -2943 2353 -2942 2387
rect -2875 2353 -2870 2387
rect -2807 2353 -2798 2387
rect -2739 2353 -2726 2387
rect -2671 2353 -2654 2387
rect -2603 2353 -2582 2387
rect -2535 2353 -2510 2387
rect -2467 2353 -2438 2387
rect -2399 2353 -2366 2387
rect -2331 2353 -2297 2387
rect -2260 2353 -2229 2387
rect -2188 2353 -2161 2387
rect -2116 2353 -2093 2387
rect -2044 2353 -2025 2387
rect -1972 2353 -1957 2387
rect -1900 2353 -1889 2387
rect -1828 2353 -1821 2387
rect -1756 2353 -1753 2387
rect -1719 2353 -1718 2387
rect -1651 2353 -1646 2387
rect -1583 2353 -1574 2387
rect -1515 2353 -1502 2387
rect -1447 2353 -1430 2387
rect -1379 2353 -1358 2387
rect -1311 2353 -1286 2387
rect -1243 2353 -1214 2387
rect -1175 2353 -1142 2387
rect -1107 2353 -1073 2387
rect -1036 2353 -1005 2387
rect -964 2353 -937 2387
rect -892 2353 -869 2387
rect -820 2353 -801 2387
rect -748 2353 -733 2387
rect -676 2353 -665 2387
rect -604 2353 -597 2387
rect -532 2353 -529 2387
rect -495 2353 -494 2387
rect -427 2353 -422 2387
rect -359 2353 -350 2387
rect -291 2353 -278 2387
rect -223 2353 -206 2387
rect -155 2353 -134 2387
rect -87 2353 -62 2387
rect -19 2353 10 2387
rect 49 2353 82 2387
rect 117 2353 151 2387
rect 188 2353 219 2387
rect 260 2353 287 2387
rect 332 2353 355 2387
rect 404 2353 423 2387
rect 476 2353 488 2387
rect -6197 2345 488 2353
rect -6119 2291 -6017 2307
rect -6085 2257 -6051 2291
rect -6119 2241 -6017 2257
rect -5819 2291 -5717 2307
rect -5785 2257 -5751 2291
rect -5819 2241 -5717 2257
rect -5519 2291 -5417 2307
rect -5485 2257 -5451 2291
rect -5519 2241 -5417 2257
rect -5343 2291 -5241 2307
rect -5309 2257 -5275 2291
rect -5343 2241 -5241 2257
rect -5043 2291 -4941 2307
rect -5009 2257 -4975 2291
rect -5043 2241 -4941 2257
rect -4743 2291 -4641 2307
rect -4709 2257 -4675 2291
rect -4743 2241 -4641 2257
rect -4567 2291 -4465 2307
rect -4533 2257 -4499 2291
rect -4567 2241 -4465 2257
rect -4267 2291 -4165 2307
rect -4233 2257 -4199 2291
rect -4267 2241 -4165 2257
rect -3667 2291 -3565 2307
rect -3633 2257 -3599 2291
rect -3667 2241 -3565 2257
rect -3491 2291 -3389 2307
rect -3457 2257 -3423 2291
rect -3491 2241 -3389 2257
rect -3191 2291 -3089 2307
rect -3157 2257 -3123 2291
rect -3191 2241 -3089 2257
rect -2891 2291 -2789 2307
rect -2857 2257 -2823 2291
rect -2891 2241 -2789 2257
rect -2715 2291 -2613 2307
rect -2681 2257 -2647 2291
rect -2715 2241 -2613 2257
rect -2415 2291 -2313 2307
rect -2381 2257 -2347 2291
rect -2415 2241 -2313 2257
rect -1814 2291 -1712 2307
rect -1780 2257 -1746 2291
rect -1814 2241 -1712 2257
rect -1638 2291 -1536 2307
rect -1604 2257 -1570 2291
rect -1638 2241 -1536 2257
rect -1338 2291 -1236 2307
rect -1304 2257 -1270 2291
rect -1338 2241 -1236 2257
rect -1038 2291 -936 2307
rect -1004 2257 -970 2291
rect -1038 2241 -936 2257
rect -862 2291 -760 2307
rect -828 2257 -794 2291
rect -862 2241 -760 2257
rect -562 2291 -460 2307
rect -528 2257 -494 2291
rect -562 2241 -460 2257
rect -6173 1795 -6139 1807
rect -6173 1723 -6139 1761
rect -6173 1651 -6139 1689
rect -6173 1605 -6139 1617
rect -6105 48 -6031 2241
rect -6103 14 -6065 48
rect -6173 -112 -6139 -74
rect -6173 -184 -6139 -146
rect -6173 -230 -6139 -218
rect -6105 -284 -6031 14
rect -5997 117 -5963 2208
rect -5873 1795 -5839 1807
rect -5873 1723 -5839 1761
rect -5873 1651 -5839 1689
rect -5873 1605 -5839 1617
rect -5805 117 -5731 2241
rect -5997 15 -5731 117
rect -5997 -250 -5963 15
rect -5873 -112 -5839 -74
rect -5873 -184 -5839 -146
rect -5873 -230 -5839 -218
rect -5805 -284 -5731 15
rect -5697 117 -5663 2208
rect -5573 1795 -5539 1807
rect -5573 1723 -5539 1761
rect -5573 1651 -5539 1689
rect -5573 1609 -5539 1617
rect -5505 117 -5431 2241
rect -5697 15 -5431 117
rect -5697 -250 -5663 15
rect -5573 -40 -5539 -37
rect -5573 -112 -5539 -74
rect -5573 -184 -5539 -146
rect -5573 -250 -5539 -218
rect -5505 -284 -5431 15
rect -5397 48 -5363 2208
rect -5397 -225 -5363 14
rect -5329 -284 -5255 2241
rect -5221 1795 -5187 1807
rect -5221 1723 -5187 1761
rect -5221 1651 -5187 1689
rect -5221 1605 -5187 1617
rect -5097 1795 -5063 1807
rect -5097 1723 -5063 1761
rect -5097 1651 -5063 1689
rect -5097 1605 -5063 1617
rect -5029 117 -4955 2241
rect -5221 48 -4955 117
rect -5187 15 -4955 48
rect -5221 -54 -5187 14
rect -5097 -112 -5063 -74
rect -5221 -250 -5187 -147
rect -5097 -184 -5063 -146
rect -5097 -230 -5063 -218
rect -5029 -284 -4955 15
rect -4921 2139 -4887 2177
rect -4921 -250 -4887 2105
rect -4797 1795 -4763 1807
rect -4797 1723 -4763 1761
rect -4797 1651 -4763 1689
rect -4797 1609 -4763 1617
rect -4729 160 -4655 2241
rect -4727 126 -4689 160
rect -4797 -40 -4763 -37
rect -4797 -112 -4763 -74
rect -4797 -184 -4763 -146
rect -4797 -250 -4763 -218
rect -4729 -284 -4655 126
rect -4621 48 -4587 2208
rect -4621 -225 -4587 14
rect -4553 1966 -4479 2241
rect -4553 1932 -4536 1966
rect -4502 1932 -4479 1966
rect -4553 1894 -4479 1932
rect -4553 1860 -4536 1894
rect -4502 1860 -4479 1894
rect -4553 -284 -4479 1860
rect -4445 1795 -4411 1807
rect -4445 1723 -4411 1761
rect -4445 1651 -4411 1689
rect -4445 1605 -4411 1617
rect -4321 1795 -4287 1807
rect -4321 1723 -4287 1761
rect -4321 1651 -4287 1689
rect -4321 1605 -4287 1617
rect -4253 117 -4179 2241
rect -4445 48 -4179 117
rect -4411 15 -4179 48
rect -4445 -54 -4411 14
rect -4321 -112 -4287 -74
rect -4445 -250 -4411 -147
rect -4321 -184 -4287 -146
rect -4321 -230 -4287 -218
rect -4253 -284 -4179 15
rect -4145 117 -4111 2208
rect -3721 1795 -3687 1807
rect -3721 1723 -3687 1761
rect -3721 1651 -3687 1689
rect -3721 1609 -3687 1617
rect -3653 117 -3579 2241
rect -4145 15 -3579 117
rect -4145 -250 -4111 15
rect -3721 -40 -3687 -37
rect -3721 -112 -3687 -74
rect -3721 -184 -3687 -146
rect -3721 -250 -3687 -218
rect -3653 -284 -3579 15
rect -3545 48 -3511 2208
rect -3545 -225 -3511 14
rect -3477 -284 -3403 2241
rect -3369 1795 -3335 1807
rect -3369 1723 -3335 1761
rect -3369 1651 -3335 1689
rect -3369 1605 -3335 1617
rect -3245 1795 -3211 1807
rect -3245 1723 -3211 1761
rect -3245 1651 -3211 1689
rect -3245 1605 -3211 1617
rect -3177 117 -3103 2241
rect -3369 48 -3103 117
rect -3335 15 -3103 48
rect -3369 -54 -3335 14
rect -3245 -112 -3211 -74
rect -3369 -250 -3335 -147
rect -3245 -184 -3211 -146
rect -3245 -230 -3211 -218
rect -3177 -284 -3103 15
rect -3069 1965 -3035 2208
rect -3069 1893 -3035 1931
rect -3069 -250 -3035 1859
rect -2945 1795 -2911 1807
rect -2945 1723 -2911 1761
rect -2945 1651 -2911 1689
rect -2945 1609 -2911 1617
rect -2877 160 -2803 2241
rect -2875 126 -2837 160
rect -2945 -40 -2911 -37
rect -2945 -112 -2911 -74
rect -2945 -184 -2911 -146
rect -2945 -250 -2911 -218
rect -2877 -284 -2803 126
rect -2769 48 -2735 2208
rect -2769 -225 -2735 14
rect -2701 2094 -2627 2241
rect -2701 2060 -2680 2094
rect -2646 2060 -2627 2094
rect -2701 2022 -2627 2060
rect -2701 1988 -2680 2022
rect -2646 1988 -2627 2022
rect -2701 -284 -2627 1988
rect -2593 1795 -2559 1807
rect -2593 1723 -2559 1761
rect -2593 1651 -2559 1689
rect -2593 1605 -2559 1617
rect -2469 1795 -2435 1807
rect -2469 1723 -2435 1761
rect -2469 1651 -2435 1689
rect -2469 1605 -2435 1617
rect -2401 117 -2327 2241
rect -2593 48 -2327 117
rect -2559 15 -2327 48
rect -2593 -54 -2559 14
rect -2469 -112 -2435 -74
rect -2593 -250 -2559 -147
rect -2469 -184 -2435 -146
rect -2469 -230 -2435 -218
rect -2401 -284 -2327 15
rect -2293 117 -2259 2208
rect -1868 1795 -1834 1807
rect -1868 1723 -1834 1761
rect -1868 1651 -1834 1689
rect -1868 1609 -1834 1617
rect -1800 117 -1726 2241
rect -2293 15 -1726 117
rect -2293 -250 -2259 15
rect -1868 -40 -1834 -37
rect -1868 -112 -1834 -74
rect -1868 -184 -1834 -146
rect -1868 -250 -1834 -218
rect -1800 -284 -1726 15
rect -1692 1494 -1658 2208
rect -1692 -225 -1658 1460
rect -1624 -284 -1550 2241
rect -1516 1795 -1482 1807
rect -1516 1723 -1482 1761
rect -1516 1651 -1482 1689
rect -1516 1605 -1482 1617
rect -1392 1795 -1358 1807
rect -1392 1723 -1358 1761
rect -1392 1651 -1358 1689
rect -1392 1605 -1358 1617
rect -1324 1494 -1250 2241
rect -1324 1460 -1305 1494
rect -1271 1460 -1250 1494
rect -1324 117 -1250 1460
rect -1516 15 -1250 117
rect -1516 -54 -1482 15
rect -1392 -112 -1358 -74
rect -1516 -250 -1482 -147
rect -1392 -184 -1358 -146
rect -1392 -230 -1358 -218
rect -1324 -284 -1250 15
rect -1216 48 -1182 2208
rect -1092 1795 -1058 1807
rect -1092 1723 -1058 1761
rect -1092 1651 -1058 1689
rect -1092 1609 -1058 1617
rect -1182 14 -1144 48
rect -1216 -250 -1182 14
rect -1092 -40 -1058 -37
rect -1092 -112 -1058 -74
rect -1092 -184 -1058 -146
rect -1092 -250 -1058 -218
rect -1024 -284 -950 2241
rect -916 48 -882 2208
rect -916 -225 -882 14
rect -848 -284 -774 2241
rect -740 1795 -706 1807
rect -740 1723 -706 1761
rect -740 1651 -706 1689
rect -740 1605 -706 1617
rect -616 1795 -582 1807
rect -616 1723 -582 1761
rect -616 1651 -582 1689
rect -616 1605 -582 1617
rect -548 117 -474 2241
rect -740 48 -474 117
rect -706 15 -474 48
rect -740 -54 -706 14
rect -616 -112 -582 -74
rect -740 -250 -706 -147
rect -616 -184 -582 -146
rect -616 -230 -582 -218
rect -548 -284 -474 15
rect -440 432 -406 2208
rect -82 1896 -48 1934
rect 270 1896 304 1934
rect -258 1723 -224 1761
rect -258 1651 -224 1689
rect 94 1723 128 1761
rect 94 1651 128 1689
rect 446 1723 480 1761
rect 446 1651 480 1689
rect -213 1527 -197 1561
rect -163 1527 -124 1561
rect -90 1527 -51 1561
rect -17 1527 22 1561
rect 56 1527 95 1561
rect 129 1527 168 1561
rect 202 1527 241 1561
rect 275 1527 313 1561
rect 347 1527 385 1561
rect 419 1527 435 1561
rect -440 360 -406 398
rect -440 -250 -406 326
rect -268 -112 -234 -74
rect -268 -184 -234 -146
rect -93 -112 -59 -74
rect -93 -184 -59 -146
rect -6119 -300 -6017 -284
rect -6085 -334 -6051 -300
rect -6119 -350 -6017 -334
rect -5819 -300 -5717 -284
rect -5785 -334 -5751 -300
rect -5819 -350 -5717 -334
rect -5519 -300 -5417 -284
rect -5343 -300 -5241 -284
rect -5043 -300 -4941 -284
rect -5485 -334 -5451 -300
rect -5309 -334 -5275 -300
rect -5009 -334 -4975 -300
rect -5519 -350 -5417 -334
rect -5343 -350 -5241 -334
rect -5043 -350 -4941 -334
rect -4743 -300 -4641 -284
rect -4709 -334 -4675 -300
rect -4743 -350 -4641 -334
rect -4567 -300 -4465 -284
rect -4533 -334 -4499 -300
rect -4567 -350 -4465 -334
rect -4267 -300 -4165 -284
rect -4233 -334 -4199 -300
rect -4267 -350 -4165 -334
rect -3667 -300 -3565 -284
rect -3491 -300 -3389 -284
rect -3191 -300 -3089 -284
rect -3633 -334 -3599 -300
rect -3457 -334 -3423 -300
rect -3157 -334 -3123 -300
rect -3667 -350 -3565 -334
rect -3491 -350 -3389 -334
rect -3191 -350 -3089 -334
rect -2891 -300 -2789 -284
rect -2857 -334 -2823 -300
rect -2891 -350 -2789 -334
rect -2715 -300 -2613 -284
rect -2681 -334 -2647 -300
rect -2715 -350 -2613 -334
rect -2415 -300 -2313 -284
rect -2381 -334 -2347 -300
rect -2415 -350 -2313 -334
rect -1814 -300 -1712 -284
rect -1638 -300 -1536 -284
rect -1338 -300 -1236 -284
rect -1038 -300 -936 -284
rect -862 -300 -760 -284
rect -562 -300 -460 -284
rect -1780 -334 -1746 -300
rect -1604 -334 -1570 -300
rect -1304 -334 -1270 -300
rect -1004 -334 -982 -300
rect -828 -334 -794 -300
rect -528 -334 -494 -300
rect -231 -324 -216 -290
rect -181 -324 -147 -290
rect -110 -324 -97 -290
rect -1814 -350 -1712 -334
rect -1638 -350 -1536 -334
rect -1338 -350 -1236 -334
rect -1038 -350 -936 -334
rect -862 -350 -760 -334
rect -562 -350 -460 -334
rect -6160 -427 -398 -419
rect -6160 -461 -6136 -427
rect -6102 -461 -6068 -427
rect -6034 -461 -6000 -427
rect -5966 -461 -5932 -427
rect -5898 -461 -5864 -427
rect -5830 -461 -5796 -427
rect -5762 -461 -5728 -427
rect -5694 -461 -5660 -427
rect -5626 -461 -5592 -427
rect -5558 -461 -5524 -427
rect -5490 -461 -5456 -427
rect -5422 -461 -5388 -427
rect -5354 -461 -5320 -427
rect -5286 -461 -5252 -427
rect -5218 -461 -5184 -427
rect -5150 -461 -5116 -427
rect -5082 -461 -5048 -427
rect -5014 -461 -4980 -427
rect -4946 -461 -4912 -427
rect -4878 -461 -4844 -427
rect -4810 -461 -4776 -427
rect -4742 -461 -4708 -427
rect -4674 -461 -4640 -427
rect -4606 -461 -4572 -427
rect -4538 -461 -4504 -427
rect -4470 -461 -4436 -427
rect -4402 -461 -4368 -427
rect -4334 -461 -4300 -427
rect -4266 -461 -4232 -427
rect -4198 -461 -4164 -427
rect -4130 -461 -4096 -427
rect -4062 -461 -4028 -427
rect -3994 -461 -3960 -427
rect -3926 -461 -3892 -427
rect -3858 -461 -3824 -427
rect -3790 -461 -3756 -427
rect -3722 -461 -3688 -427
rect -3654 -461 -3620 -427
rect -3586 -461 -3552 -427
rect -3518 -461 -3484 -427
rect -3450 -461 -3416 -427
rect -3382 -461 -3348 -427
rect -3314 -461 -3280 -427
rect -3246 -461 -3212 -427
rect -3178 -461 -3144 -427
rect -3110 -461 -3076 -427
rect -3042 -461 -3008 -427
rect -2974 -461 -2940 -427
rect -2906 -461 -2872 -427
rect -2838 -461 -2804 -427
rect -2770 -461 -2736 -427
rect -2702 -461 -2668 -427
rect -2634 -461 -2600 -427
rect -2566 -461 -2532 -427
rect -2498 -461 -2464 -427
rect -2430 -461 -2396 -427
rect -2362 -461 -2328 -427
rect -2294 -461 -2260 -427
rect -2226 -461 -2192 -427
rect -2158 -461 -2124 -427
rect -2090 -461 -2056 -427
rect -2022 -461 -1988 -427
rect -1954 -461 -1920 -427
rect -1886 -461 -1852 -427
rect -1818 -461 -1784 -427
rect -1750 -461 -1716 -427
rect -1682 -461 -1648 -427
rect -1614 -461 -1580 -427
rect -1546 -461 -1512 -427
rect -1478 -461 -1444 -427
rect -1410 -461 -1376 -427
rect -1342 -461 -1308 -427
rect -1274 -461 -1240 -427
rect -1206 -461 -1172 -427
rect -1138 -461 -1104 -427
rect -1070 -461 -1036 -427
rect -1002 -461 -968 -427
rect -934 -461 -900 -427
rect -866 -461 -832 -427
rect -798 -461 -764 -427
rect -730 -461 -696 -427
rect -662 -461 -628 -427
rect -594 -461 -560 -427
rect -526 -461 -492 -427
rect -458 -461 -398 -427
rect -6160 -469 -398 -461
rect -6001 -537 -5899 -521
rect -6585 -571 -6547 -537
rect -5967 -571 -5933 -537
rect -6669 -725 -6635 -687
rect -6669 -797 -6635 -759
rect -6597 -867 -6529 -571
rect -6001 -587 -5899 -571
rect -5701 -537 -5599 -521
rect -5667 -571 -5633 -537
rect -5701 -587 -5599 -571
rect -5401 -537 -5299 -521
rect -5225 -537 -5123 -521
rect -4925 -537 -4823 -521
rect -5367 -571 -5333 -537
rect -5191 -571 -5157 -537
rect -4891 -571 -4857 -537
rect -5401 -587 -5299 -571
rect -5225 -587 -5123 -571
rect -4925 -587 -4823 -571
rect -4749 -537 -4647 -521
rect -4715 -571 -4681 -537
rect -4749 -587 -4647 -571
rect -4449 -537 -4347 -521
rect -4415 -571 -4381 -537
rect -4449 -587 -4347 -571
rect -4149 -537 -4047 -521
rect -3973 -537 -3871 -521
rect -3673 -537 -3571 -521
rect -4115 -571 -4081 -537
rect -3939 -571 -3905 -537
rect -3639 -571 -3605 -537
rect -4149 -587 -4047 -571
rect -3973 -587 -3871 -571
rect -3673 -587 -3571 -571
rect -3497 -537 -3395 -521
rect -3463 -571 -3429 -537
rect -3497 -587 -3395 -571
rect -3197 -537 -3095 -521
rect -3163 -571 -3129 -537
rect -3197 -587 -3095 -571
rect -2897 -537 -2795 -521
rect -2721 -537 -2619 -521
rect -2421 -537 -2319 -521
rect -2863 -571 -2829 -537
rect -2687 -571 -2653 -537
rect -2387 -571 -2356 -537
rect -2897 -587 -2795 -571
rect -2721 -587 -2619 -571
rect -2421 -587 -2319 -571
rect -2245 -537 -2143 -521
rect -2211 -571 -2177 -537
rect -2245 -587 -2143 -571
rect -1945 -537 -1843 -521
rect -1911 -571 -1877 -537
rect -1945 -587 -1843 -571
rect -6055 -653 -6021 -641
rect -6493 -725 -6459 -687
rect -6493 -797 -6459 -759
rect -6055 -725 -6021 -687
rect -6055 -797 -6021 -759
rect -6633 -901 -6617 -867
rect -6583 -901 -6549 -867
rect -6515 -901 -6499 -867
rect -5987 -885 -5913 -587
rect -6597 -1089 -6529 -901
rect -5985 -919 -5947 -885
rect -6896 -1123 -6880 -1089
rect -6846 -1123 -6807 -1089
rect -6773 -1123 -6734 -1089
rect -6700 -1123 -6661 -1089
rect -6627 -1123 -6588 -1089
rect -6554 -1123 -6515 -1089
rect -6481 -1123 -6442 -1089
rect -6408 -1123 -6370 -1089
rect -6336 -1123 -6298 -1089
rect -6264 -1123 -6248 -1089
rect -6055 -1179 -6021 -1167
rect -6941 -1251 -6907 -1213
rect -6941 -1323 -6907 -1285
rect -6589 -1251 -6555 -1213
rect -6589 -1323 -6555 -1285
rect -6237 -1251 -6203 -1213
rect -6237 -1323 -6203 -1285
rect -6055 -1251 -6021 -1213
rect -6055 -1323 -6021 -1285
rect -6055 -1369 -6021 -1357
rect -6765 -1776 -6731 -1738
rect -6413 -1776 -6379 -1738
rect -5987 -1819 -5913 -919
rect -5879 -886 -5845 -621
rect -5755 -653 -5721 -641
rect -5755 -725 -5721 -687
rect -5755 -797 -5721 -759
rect -5687 -886 -5613 -587
rect -5879 -988 -5613 -886
rect -5879 -1770 -5845 -988
rect -5755 -1179 -5721 -1167
rect -5755 -1251 -5721 -1213
rect -5755 -1323 -5721 -1285
rect -5755 -1369 -5721 -1357
rect -5687 -1819 -5613 -988
rect -5579 -886 -5545 -621
rect -5455 -653 -5421 -621
rect -5455 -725 -5421 -687
rect -5455 -797 -5421 -759
rect -5455 -834 -5421 -831
rect -5387 -886 -5313 -587
rect -5579 -988 -5313 -886
rect -5579 -1770 -5545 -988
rect -5455 -1179 -5421 -1171
rect -5455 -1251 -5421 -1213
rect -5455 -1323 -5421 -1285
rect -5455 -1369 -5421 -1357
rect -5387 -1819 -5313 -988
rect -5279 -885 -5245 -646
rect -5279 -1667 -5245 -919
rect -5279 -1739 -5245 -1701
rect -5211 -1819 -5137 -587
rect -5103 -724 -5069 -621
rect -4979 -653 -4945 -621
rect -4979 -725 -4945 -687
rect -4979 -797 -4945 -759
rect -5103 -885 -5069 -817
rect -4979 -834 -4945 -831
rect -4911 -997 -4837 -587
rect -4909 -1031 -4871 -997
rect -5103 -1179 -5069 -1167
rect -5103 -1251 -5069 -1213
rect -5103 -1323 -5069 -1285
rect -5103 -1369 -5069 -1357
rect -4979 -1179 -4945 -1171
rect -4979 -1251 -4945 -1213
rect -4979 -1323 -4945 -1285
rect -4979 -1369 -4945 -1357
rect -4911 -1819 -4837 -1031
rect -4803 -885 -4769 -646
rect -4803 -1770 -4769 -919
rect -4735 -1422 -4661 -587
rect -4627 -724 -4593 -621
rect -4503 -653 -4469 -641
rect -4503 -725 -4469 -687
rect -4503 -797 -4469 -759
rect -4627 -885 -4593 -817
rect -4435 -886 -4361 -587
rect -4593 -919 -4361 -886
rect -4627 -988 -4361 -919
rect -4627 -1179 -4593 -1167
rect -4627 -1251 -4593 -1213
rect -4627 -1323 -4593 -1285
rect -4627 -1369 -4593 -1357
rect -4503 -1179 -4469 -1167
rect -4503 -1251 -4469 -1213
rect -4503 -1323 -4469 -1285
rect -4503 -1369 -4469 -1357
rect -4735 -1456 -4718 -1422
rect -4684 -1456 -4661 -1422
rect -4735 -1494 -4661 -1456
rect -4735 -1528 -4718 -1494
rect -4684 -1528 -4661 -1494
rect -4735 -1819 -4661 -1528
rect -4435 -1819 -4361 -988
rect -4327 -886 -4293 -621
rect -4203 -653 -4169 -621
rect -4203 -725 -4169 -687
rect -4203 -797 -4169 -759
rect -4203 -834 -4169 -831
rect -4135 -886 -4061 -587
rect -4327 -988 -4061 -886
rect -4327 -1770 -4293 -988
rect -4203 -1179 -4169 -1171
rect -4203 -1251 -4169 -1213
rect -4203 -1323 -4169 -1285
rect -4203 -1369 -4169 -1357
rect -4135 -1819 -4061 -988
rect -4027 -885 -3993 -646
rect -4027 -1421 -3993 -919
rect -4027 -1493 -3993 -1455
rect -4027 -1770 -3993 -1527
rect -3959 -1819 -3885 -587
rect -3851 -724 -3817 -621
rect -3727 -653 -3693 -621
rect -3727 -725 -3693 -687
rect -3727 -797 -3693 -759
rect -3851 -885 -3817 -817
rect -3727 -834 -3693 -831
rect -3659 -997 -3585 -587
rect -3657 -1031 -3619 -997
rect -3851 -1179 -3817 -1167
rect -3851 -1251 -3817 -1213
rect -3851 -1323 -3817 -1285
rect -3851 -1369 -3817 -1357
rect -3727 -1179 -3693 -1171
rect -3727 -1251 -3693 -1213
rect -3727 -1323 -3693 -1285
rect -3727 -1369 -3693 -1357
rect -3659 -1819 -3585 -1031
rect -3551 -885 -3517 -646
rect -3551 -1770 -3517 -919
rect -3483 -1550 -3409 -587
rect -3375 -724 -3341 -621
rect -3251 -653 -3217 -641
rect -3251 -725 -3217 -687
rect -3251 -797 -3217 -759
rect -3375 -885 -3341 -817
rect -3183 -886 -3109 -587
rect -3341 -919 -3109 -886
rect -3375 -988 -3109 -919
rect -3375 -1179 -3341 -1167
rect -3375 -1251 -3341 -1213
rect -3375 -1323 -3341 -1285
rect -3375 -1369 -3341 -1357
rect -3251 -1179 -3217 -1167
rect -3251 -1251 -3217 -1213
rect -3251 -1323 -3217 -1285
rect -3251 -1369 -3217 -1357
rect -3483 -1584 -3462 -1550
rect -3428 -1584 -3409 -1550
rect -3483 -1622 -3409 -1584
rect -3483 -1656 -3462 -1622
rect -3428 -1656 -3409 -1622
rect -3483 -1819 -3409 -1656
rect -3183 -1819 -3109 -988
rect -3075 -886 -3041 -621
rect -2951 -653 -2917 -621
rect -2951 -725 -2917 -687
rect -2951 -797 -2917 -759
rect -2951 -834 -2917 -831
rect -2883 -886 -2809 -587
rect -3075 -988 -2809 -886
rect -3075 -1770 -3041 -988
rect -2951 -1179 -2917 -1171
rect -2951 -1251 -2917 -1213
rect -2951 -1323 -2917 -1285
rect -2951 -1369 -2917 -1357
rect -2883 -1819 -2809 -988
rect -2775 -885 -2741 -646
rect -2775 -1770 -2741 -919
rect -2707 -1819 -2633 -587
rect -2599 -724 -2565 -621
rect -2475 -653 -2441 -621
rect -2475 -725 -2441 -687
rect -2475 -797 -2441 -759
rect -2599 -885 -2565 -817
rect -2475 -834 -2441 -831
rect -2599 -1179 -2565 -1167
rect -2599 -1251 -2565 -1213
rect -2599 -1323 -2565 -1285
rect -2599 -1369 -2565 -1357
rect -2475 -1179 -2441 -1171
rect -2475 -1251 -2441 -1213
rect -2475 -1323 -2441 -1285
rect -2475 -1369 -2441 -1357
rect -2407 -1819 -2333 -587
rect -2299 -885 -2265 -646
rect -2299 -1770 -2265 -919
rect -2231 -1819 -2157 -587
rect -2123 -724 -2089 -621
rect -1999 -653 -1965 -641
rect -1999 -725 -1965 -687
rect -1999 -797 -1965 -759
rect -2123 -885 -2089 -817
rect -1931 -886 -1857 -587
rect -2089 -919 -1857 -886
rect -2123 -988 -1857 -919
rect -2123 -1179 -2089 -1167
rect -2123 -1251 -2089 -1213
rect -2123 -1323 -2089 -1285
rect -2123 -1369 -2089 -1357
rect -1999 -1179 -1965 -1167
rect -1999 -1251 -1965 -1213
rect -1999 -1323 -1965 -1285
rect -1999 -1369 -1965 -1357
rect -1931 -1819 -1857 -988
rect -1823 -1770 -1789 -621
rect -6017 -1853 -6001 -1819
rect -5967 -1853 -5933 -1819
rect -5899 -1853 -5883 -1819
rect -5717 -1853 -5701 -1819
rect -5667 -1853 -5633 -1819
rect -5599 -1853 -5583 -1819
rect -5417 -1853 -5401 -1819
rect -5367 -1853 -5333 -1819
rect -5299 -1853 -5283 -1819
rect -5241 -1853 -5225 -1819
rect -5191 -1853 -5157 -1819
rect -5123 -1853 -5107 -1819
rect -4941 -1853 -4925 -1819
rect -4891 -1853 -4857 -1819
rect -4823 -1853 -4807 -1819
rect -4765 -1853 -4749 -1819
rect -4715 -1853 -4681 -1819
rect -4647 -1853 -4631 -1819
rect -4465 -1853 -4449 -1819
rect -4415 -1853 -4381 -1819
rect -4347 -1853 -4331 -1819
rect -4165 -1853 -4149 -1819
rect -4115 -1853 -4081 -1819
rect -4047 -1853 -4031 -1819
rect -3989 -1853 -3973 -1819
rect -3939 -1853 -3905 -1819
rect -3871 -1853 -3855 -1819
rect -3689 -1853 -3673 -1819
rect -3639 -1853 -3605 -1819
rect -3571 -1853 -3555 -1819
rect -3513 -1853 -3497 -1819
rect -3463 -1853 -3429 -1819
rect -3395 -1853 -3379 -1819
rect -3213 -1853 -3197 -1819
rect -3163 -1853 -3129 -1819
rect -3095 -1853 -3079 -1819
rect -2913 -1853 -2897 -1819
rect -2863 -1853 -2829 -1819
rect -2795 -1853 -2779 -1819
rect -2737 -1853 -2721 -1819
rect -2687 -1853 -2653 -1819
rect -2619 -1853 -2603 -1819
rect -2437 -1853 -2421 -1819
rect -2387 -1853 -2353 -1819
rect -2319 -1853 -2303 -1819
rect -2261 -1853 -2245 -1819
rect -2211 -1853 -2177 -1819
rect -2143 -1853 -2127 -1819
rect -1961 -1853 -1945 -1819
rect -1911 -1853 -1877 -1819
rect -1843 -1853 -1827 -1819
rect -6949 -1910 -1443 -1902
rect -6949 -1944 -6925 -1910
rect -6891 -1944 -6857 -1910
rect -6823 -1944 -6789 -1910
rect -6755 -1944 -6721 -1910
rect -6687 -1944 -6653 -1910
rect -6619 -1944 -6585 -1910
rect -6551 -1944 -6517 -1910
rect -6483 -1944 -6449 -1910
rect -6415 -1944 -6381 -1910
rect -6347 -1944 -6313 -1910
rect -6279 -1944 -6245 -1910
rect -6211 -1944 -6177 -1910
rect -6143 -1944 -6109 -1910
rect -6075 -1944 -6041 -1910
rect -6007 -1944 -5973 -1910
rect -5939 -1944 -5905 -1910
rect -5871 -1944 -5837 -1910
rect -5803 -1944 -5769 -1910
rect -5735 -1944 -5701 -1910
rect -5667 -1944 -5633 -1910
rect -5599 -1944 -5565 -1910
rect -5531 -1944 -5497 -1910
rect -5463 -1944 -5429 -1910
rect -5395 -1944 -5361 -1910
rect -5327 -1944 -5293 -1910
rect -5259 -1944 -5225 -1910
rect -5191 -1944 -5157 -1910
rect -5123 -1944 -5089 -1910
rect -5055 -1944 -5021 -1910
rect -4987 -1944 -4953 -1910
rect -4919 -1944 -4885 -1910
rect -4851 -1944 -4817 -1910
rect -4783 -1944 -4749 -1910
rect -4715 -1944 -4681 -1910
rect -4647 -1944 -4613 -1910
rect -4579 -1944 -4545 -1910
rect -4511 -1944 -4477 -1910
rect -4443 -1944 -4409 -1910
rect -4375 -1944 -4341 -1910
rect -4307 -1944 -4273 -1910
rect -4239 -1944 -4205 -1910
rect -4171 -1944 -4137 -1910
rect -4103 -1944 -4069 -1910
rect -4035 -1944 -4001 -1910
rect -3967 -1944 -3933 -1910
rect -3899 -1944 -3865 -1910
rect -3831 -1944 -3797 -1910
rect -3763 -1944 -3729 -1910
rect -3695 -1944 -3661 -1910
rect -3627 -1944 -3593 -1910
rect -3559 -1944 -3525 -1910
rect -3491 -1944 -3457 -1910
rect -3423 -1944 -3389 -1910
rect -3355 -1944 -3321 -1910
rect -3287 -1944 -3253 -1910
rect -3219 -1944 -3185 -1910
rect -3151 -1944 -3117 -1910
rect -3083 -1944 -3049 -1910
rect -3015 -1944 -2981 -1910
rect -2947 -1944 -2913 -1910
rect -2879 -1944 -2845 -1910
rect -2811 -1944 -2777 -1910
rect -2743 -1944 -2709 -1910
rect -2675 -1944 -2641 -1910
rect -2607 -1944 -2573 -1910
rect -2539 -1944 -2505 -1910
rect -2471 -1944 -2437 -1910
rect -2403 -1944 -2369 -1910
rect -2335 -1944 -2301 -1910
rect -2267 -1944 -2233 -1910
rect -2199 -1944 -2165 -1910
rect -2131 -1944 -2097 -1910
rect -2063 -1944 -2029 -1910
rect -1995 -1944 -1961 -1910
rect -1927 -1944 -1893 -1910
rect -1859 -1944 -1825 -1910
rect -1791 -1944 -1757 -1910
rect -1723 -1944 -1689 -1910
rect -1655 -1944 -1621 -1910
rect -1587 -1944 -1553 -1910
rect -1519 -1944 -1443 -1910
rect -6949 -1952 -1443 -1944
<< viali >>
rect -6197 2353 -6173 2387
rect -6173 2353 -6163 2387
rect -6124 2353 -6105 2387
rect -6105 2353 -6090 2387
rect -6051 2353 -6037 2387
rect -6037 2353 -6017 2387
rect -5978 2353 -5969 2387
rect -5969 2353 -5944 2387
rect -5905 2353 -5901 2387
rect -5901 2353 -5871 2387
rect -5832 2353 -5799 2387
rect -5799 2353 -5798 2387
rect -5759 2353 -5731 2387
rect -5731 2353 -5725 2387
rect -5686 2353 -5663 2387
rect -5663 2353 -5652 2387
rect -5613 2353 -5595 2387
rect -5595 2353 -5579 2387
rect -5540 2353 -5527 2387
rect -5527 2353 -5506 2387
rect -5467 2353 -5459 2387
rect -5459 2353 -5433 2387
rect -5394 2353 -5391 2387
rect -5391 2353 -5360 2387
rect -5321 2353 -5289 2387
rect -5289 2353 -5287 2387
rect -5248 2353 -5221 2387
rect -5221 2353 -5214 2387
rect -5175 2353 -5153 2387
rect -5153 2353 -5141 2387
rect -5102 2353 -5085 2387
rect -5085 2353 -5068 2387
rect -5030 2353 -5017 2387
rect -5017 2353 -4996 2387
rect -4958 2353 -4949 2387
rect -4949 2353 -4924 2387
rect -4886 2353 -4881 2387
rect -4881 2353 -4852 2387
rect -4814 2353 -4813 2387
rect -4813 2353 -4780 2387
rect -4742 2353 -4711 2387
rect -4711 2353 -4708 2387
rect -4670 2353 -4643 2387
rect -4643 2353 -4636 2387
rect -4598 2353 -4575 2387
rect -4575 2353 -4564 2387
rect -4526 2353 -4507 2387
rect -4507 2353 -4492 2387
rect -4454 2353 -4439 2387
rect -4439 2353 -4420 2387
rect -4382 2353 -4371 2387
rect -4371 2353 -4348 2387
rect -4310 2353 -4303 2387
rect -4303 2353 -4276 2387
rect -4238 2353 -4235 2387
rect -4235 2353 -4204 2387
rect -4166 2353 -4133 2387
rect -4133 2353 -4132 2387
rect -4094 2353 -4065 2387
rect -4065 2353 -4060 2387
rect -4022 2353 -3997 2387
rect -3997 2353 -3988 2387
rect -3950 2353 -3929 2387
rect -3929 2353 -3916 2387
rect -3878 2353 -3861 2387
rect -3861 2353 -3844 2387
rect -3806 2353 -3793 2387
rect -3793 2353 -3772 2387
rect -3734 2353 -3725 2387
rect -3725 2353 -3700 2387
rect -3662 2353 -3657 2387
rect -3657 2353 -3628 2387
rect -3590 2353 -3589 2387
rect -3589 2353 -3556 2387
rect -3518 2353 -3487 2387
rect -3487 2353 -3484 2387
rect -3446 2353 -3419 2387
rect -3419 2353 -3412 2387
rect -3374 2353 -3351 2387
rect -3351 2353 -3340 2387
rect -3302 2353 -3283 2387
rect -3283 2353 -3268 2387
rect -3230 2353 -3215 2387
rect -3215 2353 -3196 2387
rect -3158 2353 -3147 2387
rect -3147 2353 -3124 2387
rect -3086 2353 -3079 2387
rect -3079 2353 -3052 2387
rect -3014 2353 -3011 2387
rect -3011 2353 -2980 2387
rect -2942 2353 -2909 2387
rect -2909 2353 -2908 2387
rect -2870 2353 -2841 2387
rect -2841 2353 -2836 2387
rect -2798 2353 -2773 2387
rect -2773 2353 -2764 2387
rect -2726 2353 -2705 2387
rect -2705 2353 -2692 2387
rect -2654 2353 -2637 2387
rect -2637 2353 -2620 2387
rect -2582 2353 -2569 2387
rect -2569 2353 -2548 2387
rect -2510 2353 -2501 2387
rect -2501 2353 -2476 2387
rect -2438 2353 -2433 2387
rect -2433 2353 -2404 2387
rect -2366 2353 -2365 2387
rect -2365 2353 -2332 2387
rect -2294 2353 -2263 2387
rect -2263 2353 -2260 2387
rect -2222 2353 -2195 2387
rect -2195 2353 -2188 2387
rect -2150 2353 -2127 2387
rect -2127 2353 -2116 2387
rect -2078 2353 -2059 2387
rect -2059 2353 -2044 2387
rect -2006 2353 -1991 2387
rect -1991 2353 -1972 2387
rect -1934 2353 -1923 2387
rect -1923 2353 -1900 2387
rect -1862 2353 -1855 2387
rect -1855 2353 -1828 2387
rect -1790 2353 -1787 2387
rect -1787 2353 -1756 2387
rect -1718 2353 -1685 2387
rect -1685 2353 -1684 2387
rect -1646 2353 -1617 2387
rect -1617 2353 -1612 2387
rect -1574 2353 -1549 2387
rect -1549 2353 -1540 2387
rect -1502 2353 -1481 2387
rect -1481 2353 -1468 2387
rect -1430 2353 -1413 2387
rect -1413 2353 -1396 2387
rect -1358 2353 -1345 2387
rect -1345 2353 -1324 2387
rect -1286 2353 -1277 2387
rect -1277 2353 -1252 2387
rect -1214 2353 -1209 2387
rect -1209 2353 -1180 2387
rect -1142 2353 -1141 2387
rect -1141 2353 -1108 2387
rect -1070 2353 -1039 2387
rect -1039 2353 -1036 2387
rect -998 2353 -971 2387
rect -971 2353 -964 2387
rect -926 2353 -903 2387
rect -903 2353 -892 2387
rect -854 2353 -835 2387
rect -835 2353 -820 2387
rect -782 2353 -767 2387
rect -767 2353 -748 2387
rect -710 2353 -699 2387
rect -699 2353 -676 2387
rect -638 2353 -631 2387
rect -631 2353 -604 2387
rect -566 2353 -563 2387
rect -563 2353 -532 2387
rect -494 2353 -461 2387
rect -461 2353 -460 2387
rect -422 2353 -393 2387
rect -393 2353 -388 2387
rect -350 2353 -325 2387
rect -325 2353 -316 2387
rect -278 2353 -257 2387
rect -257 2353 -244 2387
rect -206 2353 -189 2387
rect -189 2353 -172 2387
rect -134 2353 -121 2387
rect -121 2353 -100 2387
rect -62 2353 -53 2387
rect -53 2353 -28 2387
rect 10 2353 15 2387
rect 15 2353 44 2387
rect 82 2353 83 2387
rect 83 2353 116 2387
rect 154 2353 185 2387
rect 185 2353 188 2387
rect 226 2353 253 2387
rect 253 2353 260 2387
rect 298 2353 321 2387
rect 321 2353 332 2387
rect 370 2353 389 2387
rect 389 2353 404 2387
rect 442 2353 457 2387
rect 457 2353 476 2387
rect -6173 1761 -6139 1795
rect -6173 1689 -6139 1723
rect -6173 1617 -6139 1651
rect -6137 14 -6103 48
rect -6065 14 -6031 48
rect -6173 -74 -6139 -40
rect -6173 -146 -6139 -112
rect -6173 -218 -6139 -184
rect -5873 1761 -5839 1795
rect -5873 1689 -5839 1723
rect -5873 1617 -5839 1651
rect -5873 -74 -5839 -40
rect -5873 -146 -5839 -112
rect -5873 -218 -5839 -184
rect -5573 1761 -5539 1795
rect -5573 1689 -5539 1723
rect -5573 1617 -5539 1651
rect -5573 -74 -5539 -40
rect -5573 -146 -5539 -112
rect -5573 -218 -5539 -184
rect -5397 14 -5363 48
rect -5221 1761 -5187 1795
rect -5221 1689 -5187 1723
rect -5221 1617 -5187 1651
rect -5097 1761 -5063 1795
rect -5097 1689 -5063 1723
rect -5097 1617 -5063 1651
rect -5221 14 -5187 48
rect -5097 -74 -5063 -40
rect -5097 -146 -5063 -112
rect -5097 -218 -5063 -184
rect -4921 2177 -4887 2211
rect -4921 2105 -4887 2139
rect -4797 1761 -4763 1795
rect -4797 1689 -4763 1723
rect -4797 1617 -4763 1651
rect -4761 126 -4727 160
rect -4689 126 -4655 160
rect -4797 -74 -4763 -40
rect -4797 -146 -4763 -112
rect -4797 -218 -4763 -184
rect -4621 14 -4587 48
rect -4536 1932 -4502 1966
rect -4536 1860 -4502 1894
rect -4445 1761 -4411 1795
rect -4445 1689 -4411 1723
rect -4445 1617 -4411 1651
rect -4321 1761 -4287 1795
rect -4321 1689 -4287 1723
rect -4321 1617 -4287 1651
rect -4445 14 -4411 48
rect -4321 -74 -4287 -40
rect -4321 -146 -4287 -112
rect -4321 -218 -4287 -184
rect -3721 1761 -3687 1795
rect -3721 1689 -3687 1723
rect -3721 1617 -3687 1651
rect -3721 -74 -3687 -40
rect -3721 -146 -3687 -112
rect -3721 -218 -3687 -184
rect -3545 14 -3511 48
rect -3369 1761 -3335 1795
rect -3369 1689 -3335 1723
rect -3369 1617 -3335 1651
rect -3245 1761 -3211 1795
rect -3245 1689 -3211 1723
rect -3245 1617 -3211 1651
rect -3369 14 -3335 48
rect -3245 -74 -3211 -40
rect -3245 -146 -3211 -112
rect -3245 -218 -3211 -184
rect -3069 1931 -3035 1965
rect -3069 1859 -3035 1893
rect -2945 1761 -2911 1795
rect -2945 1689 -2911 1723
rect -2945 1617 -2911 1651
rect -2909 126 -2875 160
rect -2837 126 -2803 160
rect -2945 -74 -2911 -40
rect -2945 -146 -2911 -112
rect -2945 -218 -2911 -184
rect -2769 14 -2735 48
rect -2680 2060 -2646 2094
rect -2680 1988 -2646 2022
rect -2593 1761 -2559 1795
rect -2593 1689 -2559 1723
rect -2593 1617 -2559 1651
rect -2469 1761 -2435 1795
rect -2469 1689 -2435 1723
rect -2469 1617 -2435 1651
rect -2593 14 -2559 48
rect -2469 -74 -2435 -40
rect -2469 -146 -2435 -112
rect -2469 -218 -2435 -184
rect -1868 1761 -1834 1795
rect -1868 1689 -1834 1723
rect -1868 1617 -1834 1651
rect -1868 -74 -1834 -40
rect -1868 -146 -1834 -112
rect -1868 -218 -1834 -184
rect -1692 1460 -1658 1494
rect -1516 1761 -1482 1795
rect -1516 1689 -1482 1723
rect -1516 1617 -1482 1651
rect -1392 1761 -1358 1795
rect -1392 1689 -1358 1723
rect -1392 1617 -1358 1651
rect -1305 1460 -1271 1494
rect -1392 -74 -1358 -40
rect -1392 -146 -1358 -112
rect -1392 -218 -1358 -184
rect -1092 1761 -1058 1795
rect -1092 1689 -1058 1723
rect -1092 1617 -1058 1651
rect -1216 14 -1182 48
rect -1144 14 -1110 48
rect -1092 -74 -1058 -40
rect -1092 -146 -1058 -112
rect -1092 -218 -1058 -184
rect -916 14 -882 48
rect -740 1761 -706 1795
rect -740 1689 -706 1723
rect -740 1617 -706 1651
rect -616 1761 -582 1795
rect -616 1689 -582 1723
rect -616 1617 -582 1651
rect -740 14 -706 48
rect -616 -74 -582 -40
rect -616 -146 -582 -112
rect -616 -218 -582 -184
rect -82 1934 -48 1968
rect -82 1862 -48 1896
rect 270 1934 304 1968
rect 270 1862 304 1896
rect -258 1761 -224 1795
rect -258 1689 -224 1723
rect -258 1617 -224 1651
rect 94 1761 128 1795
rect 94 1689 128 1723
rect 94 1617 128 1651
rect 446 1761 480 1795
rect 446 1689 480 1723
rect 446 1617 480 1651
rect -440 398 -406 432
rect -440 326 -406 360
rect -268 -74 -234 -40
rect -268 -146 -234 -112
rect -268 -218 -234 -184
rect -93 -74 -59 -40
rect -93 -146 -59 -112
rect -93 -218 -59 -184
rect -5344 -334 -5343 -300
rect -5343 -334 -5310 -300
rect -5272 -334 -5241 -300
rect -5241 -334 -5238 -300
rect -3494 -334 -3491 -300
rect -3491 -334 -3460 -300
rect -3422 -334 -3389 -300
rect -3389 -334 -3388 -300
rect -1640 -334 -1638 -300
rect -1638 -334 -1606 -300
rect -1568 -334 -1536 -300
rect -1536 -334 -1534 -300
rect -1054 -334 -1038 -300
rect -1038 -334 -1020 -300
rect -982 -334 -970 -300
rect -970 -334 -948 -300
rect -864 -334 -862 -300
rect -862 -334 -830 -300
rect -792 -334 -760 -300
rect -760 -334 -758 -300
rect -216 -324 -215 -290
rect -215 -324 -182 -290
rect -144 -324 -113 -290
rect -113 -324 -110 -290
rect -6619 -571 -6585 -537
rect -6547 -571 -6513 -537
rect -6669 -687 -6635 -653
rect -6669 -759 -6635 -725
rect -6669 -831 -6635 -797
rect -5226 -571 -5225 -537
rect -5225 -571 -5192 -537
rect -5154 -571 -5123 -537
rect -5123 -571 -5120 -537
rect -3976 -571 -3973 -537
rect -3973 -571 -3942 -537
rect -3904 -571 -3871 -537
rect -3871 -571 -3870 -537
rect -2723 -571 -2721 -537
rect -2721 -571 -2689 -537
rect -2651 -571 -2619 -537
rect -2619 -571 -2617 -537
rect -2428 -571 -2421 -537
rect -2421 -571 -2394 -537
rect -2356 -571 -2353 -537
rect -2353 -571 -2322 -537
rect -6493 -687 -6459 -653
rect -6493 -759 -6459 -725
rect -6493 -831 -6459 -797
rect -6055 -687 -6021 -653
rect -6055 -759 -6021 -725
rect -6055 -831 -6021 -797
rect -6019 -919 -5985 -885
rect -5947 -919 -5913 -885
rect -6941 -1213 -6907 -1179
rect -6941 -1285 -6907 -1251
rect -6941 -1357 -6907 -1323
rect -6589 -1213 -6555 -1179
rect -6589 -1285 -6555 -1251
rect -6589 -1357 -6555 -1323
rect -6237 -1213 -6203 -1179
rect -6237 -1285 -6203 -1251
rect -6237 -1357 -6203 -1323
rect -6055 -1213 -6021 -1179
rect -6055 -1285 -6021 -1251
rect -6055 -1357 -6021 -1323
rect -6765 -1738 -6731 -1704
rect -6765 -1810 -6731 -1776
rect -6413 -1738 -6379 -1704
rect -6413 -1810 -6379 -1776
rect -5755 -687 -5721 -653
rect -5755 -759 -5721 -725
rect -5755 -831 -5721 -797
rect -5755 -1213 -5721 -1179
rect -5755 -1285 -5721 -1251
rect -5755 -1357 -5721 -1323
rect -5455 -687 -5421 -653
rect -5455 -759 -5421 -725
rect -5455 -831 -5421 -797
rect -5455 -1213 -5421 -1179
rect -5455 -1285 -5421 -1251
rect -5455 -1357 -5421 -1323
rect -5279 -919 -5245 -885
rect -5279 -1701 -5245 -1667
rect -5279 -1773 -5245 -1739
rect -4979 -687 -4945 -653
rect -4979 -759 -4945 -725
rect -4979 -831 -4945 -797
rect -5103 -919 -5069 -885
rect -4943 -1031 -4909 -997
rect -4871 -1031 -4837 -997
rect -5103 -1213 -5069 -1179
rect -5103 -1285 -5069 -1251
rect -5103 -1357 -5069 -1323
rect -4979 -1213 -4945 -1179
rect -4979 -1285 -4945 -1251
rect -4979 -1357 -4945 -1323
rect -4803 -919 -4769 -885
rect -4503 -687 -4469 -653
rect -4503 -759 -4469 -725
rect -4503 -831 -4469 -797
rect -4627 -919 -4593 -885
rect -4627 -1213 -4593 -1179
rect -4627 -1285 -4593 -1251
rect -4627 -1357 -4593 -1323
rect -4503 -1213 -4469 -1179
rect -4503 -1285 -4469 -1251
rect -4503 -1357 -4469 -1323
rect -4718 -1456 -4684 -1422
rect -4718 -1528 -4684 -1494
rect -4203 -687 -4169 -653
rect -4203 -759 -4169 -725
rect -4203 -831 -4169 -797
rect -4203 -1213 -4169 -1179
rect -4203 -1285 -4169 -1251
rect -4203 -1357 -4169 -1323
rect -4027 -919 -3993 -885
rect -4027 -1455 -3993 -1421
rect -4027 -1527 -3993 -1493
rect -3727 -687 -3693 -653
rect -3727 -759 -3693 -725
rect -3727 -831 -3693 -797
rect -3851 -919 -3817 -885
rect -3691 -1031 -3657 -997
rect -3619 -1031 -3585 -997
rect -3851 -1213 -3817 -1179
rect -3851 -1285 -3817 -1251
rect -3851 -1357 -3817 -1323
rect -3727 -1213 -3693 -1179
rect -3727 -1285 -3693 -1251
rect -3727 -1357 -3693 -1323
rect -3551 -919 -3517 -885
rect -3251 -687 -3217 -653
rect -3251 -759 -3217 -725
rect -3251 -831 -3217 -797
rect -3375 -919 -3341 -885
rect -3375 -1213 -3341 -1179
rect -3375 -1285 -3341 -1251
rect -3375 -1357 -3341 -1323
rect -3251 -1213 -3217 -1179
rect -3251 -1285 -3217 -1251
rect -3251 -1357 -3217 -1323
rect -3462 -1584 -3428 -1550
rect -3462 -1656 -3428 -1622
rect -2951 -687 -2917 -653
rect -2951 -759 -2917 -725
rect -2951 -831 -2917 -797
rect -2951 -1213 -2917 -1179
rect -2951 -1285 -2917 -1251
rect -2951 -1357 -2917 -1323
rect -2775 -919 -2741 -885
rect -2475 -687 -2441 -653
rect -2475 -759 -2441 -725
rect -2475 -831 -2441 -797
rect -2599 -919 -2565 -885
rect -2599 -1213 -2565 -1179
rect -2599 -1285 -2565 -1251
rect -2599 -1357 -2565 -1323
rect -2475 -1213 -2441 -1179
rect -2475 -1285 -2441 -1251
rect -2475 -1357 -2441 -1323
rect -2299 -919 -2265 -885
rect -1999 -687 -1965 -653
rect -1999 -759 -1965 -725
rect -1999 -831 -1965 -797
rect -2123 -919 -2089 -885
rect -2123 -1213 -2089 -1179
rect -2123 -1285 -2089 -1251
rect -2123 -1357 -2089 -1323
rect -1999 -1213 -1965 -1179
rect -1999 -1285 -1965 -1251
rect -1999 -1357 -1965 -1323
<< metal1 >>
rect -6209 2387 488 2393
rect -6209 2353 -6197 2387
rect -6163 2353 -6124 2387
rect -6090 2353 -6051 2387
rect -6017 2353 -5978 2387
rect -5944 2353 -5905 2387
rect -5871 2353 -5832 2387
rect -5798 2353 -5759 2387
rect -5725 2353 -5686 2387
rect -5652 2353 -5613 2387
rect -5579 2353 -5540 2387
rect -5506 2353 -5467 2387
rect -5433 2353 -5394 2387
rect -5360 2353 -5321 2387
rect -5287 2353 -5248 2387
rect -5214 2353 -5175 2387
rect -5141 2353 -5102 2387
rect -5068 2353 -5030 2387
rect -4996 2353 -4958 2387
rect -4924 2353 -4886 2387
rect -4852 2353 -4814 2387
rect -4780 2353 -4742 2387
rect -4708 2353 -4670 2387
rect -4636 2353 -4598 2387
rect -4564 2353 -4526 2387
rect -4492 2353 -4454 2387
rect -4420 2353 -4382 2387
rect -4348 2353 -4310 2387
rect -4276 2353 -4238 2387
rect -4204 2353 -4166 2387
rect -4132 2353 -4094 2387
rect -4060 2353 -4022 2387
rect -3988 2353 -3950 2387
rect -3916 2353 -3878 2387
rect -3844 2353 -3806 2387
rect -3772 2353 -3734 2387
rect -3700 2353 -3662 2387
rect -3628 2353 -3590 2387
rect -3556 2353 -3518 2387
rect -3484 2353 -3446 2387
rect -3412 2353 -3374 2387
rect -3340 2353 -3302 2387
rect -3268 2353 -3230 2387
rect -3196 2353 -3158 2387
rect -3124 2353 -3086 2387
rect -3052 2353 -3014 2387
rect -2980 2353 -2942 2387
rect -2908 2353 -2870 2387
rect -2836 2353 -2798 2387
rect -2764 2353 -2726 2387
rect -2692 2353 -2654 2387
rect -2620 2353 -2582 2387
rect -2548 2353 -2510 2387
rect -2476 2353 -2438 2387
rect -2404 2353 -2366 2387
rect -2332 2353 -2294 2387
rect -2260 2353 -2222 2387
rect -2188 2353 -2150 2387
rect -2116 2353 -2078 2387
rect -2044 2353 -2006 2387
rect -1972 2353 -1934 2387
rect -1900 2353 -1862 2387
rect -1828 2353 -1790 2387
rect -1756 2353 -1718 2387
rect -1684 2353 -1646 2387
rect -1612 2353 -1574 2387
rect -1540 2353 -1502 2387
rect -1468 2353 -1430 2387
rect -1396 2353 -1358 2387
rect -1324 2353 -1286 2387
rect -1252 2353 -1214 2387
rect -1180 2353 -1142 2387
rect -1108 2353 -1070 2387
rect -1036 2353 -998 2387
rect -964 2353 -926 2387
rect -892 2353 -854 2387
rect -820 2353 -782 2387
rect -748 2353 -710 2387
rect -676 2353 -638 2387
rect -604 2353 -566 2387
rect -532 2353 -494 2387
rect -460 2353 -422 2387
rect -388 2353 -350 2387
rect -316 2353 -278 2387
rect -244 2353 -206 2387
rect -172 2353 -134 2387
rect -100 2353 -62 2387
rect -28 2353 10 2387
rect 44 2353 82 2387
rect 116 2353 154 2387
rect 188 2353 226 2387
rect 260 2353 298 2387
rect 332 2353 370 2387
rect 404 2353 442 2387
rect 476 2353 488 2387
rect -6209 2347 488 2353
rect -4927 2211 -4881 2223
rect -4927 2177 -4921 2211
rect -4887 2181 -4881 2211
rect -4887 2177 -1427 2181
rect -4927 2139 -1427 2177
rect -4927 2105 -4921 2139
rect -4887 2135 -1427 2139
rect -4887 2105 -4881 2135
rect -4927 2093 -4881 2105
rect -2686 2094 -2640 2106
rect -2686 2064 -2680 2094
rect -6188 2060 -2680 2064
rect -2646 2060 -2640 2094
rect -6188 2022 -2640 2060
rect -6188 2018 -2680 2022
rect -2686 1988 -2680 2018
rect -2646 1988 -2640 2022
rect -4542 1966 -4496 1978
rect -4542 1936 -4536 1966
rect -6188 1932 -4536 1936
rect -4502 1932 -4496 1966
rect -6188 1894 -4496 1932
rect -6188 1890 -4536 1894
rect -4542 1860 -4536 1890
rect -4502 1860 -4496 1894
rect -4542 1848 -4496 1860
rect -3075 1965 -3029 1977
rect -2686 1976 -2640 1988
rect -3075 1931 -3069 1965
rect -3035 1935 -3029 1965
rect -88 1973 372 1980
rect -88 1968 320 1973
rect -3035 1931 -1427 1935
rect -3075 1893 -1427 1931
rect -3075 1859 -3069 1893
rect -3035 1889 -1427 1893
rect -88 1934 -82 1968
rect -48 1934 270 1968
rect 304 1934 320 1968
rect -88 1921 320 1934
rect -88 1909 372 1921
rect -88 1896 320 1909
rect -3035 1859 -3029 1889
rect -3075 1847 -3029 1859
rect -88 1862 -82 1896
rect -48 1862 270 1896
rect 304 1862 320 1896
rect -88 1857 320 1862
rect -88 1850 372 1857
rect -6185 1795 486 1807
rect -6185 1761 -6173 1795
rect -6139 1761 -5873 1795
rect -5839 1761 -5573 1795
rect -5539 1761 -5221 1795
rect -5187 1761 -5097 1795
rect -5063 1761 -4797 1795
rect -4763 1761 -4445 1795
rect -4411 1761 -4321 1795
rect -4287 1761 -3721 1795
rect -3687 1761 -3369 1795
rect -3335 1761 -3245 1795
rect -3211 1761 -2945 1795
rect -2911 1761 -2593 1795
rect -2559 1761 -2469 1795
rect -2435 1761 -1868 1795
rect -1834 1761 -1516 1795
rect -1482 1761 -1392 1795
rect -1358 1761 -1092 1795
rect -1058 1761 -740 1795
rect -706 1761 -616 1795
rect -582 1761 -258 1795
rect -224 1761 94 1795
rect 128 1761 446 1795
rect 480 1761 486 1795
rect -6185 1723 486 1761
rect -6185 1689 -6173 1723
rect -6139 1689 -5873 1723
rect -5839 1689 -5573 1723
rect -5539 1689 -5221 1723
rect -5187 1689 -5097 1723
rect -5063 1689 -4797 1723
rect -4763 1689 -4445 1723
rect -4411 1689 -4321 1723
rect -4287 1689 -3721 1723
rect -3687 1689 -3369 1723
rect -3335 1689 -3245 1723
rect -3211 1689 -2945 1723
rect -2911 1689 -2593 1723
rect -2559 1689 -2469 1723
rect -2435 1689 -1868 1723
rect -1834 1689 -1516 1723
rect -1482 1689 -1392 1723
rect -1358 1689 -1092 1723
rect -1058 1689 -740 1723
rect -706 1689 -616 1723
rect -582 1689 -258 1723
rect -224 1689 94 1723
rect 128 1689 446 1723
rect 480 1689 486 1723
rect -6185 1651 486 1689
rect -6185 1617 -6173 1651
rect -6139 1617 -5873 1651
rect -5839 1617 -5573 1651
rect -5539 1617 -5221 1651
rect -5187 1617 -5097 1651
rect -5063 1617 -4797 1651
rect -4763 1617 -4445 1651
rect -4411 1617 -4321 1651
rect -4287 1617 -3721 1651
rect -3687 1617 -3369 1651
rect -3335 1617 -3245 1651
rect -3211 1617 -2945 1651
rect -2911 1617 -2593 1651
rect -2559 1617 -2469 1651
rect -2435 1617 -1868 1651
rect -1834 1617 -1516 1651
rect -1482 1617 -1392 1651
rect -1358 1617 -1092 1651
rect -1058 1617 -740 1651
rect -706 1617 -616 1651
rect -582 1617 -258 1651
rect -224 1617 94 1651
rect 128 1617 446 1651
rect 480 1617 486 1651
rect -6185 1605 486 1617
rect -6185 1531 -570 1605
rect -1704 1494 -1259 1500
rect -1704 1460 -1692 1494
rect -1658 1460 -1305 1494
rect -1271 1460 -1259 1494
rect -1704 1454 -1259 1460
rect -11395 621 -9201 751
rect -5946 432 -400 444
rect -5946 398 -440 432
rect -406 398 -400 432
rect -446 360 -400 398
rect -446 326 -440 360
rect -406 326 -400 360
rect -446 314 -400 326
rect -6188 160 -2791 166
rect -6188 126 -4761 160
rect -4727 126 -4689 160
rect -4655 126 -2909 160
rect -2875 126 -2837 160
rect -2803 126 -2791 160
rect -6188 120 -2791 126
rect 320 137 372 143
rect 320 73 372 85
rect -6188 48 -6019 54
rect -6188 14 -6137 48
rect -6103 14 -6065 48
rect -6031 14 -6019 48
rect -6188 8 -6019 14
rect -5409 48 -5175 54
rect -5409 14 -5397 48
rect -5363 14 -5221 48
rect -5187 14 -5175 48
rect -5409 8 -5175 14
rect -4633 48 -4399 54
rect -4633 14 -4621 48
rect -4587 14 -4445 48
rect -4411 14 -4399 48
rect -4633 8 -4399 14
rect -3557 48 -3323 54
rect -3557 14 -3545 48
rect -3511 14 -3369 48
rect -3335 14 -3323 48
rect -3557 8 -3323 14
rect -2781 48 -2547 54
rect -2781 14 -2769 48
rect -2735 14 -2593 48
rect -2559 14 -2547 48
rect -2781 8 -2547 14
rect -1228 48 -1098 54
rect -1228 14 -1216 48
rect -1182 14 -1144 48
rect -1110 14 -1098 48
rect -1228 8 -1098 14
rect -928 48 -694 54
rect -928 14 -916 48
rect -882 14 -740 48
rect -706 14 -694 48
rect 320 15 372 21
rect -928 8 -694 14
rect -6185 -40 -228 -28
rect -6185 -74 -6173 -40
rect -6139 -74 -5873 -40
rect -5839 -74 -5573 -40
rect -5539 -74 -5097 -40
rect -5063 -74 -4797 -40
rect -4763 -74 -4321 -40
rect -4287 -74 -3721 -40
rect -3687 -74 -3245 -40
rect -3211 -74 -2945 -40
rect -2911 -74 -2469 -40
rect -2435 -74 -1868 -40
rect -1834 -74 -1392 -40
rect -1358 -74 -1092 -40
rect -1058 -74 -616 -40
rect -582 -74 -268 -40
rect -234 -74 -228 -40
rect -6185 -112 -228 -74
rect -6185 -146 -6173 -112
rect -6139 -146 -5873 -112
rect -5839 -146 -5573 -112
rect -5539 -146 -5097 -112
rect -5063 -146 -4797 -112
rect -4763 -146 -4321 -112
rect -4287 -146 -3721 -112
rect -3687 -146 -3245 -112
rect -3211 -146 -2945 -112
rect -2911 -146 -2469 -112
rect -2435 -146 -1868 -112
rect -1834 -146 -1392 -112
rect -1358 -146 -1092 -112
rect -1058 -146 -616 -112
rect -582 -146 -268 -112
rect -234 -146 -228 -112
rect -6185 -184 -228 -146
rect -6185 -218 -6173 -184
rect -6139 -218 -5873 -184
rect -5839 -218 -5573 -184
rect -5539 -218 -5097 -184
rect -5063 -218 -4797 -184
rect -4763 -218 -4321 -184
rect -4287 -218 -3721 -184
rect -3687 -218 -3245 -184
rect -3211 -218 -2945 -184
rect -2911 -218 -2469 -184
rect -2435 -218 -1868 -184
rect -1834 -218 -1392 -184
rect -1358 -218 -1092 -184
rect -1058 -218 -616 -184
rect -582 -218 -268 -184
rect -234 -218 -228 -184
rect -6185 -230 -228 -218
rect -99 -40 -53 -28
rect -99 -74 -93 -40
rect -59 -74 -53 -40
rect -99 -112 -53 -74
tri 289 -98 324 -63 se
rect 324 -83 370 15
rect 324 -98 355 -83
tri 355 -98 370 -83 nw
rect -99 -146 -93 -112
rect -59 -146 -53 -112
rect -99 -184 -53 -146
tri 223 -164 289 -98 se
tri 289 -164 355 -98 nw
tri 203 -184 223 -164 se
rect -99 -218 -93 -184
rect -59 -218 223 -184
rect -99 -230 223 -218
tri 223 -230 289 -164 nw
rect -228 -290 -98 -284
rect -6182 -300 -1522 -294
rect -6182 -334 -5344 -300
rect -5310 -334 -5272 -300
rect -5238 -334 -3494 -300
rect -3460 -334 -3422 -300
rect -3388 -334 -1640 -300
rect -1606 -334 -1568 -300
rect -1534 -334 -1522 -300
rect -6182 -340 -1522 -334
rect -1066 -300 -936 -294
rect -1066 -334 -1054 -300
rect -1020 -334 -982 -300
rect -948 -334 -936 -300
rect -1066 -340 -936 -334
rect -876 -300 -746 -294
rect -876 -334 -864 -300
rect -830 -334 -792 -300
rect -758 -334 -746 -300
rect -876 -340 -746 -334
rect -228 -324 -216 -290
rect -182 -324 -144 -290
rect -110 -324 -98 -290
rect -228 -495 -98 -324
rect -6636 -537 -2605 -531
rect -6636 -571 -6619 -537
rect -6585 -571 -6547 -537
rect -6513 -571 -5226 -537
rect -5192 -571 -5154 -537
rect -5120 -571 -3976 -537
rect -3942 -571 -3904 -537
rect -3870 -571 -2723 -537
rect -2689 -571 -2651 -537
rect -2617 -571 -2605 -537
rect -6636 -577 -2605 -571
rect -2440 -537 -2310 -531
rect -2440 -571 -2428 -537
rect -2394 -571 -2356 -537
rect -2322 -571 -2310 -537
rect -2440 -577 -2310 -571
rect -6677 -647 -6625 -641
rect -6677 -716 -6625 -699
rect -6677 -785 -6625 -768
tri -12350 -831 -12339 -820 se
rect -12339 -831 -10377 -820
tri -10377 -831 -10366 -820 sw
tri -12368 -849 -12350 -831 se
rect -12350 -849 -10366 -831
rect -12728 -905 -12598 -849
tri -12404 -885 -12368 -849 se
rect -12368 -851 -10366 -849
tri -10366 -851 -10346 -831 sw
rect -6677 -843 -6625 -837
rect -6499 -653 -1959 -641
rect -6499 -687 -6493 -653
rect -6459 -687 -6055 -653
rect -6021 -687 -5755 -653
rect -5721 -687 -5455 -653
rect -5421 -687 -4979 -653
rect -4945 -687 -4503 -653
rect -4469 -687 -4203 -653
rect -4169 -687 -3727 -653
rect -3693 -687 -3251 -653
rect -3217 -687 -2951 -653
rect -2917 -687 -2475 -653
rect -2441 -687 -1999 -653
rect -1965 -687 -1959 -653
rect -6499 -725 -1959 -687
rect -6499 -759 -6493 -725
rect -6459 -759 -6055 -725
rect -6021 -759 -5755 -725
rect -5721 -759 -5455 -725
rect -5421 -759 -4979 -725
rect -4945 -759 -4503 -725
rect -4469 -759 -4203 -725
rect -4169 -759 -3727 -725
rect -3693 -759 -3251 -725
rect -3217 -759 -2951 -725
rect -2917 -759 -2475 -725
rect -2441 -759 -1999 -725
rect -1965 -759 -1959 -725
rect -6499 -797 -1959 -759
rect -6499 -831 -6493 -797
rect -6459 -831 -6055 -797
rect -6021 -831 -5755 -797
rect -5721 -831 -5455 -797
rect -5421 -831 -4979 -797
rect -4945 -831 -4503 -797
rect -4469 -831 -4203 -797
rect -4169 -831 -3727 -797
rect -3693 -831 -3251 -797
rect -3217 -831 -2951 -797
rect -2917 -831 -2475 -797
rect -2441 -831 -1999 -797
rect -1965 -831 -1959 -797
rect -6499 -843 -1959 -831
rect -12368 -866 -10346 -851
rect -12368 -885 -12338 -866
tri -12338 -885 -12319 -866 nw
tri -10397 -885 -10378 -866 ne
rect -10378 -885 -10346 -866
tri -10346 -885 -10312 -851 sw
tri -12405 -886 -12404 -885 se
rect -12404 -886 -12339 -885
tri -12339 -886 -12338 -885 nw
tri -10378 -886 -10377 -885 ne
rect -10377 -886 -10312 -885
tri -12424 -905 -12405 -886 se
rect -12405 -905 -12372 -886
rect -12728 -919 -12372 -905
tri -12372 -919 -12339 -886 nw
tri -10377 -917 -10346 -886 ne
rect -10346 -917 -10312 -886
tri -10312 -917 -10280 -885 sw
rect -10004 -917 -9874 -849
rect -9146 -917 -9016 -849
rect -6070 -885 -5901 -879
rect -8657 -917 -8651 -911
tri -10346 -919 -10344 -917 ne
rect -10344 -919 -8651 -917
rect -12728 -951 -12404 -919
tri -12404 -951 -12372 -919 nw
tri -10344 -951 -10312 -919 ne
rect -10312 -951 -8651 -919
tri -10312 -963 -10300 -951 ne
rect -10300 -963 -8651 -951
rect -8599 -963 -8587 -911
rect -8535 -963 -8529 -911
rect -6070 -919 -6019 -885
rect -5985 -919 -5947 -885
rect -5913 -919 -5901 -885
rect -6070 -925 -5901 -919
rect -5291 -885 -5057 -879
rect -5291 -919 -5279 -885
rect -5245 -919 -5103 -885
rect -5069 -919 -5057 -885
rect -5291 -925 -5057 -919
rect -4815 -885 -4581 -879
rect -4815 -919 -4803 -885
rect -4769 -919 -4627 -885
rect -4593 -919 -4581 -885
rect -4815 -925 -4581 -919
rect -4039 -885 -3805 -879
rect -4039 -919 -4027 -885
rect -3993 -919 -3851 -885
rect -3817 -919 -3805 -885
rect -4039 -925 -3805 -919
rect -3563 -885 -3329 -879
rect -3563 -919 -3551 -885
rect -3517 -919 -3375 -885
rect -3341 -919 -3329 -885
rect -3563 -925 -3329 -919
rect -2787 -885 -2553 -879
rect -2787 -919 -2775 -885
rect -2741 -919 -2599 -885
rect -2565 -919 -2553 -885
rect -2787 -925 -2553 -919
rect -2311 -885 -2077 -879
rect -2311 -919 -2299 -885
rect -2265 -919 -2123 -885
rect -2089 -919 -2077 -885
rect -2311 -925 -2077 -919
rect -6070 -997 -3573 -991
rect -6070 -1031 -4943 -997
rect -4909 -1031 -4871 -997
rect -4837 -1031 -3691 -997
rect -3657 -1031 -3619 -997
rect -3585 -1031 -3573 -997
rect -6070 -1037 -3573 -1031
rect -6947 -1179 -1449 -1167
rect -6947 -1213 -6941 -1179
rect -6907 -1213 -6589 -1179
rect -6555 -1213 -6237 -1179
rect -6203 -1213 -6055 -1179
rect -6021 -1213 -5755 -1179
rect -5721 -1213 -5455 -1179
rect -5421 -1213 -5103 -1179
rect -5069 -1213 -4979 -1179
rect -4945 -1213 -4627 -1179
rect -4593 -1213 -4503 -1179
rect -4469 -1213 -4203 -1179
rect -4169 -1213 -3851 -1179
rect -3817 -1213 -3727 -1179
rect -3693 -1213 -3375 -1179
rect -3341 -1213 -3251 -1179
rect -3217 -1213 -2951 -1179
rect -2917 -1213 -2599 -1179
rect -2565 -1213 -2475 -1179
rect -2441 -1213 -2123 -1179
rect -2089 -1213 -1999 -1179
rect -1965 -1213 -1449 -1179
rect -12406 -1279 -8954 -1233
rect -6947 -1251 -1449 -1213
rect -6947 -1285 -6941 -1251
rect -6907 -1285 -6589 -1251
rect -6555 -1285 -6237 -1251
rect -6203 -1285 -6055 -1251
rect -6021 -1285 -5755 -1251
rect -5721 -1285 -5455 -1251
rect -5421 -1285 -5103 -1251
rect -5069 -1285 -4979 -1251
rect -4945 -1285 -4627 -1251
rect -4593 -1285 -4503 -1251
rect -4469 -1285 -4203 -1251
rect -4169 -1285 -3851 -1251
rect -3817 -1285 -3727 -1251
rect -3693 -1285 -3375 -1251
rect -3341 -1285 -3251 -1251
rect -3217 -1285 -2951 -1251
rect -2917 -1285 -2599 -1251
rect -2565 -1285 -2475 -1251
rect -2441 -1285 -2123 -1251
rect -2089 -1285 -1999 -1251
rect -1965 -1285 -1449 -1251
rect -6947 -1323 -1449 -1285
rect -6947 -1357 -6941 -1323
rect -6907 -1357 -6589 -1323
rect -6555 -1357 -6237 -1323
rect -6203 -1357 -6055 -1323
rect -6021 -1357 -5755 -1323
rect -5721 -1357 -5455 -1323
rect -5421 -1357 -5103 -1323
rect -5069 -1357 -4979 -1323
rect -4945 -1357 -4627 -1323
rect -4593 -1357 -4503 -1323
rect -4469 -1357 -4203 -1323
rect -4169 -1357 -3851 -1323
rect -3817 -1357 -3727 -1323
rect -3693 -1357 -3375 -1323
rect -3341 -1357 -3251 -1323
rect -3217 -1357 -2951 -1323
rect -2917 -1357 -2599 -1323
rect -2565 -1357 -2475 -1323
rect -2441 -1357 -2123 -1323
rect -2089 -1357 -1999 -1323
rect -1965 -1357 -1449 -1323
rect -6947 -1369 -1449 -1357
rect -4724 -1422 -4678 -1410
rect -4724 -1452 -4718 -1422
rect -6070 -1456 -4718 -1452
rect -4684 -1456 -4678 -1422
rect -6070 -1494 -4678 -1456
rect -6070 -1498 -4718 -1494
rect -4724 -1528 -4718 -1498
rect -4684 -1528 -4678 -1494
rect -4724 -1540 -4678 -1528
rect -4033 -1421 -3987 -1409
rect -4033 -1455 -4027 -1421
rect -3993 -1451 -3987 -1421
rect -3993 -1455 -2510 -1451
rect -4033 -1493 -2510 -1455
rect -4033 -1527 -4027 -1493
rect -3993 -1497 -2510 -1493
rect -3993 -1527 -3987 -1497
rect -4033 -1539 -3987 -1527
rect -11676 -1550 -8162 -1544
tri -8162 -1550 -8156 -1544 sw
rect -3468 -1550 -3422 -1538
rect -11676 -1584 -8156 -1550
tri -8156 -1584 -8122 -1550 sw
rect -3468 -1580 -3462 -1550
rect -6070 -1584 -3462 -1580
rect -3428 -1584 -3422 -1550
rect -11676 -1585 -8122 -1584
tri -8122 -1585 -8121 -1584 sw
rect -11676 -1590 -8094 -1585
tri -8182 -1622 -8150 -1590 ne
rect -8150 -1622 -8094 -1590
tri -8150 -1631 -8141 -1622 ne
rect -8141 -1631 -8094 -1622
rect -6070 -1622 -3422 -1584
rect -6070 -1626 -3462 -1622
rect -5285 -1667 -5239 -1655
rect -6895 -1698 -6373 -1692
rect -6895 -1704 -6677 -1698
rect -6895 -1738 -6765 -1704
rect -6731 -1738 -6677 -1704
rect -6895 -1750 -6677 -1738
rect -6625 -1704 -6373 -1698
rect -6625 -1738 -6413 -1704
rect -6379 -1738 -6373 -1704
rect -6625 -1750 -6373 -1738
rect -6895 -1764 -6373 -1750
rect -6895 -1776 -6677 -1764
rect -6895 -1810 -6765 -1776
rect -6731 -1810 -6677 -1776
rect -6895 -1816 -6677 -1810
rect -6625 -1776 -6373 -1764
rect -6625 -1810 -6413 -1776
rect -6379 -1810 -6373 -1776
rect -5285 -1701 -5279 -1667
rect -5245 -1697 -5239 -1667
rect -3468 -1656 -3462 -1626
rect -3428 -1656 -3422 -1622
rect -3468 -1668 -3422 -1656
rect -5245 -1701 -2510 -1697
rect -5285 -1739 -2510 -1701
rect -5285 -1773 -5279 -1739
rect -5245 -1743 -2510 -1739
rect -5245 -1773 -5239 -1743
rect -5285 -1785 -5239 -1773
rect -6625 -1816 -6373 -1810
rect -6895 -1822 -6373 -1816
rect -11676 -2660 -11670 -2608
rect -11618 -2660 -11606 -2608
rect -11554 -2660 -11548 -2608
rect -11056 -2660 -11050 -2608
rect -10998 -2660 -10986 -2608
rect -10934 -2660 -10928 -2608
rect -8094 -2660 -8088 -2608
rect -8036 -2660 -8024 -2608
rect -7972 -2660 -7966 -2608
rect -7474 -2660 -7468 -2608
rect -7416 -2660 -7404 -2608
rect -7352 -2660 -7346 -2608
rect -4512 -2660 -4506 -2608
rect -4454 -2660 -4442 -2608
rect -4390 -2660 -4384 -2608
rect -3892 -2660 -3886 -2608
rect -3834 -2660 -3822 -2608
rect -3770 -2660 -3764 -2608
rect -12022 -2963 -12016 -2960
rect -12406 -3009 -12016 -2963
rect -12022 -3012 -12016 -3009
rect -11964 -3012 -11952 -2960
rect -11900 -3012 -11894 -2960
rect -10196 -3012 -10190 -2960
rect -10138 -3012 -10126 -2960
rect -10074 -3012 -10068 -2960
rect -8954 -3012 -8948 -2960
rect -8896 -3012 -8884 -2960
rect -8832 -3012 -8826 -2960
rect -6614 -3012 -6608 -2960
rect -6556 -3012 -6544 -2960
rect -6492 -3012 -6486 -2960
rect -5372 -3012 -5366 -2960
rect -5314 -3012 -5302 -2960
rect -5250 -3012 -5244 -2960
rect -3030 -3012 -3024 -2960
rect -2972 -3012 -2960 -2960
rect -2908 -3012 -2902 -2960
rect -12099 -3268 -12093 -3265
rect -12657 -3314 -12093 -3268
rect -12657 -3393 -12529 -3314
rect -12099 -3317 -12093 -3314
rect -12041 -3317 -12029 -3265
rect -11977 -3317 -11971 -3265
rect -10075 -3345 -10069 -3293
rect -10017 -3345 -10005 -3293
rect -9953 -3345 -9947 -3293
rect -10075 -3393 -9947 -3345
rect -9075 -3345 -9069 -3293
rect -9017 -3345 -9005 -3293
rect -8953 -3345 -8947 -3293
rect -9075 -3393 -8947 -3345
rect -6493 -3345 -6487 -3293
rect -6435 -3345 -6423 -3293
rect -6371 -3345 -6365 -3293
rect -6493 -3393 -6365 -3345
rect -5491 -3345 -5485 -3293
rect -5433 -3345 -5421 -3293
rect -5369 -3345 -5363 -3293
rect -5491 -3393 -5363 -3345
rect -2911 -3345 -2905 -3293
rect -2853 -3345 -2841 -3293
rect -2789 -3345 -2783 -3293
rect -2911 -3393 -2783 -3345
<< via1 >>
rect 320 1921 372 1973
rect 320 1857 372 1909
rect 320 85 372 137
rect 320 21 372 73
rect -6677 -653 -6625 -647
rect -6677 -687 -6669 -653
rect -6669 -687 -6635 -653
rect -6635 -687 -6625 -653
rect -6677 -699 -6625 -687
rect -6677 -725 -6625 -716
rect -6677 -759 -6669 -725
rect -6669 -759 -6635 -725
rect -6635 -759 -6625 -725
rect -6677 -768 -6625 -759
rect -6677 -797 -6625 -785
rect -6677 -831 -6669 -797
rect -6669 -831 -6635 -797
rect -6635 -831 -6625 -797
rect -6677 -837 -6625 -831
rect -8651 -963 -8599 -911
rect -8587 -963 -8535 -911
rect -6677 -1750 -6625 -1698
rect -6677 -1816 -6625 -1764
rect -11670 -2660 -11618 -2608
rect -11606 -2660 -11554 -2608
rect -11050 -2660 -10998 -2608
rect -10986 -2660 -10934 -2608
rect -8088 -2660 -8036 -2608
rect -8024 -2660 -7972 -2608
rect -7468 -2660 -7416 -2608
rect -7404 -2660 -7352 -2608
rect -4506 -2660 -4454 -2608
rect -4442 -2660 -4390 -2608
rect -3886 -2660 -3834 -2608
rect -3822 -2660 -3770 -2608
rect -12016 -3012 -11964 -2960
rect -11952 -3012 -11900 -2960
rect -10190 -3012 -10138 -2960
rect -10126 -3012 -10074 -2960
rect -8948 -3012 -8896 -2960
rect -8884 -3012 -8832 -2960
rect -6608 -3012 -6556 -2960
rect -6544 -3012 -6492 -2960
rect -5366 -3012 -5314 -2960
rect -5302 -3012 -5250 -2960
rect -3024 -3012 -2972 -2960
rect -2960 -3012 -2908 -2960
rect -12093 -3317 -12041 -3265
rect -12029 -3317 -11977 -3265
rect -10069 -3345 -10017 -3293
rect -10005 -3345 -9953 -3293
rect -9069 -3345 -9017 -3293
rect -9005 -3345 -8953 -3293
rect -6487 -3345 -6435 -3293
rect -6423 -3345 -6371 -3293
rect -5485 -3345 -5433 -3293
rect -5421 -3345 -5369 -3293
rect -2905 -3345 -2853 -3293
rect -2841 -3345 -2789 -3293
<< metal2 >>
rect 320 1973 372 1979
rect 320 1909 372 1921
rect 320 1851 372 1857
rect 324 143 370 1851
rect 320 137 372 143
rect 320 73 372 85
rect 320 15 372 21
rect -6677 -647 -6625 -641
rect -6677 -716 -6625 -699
rect -6677 -785 -6625 -768
rect -8657 -963 -8651 -911
rect -8599 -963 -8587 -911
rect -8535 -963 -8529 -911
rect -8597 -2266 -8545 -963
rect -6677 -1698 -6625 -837
rect -6677 -1764 -6625 -1750
tri -6719 -2244 -6677 -2202 se
rect -6677 -2224 -6625 -1816
tri -8597 -2318 -8545 -2266 ne
tri -8545 -2316 -8473 -2244 sw
tri -6751 -2276 -6719 -2244 se
rect -6719 -2276 -6677 -2244
tri -6677 -2276 -6625 -2224 nw
tri -6791 -2316 -6751 -2276 se
rect -6751 -2316 -6717 -2276
tri -6717 -2316 -6677 -2276 nw
rect -8545 -2318 -6769 -2316
tri -8545 -2368 -8495 -2318 ne
rect -8495 -2368 -6769 -2318
tri -6769 -2368 -6717 -2316 nw
rect -11676 -2660 -11670 -2608
rect -11618 -2660 -11606 -2608
rect -11554 -2660 -11050 -2608
rect -10998 -2660 -10986 -2608
rect -10934 -2660 -8088 -2608
rect -8036 -2660 -8024 -2608
rect -7972 -2660 -7468 -2608
rect -7416 -2660 -7404 -2608
rect -7352 -2660 -4506 -2608
rect -4454 -2660 -4442 -2608
rect -4390 -2660 -3886 -2608
rect -3834 -2660 -3822 -2608
rect -3770 -2660 -3764 -2608
rect -12022 -3012 -12016 -2960
rect -11964 -3012 -11952 -2960
rect -11900 -3012 -10190 -2960
rect -10138 -3012 -10126 -2960
rect -10074 -3012 -8948 -2960
rect -8896 -3012 -8884 -2960
rect -8832 -3012 -6608 -2960
rect -6556 -3012 -6544 -2960
rect -6492 -3012 -5366 -2960
rect -5314 -3012 -5302 -2960
rect -5250 -3012 -3024 -2960
rect -2972 -3012 -2960 -2960
rect -2908 -3012 -2902 -2960
rect -12099 -3317 -12093 -3265
rect -12041 -3317 -12029 -3265
rect -11977 -3293 -11971 -3265
rect -11977 -3317 -10069 -3293
rect -12099 -3345 -10069 -3317
rect -10017 -3345 -10005 -3293
rect -9953 -3345 -9069 -3293
rect -9017 -3345 -9005 -3293
rect -8953 -3345 -6487 -3293
rect -6435 -3345 -6423 -3293
rect -6371 -3345 -5485 -3293
rect -5433 -3345 -5421 -3293
rect -5369 -3345 -2905 -3293
rect -2853 -3345 -2841 -3293
rect -2789 -3345 -2158 -3293
tri -2158 -3345 -2106 -3293 sw
tri -2180 -3419 -2106 -3345 ne
tri -2106 -3419 -2032 -3345 sw
tri -2106 -3493 -2032 -3419 ne
tri -2032 -3493 -1958 -3419 sw
tri -2032 -3567 -1958 -3493 ne
tri -1958 -3542 -1909 -3493 sw
rect -1958 -3567 -1582 -3542
tri -1958 -3594 -1931 -3567 ne
rect -1931 -3594 -1582 -3567
use hvnTran_CDNS_52468879185403  hvnTran_CDNS_52468879185403_0
timestamp 1704896540
transform -1 0 -2610 0 1 -819
box -79 -26 196 226
use hvnTran_CDNS_52468879185403  hvnTran_CDNS_52468879185403_1
timestamp 1704896540
transform -1 0 -3386 0 1 -819
box -79 -26 196 226
use hvnTran_CDNS_52468879185403  hvnTran_CDNS_52468879185403_2
timestamp 1704896540
transform -1 0 -3862 0 1 -819
box -79 -26 196 226
use hvnTran_CDNS_52468879185403  hvnTran_CDNS_52468879185403_3
timestamp 1704896540
transform -1 0 -4638 0 1 -819
box -79 -26 196 226
use hvnTran_CDNS_52468879185403  hvnTran_CDNS_52468879185403_4
timestamp 1704896540
transform -1 0 -5114 0 1 -819
box -79 -26 196 226
use hvnTran_CDNS_52468879185403  hvnTran_CDNS_52468879185403_5
timestamp 1704896540
transform -1 0 -2134 0 1 -819
box -79 -26 196 226
use hvnTran_CDNS_52468879185403  hvnTran_CDNS_52468879185403_6
timestamp 1704896540
transform -1 0 -4456 0 -1 -52
box -79 -26 196 226
use hvnTran_CDNS_52468879185403  hvnTran_CDNS_52468879185403_7
timestamp 1704896540
transform -1 0 -5232 0 -1 -52
box -79 -26 196 226
use hvnTran_CDNS_52468879185403  hvnTran_CDNS_52468879185403_8
timestamp 1704896540
transform -1 0 -1527 0 -1 -52
box -79 -26 196 226
use hvnTran_CDNS_52468879185403  hvnTran_CDNS_52468879185403_9
timestamp 1704896540
transform -1 0 -2604 0 -1 -52
box -79 -26 196 226
use hvnTran_CDNS_52468879185403  hvnTran_CDNS_52468879185403_10
timestamp 1704896540
transform -1 0 -3380 0 -1 -52
box -79 -26 196 226
use hvnTran_CDNS_52468879185403  hvnTran_CDNS_52468879185403_11
timestamp 1704896540
transform -1 0 -751 0 -1 -52
box -79 -26 196 226
use hvnTran_CDNS_52468879185403  hvnTran_CDNS_52468879185403_12
timestamp 1704896540
transform 1 0 -5528 0 -1 -52
box -79 -26 196 226
use hvnTran_CDNS_52468879185403  hvnTran_CDNS_52468879185403_13
timestamp 1704896540
transform 1 0 -1823 0 -1 -52
box -79 -26 196 226
use hvnTran_CDNS_52468879185403  hvnTran_CDNS_52468879185403_14
timestamp 1704896540
transform 1 0 -2900 0 -1 -52
box -79 -26 196 226
use hvnTran_CDNS_52468879185403  hvnTran_CDNS_52468879185403_15
timestamp 1704896540
transform 1 0 -3676 0 -1 -52
box -79 -26 196 226
use hvnTran_CDNS_52468879185403  hvnTran_CDNS_52468879185403_16
timestamp 1704896540
transform 1 0 -4752 0 -1 -52
box -79 -26 196 226
use hvnTran_CDNS_52468879185403  hvnTran_CDNS_52468879185403_17
timestamp 1704896540
transform 1 0 -1047 0 -1 -52
box -79 -26 196 226
use hvnTran_CDNS_52468879185403  hvnTran_CDNS_52468879185403_18
timestamp 1704896540
transform 1 0 -2906 0 1 -819
box -79 -26 196 226
use hvnTran_CDNS_52468879185403  hvnTran_CDNS_52468879185403_19
timestamp 1704896540
transform 1 0 -3682 0 1 -819
box -79 -26 196 226
use hvnTran_CDNS_52468879185403  hvnTran_CDNS_52468879185403_20
timestamp 1704896540
transform 1 0 -4158 0 1 -819
box -79 -26 196 226
use hvnTran_CDNS_52468879185403  hvnTran_CDNS_52468879185403_21
timestamp 1704896540
transform 1 0 -4934 0 1 -819
box -79 -26 196 226
use hvnTran_CDNS_52468879185403  hvnTran_CDNS_52468879185403_22
timestamp 1704896540
transform 1 0 -5410 0 1 -819
box -79 -26 196 226
use hvnTran_CDNS_52468879185403  hvnTran_CDNS_52468879185403_23
timestamp 1704896540
transform 1 0 -2430 0 1 -819
box -79 -26 196 226
use hvnTran_CDNS_52468879185404  hvnTran_CDNS_52468879185404_0
timestamp 1704896540
transform 1 0 -4276 0 -1 -52
box -79 -26 199 226
use hvnTran_CDNS_52468879185404  hvnTran_CDNS_52468879185404_1
timestamp 1704896540
transform 1 0 -5828 0 -1 -52
box -79 -26 199 226
use hvnTran_CDNS_52468879185404  hvnTran_CDNS_52468879185404_2
timestamp 1704896540
transform 1 0 -6128 0 -1 -52
box -79 -26 199 226
use hvnTran_CDNS_52468879185404  hvnTran_CDNS_52468879185404_3
timestamp 1704896540
transform 1 0 -1347 0 -1 -52
box -79 -26 199 226
use hvnTran_CDNS_52468879185404  hvnTran_CDNS_52468879185404_4
timestamp 1704896540
transform 1 0 -2424 0 -1 -52
box -79 -26 199 226
use hvnTran_CDNS_52468879185404  hvnTran_CDNS_52468879185404_5
timestamp 1704896540
transform 1 0 -5052 0 -1 -52
box -79 -26 199 226
use hvnTran_CDNS_52468879185404  hvnTran_CDNS_52468879185404_6
timestamp 1704896540
transform 1 0 -3200 0 -1 -52
box -79 -26 199 226
use hvnTran_CDNS_52468879185404  hvnTran_CDNS_52468879185404_7
timestamp 1704896540
transform 1 0 -571 0 -1 -52
box -79 -26 199 226
use hvnTran_CDNS_52468879185404  hvnTran_CDNS_52468879185404_8
timestamp 1704896540
transform 1 0 -3206 0 1 -819
box -79 -26 199 226
use hvnTran_CDNS_52468879185404  hvnTran_CDNS_52468879185404_9
timestamp 1704896540
transform 1 0 -4458 0 1 -819
box -79 -26 199 226
use hvnTran_CDNS_52468879185404  hvnTran_CDNS_52468879185404_10
timestamp 1704896540
transform 1 0 -5710 0 1 -819
box -79 -26 199 226
use hvnTran_CDNS_52468879185404  hvnTran_CDNS_52468879185404_11
timestamp 1704896540
transform 1 0 -6010 0 1 -819
box -79 -26 199 226
use hvnTran_CDNS_52468879185404  hvnTran_CDNS_52468879185404_12
timestamp 1704896540
transform 1 0 -1954 0 1 -819
box -79 -26 199 226
use hvpTran_CDNS_52468879185405  hvpTran_CDNS_52468879185405_0
timestamp 1704896540
transform 1 0 -2906 0 -1 -1171
box -119 -66 415 666
use hvpTran_CDNS_52468879185405  hvpTran_CDNS_52468879185405_1
timestamp 1704896540
transform 1 0 -3682 0 -1 -1171
box -119 -66 415 666
use hvpTran_CDNS_52468879185405  hvpTran_CDNS_52468879185405_2
timestamp 1704896540
transform 1 0 -4158 0 -1 -1171
box -119 -66 415 666
use hvpTran_CDNS_52468879185405  hvpTran_CDNS_52468879185405_3
timestamp 1704896540
transform 1 0 -4934 0 -1 -1171
box -119 -66 415 666
use hvpTran_CDNS_52468879185405  hvpTran_CDNS_52468879185405_4
timestamp 1704896540
transform 1 0 -5410 0 -1 -1171
box -119 -66 415 666
use hvpTran_CDNS_52468879185405  hvpTran_CDNS_52468879185405_5
timestamp 1704896540
transform 1 0 -2430 0 -1 -1171
box -119 -66 415 666
use hvpTran_CDNS_52468879185405  hvpTran_CDNS_52468879185405_6
timestamp 1704896540
transform 1 0 -1823 0 1 1609
box -119 -66 415 666
use hvpTran_CDNS_52468879185405  hvpTran_CDNS_52468879185405_7
timestamp 1704896540
transform 1 0 -2900 0 1 1609
box -119 -66 415 666
use hvpTran_CDNS_52468879185405  hvpTran_CDNS_52468879185405_8
timestamp 1704896540
transform 1 0 -3676 0 1 1609
box -119 -66 415 666
use hvpTran_CDNS_52468879185405  hvpTran_CDNS_52468879185405_9
timestamp 1704896540
transform 1 0 -4752 0 1 1609
box -119 -66 415 666
use hvpTran_CDNS_52468879185405  hvpTran_CDNS_52468879185405_10
timestamp 1704896540
transform 1 0 -5528 0 1 1609
box -119 -66 415 666
use hvpTran_CDNS_52468879185405  hvpTran_CDNS_52468879185405_11
timestamp 1704896540
transform 1 0 -1047 0 1 1609
box -119 -66 415 666
use hvpTran_CDNS_52468879185406  hvpTran_CDNS_52468879185406_0
timestamp 1704896540
transform 1 0 -5710 0 -1 -1171
box -119 -66 239 666
use hvpTran_CDNS_52468879185406  hvpTran_CDNS_52468879185406_1
timestamp 1704896540
transform 1 0 -3206 0 -1 -1171
box -119 -66 239 666
use hvpTran_CDNS_52468879185406  hvpTran_CDNS_52468879185406_2
timestamp 1704896540
transform 1 0 -4458 0 -1 -1171
box -119 -66 239 666
use hvpTran_CDNS_52468879185406  hvpTran_CDNS_52468879185406_3
timestamp 1704896540
transform 1 0 -6010 0 -1 -1171
box -119 -66 239 666
use hvpTran_CDNS_52468879185406  hvpTran_CDNS_52468879185406_4
timestamp 1704896540
transform 1 0 -1954 0 -1 -1171
box -119 -66 239 666
use hvpTran_CDNS_52468879185406  hvpTran_CDNS_52468879185406_5
timestamp 1704896540
transform 1 0 -5828 0 1 1609
box -119 -66 239 666
use hvpTran_CDNS_52468879185406  hvpTran_CDNS_52468879185406_6
timestamp 1704896540
transform 1 0 -6128 0 1 1609
box -119 -66 239 666
use hvpTran_CDNS_52468879185406  hvpTran_CDNS_52468879185406_7
timestamp 1704896540
transform 1 0 -4276 0 1 1609
box -119 -66 239 666
use hvpTran_CDNS_52468879185406  hvpTran_CDNS_52468879185406_8
timestamp 1704896540
transform 1 0 -1347 0 1 1609
box -119 -66 239 666
use hvpTran_CDNS_52468879185406  hvpTran_CDNS_52468879185406_9
timestamp 1704896540
transform 1 0 -2424 0 1 1609
box -119 -66 239 666
use hvpTran_CDNS_52468879185406  hvpTran_CDNS_52468879185406_10
timestamp 1704896540
transform 1 0 -5052 0 1 1609
box -119 -66 239 666
use hvpTran_CDNS_52468879185406  hvpTran_CDNS_52468879185406_11
timestamp 1704896540
transform 1 0 -3200 0 1 1609
box -119 -66 239 666
use hvpTran_CDNS_52468879185406  hvpTran_CDNS_52468879185406_12
timestamp 1704896540
transform 1 0 -571 0 1 1609
box -119 -66 239 666
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1704896540
transform 0 -1 -1834 -1 0 -40
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_1
timestamp 1704896540
transform 0 -1 -5539 -1 0 -40
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_2
timestamp 1704896540
transform 0 -1 -5839 -1 0 -40
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_3
timestamp 1704896540
transform 0 -1 -2911 -1 0 -40
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_4
timestamp 1704896540
transform 0 -1 -6139 -1 0 -40
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_5
timestamp 1704896540
transform 0 -1 -234 -1 0 -40
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_6
timestamp 1704896540
transform 0 -1 -3687 -1 0 -40
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_7
timestamp 1704896540
transform 0 -1 -59 -1 0 -40
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_8
timestamp 1704896540
transform 0 -1 -4287 -1 0 -40
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_9
timestamp 1704896540
transform 0 -1 -4763 -1 0 -40
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_10
timestamp 1704896540
transform 0 -1 -2565 -1 0 -1179
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_11
timestamp 1704896540
transform 0 -1 -2917 -1 0 -1179
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_12
timestamp 1704896540
transform 0 -1 -3217 -1 0 -1179
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_13
timestamp 1704896540
transform 0 -1 -3341 -1 0 -1179
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_14
timestamp 1704896540
transform 0 -1 -3693 -1 0 -1179
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_15
timestamp 1704896540
transform 0 -1 -3817 -1 0 -1179
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_16
timestamp 1704896540
transform 0 -1 -4169 -1 0 -1179
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_17
timestamp 1704896540
transform 0 -1 -4469 -1 0 -1179
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_18
timestamp 1704896540
transform 0 -1 -4593 -1 0 -1179
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_19
timestamp 1704896540
transform 0 -1 -4945 -1 0 -1179
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_20
timestamp 1704896540
transform 0 -1 -5069 -1 0 -1179
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_21
timestamp 1704896540
transform 0 -1 -5421 -1 0 -1179
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_22
timestamp 1704896540
transform 0 -1 -5721 -1 0 -1179
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_23
timestamp 1704896540
transform 0 -1 -6021 -1 0 -1179
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_24
timestamp 1704896540
transform 0 -1 -1358 -1 0 -40
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_25
timestamp 1704896540
transform 0 -1 -2435 -1 0 -40
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_26
timestamp 1704896540
transform 0 -1 -5063 -1 0 -40
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_27
timestamp 1704896540
transform 0 -1 -3211 -1 0 -40
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_28
timestamp 1704896540
transform 0 -1 -2441 -1 0 -1179
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_29
timestamp 1704896540
transform 0 -1 -2089 -1 0 -1179
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_30
timestamp 1704896540
transform 0 -1 -1965 -1 0 -1179
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_31
timestamp 1704896540
transform 0 -1 -582 -1 0 -40
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_32
timestamp 1704896540
transform 0 -1 -1058 -1 0 -40
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_33
timestamp 1704896540
transform 0 -1 -6203 -1 0 -1179
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_34
timestamp 1704896540
transform 0 -1 -6555 -1 0 -1179
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_35
timestamp 1704896540
transform 0 -1 -6907 -1 0 -1179
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_36
timestamp 1704896540
transform 0 -1 -5187 1 0 1617
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_37
timestamp 1704896540
transform 0 -1 -1834 1 0 1617
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_38
timestamp 1704896540
transform 0 -1 -1482 1 0 1617
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_39
timestamp 1704896540
transform 0 -1 -2559 1 0 1617
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_40
timestamp 1704896540
transform 0 -1 -5539 1 0 1617
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_41
timestamp 1704896540
transform 0 -1 -2911 1 0 1617
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_42
timestamp 1704896540
transform 0 -1 -5839 1 0 1617
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_43
timestamp 1704896540
transform 0 -1 -6139 1 0 1617
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_44
timestamp 1704896540
transform 0 -1 -3335 1 0 1617
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_45
timestamp 1704896540
transform 0 -1 -3687 1 0 1617
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_46
timestamp 1704896540
transform 0 -1 -4287 1 0 1617
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_47
timestamp 1704896540
transform 0 -1 -4411 1 0 1617
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_48
timestamp 1704896540
transform 0 -1 -4763 1 0 1617
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_49
timestamp 1704896540
transform 0 -1 -2917 1 0 -831
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_50
timestamp 1704896540
transform 0 -1 -3217 1 0 -831
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_51
timestamp 1704896540
transform 0 -1 -3693 1 0 -831
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_52
timestamp 1704896540
transform 0 -1 -4169 1 0 -831
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_53
timestamp 1704896540
transform 0 -1 -4469 1 0 -831
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_54
timestamp 1704896540
transform 0 -1 -4945 1 0 -831
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_55
timestamp 1704896540
transform 0 -1 -5421 1 0 -831
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_56
timestamp 1704896540
transform 0 -1 -5721 1 0 -831
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_57
timestamp 1704896540
transform 0 -1 -6021 1 0 -831
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_58
timestamp 1704896540
transform 0 -1 -1358 1 0 1617
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_59
timestamp 1704896540
transform 0 -1 -2435 1 0 1617
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_60
timestamp 1704896540
transform 0 -1 -5063 1 0 1617
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_61
timestamp 1704896540
transform 0 -1 -3211 1 0 1617
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_62
timestamp 1704896540
transform 0 -1 -2441 1 0 -831
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_63
timestamp 1704896540
transform 0 -1 -1965 1 0 -831
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_64
timestamp 1704896540
transform 0 -1 -1058 1 0 1617
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_65
timestamp 1704896540
transform 0 -1 -706 1 0 1617
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_66
timestamp 1704896540
transform 0 -1 -582 1 0 1617
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_67
timestamp 1704896540
transform 0 -1 -6459 1 0 -831
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_68
timestamp 1704896540
transform 0 -1 -6635 1 0 -831
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_0
timestamp 1704896540
transform 1 0 -5221 0 -1 48
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_1
timestamp 1704896540
transform 1 0 -5397 0 -1 48
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_2
timestamp 1704896540
transform 1 0 -4445 0 -1 48
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_3
timestamp 1704896540
transform 1 0 -4621 0 -1 48
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_4
timestamp 1704896540
transform 1 0 -2769 0 -1 48
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_5
timestamp 1704896540
transform 1 0 -3369 0 -1 48
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_6
timestamp 1704896540
transform 1 0 -2593 0 -1 48
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_7
timestamp 1704896540
transform 1 0 -3545 0 -1 48
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_8
timestamp 1704896540
transform 1 0 -1305 0 -1 1494
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_9
timestamp 1704896540
transform 1 0 -1692 0 -1 1494
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_10
timestamp 1704896540
transform 1 0 -916 0 -1 48
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_11
timestamp 1704896540
transform 1 0 -740 0 -1 48
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_12
timestamp 1704896540
transform 1 0 -3551 0 1 -919
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_13
timestamp 1704896540
transform 1 0 -3375 0 1 -919
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_14
timestamp 1704896540
transform 1 0 -2775 0 1 -919
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_15
timestamp 1704896540
transform 1 0 -2599 0 1 -919
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_16
timestamp 1704896540
transform 1 0 -4027 0 1 -919
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_17
timestamp 1704896540
transform 1 0 -3851 0 1 -919
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_18
timestamp 1704896540
transform 1 0 -4803 0 1 -919
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_19
timestamp 1704896540
transform 1 0 -4627 0 1 -919
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_20
timestamp 1704896540
transform 1 0 -5279 0 1 -919
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_21
timestamp 1704896540
transform 1 0 -5103 0 1 -919
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_22
timestamp 1704896540
transform 1 0 -2123 0 1 -919
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_23
timestamp 1704896540
transform 1 0 -2299 0 1 -919
box 0 0 1 1
use nfet_CDNS_52468879185797  nfet_CDNS_52468879185797_0
timestamp 1704896540
transform 1 0 -6624 0 -1 -619
box -79 -32 199 232
use nfet_CDNS_52468879185797  nfet_CDNS_52468879185797_1
timestamp 1704896540
transform 1 0 -224 0 -1 -42
box -79 -32 199 232
use pfet_CDNS_52468879185917  pfet_CDNS_52468879185917_0
timestamp 1704896540
transform 1 0 -213 0 -1 2209
box -119 -66 767 666
use pfet_CDNS_52468879185917  pfet_CDNS_52468879185917_1
timestamp 1704896540
transform 1 0 -6896 0 1 -1771
box -119 -66 767 666
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_0
timestamp 1704896540
transform -1 0 -4149 0 1 -350
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_1
timestamp 1704896540
transform -1 0 -5701 0 1 -350
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_2
timestamp 1704896540
transform -1 0 -6001 0 1 -350
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_3
timestamp 1704896540
transform -1 0 -1220 0 1 -350
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_4
timestamp 1704896540
transform -1 0 -2297 0 1 -350
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_5
timestamp 1704896540
transform -1 0 -4925 0 1 -350
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_6
timestamp 1704896540
transform -1 0 -3073 0 1 -350
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_7
timestamp 1704896540
transform -1 0 -444 0 1 -350
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_8
timestamp 1704896540
transform -1 0 -4149 0 -1 2307
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_9
timestamp 1704896540
transform -1 0 -5701 0 -1 2307
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_10
timestamp 1704896540
transform -1 0 -6001 0 -1 2307
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_11
timestamp 1704896540
transform -1 0 -3079 0 -1 -521
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_12
timestamp 1704896540
transform -1 0 -4331 0 -1 -521
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_13
timestamp 1704896540
transform -1 0 -5583 0 -1 -521
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_14
timestamp 1704896540
transform -1 0 -5883 0 -1 -521
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_15
timestamp 1704896540
transform -1 0 -1220 0 -1 2307
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_16
timestamp 1704896540
transform -1 0 -2297 0 -1 2307
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_17
timestamp 1704896540
transform -1 0 -4925 0 -1 2307
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_18
timestamp 1704896540
transform -1 0 -3073 0 -1 2307
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_19
timestamp 1704896540
transform -1 0 -1827 0 -1 -521
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_20
timestamp 1704896540
transform -1 0 -444 0 -1 2307
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_21
timestamp 1704896540
transform 1 0 -3507 0 -1 2307
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_22
timestamp 1704896540
transform 1 0 -3683 0 -1 2307
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_23
timestamp 1704896540
transform 1 0 -5359 0 -1 2307
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_24
timestamp 1704896540
transform 1 0 -5535 0 -1 2307
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_25
timestamp 1704896540
transform 1 0 -2731 0 -1 2307
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_26
timestamp 1704896540
transform 1 0 -1830 0 -1 2307
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_27
timestamp 1704896540
transform 1 0 -2907 0 -1 2307
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_28
timestamp 1704896540
transform 1 0 -1654 0 -1 2307
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_29
timestamp 1704896540
transform 1 0 -4583 0 -1 2307
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_30
timestamp 1704896540
transform 1 0 -4759 0 -1 2307
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_31
timestamp 1704896540
transform 1 0 -2913 0 -1 -521
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_32
timestamp 1704896540
transform 1 0 -2737 0 -1 -521
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_33
timestamp 1704896540
transform 1 0 -3689 0 -1 -521
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_34
timestamp 1704896540
transform 1 0 -3513 0 -1 -521
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_35
timestamp 1704896540
transform 1 0 -4165 0 -1 -521
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_36
timestamp 1704896540
transform 1 0 -3989 0 -1 -521
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_37
timestamp 1704896540
transform 1 0 -4941 0 -1 -521
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_38
timestamp 1704896540
transform 1 0 -4765 0 -1 -521
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_39
timestamp 1704896540
transform 1 0 -5417 0 -1 -521
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_40
timestamp 1704896540
transform 1 0 -5241 0 -1 -521
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_41
timestamp 1704896540
transform 1 0 -2261 0 -1 -521
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_42
timestamp 1704896540
transform 1 0 -2437 0 -1 -521
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_43
timestamp 1704896540
transform 1 0 -1054 0 -1 2307
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_44
timestamp 1704896540
transform 1 0 -878 0 -1 2307
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_45
timestamp 1704896540
transform 1 0 -5359 0 1 -350
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_46
timestamp 1704896540
transform 1 0 -2907 0 1 -350
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_47
timestamp 1704896540
transform 1 0 -2731 0 1 -350
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_48
timestamp 1704896540
transform 1 0 -4759 0 1 -350
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_49
timestamp 1704896540
transform 1 0 -1654 0 1 -350
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_50
timestamp 1704896540
transform 1 0 -4583 0 1 -350
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_51
timestamp 1704896540
transform 1 0 -1830 0 1 -350
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_52
timestamp 1704896540
transform 1 0 -3683 0 1 -350
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_53
timestamp 1704896540
transform 1 0 -3507 0 1 -350
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_54
timestamp 1704896540
transform 1 0 -5535 0 1 -350
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_55
timestamp 1704896540
transform 1 0 -1054 0 1 -350
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_56
timestamp 1704896540
transform 1 0 -878 0 1 -350
box 0 0 1 1
use PYL1_CDNS_52468879185123  PYL1_CDNS_52468879185123_0
timestamp 1704896540
transform -1 0 -3079 0 1 -1869
box 0 0 1 1
use PYL1_CDNS_52468879185123  PYL1_CDNS_52468879185123_1
timestamp 1704896540
transform -1 0 -4331 0 1 -1869
box 0 0 1 1
use PYL1_CDNS_52468879185123  PYL1_CDNS_52468879185123_2
timestamp 1704896540
transform -1 0 -5583 0 1 -1869
box 0 0 1 1
use PYL1_CDNS_52468879185123  PYL1_CDNS_52468879185123_3
timestamp 1704896540
transform -1 0 -5883 0 1 -1869
box 0 0 1 1
use PYL1_CDNS_52468879185123  PYL1_CDNS_52468879185123_4
timestamp 1704896540
transform -1 0 -1827 0 1 -1869
box 0 0 1 1
use PYL1_CDNS_52468879185123  PYL1_CDNS_52468879185123_5
timestamp 1704896540
transform 1 0 -2737 0 1 -1869
box 0 0 1 1
use PYL1_CDNS_52468879185123  PYL1_CDNS_52468879185123_6
timestamp 1704896540
transform 1 0 -2913 0 1 -1869
box 0 0 1 1
use PYL1_CDNS_52468879185123  PYL1_CDNS_52468879185123_7
timestamp 1704896540
transform 1 0 -3513 0 1 -1869
box 0 0 1 1
use PYL1_CDNS_52468879185123  PYL1_CDNS_52468879185123_8
timestamp 1704896540
transform 1 0 -3689 0 1 -1869
box 0 0 1 1
use PYL1_CDNS_52468879185123  PYL1_CDNS_52468879185123_9
timestamp 1704896540
transform 1 0 -3989 0 1 -1869
box 0 0 1 1
use PYL1_CDNS_52468879185123  PYL1_CDNS_52468879185123_10
timestamp 1704896540
transform 1 0 -4165 0 1 -1869
box 0 0 1 1
use PYL1_CDNS_52468879185123  PYL1_CDNS_52468879185123_11
timestamp 1704896540
transform 1 0 -4765 0 1 -1869
box 0 0 1 1
use PYL1_CDNS_52468879185123  PYL1_CDNS_52468879185123_12
timestamp 1704896540
transform 1 0 -4941 0 1 -1869
box 0 0 1 1
use PYL1_CDNS_52468879185123  PYL1_CDNS_52468879185123_13
timestamp 1704896540
transform 1 0 -5241 0 1 -1869
box 0 0 1 1
use PYL1_CDNS_52468879185123  PYL1_CDNS_52468879185123_14
timestamp 1704896540
transform 1 0 -5417 0 1 -1869
box 0 0 1 1
use PYL1_CDNS_52468879185123  PYL1_CDNS_52468879185123_15
timestamp 1704896540
transform 1 0 -2437 0 1 -1869
box 0 0 1 1
use PYL1_CDNS_52468879185123  PYL1_CDNS_52468879185123_16
timestamp 1704896540
transform 1 0 -2261 0 1 -1869
box 0 0 1 1
use sky130_fd_io__refgen_ctl_vdda_ls  sky130_fd_io__refgen_ctl_vdda_ls_0
timestamp 1704896540
transform -1 0 -9555 0 1 -6427
box -336 -32 2037 4597
use sky130_fd_io__refgen_ctl_vdda_ls  sky130_fd_io__refgen_ctl_vdda_ls_1
timestamp 1704896540
transform -1 0 -5973 0 1 -6427
box -336 -32 2037 4597
use sky130_fd_io__refgen_ctl_vdda_ls  sky130_fd_io__refgen_ctl_vdda_ls_2
timestamp 1704896540
transform -1 0 -2391 0 1 -6427
box -336 -32 2037 4597
use sky130_fd_io__refgen_ctl_vdda_ls  sky130_fd_io__refgen_ctl_vdda_ls_3
timestamp 1704896540
transform 1 0 -13047 0 1 -6427
box -336 -32 2037 4597
use sky130_fd_io__refgen_ctl_vdda_ls  sky130_fd_io__refgen_ctl_vdda_ls_4
timestamp 1704896540
transform 1 0 -9465 0 1 -6427
box -336 -32 2037 4597
use sky130_fd_io__refgen_ctl_vdda_ls  sky130_fd_io__refgen_ctl_vdda_ls_5
timestamp 1704896540
transform 1 0 -5883 0 1 -6427
box -336 -32 2037 4597
use sky130_fd_io__refgen_ctl_vdda_ls_vdda  sky130_fd_io__refgen_ctl_vdda_ls_vdda_0
timestamp 1704896540
transform -1 0 -9555 0 -1 2185
box -336 1103 2037 4597
use sky130_fd_io__refgen_ctl_vdda_ls_vdda  sky130_fd_io__refgen_ctl_vdda_ls_vdda_1
timestamp 1704896540
transform 1 0 -13047 0 -1 2185
box -336 1103 2037 4597
use sky130_fd_io__refgen_ctl_vdda_ls_vdda  sky130_fd_io__refgen_ctl_vdda_ls_vdda_2
timestamp 1704896540
transform 1 0 -9465 0 -1 2185
box -336 1103 2037 4597
<< labels >>
flabel comment s -5903 -1606 -5903 -1606 0 FreeSans 400 0 0 0 vref_sel0_vdda
flabel comment s -5903 -1478 -5903 -1478 0 FreeSans 400 0 0 0 vref_sel0_vdda_n
flabel comment s -5932 -1016 -5932 -1016 0 FreeSans 400 0 0 0 vref_sel1_vdda
flabel comment s -5951 -908 -5951 -908 0 FreeSans 400 0 0 0 vref_sel1_vdda_n
flabel comment s -5951 -559 -5951 -559 0 FreeSans 400 0 0 0 enable_vdda_h
flabel comment s -2655 -1726 -2655 -1726 0 FreeSans 400 0 0 0 sel_vdda_vref
flabel comment s -2774 -1481 -2774 -1481 0 FreeSans 400 0 0 0 sel_vdda_amuxbusa
flabel comment s -2774 -907 -2774 -907 0 FreeSans 400 0 0 0 sel_vdda_amuxbusb
flabel comment s -5927 43 -5927 43 0 FreeSans 400 0 0 0 vref_sel1_vddio_n
flabel comment s -5879 2040 -5879 2040 0 FreeSans 400 0 0 0 vref_sel0_vddio
flabel comment s -5879 1912 -5879 1912 0 FreeSans 400 0 0 0 vref_sel0_vddio_n
flabel comment s -5908 151 -5908 151 0 FreeSans 400 0 0 0 vref_sel1_vddio
flabel comment s -5927 -306 -5927 -306 0 FreeSans 400 0 0 0 enable_vswitch_h
flabel comment s -1430 2160 -1430 2160 0 FreeSans 400 0 0 0 sel_vddio_vref
flabel comment s -1549 1915 -1549 1915 0 FreeSans 400 0 0 0 sel_vddio_amuxbusa
flabel comment s -1227 42 -1227 42 0 FreeSans 400 0 0 0 sel_vddio_amuxbusb
<< properties >>
string GDS_END 80818612
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 80735712
string path 8.650 0.375 8.650 3.575 
<< end >>
