magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< pwell >>
rect 82 3520 202 3524
rect 1234 3520 1354 3524
rect 82 8 252 3520
rect 1184 8 1354 3520
rect 82 4 202 8
rect 1234 4 1354 8
<< mvndiff >>
rect 108 3494 176 3498
rect 1260 3494 1328 3498
rect 108 3482 226 3494
rect 108 3448 116 3482
rect 150 3448 184 3482
rect 218 3448 226 3482
rect 108 3436 226 3448
rect 1210 3482 1328 3494
rect 1210 3448 1218 3482
rect 1252 3448 1286 3482
rect 1320 3448 1328 3482
rect 1210 3436 1328 3448
rect 108 3432 176 3436
rect 1260 3432 1328 3436
rect 108 3368 176 3372
rect 1260 3368 1328 3372
rect 108 3356 226 3368
rect 108 3322 116 3356
rect 150 3322 184 3356
rect 218 3322 226 3356
rect 108 3310 226 3322
rect 1210 3356 1328 3368
rect 1210 3322 1218 3356
rect 1252 3322 1286 3356
rect 1320 3322 1328 3356
rect 1210 3310 1328 3322
rect 108 3306 176 3310
rect 1260 3306 1328 3310
rect 108 3242 176 3246
rect 1260 3242 1328 3246
rect 108 3230 226 3242
rect 108 3196 116 3230
rect 150 3196 184 3230
rect 218 3196 226 3230
rect 108 3184 226 3196
rect 1210 3230 1328 3242
rect 1210 3196 1218 3230
rect 1252 3196 1286 3230
rect 1320 3196 1328 3230
rect 1210 3184 1328 3196
rect 108 3180 176 3184
rect 1260 3180 1328 3184
rect 108 3116 176 3120
rect 1260 3116 1328 3120
rect 108 3104 226 3116
rect 108 3070 116 3104
rect 150 3070 184 3104
rect 218 3070 226 3104
rect 108 3058 226 3070
rect 1210 3104 1328 3116
rect 1210 3070 1218 3104
rect 1252 3070 1286 3104
rect 1320 3070 1328 3104
rect 1210 3058 1328 3070
rect 108 3054 176 3058
rect 1260 3054 1328 3058
rect 108 2990 176 2994
rect 1260 2990 1328 2994
rect 108 2978 226 2990
rect 108 2944 116 2978
rect 150 2944 184 2978
rect 218 2944 226 2978
rect 108 2932 226 2944
rect 1210 2978 1328 2990
rect 1210 2944 1218 2978
rect 1252 2944 1286 2978
rect 1320 2944 1328 2978
rect 1210 2932 1328 2944
rect 108 2928 176 2932
rect 1260 2928 1328 2932
rect 108 2864 176 2868
rect 1260 2864 1328 2868
rect 108 2852 226 2864
rect 108 2818 116 2852
rect 150 2818 184 2852
rect 218 2818 226 2852
rect 108 2806 226 2818
rect 1210 2852 1328 2864
rect 1210 2818 1218 2852
rect 1252 2818 1286 2852
rect 1320 2818 1328 2852
rect 1210 2806 1328 2818
rect 108 2802 176 2806
rect 1260 2802 1328 2806
rect 108 2738 176 2742
rect 1260 2738 1328 2742
rect 108 2726 226 2738
rect 108 2692 116 2726
rect 150 2692 184 2726
rect 218 2692 226 2726
rect 108 2680 226 2692
rect 1210 2726 1328 2738
rect 1210 2692 1218 2726
rect 1252 2692 1286 2726
rect 1320 2692 1328 2726
rect 1210 2680 1328 2692
rect 108 2676 176 2680
rect 1260 2676 1328 2680
rect 108 2612 176 2616
rect 1260 2612 1328 2616
rect 108 2600 226 2612
rect 108 2566 116 2600
rect 150 2566 184 2600
rect 218 2566 226 2600
rect 108 2554 226 2566
rect 1210 2600 1328 2612
rect 1210 2566 1218 2600
rect 1252 2566 1286 2600
rect 1320 2566 1328 2600
rect 1210 2554 1328 2566
rect 108 2550 176 2554
rect 1260 2550 1328 2554
rect 108 2486 176 2490
rect 1260 2486 1328 2490
rect 108 2474 226 2486
rect 108 2440 116 2474
rect 150 2440 184 2474
rect 218 2440 226 2474
rect 108 2428 226 2440
rect 1210 2474 1328 2486
rect 1210 2440 1218 2474
rect 1252 2440 1286 2474
rect 1320 2440 1328 2474
rect 1210 2428 1328 2440
rect 108 2424 176 2428
rect 1260 2424 1328 2428
rect 108 2360 176 2364
rect 1260 2360 1328 2364
rect 108 2348 226 2360
rect 108 2314 116 2348
rect 150 2314 184 2348
rect 218 2314 226 2348
rect 108 2302 226 2314
rect 1210 2348 1328 2360
rect 1210 2314 1218 2348
rect 1252 2314 1286 2348
rect 1320 2314 1328 2348
rect 1210 2302 1328 2314
rect 108 2298 176 2302
rect 1260 2298 1328 2302
rect 108 2234 176 2238
rect 1260 2234 1328 2238
rect 108 2222 226 2234
rect 108 2188 116 2222
rect 150 2188 184 2222
rect 218 2188 226 2222
rect 108 2176 226 2188
rect 1210 2222 1328 2234
rect 1210 2188 1218 2222
rect 1252 2188 1286 2222
rect 1320 2188 1328 2222
rect 1210 2176 1328 2188
rect 108 2172 176 2176
rect 1260 2172 1328 2176
rect 108 2108 176 2112
rect 1260 2108 1328 2112
rect 108 2096 226 2108
rect 108 2062 116 2096
rect 150 2062 184 2096
rect 218 2062 226 2096
rect 108 2050 226 2062
rect 1210 2096 1328 2108
rect 1210 2062 1218 2096
rect 1252 2062 1286 2096
rect 1320 2062 1328 2096
rect 1210 2050 1328 2062
rect 108 2046 176 2050
rect 1260 2046 1328 2050
rect 108 1982 176 1986
rect 1260 1982 1328 1986
rect 108 1970 226 1982
rect 108 1936 116 1970
rect 150 1936 184 1970
rect 218 1936 226 1970
rect 108 1924 226 1936
rect 1210 1970 1328 1982
rect 1210 1936 1218 1970
rect 1252 1936 1286 1970
rect 1320 1936 1328 1970
rect 1210 1924 1328 1936
rect 108 1920 176 1924
rect 1260 1920 1328 1924
rect 108 1856 176 1860
rect 1260 1856 1328 1860
rect 108 1844 226 1856
rect 108 1810 116 1844
rect 150 1810 184 1844
rect 218 1810 226 1844
rect 108 1798 226 1810
rect 1210 1844 1328 1856
rect 1210 1810 1218 1844
rect 1252 1810 1286 1844
rect 1320 1810 1328 1844
rect 1210 1798 1328 1810
rect 108 1794 176 1798
rect 1260 1794 1328 1798
rect 108 1730 176 1734
rect 1260 1730 1328 1734
rect 108 1718 226 1730
rect 108 1684 116 1718
rect 150 1684 184 1718
rect 218 1684 226 1718
rect 108 1672 226 1684
rect 1210 1718 1328 1730
rect 1210 1684 1218 1718
rect 1252 1684 1286 1718
rect 1320 1684 1328 1718
rect 1210 1672 1328 1684
rect 108 1668 176 1672
rect 1260 1668 1328 1672
rect 108 1604 176 1608
rect 1260 1604 1328 1608
rect 108 1592 226 1604
rect 108 1558 116 1592
rect 150 1558 184 1592
rect 218 1558 226 1592
rect 108 1546 226 1558
rect 1210 1592 1328 1604
rect 1210 1558 1218 1592
rect 1252 1558 1286 1592
rect 1320 1558 1328 1592
rect 1210 1546 1328 1558
rect 108 1542 176 1546
rect 1260 1542 1328 1546
rect 108 1478 176 1482
rect 1260 1478 1328 1482
rect 108 1466 226 1478
rect 108 1432 116 1466
rect 150 1432 184 1466
rect 218 1432 226 1466
rect 108 1420 226 1432
rect 1210 1466 1328 1478
rect 1210 1432 1218 1466
rect 1252 1432 1286 1466
rect 1320 1432 1328 1466
rect 1210 1420 1328 1432
rect 108 1416 176 1420
rect 1260 1416 1328 1420
rect 108 1352 176 1356
rect 1260 1352 1328 1356
rect 108 1340 226 1352
rect 108 1306 116 1340
rect 150 1306 184 1340
rect 218 1306 226 1340
rect 108 1294 226 1306
rect 1210 1340 1328 1352
rect 1210 1306 1218 1340
rect 1252 1306 1286 1340
rect 1320 1306 1328 1340
rect 1210 1294 1328 1306
rect 108 1290 176 1294
rect 1260 1290 1328 1294
rect 108 1226 176 1230
rect 1260 1226 1328 1230
rect 108 1214 226 1226
rect 108 1180 116 1214
rect 150 1180 184 1214
rect 218 1180 226 1214
rect 108 1168 226 1180
rect 1210 1214 1328 1226
rect 1210 1180 1218 1214
rect 1252 1180 1286 1214
rect 1320 1180 1328 1214
rect 1210 1168 1328 1180
rect 108 1164 176 1168
rect 1260 1164 1328 1168
rect 108 1100 176 1104
rect 1260 1100 1328 1104
rect 108 1088 226 1100
rect 108 1054 116 1088
rect 150 1054 184 1088
rect 218 1054 226 1088
rect 108 1042 226 1054
rect 1210 1088 1328 1100
rect 1210 1054 1218 1088
rect 1252 1054 1286 1088
rect 1320 1054 1328 1088
rect 1210 1042 1328 1054
rect 108 1038 176 1042
rect 1260 1038 1328 1042
rect 108 974 176 978
rect 1260 974 1328 978
rect 108 962 226 974
rect 108 928 116 962
rect 150 928 184 962
rect 218 928 226 962
rect 108 916 226 928
rect 1210 962 1328 974
rect 1210 928 1218 962
rect 1252 928 1286 962
rect 1320 928 1328 962
rect 1210 916 1328 928
rect 108 912 176 916
rect 1260 912 1328 916
rect 108 848 176 852
rect 1260 848 1328 852
rect 108 836 226 848
rect 108 802 116 836
rect 150 802 184 836
rect 218 802 226 836
rect 108 790 226 802
rect 1210 836 1328 848
rect 1210 802 1218 836
rect 1252 802 1286 836
rect 1320 802 1328 836
rect 1210 790 1328 802
rect 108 786 176 790
rect 1260 786 1328 790
rect 108 722 176 726
rect 1260 722 1328 726
rect 108 710 226 722
rect 108 676 116 710
rect 150 676 184 710
rect 218 676 226 710
rect 108 664 226 676
rect 1210 710 1328 722
rect 1210 676 1218 710
rect 1252 676 1286 710
rect 1320 676 1328 710
rect 1210 664 1328 676
rect 108 660 176 664
rect 1260 660 1328 664
rect 108 596 176 600
rect 1260 596 1328 600
rect 108 584 226 596
rect 108 550 116 584
rect 150 550 184 584
rect 218 550 226 584
rect 108 538 226 550
rect 1210 584 1328 596
rect 1210 550 1218 584
rect 1252 550 1286 584
rect 1320 550 1328 584
rect 1210 538 1328 550
rect 108 534 176 538
rect 1260 534 1328 538
rect 108 470 176 474
rect 1260 470 1328 474
rect 108 458 226 470
rect 108 424 116 458
rect 150 424 184 458
rect 218 424 226 458
rect 108 412 226 424
rect 1210 458 1328 470
rect 1210 424 1218 458
rect 1252 424 1286 458
rect 1320 424 1328 458
rect 1210 412 1328 424
rect 108 408 176 412
rect 1260 408 1328 412
rect 108 344 176 348
rect 1260 344 1328 348
rect 108 332 226 344
rect 108 298 116 332
rect 150 298 184 332
rect 218 298 226 332
rect 108 286 226 298
rect 1210 332 1328 344
rect 1210 298 1218 332
rect 1252 298 1286 332
rect 1320 298 1328 332
rect 1210 286 1328 298
rect 108 282 176 286
rect 1260 282 1328 286
rect 108 218 176 222
rect 1260 218 1328 222
rect 108 206 226 218
rect 108 172 116 206
rect 150 172 184 206
rect 218 172 226 206
rect 108 160 226 172
rect 1210 206 1328 218
rect 1210 172 1218 206
rect 1252 172 1286 206
rect 1320 172 1328 206
rect 1210 160 1328 172
rect 108 156 176 160
rect 1260 156 1328 160
rect 108 92 176 96
rect 1260 92 1328 96
rect 108 80 226 92
rect 108 46 116 80
rect 150 46 184 80
rect 218 46 226 80
rect 108 34 226 46
rect 1210 80 1328 92
rect 1210 46 1218 80
rect 1252 46 1286 80
rect 1320 46 1328 80
rect 1210 34 1328 46
rect 108 30 176 34
rect 1260 30 1328 34
<< ndiffc >>
rect 184 3448 218 3482
rect 1218 3448 1252 3482
rect 184 3322 218 3356
rect 1218 3322 1252 3356
rect 184 3196 218 3230
rect 1218 3196 1252 3230
rect 184 3070 218 3104
rect 1218 3070 1252 3104
rect 184 2944 218 2978
rect 1218 2944 1252 2978
rect 184 2818 218 2852
rect 1218 2818 1252 2852
rect 184 2692 218 2726
rect 1218 2692 1252 2726
rect 184 2566 218 2600
rect 1218 2566 1252 2600
rect 184 2440 218 2474
rect 1218 2440 1252 2474
rect 184 2314 218 2348
rect 1218 2314 1252 2348
rect 184 2188 218 2222
rect 1218 2188 1252 2222
rect 184 2062 218 2096
rect 1218 2062 1252 2096
rect 184 1936 218 1970
rect 1218 1936 1252 1970
rect 184 1810 218 1844
rect 1218 1810 1252 1844
rect 184 1684 218 1718
rect 1218 1684 1252 1718
rect 184 1558 218 1592
rect 1218 1558 1252 1592
rect 184 1432 218 1466
rect 1218 1432 1252 1466
rect 184 1306 218 1340
rect 1218 1306 1252 1340
rect 184 1180 218 1214
rect 1218 1180 1252 1214
rect 184 1054 218 1088
rect 1218 1054 1252 1088
rect 184 928 218 962
rect 1218 928 1252 962
rect 184 802 218 836
rect 1218 802 1252 836
rect 184 676 218 710
rect 1218 676 1252 710
rect 184 550 218 584
rect 1218 550 1252 584
rect 184 424 218 458
rect 1218 424 1252 458
rect 184 298 218 332
rect 1218 298 1252 332
rect 184 172 218 206
rect 1218 172 1252 206
rect 184 46 218 80
rect 1218 46 1252 80
<< mvndiffc >>
rect 116 3448 150 3482
rect 1286 3448 1320 3482
rect 116 3322 150 3356
rect 1286 3322 1320 3356
rect 116 3196 150 3230
rect 1286 3196 1320 3230
rect 116 3070 150 3104
rect 1286 3070 1320 3104
rect 116 2944 150 2978
rect 1286 2944 1320 2978
rect 116 2818 150 2852
rect 1286 2818 1320 2852
rect 116 2692 150 2726
rect 1286 2692 1320 2726
rect 116 2566 150 2600
rect 1286 2566 1320 2600
rect 116 2440 150 2474
rect 1286 2440 1320 2474
rect 116 2314 150 2348
rect 1286 2314 1320 2348
rect 116 2188 150 2222
rect 1286 2188 1320 2222
rect 116 2062 150 2096
rect 1286 2062 1320 2096
rect 116 1936 150 1970
rect 1286 1936 1320 1970
rect 116 1810 150 1844
rect 1286 1810 1320 1844
rect 116 1684 150 1718
rect 1286 1684 1320 1718
rect 116 1558 150 1592
rect 1286 1558 1320 1592
rect 116 1432 150 1466
rect 1286 1432 1320 1466
rect 116 1306 150 1340
rect 1286 1306 1320 1340
rect 116 1180 150 1214
rect 1286 1180 1320 1214
rect 116 1054 150 1088
rect 1286 1054 1320 1088
rect 116 928 150 962
rect 1286 928 1320 962
rect 116 802 150 836
rect 1286 802 1320 836
rect 116 676 150 710
rect 1286 676 1320 710
rect 116 550 150 584
rect 1286 550 1320 584
rect 116 424 150 458
rect 1286 424 1320 458
rect 116 298 150 332
rect 1286 298 1320 332
rect 116 172 150 206
rect 1286 172 1320 206
rect 116 46 150 80
rect 1286 46 1320 80
<< locali >>
rect 116 3482 218 3498
rect 1218 3482 1320 3498
rect 158 3448 196 3482
rect 1218 3448 1286 3482
rect 116 3432 218 3448
rect 116 3356 218 3372
rect 150 3322 218 3356
rect 116 3230 218 3322
rect 1218 3356 1320 3448
rect 1218 3322 1286 3356
rect 1218 3306 1320 3322
rect 150 3196 218 3230
rect 116 3180 218 3196
rect 1218 3230 1320 3246
rect 1218 3196 1286 3230
rect 116 3104 218 3120
rect 150 3070 218 3104
rect 116 2978 218 3070
rect 1218 3104 1320 3196
rect 1218 3070 1286 3104
rect 1218 3054 1320 3070
rect 150 2944 218 2978
rect 116 2928 218 2944
rect 1218 2978 1320 2994
rect 1218 2944 1286 2978
rect 116 2852 218 2868
rect 150 2818 218 2852
rect 116 2726 218 2818
rect 1218 2852 1320 2944
rect 1218 2818 1286 2852
rect 1218 2802 1320 2818
rect 150 2692 218 2726
rect 116 2676 218 2692
rect 1218 2726 1320 2742
rect 1218 2692 1286 2726
rect 1218 2658 1252 2692
rect 1286 2658 1320 2692
rect 1218 2620 1320 2658
rect 116 2600 218 2616
rect 150 2566 218 2600
rect 116 2474 218 2566
rect 1218 2586 1252 2620
rect 1286 2600 1320 2620
rect 1218 2566 1286 2586
rect 1218 2550 1320 2566
rect 150 2440 218 2474
rect 116 2424 218 2440
rect 1218 2474 1320 2490
rect 1218 2440 1286 2474
rect 116 2348 218 2364
rect 150 2314 218 2348
rect 116 2222 218 2314
rect 1218 2348 1320 2440
rect 1218 2314 1286 2348
rect 1218 2298 1320 2314
rect 150 2188 218 2222
rect 116 2172 218 2188
rect 1218 2222 1320 2238
rect 1218 2188 1286 2222
rect 116 2096 218 2112
rect 150 2062 218 2096
rect 116 1970 218 2062
rect 1218 2096 1320 2188
rect 1218 2062 1286 2096
rect 1218 2046 1320 2062
rect 150 1936 218 1970
rect 116 1920 218 1936
rect 1218 1970 1320 1986
rect 1218 1936 1286 1970
rect 116 1844 218 1860
rect 150 1810 218 1844
rect 116 1784 218 1810
rect 1218 1844 1320 1936
rect 1218 1810 1286 1844
rect 1218 1794 1320 1810
rect 116 1750 124 1784
rect 158 1750 196 1784
rect 116 1718 218 1750
rect 150 1684 218 1718
rect 116 1668 218 1684
rect 1218 1718 1320 1734
rect 1218 1684 1286 1718
rect 116 1592 218 1608
rect 150 1558 218 1592
rect 116 1466 218 1558
rect 1218 1592 1320 1684
rect 1218 1558 1286 1592
rect 1218 1542 1320 1558
rect 150 1432 218 1466
rect 116 1416 218 1432
rect 1218 1466 1320 1482
rect 1218 1432 1286 1466
rect 116 1340 218 1356
rect 150 1306 218 1340
rect 116 1214 218 1306
rect 1218 1340 1320 1432
rect 1218 1306 1286 1340
rect 1218 1290 1320 1306
rect 150 1180 218 1214
rect 116 1164 218 1180
rect 1218 1214 1320 1230
rect 1218 1180 1286 1214
rect 116 1088 218 1104
rect 150 1054 218 1088
rect 116 962 218 1054
rect 1218 1088 1320 1180
rect 1218 1054 1286 1088
rect 1218 1038 1320 1054
rect 150 928 218 962
rect 116 912 218 928
rect 1218 962 1320 978
rect 1218 937 1286 962
rect 1218 903 1252 937
rect 1286 903 1320 928
rect 1218 865 1320 903
rect 116 836 218 852
rect 150 802 218 836
rect 116 710 218 802
rect 1218 831 1252 865
rect 1286 836 1320 865
rect 1218 802 1286 831
rect 1218 786 1320 802
rect 150 676 218 710
rect 116 660 218 676
rect 1218 710 1320 726
rect 1218 676 1286 710
rect 116 584 218 600
rect 150 550 218 584
rect 116 458 218 550
rect 1218 584 1320 676
rect 1218 550 1286 584
rect 1218 534 1320 550
rect 150 424 218 458
rect 116 408 218 424
rect 1218 458 1320 474
rect 1218 424 1286 458
rect 116 332 218 348
rect 150 298 218 332
rect 116 206 218 298
rect 1218 332 1320 424
rect 1218 298 1286 332
rect 1218 282 1320 298
rect 150 172 218 206
rect 116 156 218 172
rect 1218 206 1320 222
rect 1218 172 1286 206
rect 116 80 218 96
rect 1218 80 1320 172
rect 158 46 196 80
rect 1218 46 1286 80
rect 116 30 218 46
rect 1218 30 1320 46
<< viali >>
rect 124 3448 150 3482
rect 150 3448 158 3482
rect 196 3448 230 3482
rect 1252 2658 1286 2692
rect 1252 2586 1286 2620
rect 124 1750 158 1784
rect 196 1750 230 1784
rect 1252 903 1286 937
rect 1252 831 1286 865
rect 124 46 150 80
rect 150 46 158 80
rect 196 46 230 80
<< metal1 >>
rect 108 3492 236 3494
rect 108 3440 114 3492
rect 166 3440 178 3492
rect 230 3440 236 3492
rect 1200 3440 1206 3492
rect 1258 3440 1270 3492
rect 1322 3440 1328 3492
rect 108 3436 236 3440
tri 1221 3436 1225 3440 ne
rect 1225 3436 1292 3440
tri 1225 3415 1246 3436 ne
rect 1246 2789 1292 3436
tri 1292 3415 1317 3440 nw
rect 1247 2787 1291 2788
rect 1247 2750 1291 2751
rect 1246 2692 1292 2749
rect 1246 2658 1252 2692
rect 1286 2658 1292 2692
rect 1246 2620 1292 2658
rect 1246 2586 1252 2620
rect 1286 2586 1292 2620
rect 1246 2538 1292 2586
rect 1247 2536 1291 2537
rect 1247 2499 1291 2500
tri 1225 1796 1246 1817 se
rect 1246 1796 1292 2498
rect 108 1792 236 1796
tri 1221 1792 1225 1796 se
rect 1225 1792 1292 1796
tri 1292 1792 1317 1817 sw
rect 108 1740 114 1792
rect 166 1740 178 1792
rect 230 1740 236 1792
rect 1200 1740 1206 1792
rect 1258 1740 1270 1792
rect 1322 1740 1328 1792
rect 108 1738 236 1740
tri 1221 1738 1223 1740 ne
rect 1223 1738 1292 1740
tri 1223 1715 1246 1738 ne
rect 1246 1530 1292 1738
tri 1292 1715 1317 1740 nw
rect 1247 1528 1291 1529
rect 1246 1492 1292 1528
rect 1247 1491 1291 1492
rect 1246 937 1292 1490
rect 1246 903 1252 937
rect 1286 903 1292 937
rect 1246 865 1292 903
rect 1246 831 1252 865
rect 1286 831 1292 865
rect 1246 780 1292 831
rect 1247 778 1291 779
rect 1246 742 1292 778
rect 1247 741 1291 742
tri 1225 92 1246 113 se
rect 1246 92 1292 740
rect 108 88 236 92
tri 1221 88 1225 92 se
rect 1225 88 1292 92
tri 1292 88 1317 113 sw
rect 108 36 114 88
rect 166 36 178 88
rect 230 36 236 88
rect 1200 36 1206 88
rect 1258 36 1270 88
rect 1322 36 1328 88
rect 108 34 236 36
<< rmetal1 >>
rect 1246 2788 1292 2789
rect 1246 2787 1247 2788
rect 1291 2787 1292 2788
rect 1246 2750 1247 2751
rect 1291 2750 1292 2751
rect 1246 2749 1292 2750
rect 1246 2537 1292 2538
rect 1246 2536 1247 2537
rect 1291 2536 1292 2537
rect 1246 2499 1247 2500
rect 1291 2499 1292 2500
rect 1246 2498 1292 2499
rect 1246 1529 1292 1530
rect 1246 1528 1247 1529
rect 1291 1528 1292 1529
rect 1246 1491 1247 1492
rect 1291 1491 1292 1492
rect 1246 1490 1292 1491
rect 1246 779 1292 780
rect 1246 778 1247 779
rect 1291 778 1292 779
rect 1246 741 1247 742
rect 1291 741 1292 742
rect 1246 740 1292 741
<< via1 >>
rect 114 3482 166 3492
rect 114 3448 124 3482
rect 124 3448 158 3482
rect 158 3448 166 3482
rect 114 3440 166 3448
rect 178 3482 230 3492
rect 178 3448 196 3482
rect 196 3448 230 3482
rect 178 3440 230 3448
rect 1206 3440 1258 3492
rect 1270 3440 1322 3492
rect 114 1784 166 1792
rect 114 1750 124 1784
rect 124 1750 158 1784
rect 158 1750 166 1784
rect 114 1740 166 1750
rect 178 1784 230 1792
rect 178 1750 196 1784
rect 196 1750 230 1784
rect 178 1740 230 1750
rect 1206 1740 1258 1792
rect 1270 1740 1322 1792
rect 114 80 166 88
rect 114 46 124 80
rect 124 46 158 80
rect 158 46 166 80
rect 114 36 166 46
rect 178 80 230 88
rect 178 46 196 80
rect 196 46 230 80
rect 178 36 230 46
rect 1206 36 1258 88
rect 1270 36 1322 88
<< metal2 >>
rect 108 3440 114 3492
rect 166 3440 178 3492
rect 230 3440 1206 3492
rect 1258 3440 1270 3492
rect 1322 3440 1328 3492
rect 108 1740 114 1792
rect 166 1740 178 1792
rect 230 1740 1206 1792
rect 1258 1740 1270 1792
rect 1322 1740 1328 1792
rect 108 36 114 88
rect 166 36 178 88
rect 230 36 1206 88
rect 1258 36 1270 88
rect 1322 36 1328 88
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_0
timestamp 1704896540
transform -1 0 226 0 1 3310
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_1
timestamp 1704896540
transform -1 0 226 0 1 3184
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_2
timestamp 1704896540
transform -1 0 226 0 1 3058
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_3
timestamp 1704896540
transform -1 0 226 0 1 2932
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_4
timestamp 1704896540
transform -1 0 226 0 1 2806
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_5
timestamp 1704896540
transform -1 0 226 0 1 2680
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_6
timestamp 1704896540
transform -1 0 226 0 1 1672
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_7
timestamp 1704896540
transform -1 0 226 0 1 1546
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_8
timestamp 1704896540
transform -1 0 226 0 1 1420
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_9
timestamp 1704896540
transform -1 0 226 0 1 1294
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_10
timestamp 1704896540
transform -1 0 226 0 1 1168
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_11
timestamp 1704896540
transform -1 0 226 0 1 1042
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_12
timestamp 1704896540
transform -1 0 226 0 1 916
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_13
timestamp 1704896540
transform -1 0 226 0 1 3436
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_14
timestamp 1704896540
transform -1 0 226 0 -1 1856
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_15
timestamp 1704896540
transform -1 0 226 0 -1 1982
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_16
timestamp 1704896540
transform -1 0 226 0 -1 2108
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_17
timestamp 1704896540
transform -1 0 226 0 -1 2234
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_18
timestamp 1704896540
transform -1 0 226 0 -1 2360
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_19
timestamp 1704896540
transform -1 0 226 0 -1 2486
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_20
timestamp 1704896540
transform -1 0 226 0 -1 2612
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_21
timestamp 1704896540
transform -1 0 226 0 -1 92
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_22
timestamp 1704896540
transform -1 0 226 0 -1 218
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_23
timestamp 1704896540
transform -1 0 226 0 -1 344
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_24
timestamp 1704896540
transform -1 0 226 0 -1 470
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_25
timestamp 1704896540
transform -1 0 226 0 -1 596
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_26
timestamp 1704896540
transform -1 0 226 0 -1 722
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_27
timestamp 1704896540
transform -1 0 226 0 -1 848
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_28
timestamp 1704896540
transform 1 0 1210 0 -1 1856
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_29
timestamp 1704896540
transform 1 0 1210 0 -1 1982
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_30
timestamp 1704896540
transform 1 0 1210 0 -1 2108
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_31
timestamp 1704896540
transform 1 0 1210 0 -1 2234
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_32
timestamp 1704896540
transform 1 0 1210 0 -1 2360
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_33
timestamp 1704896540
transform 1 0 1210 0 -1 2486
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_34
timestamp 1704896540
transform 1 0 1210 0 -1 2612
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_35
timestamp 1704896540
transform 1 0 1210 0 -1 92
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_36
timestamp 1704896540
transform 1 0 1210 0 -1 218
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_37
timestamp 1704896540
transform 1 0 1210 0 -1 344
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_38
timestamp 1704896540
transform 1 0 1210 0 -1 470
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_39
timestamp 1704896540
transform 1 0 1210 0 -1 596
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_40
timestamp 1704896540
transform 1 0 1210 0 -1 722
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_41
timestamp 1704896540
transform 1 0 1210 0 -1 848
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_42
timestamp 1704896540
transform 1 0 1210 0 1 3436
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_43
timestamp 1704896540
transform 1 0 1210 0 1 3310
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_44
timestamp 1704896540
transform 1 0 1210 0 1 3184
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_45
timestamp 1704896540
transform 1 0 1210 0 1 3058
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_46
timestamp 1704896540
transform 1 0 1210 0 1 2932
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_47
timestamp 1704896540
transform 1 0 1210 0 1 2806
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_48
timestamp 1704896540
transform 1 0 1210 0 1 2680
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_49
timestamp 1704896540
transform 1 0 1210 0 1 1672
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_50
timestamp 1704896540
transform 1 0 1210 0 1 1546
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_51
timestamp 1704896540
transform 1 0 1210 0 1 1420
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_52
timestamp 1704896540
transform 1 0 1210 0 1 1294
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_53
timestamp 1704896540
transform 1 0 1210 0 1 1168
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_54
timestamp 1704896540
transform 1 0 1210 0 1 1042
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_55
timestamp 1704896540
transform 1 0 1210 0 1 916
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_0
timestamp 1704896540
transform 0 1 124 -1 0 1784
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_1
timestamp 1704896540
transform 0 1 124 -1 0 80
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_2
timestamp 1704896540
transform 0 1 124 1 0 3448
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1704896540
transform 0 -1 1286 1 0 2586
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1704896540
transform 0 -1 1286 1 0 831
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1704896540
transform 1 0 108 0 -1 1792
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_1
timestamp 1704896540
transform 1 0 1200 0 -1 1792
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_2
timestamp 1704896540
transform 1 0 108 0 -1 88
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_3
timestamp 1704896540
transform 1 0 1200 0 -1 88
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_4
timestamp 1704896540
transform 1 0 1200 0 1 3440
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_5
timestamp 1704896540
transform 1 0 108 0 1 3440
box 0 0 1 1
use nDFres_CDNS_524688791851622  nDFres_CDNS_524688791851622_0
timestamp 1704896540
transform -1 0 1218 0 1 2802
box -68 -26 1068 92
use nDFres_CDNS_524688791851622  nDFres_CDNS_524688791851622_1
timestamp 1704896540
transform -1 0 1218 0 1 1038
box -68 -26 1068 92
use nDFres_CDNS_524688791851622  nDFres_CDNS_524688791851622_2
timestamp 1704896540
transform -1 0 1218 0 1 3054
box -68 -26 1068 92
use nDFres_CDNS_524688791851622  nDFres_CDNS_524688791851622_3
timestamp 1704896540
transform -1 0 1218 0 1 1290
box -68 -26 1068 92
use nDFres_CDNS_524688791851622  nDFres_CDNS_524688791851622_4
timestamp 1704896540
transform -1 0 1218 0 1 3306
box -68 -26 1068 92
use nDFres_CDNS_524688791851622  nDFres_CDNS_524688791851622_5
timestamp 1704896540
transform -1 0 1218 0 1 1542
box -68 -26 1068 92
use nDFres_CDNS_524688791851622  nDFres_CDNS_524688791851622_6
timestamp 1704896540
transform -1 0 1218 0 -1 2490
box -68 -26 1068 92
use nDFres_CDNS_524688791851622  nDFres_CDNS_524688791851622_7
timestamp 1704896540
transform -1 0 1218 0 -1 726
box -68 -26 1068 92
use nDFres_CDNS_524688791851622  nDFres_CDNS_524688791851622_8
timestamp 1704896540
transform -1 0 1218 0 -1 2238
box -68 -26 1068 92
use nDFres_CDNS_524688791851622  nDFres_CDNS_524688791851622_9
timestamp 1704896540
transform -1 0 1218 0 -1 474
box -68 -26 1068 92
use nDFres_CDNS_524688791851622  nDFres_CDNS_524688791851622_10
timestamp 1704896540
transform -1 0 1218 0 -1 1986
box -68 -26 1068 92
use nDFres_CDNS_524688791851622  nDFres_CDNS_524688791851622_11
timestamp 1704896540
transform -1 0 1218 0 -1 222
box -68 -26 1068 92
use nDFres_CDNS_524688791851622  nDFres_CDNS_524688791851622_12
timestamp 1704896540
transform 1 0 218 0 -1 2616
box -68 -26 1068 92
use nDFres_CDNS_524688791851622  nDFres_CDNS_524688791851622_13
timestamp 1704896540
transform 1 0 218 0 -1 852
box -68 -26 1068 92
use nDFres_CDNS_524688791851622  nDFres_CDNS_524688791851622_14
timestamp 1704896540
transform 1 0 218 0 -1 2364
box -68 -26 1068 92
use nDFres_CDNS_524688791851622  nDFres_CDNS_524688791851622_15
timestamp 1704896540
transform 1 0 218 0 -1 600
box -68 -26 1068 92
use nDFres_CDNS_524688791851622  nDFres_CDNS_524688791851622_16
timestamp 1704896540
transform 1 0 218 0 -1 2112
box -68 -26 1068 92
use nDFres_CDNS_524688791851622  nDFres_CDNS_524688791851622_17
timestamp 1704896540
transform 1 0 218 0 -1 348
box -68 -26 1068 92
use nDFres_CDNS_524688791851622  nDFres_CDNS_524688791851622_18
timestamp 1704896540
transform 1 0 218 0 -1 1860
box -68 -26 1068 92
use nDFres_CDNS_524688791851622  nDFres_CDNS_524688791851622_19
timestamp 1704896540
transform 1 0 218 0 -1 96
box -68 -26 1068 92
use nDFres_CDNS_524688791851622  nDFres_CDNS_524688791851622_20
timestamp 1704896540
transform 1 0 218 0 1 2676
box -68 -26 1068 92
use nDFres_CDNS_524688791851622  nDFres_CDNS_524688791851622_21
timestamp 1704896540
transform 1 0 218 0 1 912
box -68 -26 1068 92
use nDFres_CDNS_524688791851622  nDFres_CDNS_524688791851622_22
timestamp 1704896540
transform 1 0 218 0 1 2928
box -68 -26 1068 92
use nDFres_CDNS_524688791851622  nDFres_CDNS_524688791851622_23
timestamp 1704896540
transform 1 0 218 0 1 1164
box -68 -26 1068 92
use nDFres_CDNS_524688791851622  nDFres_CDNS_524688791851622_24
timestamp 1704896540
transform 1 0 218 0 1 3180
box -68 -26 1068 92
use nDFres_CDNS_524688791851622  nDFres_CDNS_524688791851622_25
timestamp 1704896540
transform 1 0 218 0 1 1416
box -68 -26 1068 92
use nDFres_CDNS_524688791851622  nDFres_CDNS_524688791851622_26
timestamp 1704896540
transform 1 0 218 0 1 3432
box -68 -26 1068 92
use nDFres_CDNS_524688791851622  nDFres_CDNS_524688791851622_27
timestamp 1704896540
transform 1 0 218 0 1 1668
box -68 -26 1068 92
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851293  sky130_fd_io__sio_tk_em1o_CDNS_524688791851293_0
timestamp 1704896540
transform 0 1 1246 -1 0 2590
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851293  sky130_fd_io__sio_tk_em1o_CDNS_524688791851293_1
timestamp 1704896540
transform 0 -1 1292 1 0 2697
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851295  sky130_fd_io__sio_tk_em1s_CDNS_524688791851295_0
timestamp 1704896540
transform 0 1 1246 -1 0 832
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851295  sky130_fd_io__sio_tk_em1s_CDNS_524688791851295_1
timestamp 1704896540
transform 0 -1 1292 1 0 1438
box 0 0 1 1
<< labels >>
flabel metal1 s 108 34 236 92 3 FreeSans 600 0 0 0 r2
port 2 nsew
flabel metal1 s 108 3436 236 3494 3 FreeSans 600 0 0 0 r1
port 1 nsew
<< properties >>
string GDS_END 96461006
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 96448168
<< end >>
