magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< pwell >>
rect -26 -26 176 626
<< scnmos >>
rect 60 0 90 600
<< ndiff >>
rect 0 317 60 600
rect 0 283 8 317
rect 42 283 60 317
rect 0 0 60 283
rect 90 317 150 600
rect 90 283 108 317
rect 142 283 150 317
rect 90 0 150 283
<< ndiffc >>
rect 8 283 42 317
rect 108 283 142 317
<< poly >>
rect 60 600 90 626
rect 60 -26 90 0
<< locali >>
rect 8 317 42 333
rect 8 267 42 283
rect 108 317 142 333
rect 108 267 142 283
use contact_17  contact_17_0
timestamp 1704896540
transform 1 0 100 0 1 267
box 0 0 1 1
use contact_17  contact_17_1
timestamp 1704896540
transform 1 0 0 0 1 267
box 0 0 1 1
<< labels >>
rlabel locali s 125 300 125 300 4 D
port 1 nsew
rlabel locali s 25 300 25 300 4 S
port 2 nsew
rlabel poly s 75 300 75 300 4 G
port 3 nsew
<< properties >>
string FIXED_BBOX -25 -26 175 626
string GDS_END 33512
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 32760
<< end >>
