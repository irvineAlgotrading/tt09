magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 1 21 879 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 331 47 361 177
rect 519 47 549 177
rect 603 47 633 177
rect 687 47 717 177
rect 771 47 801 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 331 297 361 497
rect 519 297 549 497
rect 603 297 633 497
rect 687 297 717 497
rect 771 297 801 497
<< ndiff >>
rect 27 131 79 177
rect 27 97 35 131
rect 69 97 79 131
rect 27 47 79 97
rect 109 97 163 177
rect 109 63 119 97
rect 153 63 163 97
rect 109 47 163 63
rect 193 131 247 177
rect 193 97 203 131
rect 237 97 247 131
rect 193 47 247 97
rect 277 169 331 177
rect 277 135 287 169
rect 321 135 331 169
rect 277 47 331 135
rect 361 101 413 177
rect 361 67 371 101
rect 405 67 413 101
rect 361 47 413 67
rect 467 101 519 177
rect 467 67 475 101
rect 509 67 519 101
rect 467 47 519 67
rect 549 169 603 177
rect 549 135 559 169
rect 593 135 603 169
rect 549 47 603 135
rect 633 131 687 177
rect 633 97 643 131
rect 677 97 687 131
rect 633 47 687 97
rect 717 97 771 177
rect 717 63 727 97
rect 761 63 771 97
rect 717 47 771 63
rect 801 131 853 177
rect 801 97 811 131
rect 845 97 853 131
rect 801 47 853 97
<< pdiff >>
rect 27 445 79 497
rect 27 411 35 445
rect 69 411 79 445
rect 27 377 79 411
rect 27 343 35 377
rect 69 343 79 377
rect 27 297 79 343
rect 109 485 163 497
rect 109 451 119 485
rect 153 451 163 485
rect 109 417 163 451
rect 109 383 119 417
rect 153 383 163 417
rect 109 297 163 383
rect 193 417 247 497
rect 193 383 203 417
rect 237 383 247 417
rect 193 349 247 383
rect 193 315 203 349
rect 237 315 247 349
rect 193 297 247 315
rect 277 485 331 497
rect 277 451 287 485
rect 321 451 331 485
rect 277 417 331 451
rect 277 383 287 417
rect 321 383 331 417
rect 277 297 331 383
rect 361 417 413 497
rect 361 383 371 417
rect 405 383 413 417
rect 361 349 413 383
rect 361 315 371 349
rect 405 315 413 349
rect 361 297 413 315
rect 467 485 519 497
rect 467 451 475 485
rect 509 451 519 485
rect 467 417 519 451
rect 467 383 475 417
rect 509 383 519 417
rect 467 349 519 383
rect 467 315 475 349
rect 509 315 519 349
rect 467 297 519 315
rect 549 485 603 497
rect 549 451 559 485
rect 593 451 603 485
rect 549 417 603 451
rect 549 383 559 417
rect 593 383 603 417
rect 549 297 603 383
rect 633 485 687 497
rect 633 451 643 485
rect 677 451 687 485
rect 633 417 687 451
rect 633 383 643 417
rect 677 383 687 417
rect 633 349 687 383
rect 633 315 643 349
rect 677 315 687 349
rect 633 297 687 315
rect 717 485 771 497
rect 717 451 727 485
rect 761 451 771 485
rect 717 417 771 451
rect 717 383 727 417
rect 761 383 771 417
rect 717 297 771 383
rect 801 485 853 497
rect 801 451 811 485
rect 845 451 853 485
rect 801 417 853 451
rect 801 383 811 417
rect 845 383 853 417
rect 801 349 853 383
rect 801 315 811 349
rect 845 315 853 349
rect 801 297 853 315
<< ndiffc >>
rect 35 97 69 131
rect 119 63 153 97
rect 203 97 237 131
rect 287 135 321 169
rect 371 67 405 101
rect 475 67 509 101
rect 559 135 593 169
rect 643 97 677 131
rect 727 63 761 97
rect 811 97 845 131
<< pdiffc >>
rect 35 411 69 445
rect 35 343 69 377
rect 119 451 153 485
rect 119 383 153 417
rect 203 383 237 417
rect 203 315 237 349
rect 287 451 321 485
rect 287 383 321 417
rect 371 383 405 417
rect 371 315 405 349
rect 475 451 509 485
rect 475 383 509 417
rect 475 315 509 349
rect 559 451 593 485
rect 559 383 593 417
rect 643 451 677 485
rect 643 383 677 417
rect 643 315 677 349
rect 727 451 761 485
rect 727 383 761 417
rect 811 451 845 485
rect 811 383 845 417
rect 811 315 845 349
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 331 497 361 523
rect 519 497 549 523
rect 603 497 633 523
rect 687 497 717 523
rect 771 497 801 523
rect 79 265 109 297
rect 163 265 193 297
rect 55 249 193 265
rect 55 215 65 249
rect 99 215 193 249
rect 55 199 193 215
rect 79 177 109 199
rect 163 177 193 199
rect 247 265 277 297
rect 331 265 361 297
rect 519 265 549 297
rect 603 265 633 297
rect 247 249 361 265
rect 247 215 263 249
rect 297 215 361 249
rect 247 199 361 215
rect 495 249 633 265
rect 495 215 505 249
rect 539 215 633 249
rect 495 199 633 215
rect 247 177 277 199
rect 331 177 361 199
rect 519 177 549 199
rect 603 177 633 199
rect 687 265 717 297
rect 771 265 801 297
rect 687 249 801 265
rect 687 215 703 249
rect 737 215 801 249
rect 687 199 801 215
rect 687 177 717 199
rect 771 177 801 199
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 331 21 361 47
rect 519 21 549 47
rect 603 21 633 47
rect 687 21 717 47
rect 771 21 801 47
<< polycont >>
rect 65 215 99 249
rect 263 215 297 249
rect 505 215 539 249
rect 703 215 737 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 19 445 69 493
rect 19 411 35 445
rect 19 377 69 411
rect 19 343 35 377
rect 103 485 525 493
rect 103 451 119 485
rect 153 459 287 485
rect 103 417 153 451
rect 321 459 475 485
rect 103 383 119 417
rect 103 365 153 383
rect 187 417 253 425
rect 187 383 203 417
rect 237 383 253 417
rect 19 331 69 343
rect 187 349 253 383
rect 287 417 321 451
rect 509 451 525 485
rect 287 365 321 383
rect 355 417 432 425
rect 355 383 371 417
rect 405 383 432 417
rect 187 331 203 349
rect 19 315 203 331
rect 237 331 253 349
rect 355 349 432 383
rect 355 331 371 349
rect 237 315 371 331
rect 405 315 432 349
rect 19 297 432 315
rect 475 417 525 451
rect 509 383 525 417
rect 475 349 525 383
rect 559 485 593 527
rect 559 417 593 451
rect 559 365 593 383
rect 627 485 693 493
rect 627 451 643 485
rect 677 451 693 485
rect 627 417 693 451
rect 627 383 643 417
rect 677 383 693 417
rect 509 331 525 349
rect 627 349 693 383
rect 727 485 761 527
rect 727 417 761 451
rect 727 365 761 383
rect 795 485 861 493
rect 795 451 811 485
rect 845 451 861 485
rect 795 417 861 451
rect 795 383 811 417
rect 845 383 861 417
rect 627 331 643 349
rect 509 315 643 331
rect 677 331 693 349
rect 795 349 861 383
rect 795 331 811 349
rect 677 315 811 331
rect 845 315 861 349
rect 475 297 861 315
rect 30 249 156 255
rect 30 215 65 249
rect 99 215 156 249
rect 214 249 340 255
rect 214 215 263 249
rect 297 215 340 249
rect 19 136 237 170
rect 374 169 432 297
rect 489 249 620 255
rect 489 215 505 249
rect 539 215 620 249
rect 678 249 900 255
rect 678 215 703 249
rect 737 215 900 249
rect 19 131 69 136
rect 19 97 35 131
rect 203 131 237 136
rect 271 135 287 169
rect 321 135 559 169
rect 593 135 609 169
rect 643 136 875 170
rect 19 51 69 97
rect 103 97 169 102
rect 103 63 119 97
rect 153 63 169 97
rect 103 17 169 63
rect 643 131 677 136
rect 237 97 371 101
rect 203 67 371 97
rect 405 67 421 101
rect 203 51 421 67
rect 459 67 475 101
rect 509 97 643 101
rect 811 131 875 136
rect 509 67 677 97
rect 459 51 677 67
rect 711 97 777 102
rect 711 63 727 97
rect 761 63 777 97
rect 711 17 777 63
rect 845 97 875 131
rect 811 51 875 97
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
flabel locali s 494 221 528 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 586 221 620 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 678 221 712 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 770 221 804 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 306 221 340 255 0 FreeSans 200 0 0 0 B1
port 3 nsew signal input
flabel locali s 122 221 156 255 0 FreeSans 200 0 0 0 B2
port 4 nsew signal input
flabel locali s 398 153 432 187 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 398 221 432 255 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 398 357 432 391 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 398 289 432 323 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 122 527 156 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel locali s 122 -17 156 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 B2
port 4 nsew signal input
flabel locali s 214 221 248 255 0 FreeSans 200 0 0 0 B1
port 3 nsew signal input
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 a22oi_2
rlabel metal1 s 0 -48 920 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 920 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 920 544
string GDS_END 4051862
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 4043376
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 13.600 23.000 13.600 
<< end >>
