magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -119 -66 1719 1466
<< mvpmos >>
rect 0 0 1600 1400
<< mvpdiff >>
rect -50 0 0 1400
rect 1600 0 1650 1400
<< poly >>
rect 0 1400 1600 1426
rect 0 -26 1600 0
<< locali >>
rect -45 -4 -11 1354
rect 1611 -4 1645 1354
use DFL1sd_CDNS_52468879185620  DFL1sd_CDNS_52468879185620_0
timestamp 1704896540
transform 1 0 1600 0 1 0
box -36 -36 89 1436
use hvDFL1sd_CDNS_5246887918573  hvDFL1sd_CDNS_5246887918573_0
timestamp 1704896540
transform -1 0 0 0 1 0
box -36 -36 89 1436
<< labels >>
flabel comment s -28 675 -28 675 0 FreeSans 300 0 0 0 S
flabel comment s 1628 675 1628 675 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 96468948
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 96467932
<< end >>
