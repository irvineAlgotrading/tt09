magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< dnwell >>
rect 4927 3772 308245 36105
<< nwell >>
rect 303230 39610 311106 39640
rect 0 31750 311106 39610
rect 0 7206 7829 31750
rect 303230 7206 311106 31750
rect 0 0 311106 7206
rect 303230 -3184 311106 -3154
rect 0 -42794 311106 -3184
<< pwell >>
rect 11759 17686 13156 19032
<< psubdiff >>
rect 11785 18533 13130 19006
rect 11785 18499 12218 18533
rect 12252 18499 13130 18533
rect 11785 17712 13130 18499
<< nsubdiff >>
rect 1592 2125 2937 2598
rect 1592 2091 2025 2125
rect 2059 2091 2937 2125
rect 1592 1304 2937 2091
rect 1592 -40669 2937 -40196
rect 1592 -40703 2025 -40669
rect 2059 -40703 2937 -40669
rect 1592 -41490 2937 -40703
<< psubdiffcont >>
rect 12218 18499 12252 18533
<< nsubdiffcont >>
rect 2025 2091 2059 2125
rect 2025 -40703 2059 -40669
<< locali >>
rect 12028 18533 12590 18733
rect 12028 18499 12218 18533
rect 12252 18499 12590 18533
rect 12028 18138 12590 18499
rect 1835 2125 2397 2325
rect 1835 2091 2025 2125
rect 2059 2091 2397 2125
rect 1835 1730 2397 2091
rect 1835 -40669 2397 -40469
rect 1835 -40703 2025 -40669
rect 2059 -40703 2397 -40669
rect 1835 -41064 2397 -40703
<< metal1 >>
rect 16968 20613 19467 20671
rect 16968 20239 17042 20613
rect 14436 20181 17042 20239
rect 14436 20157 14510 20181
rect 13652 20097 14510 20157
rect 13652 19853 19553 19913
rect 16941 -24022 17447 -23964
rect 16941 -24371 17010 -24022
rect 15875 -24429 17010 -24371
rect 15875 -24631 15944 -24429
rect 14089 -24689 15944 -24631
rect 14089 -24803 14158 -24689
rect 13326 -24861 14158 -24803
rect 13326 -25191 17491 -25131
<< metal2 >>
rect 17166 20562 17858 20575
rect 17166 20506 17177 20562
rect 17233 20531 17858 20562
rect 17233 20506 17777 20531
rect 17166 20475 17777 20506
rect 17833 20475 17858 20531
rect 17166 20430 17858 20475
rect 13652 20056 15260 20062
rect 13652 20000 15189 20056
rect 15245 20000 15260 20056
rect 13652 19993 15260 20000
rect 17061 -24190 17408 -24062
rect 17061 -24486 17170 -24190
rect 16068 -24614 17170 -24486
rect 14225 -24775 15017 -24733
rect 14225 -24831 14913 -24775
rect 14969 -24831 15017 -24775
rect 14225 -24861 15017 -24831
rect 16068 -24775 16177 -24614
rect 16068 -24831 16098 -24775
rect 16154 -24831 16177 -24775
rect 14225 -24918 14298 -24861
rect 16068 -24862 16177 -24831
rect 13327 -25046 14298 -24918
<< via2 >>
rect 17177 20506 17233 20562
rect 17777 20475 17833 20531
rect 15189 20000 15245 20056
rect 14913 -24831 14969 -24775
rect 16098 -24831 16154 -24775
<< metal3 >>
rect 17166 20562 17244 20575
rect 17166 20506 17177 20562
rect 17233 20506 17244 20562
rect 17166 20137 17244 20506
rect 17756 20531 19477 20575
rect 17756 20475 17777 20531
rect 17833 20475 19477 20531
rect 17756 20415 19477 20475
rect 15179 20056 17244 20137
rect 15179 20000 15189 20056
rect 15245 20000 17244 20056
rect 15179 19993 17244 20000
rect 14892 -24775 16177 -24733
rect 14892 -24831 14913 -24775
rect 14969 -24831 16098 -24775
rect 16154 -24831 16177 -24775
rect 14892 -24862 16177 -24831
use sky130_fd_pr__rf_nfet_01v8_lvt_aF02W0p42L0p15  sky130_fd_pr__rf_nfet_01v8_lvt_aF02W0p42L0p15_0
timestamp 1704896540
transform 1 0 13768 0 1 19942
box 10 -89 290 217
use sky130_fd_pr__rf_nfet_01v8_lvt_aF02W0p84L0p15  sky130_fd_pr__rf_nfet_01v8_lvt_aF02W0p84L0p15_0
timestamp 1704896540
transform 1 0 14792 0 1 19942
box 10 -89 290 301
use sky130_fd_pr__rf_nfet_01v8_lvt_aF02W3p00L0p15  sky130_fd_pr__rf_nfet_01v8_lvt_aF02W3p00L0p15_0
timestamp 1704896540
transform 1 0 17280 0 1 19942
box 10 -89 290 733
use sky130_fd_pr__rf_nfet_01v8_lvt_aF04W0p84L0p15  sky130_fd_pr__rf_nfet_01v8_lvt_aF04W0p84L0p15_0
timestamp 1704896540
transform 1 0 15336 0 1 19942
box 10 -89 462 301
use sky130_fd_pr__rf_nfet_01v8_lvt_aF04W3p00L0p15  sky130_fd_pr__rf_nfet_01v8_lvt_aF04W3p00L0p15_0
timestamp 1704896540
transform 1 0 17978 0 1 19942
box 10 -89 462 733
use sky130_fd_pr__rf_nfet_01v8_lvt_aF08W0p84L0p15  sky130_fd_pr__rf_nfet_01v8_lvt_aF08W0p84L0p15_0
timestamp 1704896540
transform 1 0 15979 0 1 19942
box 10 -89 806 301
use sky130_fd_pr__rf_nfet_01v8_lvt_aF08W3p00L0p15  sky130_fd_pr__rf_nfet_01v8_lvt_aF08W3p00L0p15_0
timestamp 1704896540
transform 1 0 18778 0 1 19942
box 10 -89 806 733
use sky130_fd_pr__rf_pfet_01v8_aF02W0p84L0p15  sky130_fd_pr__rf_pfet_01v8_aF02W0p84L0p15_0
timestamp 1704896540
transform 1 0 13567 0 1 -25102
box 0 -89 300 303
use sky130_fd_pr__rf_pfet_01v8_aF02W1p68L0p15  sky130_fd_pr__rf_pfet_01v8_aF02W1p68L0p15_0
timestamp 1704896540
transform 1 0 14343 0 1 -25102
box 0 -89 294 475
use sky130_fd_pr__rf_pfet_01v8_aF02W3p00L0p15  sky130_fd_pr__rf_pfet_01v8_aF02W3p00L0p15_0
timestamp 1704896540
transform 1 0 16352 0 1 -25102
box 0 -89 294 735
use sky130_fd_pr__rf_pfet_01v8_aF02W5p00L0p15  sky130_fd_pr__rf_pfet_01v8_aF02W5p00L0p15_0
timestamp 1704896540
transform 1 0 17235 0 1 -25094
box 0 -97 294 1134
use sky130_fd_pr__rf_pfet_01v8_aF04W1p68L0p15  sky130_fd_pr__rf_pfet_01v8_aF04W1p68L0p15_0
timestamp 1704896540
transform 1 0 15125 0 1 -25102
box 0 -89 466 471
<< labels >>
flabel comment s 9976 31045 9976 31045 0 FreeSans 1600 0 0 0 condiode
flabel locali s 12401 18220 12529 18665 0 FreeSans 54 0 0 0 VGND
port 2 nsew
flabel locali s 2191 1808 2304 2253 0 FreeSans 54 0 0 0 NWELL
port 3 nsew
flabel locali s 2209 -40991 2318 -40518 0 FreeSans 54 0 0 0 B_P
port 4 nsew
flabel metal2 s 13652 19993 13673 20062 0 FreeSans 400 0 0 0 VPWR
port 5 nsew
flabel metal2 s 13327 -25046 13331 -24918 0 FreeSans 400 0 0 0 D_P
port 6 nsew
flabel metal1 s 13652 19853 13658 19913 0 FreeSans 400 0 0 0 S
port 7 nsew
flabel metal1 s 13326 -24861 13328 -24803 0 FreeSans 400 0 0 0 G_P
port 8 nsew
flabel metal1 s 13326 -25191 13330 -25131 0 FreeSans 400 0 0 0 S_P
port 9 nsew
flabel metal1 s 13652 20097 13674 20157 0 FreeSans 400 0 0 0 G
port 10 nsew
<< properties >>
string GDS_END 10521924
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 10516786
<< end >>
