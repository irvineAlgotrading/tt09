magic
tech sky130A
magscale 1 2
timestamp 1704896540
use sky130_fd_pr__hvdfl1sd__example_55959141808370  sky130_fd_pr__hvdfl1sd__example_55959141808370_0
timestamp 1704896540
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808370  sky130_fd_pr__hvdfl1sd__example_55959141808370_1
timestamp 1704896540
transform 1 0 120 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 16742572
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 16741518
<< end >>
