magic
tech sky130A
timestamp 1704896540
<< metal1 >>
rect 0 0 3 58
rect 381 0 384 58
<< via1 >>
rect 3 0 381 58
<< metal2 >>
rect 0 0 3 58
rect 381 0 384 58
<< properties >>
string GDS_END 94174968
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 94173300
<< end >>
