magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect 22 2201 6234 2367
rect 22 1127 188 2201
rect 2940 1139 3204 1140
rect 4650 1139 5597 1140
rect 6068 1139 6234 2201
rect 1214 973 6234 1139
rect 4650 972 5163 973
<< pwell >>
rect -124 496 128 1067
rect 42 231 128 496
rect 5708 231 5794 905
rect 42 145 5794 231
<< psubdiff >>
rect -98 1017 102 1041
rect -98 983 68 1017
rect -98 945 102 983
rect -98 911 68 945
rect -98 873 102 911
rect -98 839 68 873
rect -98 801 102 839
rect -98 767 68 801
rect -98 729 102 767
rect -98 695 68 729
rect -98 658 102 695
rect -98 624 68 658
rect -98 587 102 624
rect -98 553 68 587
rect -98 522 102 553
rect 68 516 102 522
rect 68 445 102 482
rect 68 374 102 411
rect 68 303 102 340
rect 68 205 102 269
rect 5734 855 5768 879
rect 5734 781 5768 821
rect 5734 707 5768 747
rect 5734 633 5768 673
rect 5734 559 5768 599
rect 5734 485 5768 525
rect 5734 411 5768 451
rect 5734 337 5768 377
rect 5734 205 5768 303
rect 68 171 92 205
rect 126 171 161 205
rect 195 171 230 205
rect 264 171 299 205
rect 333 171 368 205
rect 402 171 437 205
rect 471 171 506 205
rect 540 171 575 205
rect 609 171 644 205
rect 678 171 713 205
rect 747 171 782 205
rect 816 171 851 205
rect 885 171 920 205
rect 954 171 989 205
rect 1023 171 1058 205
rect 1092 171 1127 205
rect 1161 171 1196 205
rect 1230 171 1265 205
rect 1299 171 1334 205
rect 1368 171 1403 205
rect 1437 171 1472 205
rect 1506 171 1541 205
rect 1575 171 1610 205
rect 1644 171 1679 205
rect 1713 171 1748 205
rect 1782 171 1817 205
rect 1851 171 1886 205
rect 1920 171 1955 205
rect 1989 171 2024 205
rect 2058 171 2093 205
rect 2127 171 2162 205
rect 2196 171 2231 205
rect 2265 171 2300 205
rect 2334 171 2369 205
rect 2403 171 2438 205
rect 2472 171 2507 205
rect 2541 171 2576 205
rect 2610 171 2645 205
rect 2679 171 2714 205
rect 2748 171 2783 205
rect 2817 171 2852 205
rect 2886 171 2921 205
rect 2955 171 2990 205
rect 3024 171 3058 205
rect 3092 171 3126 205
rect 3160 171 3194 205
rect 3228 171 3262 205
rect 3296 171 3330 205
rect 3364 171 3398 205
rect 3432 171 3466 205
rect 3500 171 3534 205
rect 3568 171 3602 205
rect 3636 171 3670 205
rect 3704 171 3738 205
rect 3772 171 3806 205
rect 3840 171 3874 205
rect 3908 171 3942 205
rect 3976 171 4010 205
rect 4044 171 4078 205
rect 4112 171 4146 205
rect 4180 171 4214 205
rect 4248 171 4282 205
rect 4316 171 4350 205
rect 4384 171 4418 205
rect 4452 171 4486 205
rect 4520 171 4554 205
rect 4588 171 4622 205
rect 4656 171 4690 205
rect 4724 171 4758 205
rect 4792 171 4826 205
rect 4860 171 4894 205
rect 4928 171 4962 205
rect 4996 171 5030 205
rect 5064 171 5098 205
rect 5132 171 5166 205
rect 5200 171 5234 205
rect 5268 171 5302 205
rect 5336 171 5370 205
rect 5404 171 5438 205
rect 5472 171 5506 205
rect 5540 171 5574 205
rect 5608 171 5642 205
rect 5676 171 5710 205
rect 5744 171 5768 205
<< mvnsubdiff >>
rect 88 2267 112 2301
rect 146 2267 181 2301
rect 215 2267 250 2301
rect 284 2267 319 2301
rect 353 2267 388 2301
rect 422 2267 457 2301
rect 491 2267 526 2301
rect 560 2267 595 2301
rect 629 2267 664 2301
rect 698 2267 733 2301
rect 767 2267 802 2301
rect 836 2267 871 2301
rect 905 2267 940 2301
rect 974 2267 1009 2301
rect 1043 2267 1078 2301
rect 1112 2267 1146 2301
rect 1180 2267 1214 2301
rect 1248 2267 1282 2301
rect 1316 2267 1350 2301
rect 1384 2267 1418 2301
rect 1452 2267 1486 2301
rect 1520 2267 1554 2301
rect 1588 2267 1622 2301
rect 1656 2267 1690 2301
rect 1724 2267 1758 2301
rect 1792 2267 1826 2301
rect 1860 2267 1894 2301
rect 1928 2267 1962 2301
rect 1996 2267 2030 2301
rect 2064 2267 2098 2301
rect 2132 2267 2166 2301
rect 2200 2267 2234 2301
rect 2268 2267 2302 2301
rect 2336 2267 2370 2301
rect 2404 2267 2438 2301
rect 2472 2267 2506 2301
rect 2540 2267 2574 2301
rect 2608 2267 2642 2301
rect 2676 2267 2710 2301
rect 2744 2267 2778 2301
rect 2812 2267 2846 2301
rect 2880 2267 2914 2301
rect 2948 2267 2982 2301
rect 3016 2267 3050 2301
rect 3084 2267 3118 2301
rect 3152 2267 3186 2301
rect 3220 2267 3254 2301
rect 3288 2267 3322 2301
rect 3356 2267 3390 2301
rect 3424 2267 3458 2301
rect 3492 2267 3526 2301
rect 3560 2267 3594 2301
rect 3628 2267 3662 2301
rect 3696 2267 3730 2301
rect 3764 2267 3798 2301
rect 3832 2267 3866 2301
rect 3900 2267 3934 2301
rect 3968 2267 4002 2301
rect 4036 2267 4070 2301
rect 4104 2267 4138 2301
rect 4172 2267 4206 2301
rect 4240 2267 4274 2301
rect 4308 2267 4342 2301
rect 4376 2267 4410 2301
rect 4444 2267 4478 2301
rect 4512 2267 4546 2301
rect 4580 2267 4614 2301
rect 4648 2267 4682 2301
rect 4716 2267 4750 2301
rect 4784 2267 4818 2301
rect 4852 2267 4886 2301
rect 4920 2267 4954 2301
rect 4988 2267 5022 2301
rect 5056 2267 5090 2301
rect 5124 2267 5158 2301
rect 5192 2267 5226 2301
rect 5260 2267 5294 2301
rect 5328 2267 5362 2301
rect 5396 2267 5430 2301
rect 5464 2267 5498 2301
rect 5532 2267 5566 2301
rect 5600 2267 5634 2301
rect 5668 2267 5702 2301
rect 5736 2267 5770 2301
rect 5804 2267 5838 2301
rect 5872 2267 5906 2301
rect 5940 2267 5974 2301
rect 6008 2267 6042 2301
rect 6076 2277 6168 2301
rect 6076 2267 6134 2277
rect 88 2191 122 2267
rect 88 2118 122 2157
rect 88 2045 122 2084
rect 88 1972 122 2011
rect 88 1899 122 1938
rect 88 1827 122 1865
rect 88 1755 122 1793
rect 88 1683 122 1721
rect 88 1611 122 1649
rect 88 1539 122 1577
rect 88 1467 122 1505
rect 88 1395 122 1433
rect 88 1323 122 1361
rect 88 1251 122 1289
rect 88 1193 122 1217
rect 6134 2208 6168 2243
rect 6134 2139 6168 2174
rect 6134 2070 6168 2105
rect 6134 2001 6168 2036
rect 6134 1932 6168 1967
rect 6134 1863 6168 1898
rect 6134 1795 6168 1829
rect 6134 1727 6168 1761
rect 6134 1659 6168 1693
rect 6134 1591 6168 1625
rect 6134 1523 6168 1557
rect 6134 1455 6168 1489
rect 6134 1387 6168 1421
rect 6134 1319 6168 1353
rect 6134 1251 6168 1285
rect 1280 1039 1304 1073
rect 1338 1039 1373 1073
rect 1407 1039 1442 1073
rect 1476 1039 1511 1073
rect 1545 1039 1580 1073
rect 1614 1039 1649 1073
rect 1683 1039 1718 1073
rect 1752 1039 1787 1073
rect 1821 1039 1856 1073
rect 1890 1039 1925 1073
rect 1959 1039 1994 1073
rect 2028 1039 2063 1073
rect 2097 1039 2132 1073
rect 2166 1039 2201 1073
rect 2235 1039 2270 1073
rect 2304 1039 2339 1073
rect 2373 1039 2408 1073
rect 2442 1039 2477 1073
rect 2511 1039 2546 1073
rect 2580 1039 2615 1073
rect 2649 1039 2683 1073
rect 2717 1039 2751 1073
rect 2785 1039 2819 1073
rect 2853 1039 2877 1073
rect 3270 1039 3294 1073
rect 3328 1039 3363 1073
rect 3397 1039 3432 1073
rect 3466 1039 3501 1073
rect 3535 1039 3570 1073
rect 3604 1039 3639 1073
rect 3673 1039 3708 1073
rect 3742 1039 3777 1073
rect 3811 1039 3846 1073
rect 3880 1039 3914 1073
rect 3948 1039 3982 1073
rect 4016 1039 4050 1073
rect 4084 1039 4118 1073
rect 4152 1039 4186 1073
rect 4220 1039 4254 1073
rect 4288 1039 4322 1073
rect 4356 1039 4390 1073
rect 4424 1039 4458 1073
rect 4492 1039 4526 1073
rect 4560 1039 4584 1073
rect 6134 1073 6168 1217
rect 5663 1039 5687 1073
rect 5721 1039 5758 1073
rect 5792 1039 5829 1073
rect 5863 1039 5900 1073
rect 5934 1039 5970 1073
rect 6004 1039 6040 1073
rect 6074 1039 6110 1073
rect 6144 1039 6168 1073
<< psubdiffcont >>
rect 68 983 102 1017
rect 68 911 102 945
rect 68 839 102 873
rect 68 767 102 801
rect 68 695 102 729
rect 68 624 102 658
rect 68 553 102 587
rect 68 482 102 516
rect 68 411 102 445
rect 68 340 102 374
rect 68 269 102 303
rect 5734 821 5768 855
rect 5734 747 5768 781
rect 5734 673 5768 707
rect 5734 599 5768 633
rect 5734 525 5768 559
rect 5734 451 5768 485
rect 5734 377 5768 411
rect 5734 303 5768 337
rect 92 171 126 205
rect 161 171 195 205
rect 230 171 264 205
rect 299 171 333 205
rect 368 171 402 205
rect 437 171 471 205
rect 506 171 540 205
rect 575 171 609 205
rect 644 171 678 205
rect 713 171 747 205
rect 782 171 816 205
rect 851 171 885 205
rect 920 171 954 205
rect 989 171 1023 205
rect 1058 171 1092 205
rect 1127 171 1161 205
rect 1196 171 1230 205
rect 1265 171 1299 205
rect 1334 171 1368 205
rect 1403 171 1437 205
rect 1472 171 1506 205
rect 1541 171 1575 205
rect 1610 171 1644 205
rect 1679 171 1713 205
rect 1748 171 1782 205
rect 1817 171 1851 205
rect 1886 171 1920 205
rect 1955 171 1989 205
rect 2024 171 2058 205
rect 2093 171 2127 205
rect 2162 171 2196 205
rect 2231 171 2265 205
rect 2300 171 2334 205
rect 2369 171 2403 205
rect 2438 171 2472 205
rect 2507 171 2541 205
rect 2576 171 2610 205
rect 2645 171 2679 205
rect 2714 171 2748 205
rect 2783 171 2817 205
rect 2852 171 2886 205
rect 2921 171 2955 205
rect 2990 171 3024 205
rect 3058 171 3092 205
rect 3126 171 3160 205
rect 3194 171 3228 205
rect 3262 171 3296 205
rect 3330 171 3364 205
rect 3398 171 3432 205
rect 3466 171 3500 205
rect 3534 171 3568 205
rect 3602 171 3636 205
rect 3670 171 3704 205
rect 3738 171 3772 205
rect 3806 171 3840 205
rect 3874 171 3908 205
rect 3942 171 3976 205
rect 4010 171 4044 205
rect 4078 171 4112 205
rect 4146 171 4180 205
rect 4214 171 4248 205
rect 4282 171 4316 205
rect 4350 171 4384 205
rect 4418 171 4452 205
rect 4486 171 4520 205
rect 4554 171 4588 205
rect 4622 171 4656 205
rect 4690 171 4724 205
rect 4758 171 4792 205
rect 4826 171 4860 205
rect 4894 171 4928 205
rect 4962 171 4996 205
rect 5030 171 5064 205
rect 5098 171 5132 205
rect 5166 171 5200 205
rect 5234 171 5268 205
rect 5302 171 5336 205
rect 5370 171 5404 205
rect 5438 171 5472 205
rect 5506 171 5540 205
rect 5574 171 5608 205
rect 5642 171 5676 205
rect 5710 171 5744 205
<< mvnsubdiffcont >>
rect 112 2267 146 2301
rect 181 2267 215 2301
rect 250 2267 284 2301
rect 319 2267 353 2301
rect 388 2267 422 2301
rect 457 2267 491 2301
rect 526 2267 560 2301
rect 595 2267 629 2301
rect 664 2267 698 2301
rect 733 2267 767 2301
rect 802 2267 836 2301
rect 871 2267 905 2301
rect 940 2267 974 2301
rect 1009 2267 1043 2301
rect 1078 2267 1112 2301
rect 1146 2267 1180 2301
rect 1214 2267 1248 2301
rect 1282 2267 1316 2301
rect 1350 2267 1384 2301
rect 1418 2267 1452 2301
rect 1486 2267 1520 2301
rect 1554 2267 1588 2301
rect 1622 2267 1656 2301
rect 1690 2267 1724 2301
rect 1758 2267 1792 2301
rect 1826 2267 1860 2301
rect 1894 2267 1928 2301
rect 1962 2267 1996 2301
rect 2030 2267 2064 2301
rect 2098 2267 2132 2301
rect 2166 2267 2200 2301
rect 2234 2267 2268 2301
rect 2302 2267 2336 2301
rect 2370 2267 2404 2301
rect 2438 2267 2472 2301
rect 2506 2267 2540 2301
rect 2574 2267 2608 2301
rect 2642 2267 2676 2301
rect 2710 2267 2744 2301
rect 2778 2267 2812 2301
rect 2846 2267 2880 2301
rect 2914 2267 2948 2301
rect 2982 2267 3016 2301
rect 3050 2267 3084 2301
rect 3118 2267 3152 2301
rect 3186 2267 3220 2301
rect 3254 2267 3288 2301
rect 3322 2267 3356 2301
rect 3390 2267 3424 2301
rect 3458 2267 3492 2301
rect 3526 2267 3560 2301
rect 3594 2267 3628 2301
rect 3662 2267 3696 2301
rect 3730 2267 3764 2301
rect 3798 2267 3832 2301
rect 3866 2267 3900 2301
rect 3934 2267 3968 2301
rect 4002 2267 4036 2301
rect 4070 2267 4104 2301
rect 4138 2267 4172 2301
rect 4206 2267 4240 2301
rect 4274 2267 4308 2301
rect 4342 2267 4376 2301
rect 4410 2267 4444 2301
rect 4478 2267 4512 2301
rect 4546 2267 4580 2301
rect 4614 2267 4648 2301
rect 4682 2267 4716 2301
rect 4750 2267 4784 2301
rect 4818 2267 4852 2301
rect 4886 2267 4920 2301
rect 4954 2267 4988 2301
rect 5022 2267 5056 2301
rect 5090 2267 5124 2301
rect 5158 2267 5192 2301
rect 5226 2267 5260 2301
rect 5294 2267 5328 2301
rect 5362 2267 5396 2301
rect 5430 2267 5464 2301
rect 5498 2267 5532 2301
rect 5566 2267 5600 2301
rect 5634 2267 5668 2301
rect 5702 2267 5736 2301
rect 5770 2267 5804 2301
rect 5838 2267 5872 2301
rect 5906 2267 5940 2301
rect 5974 2267 6008 2301
rect 6042 2267 6076 2301
rect 88 2157 122 2191
rect 88 2084 122 2118
rect 88 2011 122 2045
rect 88 1938 122 1972
rect 88 1865 122 1899
rect 88 1793 122 1827
rect 88 1721 122 1755
rect 88 1649 122 1683
rect 88 1577 122 1611
rect 88 1505 122 1539
rect 88 1433 122 1467
rect 88 1361 122 1395
rect 88 1289 122 1323
rect 88 1217 122 1251
rect 6134 2243 6168 2277
rect 6134 2174 6168 2208
rect 6134 2105 6168 2139
rect 6134 2036 6168 2070
rect 6134 1967 6168 2001
rect 6134 1898 6168 1932
rect 6134 1829 6168 1863
rect 6134 1761 6168 1795
rect 6134 1693 6168 1727
rect 6134 1625 6168 1659
rect 6134 1557 6168 1591
rect 6134 1489 6168 1523
rect 6134 1421 6168 1455
rect 6134 1353 6168 1387
rect 6134 1285 6168 1319
rect 6134 1217 6168 1251
rect 1304 1039 1338 1073
rect 1373 1039 1407 1073
rect 1442 1039 1476 1073
rect 1511 1039 1545 1073
rect 1580 1039 1614 1073
rect 1649 1039 1683 1073
rect 1718 1039 1752 1073
rect 1787 1039 1821 1073
rect 1856 1039 1890 1073
rect 1925 1039 1959 1073
rect 1994 1039 2028 1073
rect 2063 1039 2097 1073
rect 2132 1039 2166 1073
rect 2201 1039 2235 1073
rect 2270 1039 2304 1073
rect 2339 1039 2373 1073
rect 2408 1039 2442 1073
rect 2477 1039 2511 1073
rect 2546 1039 2580 1073
rect 2615 1039 2649 1073
rect 2683 1039 2717 1073
rect 2751 1039 2785 1073
rect 2819 1039 2853 1073
rect 3294 1039 3328 1073
rect 3363 1039 3397 1073
rect 3432 1039 3466 1073
rect 3501 1039 3535 1073
rect 3570 1039 3604 1073
rect 3639 1039 3673 1073
rect 3708 1039 3742 1073
rect 3777 1039 3811 1073
rect 3846 1039 3880 1073
rect 3914 1039 3948 1073
rect 3982 1039 4016 1073
rect 4050 1039 4084 1073
rect 4118 1039 4152 1073
rect 4186 1039 4220 1073
rect 4254 1039 4288 1073
rect 4322 1039 4356 1073
rect 4390 1039 4424 1073
rect 4458 1039 4492 1073
rect 4526 1039 4560 1073
rect 5687 1039 5721 1073
rect 5758 1039 5792 1073
rect 5829 1039 5863 1073
rect 5900 1039 5934 1073
rect 5970 1039 6004 1073
rect 6040 1039 6074 1073
rect 6110 1039 6144 1073
<< poly >>
rect 249 1145 349 1167
rect 249 1111 296 1145
rect 330 1111 349 1145
rect 249 1077 349 1111
rect 249 1043 296 1077
rect 330 1043 349 1077
rect 249 905 349 1043
rect 405 1142 505 1167
rect 405 1108 436 1142
rect 470 1108 505 1142
rect 405 1074 505 1108
rect 405 1040 436 1074
rect 470 1040 505 1074
rect 405 1006 505 1040
rect 405 972 436 1006
rect 470 972 505 1006
rect 405 905 505 972
rect 691 1129 791 1167
rect 691 1095 720 1129
rect 754 1095 791 1129
rect 691 1061 791 1095
rect 691 1027 720 1061
rect 754 1027 791 1061
rect 691 905 791 1027
rect 867 1129 947 1167
rect 867 1095 890 1129
rect 924 1095 947 1129
rect 867 1061 947 1095
rect 867 1027 890 1061
rect 924 1027 947 1061
rect 1003 1145 1103 1170
rect 1003 1111 1036 1145
rect 1070 1111 1103 1145
rect 1003 1077 1103 1111
rect 1003 1043 1036 1077
rect 1070 1043 1103 1077
rect 1003 1027 1103 1043
rect 1159 1145 1259 1167
rect 1159 1111 1175 1145
rect 1209 1111 1259 1145
rect 1159 1077 1259 1111
rect 1425 1095 2305 1167
rect 2361 1095 3241 1167
rect 3297 1095 4773 1167
rect 4815 1095 5385 1167
rect 1159 1043 1175 1077
rect 1209 1043 1259 1077
rect 1159 1027 1259 1043
rect 2899 1057 3241 1095
rect 867 985 947 1027
rect 2899 1023 2919 1057
rect 2953 1023 2987 1057
rect 3021 1023 3055 1057
rect 3089 1023 3123 1057
rect 3157 1023 3191 1057
rect 3225 1023 3241 1057
rect 4607 1053 4773 1095
rect 867 905 1515 985
rect 2899 977 3241 1023
rect 1681 961 1977 977
rect 1681 927 1717 961
rect 1751 927 1785 961
rect 1819 927 1853 961
rect 1887 927 1921 961
rect 1955 927 1977 961
rect 1681 905 1977 927
rect 2033 961 2329 977
rect 2033 927 2064 961
rect 2098 927 2132 961
rect 2166 927 2200 961
rect 2234 927 2268 961
rect 2302 927 2329 961
rect 2033 905 2329 927
rect 2495 905 3495 977
rect 3551 905 4551 977
rect 4607 905 4903 1053
rect 4959 1019 5385 1095
rect 5439 1095 6007 1167
rect 5439 1077 5641 1095
rect 5439 1043 5455 1077
rect 5489 1043 5523 1077
rect 5557 1043 5591 1077
rect 5625 1043 5641 1077
rect 4959 905 5255 1019
rect 5439 977 5641 1043
rect 5311 961 5641 977
rect 5311 927 5338 961
rect 5372 927 5406 961
rect 5440 927 5474 961
rect 5508 927 5542 961
rect 5576 927 5641 961
rect 5311 905 5641 927
<< polycont >>
rect 296 1111 330 1145
rect 296 1043 330 1077
rect 436 1108 470 1142
rect 436 1040 470 1074
rect 436 972 470 1006
rect 720 1095 754 1129
rect 720 1027 754 1061
rect 890 1095 924 1129
rect 890 1027 924 1061
rect 1036 1111 1070 1145
rect 1036 1043 1070 1077
rect 1175 1111 1209 1145
rect 1175 1043 1209 1077
rect 2919 1023 2953 1057
rect 2987 1023 3021 1057
rect 3055 1023 3089 1057
rect 3123 1023 3157 1057
rect 3191 1023 3225 1057
rect 1717 927 1751 961
rect 1785 927 1819 961
rect 1853 927 1887 961
rect 1921 927 1955 961
rect 2064 927 2098 961
rect 2132 927 2166 961
rect 2200 927 2234 961
rect 2268 927 2302 961
rect 5455 1043 5489 1077
rect 5523 1043 5557 1077
rect 5591 1043 5625 1077
rect 5338 927 5372 961
rect 5406 927 5440 961
rect 5474 927 5508 961
rect 5542 927 5576 961
<< locali >>
rect 88 2267 112 2301
rect 146 2267 181 2301
rect 215 2267 250 2301
rect 284 2267 319 2301
rect 353 2267 388 2301
rect 422 2267 457 2301
rect 491 2267 526 2301
rect 560 2267 595 2301
rect 629 2267 664 2301
rect 698 2267 733 2301
rect 767 2267 802 2301
rect 836 2267 871 2301
rect 905 2267 940 2301
rect 974 2267 1009 2301
rect 1043 2267 1078 2301
rect 1112 2267 1146 2301
rect 1180 2267 1214 2301
rect 1248 2267 1282 2301
rect 1316 2267 1350 2301
rect 1384 2267 1418 2301
rect 1452 2267 1486 2301
rect 1520 2267 1554 2301
rect 1588 2267 1622 2301
rect 1656 2267 1690 2301
rect 1724 2267 1758 2301
rect 1792 2267 1826 2301
rect 1860 2267 1894 2301
rect 1928 2267 1962 2301
rect 1996 2267 2030 2301
rect 2064 2267 2098 2301
rect 2132 2267 2166 2301
rect 2200 2267 2234 2301
rect 2268 2267 2302 2301
rect 2336 2267 2370 2301
rect 2404 2267 2438 2301
rect 2472 2267 2506 2301
rect 2540 2267 2574 2301
rect 2608 2267 2642 2301
rect 2676 2267 2710 2301
rect 2744 2267 2778 2301
rect 2812 2267 2846 2301
rect 2880 2267 2914 2301
rect 2948 2267 2982 2301
rect 3016 2267 3050 2301
rect 3084 2267 3118 2301
rect 3152 2267 3186 2301
rect 3220 2267 3254 2301
rect 3288 2267 3322 2301
rect 3356 2267 3390 2301
rect 3424 2267 3458 2301
rect 3492 2267 3526 2301
rect 3560 2267 3594 2301
rect 3628 2267 3662 2301
rect 3696 2267 3730 2301
rect 3764 2267 3798 2301
rect 3832 2267 3866 2301
rect 3900 2267 3934 2301
rect 3968 2267 4002 2301
rect 4036 2267 4070 2301
rect 4104 2267 4138 2301
rect 4172 2267 4206 2301
rect 4240 2267 4274 2301
rect 88 2191 122 2267
rect 88 2118 122 2157
rect 88 2045 122 2084
rect 88 1972 122 2011
rect 88 1899 122 1938
rect 88 1827 122 1840
rect 88 1755 122 1768
rect 88 1683 122 1696
rect 88 1611 122 1649
rect 88 1539 122 1577
rect 88 1467 122 1505
rect 88 1395 122 1433
rect 88 1323 122 1361
rect 88 1251 122 1289
rect 88 1193 122 1217
rect -98 1017 102 1041
rect -98 983 68 1017
rect -98 945 102 983
rect -98 911 68 945
rect -98 873 102 911
rect -98 839 68 873
rect -98 801 102 839
rect -98 767 68 801
rect -98 729 102 767
rect -98 695 68 729
rect -98 658 102 695
rect -98 624 68 658
rect -98 587 102 624
rect -98 553 68 587
rect -98 522 102 553
rect 68 516 102 522
rect 68 445 102 482
rect 68 381 102 411
rect 68 309 102 340
rect 184 993 238 2197
rect 360 2169 394 2267
rect 360 1802 394 1840
rect 360 1730 394 1768
rect 516 1228 570 2197
rect 498 1194 536 1228
rect 296 1145 330 1161
rect 436 1154 470 1158
rect 410 1142 448 1154
rect 410 1120 436 1142
rect 296 1077 330 1111
rect 296 1027 330 1043
rect 436 1074 470 1108
rect 436 1006 470 1040
rect 184 972 436 993
rect 184 933 470 972
rect 184 275 238 933
rect 360 309 394 347
rect 516 275 570 1194
rect 622 1213 680 2197
rect 802 2150 836 2267
rect 1114 2150 1148 2267
rect 1380 2194 1414 2267
rect 1692 2194 1726 2267
rect 2004 2190 2038 2267
rect 2316 2190 2350 2267
rect 2628 2190 2662 2267
rect 2940 2183 2974 2267
rect 3252 2183 3286 2267
rect 3604 2183 3638 2267
rect 3956 2183 3990 2267
rect 4308 2181 4342 2301
rect 4376 2267 4410 2301
rect 4444 2267 4478 2301
rect 4512 2267 4546 2301
rect 4580 2267 4614 2301
rect 4648 2267 4682 2301
rect 4716 2267 4750 2301
rect 4784 2267 4818 2301
rect 4852 2267 4886 2301
rect 4920 2267 4954 2301
rect 4988 2267 5022 2301
rect 5056 2267 5090 2301
rect 5124 2267 5158 2301
rect 5192 2267 5226 2301
rect 5260 2267 5294 2301
rect 5328 2267 5362 2301
rect 5396 2267 5430 2301
rect 5464 2267 5498 2301
rect 5532 2267 5566 2301
rect 5600 2267 5634 2301
rect 5668 2267 5702 2301
rect 5736 2267 5770 2301
rect 5804 2267 5838 2301
rect 5872 2267 5906 2301
rect 5940 2267 5974 2301
rect 6008 2267 6042 2301
rect 6076 2277 6168 2301
rect 6076 2267 6134 2277
rect 4660 2166 4694 2267
rect 6134 2208 6168 2243
rect 6134 2139 6168 2174
rect 6134 2070 6168 2105
rect 6134 2001 6168 2036
rect 6134 1932 6168 1967
rect 6134 1874 6168 1898
rect 802 1802 836 1840
rect 802 1730 836 1768
rect 1114 1802 1148 1840
rect 1114 1730 1148 1768
rect 1380 1802 1414 1840
rect 1380 1730 1414 1768
rect 1692 1802 1726 1840
rect 1692 1730 1726 1768
rect 2004 1802 2038 1840
rect 2004 1730 2038 1768
rect 2316 1802 2350 1840
rect 2316 1730 2350 1768
rect 2628 1802 2662 1840
rect 2628 1730 2662 1768
rect 2940 1802 2974 1840
rect 2940 1730 2974 1768
rect 3252 1802 3286 1840
rect 3252 1730 3286 1768
rect 3604 1802 3638 1840
rect 3604 1730 3638 1768
rect 3956 1802 3990 1840
rect 3956 1730 3990 1768
rect 4308 1802 4342 1840
rect 4308 1730 4342 1768
rect 4660 1802 4694 1840
rect 4660 1730 4694 1768
rect 6134 1802 6168 1829
rect 6134 1730 6168 1761
rect 6134 1659 6168 1693
rect 2470 1613 2508 1647
rect 2782 1613 2820 1647
rect 3058 1613 3096 1647
rect 3424 1616 3462 1650
rect 3776 1616 3814 1650
rect 4128 1616 4166 1650
rect 4480 1616 4518 1650
rect 4922 1616 4960 1650
rect 5234 1616 5272 1650
rect 6134 1591 6168 1625
rect 5550 1533 5588 1567
rect 5862 1533 5900 1567
rect 6134 1523 6168 1557
rect 1532 1456 1570 1490
rect 1848 1456 1886 1490
rect 2160 1453 2198 1487
rect 4804 1456 4842 1490
rect 5078 1456 5116 1490
rect 5390 1456 5428 1490
rect 5703 1456 5741 1490
rect 5980 1456 6018 1490
rect 6134 1455 6168 1489
rect 958 1358 996 1392
rect 1232 1358 1270 1392
rect 6134 1387 6168 1421
rect 6134 1319 6168 1353
rect 6134 1251 6168 1285
rect 622 1179 1070 1213
rect 622 913 680 1179
rect 1036 1145 1070 1179
rect 720 1129 754 1145
rect 720 1061 754 1095
rect 720 1011 754 1027
rect 890 1073 924 1095
rect 1036 1077 1070 1111
rect 1036 1027 1070 1039
rect 1175 1145 1209 1161
rect 1175 1077 1209 1111
rect 1270 1145 1304 1247
rect 1270 1108 1467 1145
rect 1280 1039 1304 1073
rect 1338 1039 1373 1073
rect 1407 1039 1442 1073
rect 1476 1039 1511 1073
rect 1545 1039 1580 1073
rect 1614 1039 1649 1073
rect 1683 1039 1718 1073
rect 1752 1039 1787 1073
rect 1821 1039 1856 1073
rect 1890 1039 1925 1073
rect 1959 1039 1994 1073
rect 2028 1039 2063 1073
rect 2097 1039 2132 1073
rect 2166 1039 2201 1073
rect 2235 1039 2270 1073
rect 2304 1039 2339 1073
rect 2373 1039 2408 1073
rect 2442 1039 2477 1073
rect 2511 1039 2546 1073
rect 2580 1039 2615 1073
rect 2649 1039 2683 1073
rect 2717 1039 2751 1073
rect 2785 1039 2819 1073
rect 2853 1039 2877 1073
rect 2919 1057 3225 1145
rect 1175 1027 1209 1039
rect 890 948 924 1027
rect 2953 1023 2987 1057
rect 3021 1023 3055 1057
rect 3089 1023 3123 1057
rect 3157 1023 3191 1057
rect 3270 1039 3294 1073
rect 3328 1039 3363 1073
rect 3397 1039 3432 1073
rect 3466 1039 3501 1073
rect 3535 1039 3570 1073
rect 3604 1039 3639 1073
rect 3673 1039 3708 1073
rect 3742 1039 3777 1073
rect 3811 1039 3846 1073
rect 3880 1039 3914 1073
rect 3948 1039 3982 1073
rect 4016 1039 4050 1073
rect 4084 1039 4118 1073
rect 4152 1039 4186 1073
rect 4220 1039 4254 1073
rect 4288 1039 4322 1073
rect 4356 1039 4390 1073
rect 4424 1039 4458 1073
rect 4492 1039 4526 1073
rect 4560 1039 4584 1073
rect 4618 1029 4759 1111
rect 1701 954 1705 988
rect 1739 961 1777 988
rect 1811 961 1849 988
rect 1883 961 1921 988
rect 1751 954 1777 961
rect 1819 954 1849 961
rect 1701 927 1717 954
rect 1751 927 1785 954
rect 1819 927 1853 954
rect 1887 927 1921 961
rect 1955 927 1971 988
rect 2048 927 2064 961
rect 2098 927 2132 961
rect 2166 927 2200 961
rect 2234 927 2268 961
rect 2302 927 2318 961
rect 2919 944 3225 1023
rect 4970 961 5240 1145
rect 5455 1077 5625 1145
rect 5947 1111 5997 1145
rect 5489 1043 5523 1077
rect 5557 1043 5591 1077
rect 6134 1073 6168 1217
rect 5455 961 5625 1043
rect 5663 1062 5687 1073
rect 5721 1062 5758 1073
rect 5792 1062 5829 1073
rect 5863 1062 5900 1073
rect 5934 1062 5970 1073
rect 5721 1039 5735 1062
rect 5792 1039 5807 1062
rect 5863 1039 5879 1062
rect 5934 1039 5951 1062
rect 6004 1039 6040 1073
rect 6074 1039 6110 1073
rect 6144 1039 6168 1073
rect 5697 1028 5735 1039
rect 5769 1028 5807 1039
rect 5841 1028 5879 1039
rect 5913 1028 5951 1039
rect 4970 927 4978 961
rect 5012 927 5050 961
rect 5084 927 5122 961
rect 5156 927 5194 961
rect 5228 927 5240 961
rect 5322 927 5338 961
rect 5372 927 5406 961
rect 5440 927 5474 961
rect 5508 927 5542 961
rect 5576 927 5625 961
rect 2048 913 2318 927
rect 656 879 694 913
rect 2048 879 2052 913
rect 2086 879 2124 913
rect 2158 879 2196 913
rect 2230 879 2268 913
rect 2302 879 2318 913
rect 622 275 680 879
rect 5734 855 5768 879
rect 2166 799 2204 833
rect 3682 765 3720 799
rect 4033 765 4071 799
rect 4386 765 4424 799
rect 5734 781 5768 821
rect 4738 691 4776 725
rect 5090 691 5128 725
rect 5442 691 5480 725
rect 5734 707 5768 747
rect 5734 633 5768 673
rect 1032 527 1070 561
rect 1312 527 1350 561
rect 1809 527 1847 561
rect 5734 559 5768 599
rect 1670 453 1708 487
rect 1988 453 2026 487
rect 2302 453 2340 487
rect 2626 453 2664 487
rect 2977 453 3015 487
rect 3330 453 3368 487
rect 5734 485 5768 525
rect 5734 411 5768 451
rect 822 309 856 347
rect 1174 309 1208 347
rect 1526 309 1560 347
rect 2450 309 2484 347
rect 2802 309 2836 347
rect 3154 309 3188 347
rect 3506 309 3540 347
rect 3858 309 3892 347
rect 4210 309 4244 347
rect 4562 309 4596 347
rect 4914 309 4948 347
rect 5266 309 5300 347
rect 5618 309 5652 347
rect 5734 337 5768 347
rect 68 205 102 269
rect 5734 205 5768 275
rect 68 171 92 205
rect 126 171 161 205
rect 195 171 230 205
rect 264 171 299 205
rect 333 171 368 205
rect 402 171 437 205
rect 471 171 506 205
rect 540 171 575 205
rect 609 171 644 205
rect 678 171 713 205
rect 747 171 782 205
rect 816 171 851 205
rect 885 171 920 205
rect 954 171 989 205
rect 1023 171 1058 205
rect 1092 171 1127 205
rect 1161 171 1196 205
rect 1230 171 1265 205
rect 1299 171 1334 205
rect 1368 171 1403 205
rect 1437 171 1472 205
rect 1506 171 1541 205
rect 1575 171 1610 205
rect 1644 171 1679 205
rect 1713 171 1748 205
rect 1782 171 1817 205
rect 1851 171 1886 205
rect 1920 171 1955 205
rect 1989 171 2024 205
rect 2058 171 2093 205
rect 2127 171 2162 205
rect 2196 171 2231 205
rect 2265 171 2300 205
rect 2334 171 2369 205
rect 2403 171 2438 205
rect 2472 171 2507 205
rect 2541 171 2576 205
rect 2610 171 2645 205
rect 2679 171 2714 205
rect 2748 171 2783 205
rect 2817 171 2852 205
rect 2886 171 2921 205
rect 2955 171 2990 205
rect 3024 171 3058 205
rect 3092 171 3126 205
rect 3160 171 3194 205
rect 3228 171 3262 205
rect 3296 171 3330 205
rect 3364 171 3398 205
rect 3432 171 3466 205
rect 3500 171 3534 205
rect 3568 171 3602 205
rect 3636 171 3670 205
rect 3704 171 3738 205
rect 3772 171 3806 205
rect 3840 171 3874 205
rect 3908 171 3942 205
rect 3976 171 4010 205
rect 4044 171 4078 205
rect 4112 171 4146 205
rect 4180 171 4214 205
rect 4248 171 4282 205
rect 4316 171 4350 205
rect 4384 171 4418 205
rect 4452 171 4486 205
rect 4520 171 4554 205
rect 4588 171 4622 205
rect 4656 171 4690 205
rect 4724 171 4758 205
rect 4792 171 4826 205
rect 4860 171 4894 205
rect 4928 171 4962 205
rect 4996 171 5030 205
rect 5064 171 5098 205
rect 5132 171 5166 205
rect 5200 171 5234 205
rect 5268 171 5302 205
rect 5336 171 5370 205
rect 5404 171 5438 205
rect 5472 171 5506 205
rect 5540 171 5574 205
rect 5608 171 5642 205
rect 5676 171 5710 205
rect 5744 171 5768 205
<< viali >>
rect 88 1865 122 1874
rect 88 1840 122 1865
rect 88 1793 122 1802
rect 88 1768 122 1793
rect 88 1721 122 1730
rect 88 1696 122 1721
rect 68 374 102 381
rect 68 347 102 374
rect 68 303 102 309
rect 68 275 102 303
rect 360 1840 394 1874
rect 360 1768 394 1802
rect 360 1696 394 1730
rect 464 1194 498 1228
rect 536 1194 570 1228
rect 376 1120 410 1154
rect 448 1142 482 1154
rect 448 1120 470 1142
rect 470 1120 482 1142
rect 360 347 394 381
rect 360 275 394 309
rect 802 1840 836 1874
rect 802 1768 836 1802
rect 802 1696 836 1730
rect 1114 1840 1148 1874
rect 1114 1768 1148 1802
rect 1114 1696 1148 1730
rect 1380 1840 1414 1874
rect 1380 1768 1414 1802
rect 1380 1696 1414 1730
rect 1692 1840 1726 1874
rect 1692 1768 1726 1802
rect 1692 1696 1726 1730
rect 2004 1840 2038 1874
rect 2004 1768 2038 1802
rect 2004 1696 2038 1730
rect 2316 1840 2350 1874
rect 2316 1768 2350 1802
rect 2316 1696 2350 1730
rect 2628 1840 2662 1874
rect 2628 1768 2662 1802
rect 2628 1696 2662 1730
rect 2940 1840 2974 1874
rect 2940 1768 2974 1802
rect 2940 1696 2974 1730
rect 3252 1840 3286 1874
rect 3252 1768 3286 1802
rect 3252 1696 3286 1730
rect 3604 1840 3638 1874
rect 3604 1768 3638 1802
rect 3604 1696 3638 1730
rect 3956 1840 3990 1874
rect 3956 1768 3990 1802
rect 3956 1696 3990 1730
rect 4308 1840 4342 1874
rect 4308 1768 4342 1802
rect 4308 1696 4342 1730
rect 4660 1840 4694 1874
rect 4660 1768 4694 1802
rect 4660 1696 4694 1730
rect 6134 1863 6168 1874
rect 6134 1840 6168 1863
rect 6134 1795 6168 1802
rect 6134 1768 6168 1795
rect 6134 1727 6168 1730
rect 6134 1696 6168 1727
rect 2436 1613 2470 1647
rect 2508 1613 2542 1647
rect 2748 1613 2782 1647
rect 2820 1613 2854 1647
rect 3024 1613 3058 1647
rect 3096 1613 3130 1647
rect 3390 1616 3424 1650
rect 3462 1616 3496 1650
rect 3742 1616 3776 1650
rect 3814 1616 3848 1650
rect 4094 1616 4128 1650
rect 4166 1616 4200 1650
rect 4446 1616 4480 1650
rect 4518 1616 4552 1650
rect 4888 1616 4922 1650
rect 4960 1616 4994 1650
rect 5200 1616 5234 1650
rect 5272 1616 5306 1650
rect 5516 1533 5550 1567
rect 5588 1533 5622 1567
rect 5828 1533 5862 1567
rect 5900 1533 5934 1567
rect 1498 1456 1532 1490
rect 1570 1456 1604 1490
rect 1814 1456 1848 1490
rect 1886 1456 1920 1490
rect 2126 1453 2160 1487
rect 2198 1453 2232 1487
rect 4770 1456 4804 1490
rect 4842 1456 4876 1490
rect 5044 1456 5078 1490
rect 5116 1456 5150 1490
rect 5356 1456 5390 1490
rect 5428 1456 5462 1490
rect 5669 1456 5703 1490
rect 5741 1456 5775 1490
rect 5946 1456 5980 1490
rect 6018 1456 6052 1490
rect 924 1358 958 1392
rect 996 1358 1030 1392
rect 1198 1358 1232 1392
rect 1270 1358 1304 1392
rect 890 1129 924 1145
rect 890 1111 924 1129
rect 890 1061 924 1073
rect 890 1039 924 1061
rect 1036 1111 1070 1145
rect 1036 1043 1070 1073
rect 1036 1039 1070 1043
rect 1175 1111 1209 1145
rect 1175 1043 1209 1073
rect 1175 1039 1209 1043
rect 1705 961 1739 988
rect 1777 961 1811 988
rect 1849 961 1883 988
rect 1921 961 1955 988
rect 1705 954 1717 961
rect 1717 954 1739 961
rect 1777 954 1785 961
rect 1785 954 1811 961
rect 1849 954 1853 961
rect 1853 954 1883 961
rect 1921 954 1955 961
rect 5663 1039 5687 1062
rect 5687 1039 5697 1062
rect 5735 1039 5758 1062
rect 5758 1039 5769 1062
rect 5807 1039 5829 1062
rect 5829 1039 5841 1062
rect 5879 1039 5900 1062
rect 5900 1039 5913 1062
rect 5951 1039 5970 1062
rect 5970 1039 5985 1062
rect 5663 1028 5697 1039
rect 5735 1028 5769 1039
rect 5807 1028 5841 1039
rect 5879 1028 5913 1039
rect 5951 1028 5985 1039
rect 4978 927 5012 961
rect 5050 927 5084 961
rect 5122 927 5156 961
rect 5194 927 5228 961
rect 622 879 656 913
rect 694 879 728 913
rect 2052 879 2086 913
rect 2124 879 2158 913
rect 2196 879 2230 913
rect 2268 879 2302 913
rect 2132 799 2166 833
rect 2204 799 2238 833
rect 3648 765 3682 799
rect 3720 765 3754 799
rect 3999 765 4033 799
rect 4071 765 4105 799
rect 4352 765 4386 799
rect 4424 765 4458 799
rect 4704 691 4738 725
rect 4776 691 4810 725
rect 5056 691 5090 725
rect 5128 691 5162 725
rect 5408 691 5442 725
rect 5480 691 5514 725
rect 998 527 1032 561
rect 1070 527 1104 561
rect 1278 527 1312 561
rect 1350 527 1384 561
rect 1775 527 1809 561
rect 1847 527 1881 561
rect 1636 453 1670 487
rect 1708 453 1742 487
rect 1954 453 1988 487
rect 2026 453 2060 487
rect 2268 453 2302 487
rect 2340 453 2374 487
rect 2592 453 2626 487
rect 2664 453 2698 487
rect 2943 453 2977 487
rect 3015 453 3049 487
rect 3296 453 3330 487
rect 3368 453 3402 487
rect 822 347 856 381
rect 822 275 856 309
rect 1174 347 1208 381
rect 1174 275 1208 309
rect 1526 347 1560 381
rect 1526 275 1560 309
rect 2450 347 2484 381
rect 2450 275 2484 309
rect 2802 347 2836 381
rect 2802 275 2836 309
rect 3154 347 3188 381
rect 3154 275 3188 309
rect 3506 347 3540 381
rect 3506 275 3540 309
rect 3858 347 3892 381
rect 3858 275 3892 309
rect 4210 347 4244 381
rect 4210 275 4244 309
rect 4562 347 4596 381
rect 4562 275 4596 309
rect 4914 347 4948 381
rect 4914 275 4948 309
rect 5266 347 5300 381
rect 5266 275 5300 309
rect 5618 347 5652 381
rect 5618 275 5652 309
rect 5734 377 5768 381
rect 5734 347 5768 377
rect 5734 303 5768 309
rect 5734 275 5768 303
<< metal1 >>
rect 82 1874 6234 1886
rect 82 1840 88 1874
rect 122 1840 360 1874
rect 394 1840 802 1874
rect 836 1840 1114 1874
rect 1148 1840 1380 1874
rect 1414 1840 1692 1874
rect 1726 1840 2004 1874
rect 2038 1840 2316 1874
rect 2350 1840 2628 1874
rect 2662 1840 2940 1874
rect 2974 1840 3252 1874
rect 3286 1840 3604 1874
rect 3638 1840 3956 1874
rect 3990 1840 4308 1874
rect 4342 1840 4660 1874
rect 4694 1840 6134 1874
rect 6168 1840 6234 1874
rect 82 1802 6234 1840
rect 82 1768 88 1802
rect 122 1768 360 1802
rect 394 1768 802 1802
rect 836 1768 1114 1802
rect 1148 1768 1380 1802
rect 1414 1768 1692 1802
rect 1726 1768 2004 1802
rect 2038 1768 2316 1802
rect 2350 1768 2628 1802
rect 2662 1768 2940 1802
rect 2974 1768 3252 1802
rect 3286 1768 3604 1802
rect 3638 1768 3956 1802
rect 3990 1768 4308 1802
rect 4342 1768 4660 1802
rect 4694 1768 6134 1802
rect 6168 1768 6234 1802
rect 82 1730 6234 1768
rect 82 1696 88 1730
rect 122 1696 360 1730
rect 394 1696 802 1730
rect 836 1696 1114 1730
rect 1148 1696 1380 1730
rect 1414 1696 1692 1730
rect 1726 1696 2004 1730
rect 2038 1696 2316 1730
rect 2350 1696 2628 1730
rect 2662 1696 2940 1730
rect 2974 1696 3252 1730
rect 3286 1696 3604 1730
rect 3638 1696 3956 1730
rect 3990 1696 4308 1730
rect 4342 1696 4660 1730
rect 4694 1696 6134 1730
rect 6168 1696 6234 1730
rect 82 1684 6234 1696
rect 1163 1604 1169 1656
rect 1221 1604 1233 1656
rect 1285 1604 2420 1656
rect 2472 1604 2484 1656
rect 2536 1647 3142 1656
rect 2542 1613 2748 1647
rect 2782 1613 2820 1647
rect 2854 1613 3024 1647
rect 3058 1613 3096 1647
rect 3130 1613 3142 1647
rect 2536 1604 3142 1613
rect 3378 1650 5318 1656
rect 3378 1616 3390 1650
rect 3424 1616 3462 1650
rect 3496 1616 3742 1650
rect 3776 1616 3814 1650
rect 3848 1616 4094 1650
rect 4128 1616 4166 1650
rect 4200 1616 4446 1650
rect 4480 1616 4518 1650
rect 4552 1616 4888 1650
rect 4922 1616 4960 1650
rect 4994 1616 5200 1650
rect 5234 1616 5272 1650
rect 5306 1616 5318 1650
rect 3378 1610 5318 1616
rect 2570 1524 2576 1576
rect 2628 1524 2640 1576
rect 2692 1524 5138 1576
rect 5190 1524 5202 1576
rect 5254 1567 5946 1576
rect 5254 1533 5516 1567
rect 5550 1533 5588 1567
rect 5622 1533 5828 1567
rect 5862 1533 5900 1567
rect 5934 1533 5946 1567
rect 5254 1524 5946 1533
rect 1486 1490 4647 1496
tri 4647 1490 4653 1496 sw
rect 4758 1490 6064 1496
rect 1486 1456 1498 1490
rect 1532 1456 1570 1490
rect 1604 1456 1814 1490
rect 1848 1456 1886 1490
rect 1920 1487 4653 1490
rect 1920 1456 2126 1487
rect 1486 1453 2126 1456
rect 2160 1453 2198 1487
rect 2232 1481 4653 1487
tri 4653 1481 4662 1490 sw
rect 2232 1456 4662 1481
tri 4662 1456 4687 1481 sw
rect 4758 1456 4770 1490
rect 4804 1456 4842 1490
rect 4876 1456 5044 1490
rect 5078 1456 5116 1490
rect 5150 1456 5356 1490
rect 5390 1456 5428 1490
rect 5462 1456 5669 1490
rect 5703 1456 5741 1490
rect 5775 1456 5946 1490
rect 5980 1456 6018 1490
rect 6052 1456 6064 1490
rect 2232 1453 4687 1456
rect 1486 1444 4687 1453
tri 4625 1407 4662 1444 ne
rect 4662 1407 4687 1444
tri 4687 1407 4736 1456 sw
rect 4758 1450 6064 1456
tri 4662 1398 4671 1407 ne
rect 4671 1398 4982 1407
rect 912 1392 1316 1398
rect 912 1358 924 1392
rect 958 1358 996 1392
rect 1030 1358 1198 1392
rect 1232 1358 1270 1392
rect 1304 1358 1316 1392
rect 912 1346 1316 1358
tri 4671 1355 4714 1398 ne
rect 4714 1355 4982 1398
rect 5034 1355 5046 1407
rect 5098 1355 5104 1407
rect 452 1228 4764 1234
rect 452 1194 464 1228
rect 498 1194 536 1228
rect 570 1194 4764 1228
rect 452 1188 4764 1194
tri 3313 1163 3338 1188 ne
rect 364 1154 930 1160
rect 364 1120 376 1154
rect 410 1120 448 1154
rect 482 1145 930 1154
rect 482 1120 890 1145
rect 364 1114 890 1120
tri 859 1111 862 1114 ne
rect 862 1111 890 1114
rect 924 1111 930 1145
tri 862 1089 884 1111 ne
rect 884 1073 930 1111
rect 884 1039 890 1073
rect 924 1039 930 1073
rect 884 1027 930 1039
rect 1030 1145 1076 1157
rect 1030 1111 1036 1145
rect 1070 1111 1076 1145
rect 1030 1073 1076 1111
rect 1030 1039 1036 1073
rect 1070 1039 1076 1073
tri 1013 927 1030 944 se
rect 1030 927 1076 1039
rect 1163 1151 1215 1157
rect 1163 1087 1215 1099
rect 1350 1096 1356 1148
rect 1408 1096 1420 1148
rect 1472 1096 2293 1148
rect 2375 1096 2576 1148
rect 2628 1096 2640 1148
rect 2692 1096 3225 1148
rect 3338 1096 4764 1188
rect 4819 1096 4982 1148
rect 5034 1096 5046 1148
rect 5098 1096 5381 1148
rect 1163 1023 1215 1035
rect 1279 1062 5997 1068
rect 1279 1028 5663 1062
rect 5697 1028 5735 1062
rect 5769 1028 5807 1062
rect 5841 1028 5879 1062
rect 5913 1028 5951 1062
rect 5985 1028 5997 1062
rect 1279 1022 5997 1028
tri 1215 994 1240 1019 sw
rect 1215 988 1967 994
rect 1215 971 1705 988
rect 1163 954 1705 971
rect 1739 954 1777 988
rect 1811 954 1849 988
rect 1883 954 1921 988
rect 1955 954 1967 988
tri 2447 961 2453 967 se
rect 2453 961 4505 967
rect 1163 948 1967 954
tri 2434 948 2447 961 se
rect 2447 948 4505 961
tri 2430 944 2434 948 se
rect 2434 944 4505 948
tri 1076 927 1093 944 sw
tri 2413 927 2430 944 se
rect 2430 927 4505 944
tri 1005 919 1013 927 se
rect 1013 919 1093 927
tri 1093 919 1101 927 sw
tri 2405 919 2413 927 se
rect 2413 919 4505 927
rect 610 913 2314 919
rect 610 879 622 913
rect 656 879 694 913
rect 728 879 2052 913
rect 2086 879 2124 913
rect 2158 879 2196 913
rect 2230 879 2268 913
rect 2302 879 2314 913
tri 2379 893 2405 919 se
rect 2405 915 4505 919
rect 4966 961 4982 967
rect 4966 927 4978 961
rect 4966 915 4982 927
rect 5034 915 5046 967
rect 5098 961 5240 967
rect 5098 927 5122 961
rect 5156 927 5194 961
rect 5228 927 5240 961
rect 5098 915 5240 927
rect 2405 893 2453 915
tri 2453 893 2475 915 nw
rect 610 873 2314 879
tri 2359 873 2379 893 se
rect 2379 873 2405 893
tri 2331 845 2359 873 se
rect 2359 845 2405 873
tri 2405 845 2453 893 nw
rect 1350 793 1356 845
rect 1408 793 1420 845
rect 1472 833 2359 845
rect 1472 799 2132 833
rect 2166 799 2204 833
rect 2238 799 2359 833
tri 2359 799 2405 845 nw
rect 3636 799 4982 811
rect 1472 793 2353 799
tri 2353 793 2359 799 nw
rect 3636 765 3648 799
rect 3682 765 3720 799
rect 3754 765 3999 799
rect 4033 765 4071 799
rect 4105 765 4352 799
rect 4386 765 4424 799
rect 4458 765 4982 799
rect 3636 759 4982 765
rect 5034 759 5046 811
rect 5098 759 5104 811
rect 4692 725 5138 731
rect 4692 691 4704 725
rect 4738 691 4776 725
rect 4810 691 5056 725
rect 5090 691 5128 725
rect 4692 679 5138 691
rect 5190 679 5202 731
rect 5254 725 5526 731
rect 5254 691 5408 725
rect 5442 691 5480 725
rect 5514 691 5526 725
rect 5254 679 5526 691
rect -119 462 86 674
rect 986 561 1893 567
rect 986 527 998 561
rect 1032 527 1070 561
rect 1104 527 1278 561
rect 1312 527 1350 561
rect 1384 527 1775 561
rect 1809 527 1847 561
rect 1881 527 1893 561
rect 986 521 1893 527
rect 1624 487 2386 493
rect 1624 453 1636 487
rect 1670 453 1708 487
rect 1742 453 1954 487
rect 1988 453 2026 487
rect 2060 453 2268 487
rect 2302 453 2340 487
rect 2374 453 2386 487
rect 1624 447 2386 453
rect 2414 447 2420 499
rect 2472 447 2484 499
rect 2536 487 3414 499
rect 2536 453 2592 487
rect 2626 453 2664 487
rect 2698 453 2943 487
rect 2977 453 3015 487
rect 3049 453 3296 487
rect 3330 453 3368 487
rect 3402 453 3414 487
rect 2536 447 3414 453
rect -22 381 5794 419
rect -22 347 68 381
rect 102 347 360 381
rect 394 347 822 381
rect 856 347 1174 381
rect 1208 347 1526 381
rect 1560 347 2450 381
rect 2484 347 2802 381
rect 2836 347 3154 381
rect 3188 347 3506 381
rect 3540 347 3858 381
rect 3892 347 4210 381
rect 4244 347 4562 381
rect 4596 347 4914 381
rect 4948 347 5266 381
rect 5300 347 5618 381
rect 5652 347 5734 381
rect 5768 347 5794 381
rect -22 309 5794 347
rect -22 275 68 309
rect 102 275 360 309
rect 394 275 822 309
rect 856 275 1174 309
rect 1208 275 1526 309
rect 1560 275 2450 309
rect 2484 275 2802 309
rect 2836 275 3154 309
rect 3188 275 3506 309
rect 3540 275 3858 309
rect 3892 275 4210 309
rect 4244 275 4562 309
rect 4596 275 4914 309
rect 4948 275 5266 309
rect 5300 275 5618 309
rect 5652 275 5734 309
rect 5768 275 5794 309
rect -22 217 5794 275
<< via1 >>
rect 1169 1604 1221 1656
rect 1233 1604 1285 1656
rect 2420 1647 2472 1656
rect 2420 1613 2436 1647
rect 2436 1613 2470 1647
rect 2470 1613 2472 1647
rect 2420 1604 2472 1613
rect 2484 1647 2536 1656
rect 2484 1613 2508 1647
rect 2508 1613 2536 1647
rect 2484 1604 2536 1613
rect 2576 1524 2628 1576
rect 2640 1524 2692 1576
rect 5138 1524 5190 1576
rect 5202 1524 5254 1576
rect 4982 1355 5034 1407
rect 5046 1355 5098 1407
rect 1163 1145 1215 1151
rect 1163 1111 1175 1145
rect 1175 1111 1209 1145
rect 1209 1111 1215 1145
rect 1163 1099 1215 1111
rect 1356 1096 1408 1148
rect 1420 1096 1472 1148
rect 2576 1096 2628 1148
rect 2640 1096 2692 1148
rect 4982 1096 5034 1148
rect 5046 1096 5098 1148
rect 1163 1073 1215 1087
rect 1163 1039 1175 1073
rect 1175 1039 1209 1073
rect 1209 1039 1215 1073
rect 1163 1035 1215 1039
rect 1163 971 1215 1023
rect 4982 961 5034 967
rect 4982 927 5012 961
rect 5012 927 5034 961
rect 4982 915 5034 927
rect 5046 961 5098 967
rect 5046 927 5050 961
rect 5050 927 5084 961
rect 5084 927 5098 961
rect 5046 915 5098 927
rect 1356 793 1408 845
rect 1420 793 1472 845
rect 4982 759 5034 811
rect 5046 759 5098 811
rect 5138 725 5190 731
rect 5138 691 5162 725
rect 5162 691 5190 725
rect 5138 679 5190 691
rect 5202 679 5254 731
rect 2420 447 2472 499
rect 2484 447 2536 499
<< metal2 >>
rect 1163 1604 1169 1656
rect 1221 1604 1233 1656
rect 1285 1604 1291 1656
rect 2414 1604 2420 1656
rect 2472 1604 2484 1656
rect 2536 1604 2542 1656
rect 1163 1151 1215 1604
tri 1215 1579 1240 1604 nw
rect 1163 1087 1215 1099
rect 1163 1023 1215 1035
rect 1163 965 1215 971
rect 1350 1096 1356 1148
rect 1408 1096 1420 1148
rect 1472 1096 1478 1148
rect 1350 845 1478 1096
rect 1350 793 1356 845
rect 1408 793 1420 845
rect 1472 793 1478 845
rect -72 503 -38 537
rect 2414 499 2542 1604
rect 2570 1524 2576 1576
rect 2628 1524 2640 1576
rect 2692 1524 2698 1576
rect 2570 1148 2698 1524
rect 5132 1524 5138 1576
rect 5190 1524 5202 1576
rect 5254 1524 5260 1576
rect 2570 1096 2576 1148
rect 2628 1096 2640 1148
rect 2692 1096 2698 1148
rect 4976 1355 4982 1407
rect 5034 1355 5046 1407
rect 5098 1355 5104 1407
rect 4976 1148 5104 1355
rect 4976 1096 4982 1148
rect 5034 1096 5046 1148
rect 5098 1096 5104 1148
rect 4976 967 5104 1096
rect 4976 915 4982 967
rect 5034 915 5046 967
rect 5098 915 5104 967
rect 4976 811 5104 915
rect 4976 759 4982 811
rect 5034 759 5046 811
rect 5098 759 5104 811
rect 5132 731 5260 1524
rect 5132 679 5138 731
rect 5190 679 5202 731
rect 5254 679 5260 731
rect 2414 447 2420 499
rect 2472 447 2484 499
rect 2536 447 2542 499
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1704896540
transform 0 -1 1209 -1 0 1145
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1704896540
transform 0 -1 1070 -1 0 1145
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1704896540
transform 0 -1 856 -1 0 381
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1704896540
transform 0 -1 102 -1 0 381
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_4
timestamp 1704896540
transform 0 -1 5768 -1 0 381
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_5
timestamp 1704896540
transform 0 -1 394 -1 0 381
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_6
timestamp 1704896540
transform 0 -1 924 -1 0 1145
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_7
timestamp 1704896540
transform 0 -1 2484 -1 0 381
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_8
timestamp 1704896540
transform 0 -1 1560 -1 0 381
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_9
timestamp 1704896540
transform 0 -1 1208 -1 0 381
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_10
timestamp 1704896540
transform 0 -1 2836 -1 0 381
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_11
timestamp 1704896540
transform 0 -1 3188 -1 0 381
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_12
timestamp 1704896540
transform 0 -1 3540 -1 0 381
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_13
timestamp 1704896540
transform 0 -1 3892 -1 0 381
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_14
timestamp 1704896540
transform 0 -1 4244 -1 0 381
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_15
timestamp 1704896540
transform 0 -1 4596 -1 0 381
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_16
timestamp 1704896540
transform 0 -1 4948 -1 0 381
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_17
timestamp 1704896540
transform 0 -1 5300 -1 0 381
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_18
timestamp 1704896540
transform 0 -1 5652 -1 0 381
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_19
timestamp 1704896540
transform -1 0 6052 0 1 1456
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_20
timestamp 1704896540
transform -1 0 5514 0 1 691
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_21
timestamp 1704896540
transform -1 0 5162 0 1 691
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_22
timestamp 1704896540
transform -1 0 4810 0 1 691
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_23
timestamp 1704896540
transform -1 0 570 0 1 1194
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_24
timestamp 1704896540
transform -1 0 3496 0 1 1616
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_25
timestamp 1704896540
transform -1 0 3848 0 1 1616
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_26
timestamp 1704896540
transform -1 0 4200 0 1 1616
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_27
timestamp 1704896540
transform -1 0 4552 0 1 1616
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_28
timestamp 1704896540
transform -1 0 5306 0 1 1616
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_29
timestamp 1704896540
transform -1 0 4994 0 1 1616
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_30
timestamp 1704896540
transform -1 0 4876 0 1 1456
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_31
timestamp 1704896540
transform -1 0 5150 0 1 1456
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_32
timestamp 1704896540
transform -1 0 5462 0 1 1456
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_33
timestamp 1704896540
transform -1 0 1304 0 1 1358
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_34
timestamp 1704896540
transform -1 0 1030 0 1 1358
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_35
timestamp 1704896540
transform -1 0 2232 0 1 1453
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_36
timestamp 1704896540
transform -1 0 2374 0 1 453
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_37
timestamp 1704896540
transform -1 0 2060 0 1 453
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_38
timestamp 1704896540
transform -1 0 1742 0 1 453
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_39
timestamp 1704896540
transform -1 0 2238 0 1 799
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_40
timestamp 1704896540
transform -1 0 2854 0 1 1613
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_41
timestamp 1704896540
transform -1 0 5934 0 1 1533
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_42
timestamp 1704896540
transform -1 0 5622 0 1 1533
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_43
timestamp 1704896540
transform -1 0 3130 0 1 1613
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_44
timestamp 1704896540
transform -1 0 2542 0 1 1613
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_45
timestamp 1704896540
transform -1 0 1920 0 1 1456
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_46
timestamp 1704896540
transform -1 0 1604 0 1 1456
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_47
timestamp 1704896540
transform -1 0 1881 0 1 527
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_48
timestamp 1704896540
transform -1 0 1104 0 1 527
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_49
timestamp 1704896540
transform -1 0 5775 0 1 1456
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_50
timestamp 1704896540
transform -1 0 482 0 1 1120
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_51
timestamp 1704896540
transform -1 0 1384 0 1 527
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_52
timestamp 1704896540
transform 1 0 622 0 1 879
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_53
timestamp 1704896540
transform 1 0 2943 0 1 453
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_54
timestamp 1704896540
transform 1 0 2592 0 1 453
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_55
timestamp 1704896540
transform 1 0 3296 0 1 453
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_56
timestamp 1704896540
transform 1 0 4352 0 1 765
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_57
timestamp 1704896540
transform 1 0 3999 0 1 765
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_58
timestamp 1704896540
transform 1 0 3648 0 1 765
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1704896540
transform 0 -1 122 1 0 1696
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_1
timestamp 1704896540
transform 0 -1 4694 1 0 1696
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_2
timestamp 1704896540
transform 0 -1 4342 1 0 1696
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_3
timestamp 1704896540
transform 0 -1 3990 1 0 1696
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_4
timestamp 1704896540
transform 0 -1 2662 1 0 1696
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_5
timestamp 1704896540
transform 0 -1 2974 1 0 1696
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_6
timestamp 1704896540
transform 0 -1 3286 1 0 1696
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_7
timestamp 1704896540
transform 0 -1 3638 1 0 1696
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_8
timestamp 1704896540
transform 0 -1 2350 1 0 1696
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_9
timestamp 1704896540
transform 0 -1 2038 1 0 1696
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_10
timestamp 1704896540
transform 0 -1 1726 1 0 1696
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_11
timestamp 1704896540
transform 0 -1 1414 1 0 1696
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_12
timestamp 1704896540
transform 0 -1 1148 1 0 1696
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_13
timestamp 1704896540
transform 0 -1 836 1 0 1696
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_14
timestamp 1704896540
transform 0 -1 394 1 0 1696
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_15
timestamp 1704896540
transform 0 -1 6168 1 0 1696
box 0 0 1 1
use L1M1_CDNS_52468879185191  L1M1_CDNS_52468879185191_0
timestamp 1704896540
transform -1 0 3213 0 1 1108
box -12 -6 838 40
use L1M1_CDNS_52468879185191  L1M1_CDNS_52468879185191_1
timestamp 1704896540
transform 1 0 1455 0 1 1108
box -12 -6 838 40
use L1M1_CDNS_52468879185193  L1M1_CDNS_52468879185193_0
timestamp 1704896540
transform 1 0 5663 0 1 1028
box 0 0 1 1
use L1M1_CDNS_52468879185195  L1M1_CDNS_52468879185195_0
timestamp 1704896540
transform 1 0 4831 0 1 1108
box -12 -6 550 40
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_0
timestamp 1704896540
transform -1 0 2302 0 1 879
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_1
timestamp 1704896540
transform -1 0 1955 0 1 954
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_2
timestamp 1704896540
transform -1 0 5228 0 1 927
box 0 0 1 1
use L1M1_CDNS_52468879185302  L1M1_CDNS_52468879185302_0
timestamp 1704896540
transform 0 1 -98 -1 0 822
box -12 -6 262 184
use L1M1_CDNS_52468879185307  L1M1_CDNS_52468879185307_0
timestamp 1704896540
transform 1 0 3350 0 1 1108
box -12 -6 1414 40
use L1M1_CDNS_52468879185336  L1M1_CDNS_52468879185336_0
timestamp 1704896540
transform 1 0 1289 0 1 1028
box -12 -6 1558 40
use L1M1_CDNS_52468879185381  L1M1_CDNS_52468879185381_0
timestamp 1704896540
transform -1 0 4493 0 1 927
box -12 -6 910 40
use L1M1_CDNS_52468879185448  L1M1_CDNS_52468879185448_0
timestamp 1704896540
transform 1 0 3298 0 1 1028
box -12 -6 1270 40
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1704896540
transform -1 0 2698 0 1 1524
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_1
timestamp 1704896540
transform -1 0 5104 0 1 1096
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_2
timestamp 1704896540
transform -1 0 5104 0 1 915
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_3
timestamp 1704896540
transform -1 0 5104 0 1 759
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_4
timestamp 1704896540
transform -1 0 2698 0 -1 1148
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_5
timestamp 1704896540
transform 1 0 1350 0 -1 1148
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_6
timestamp 1704896540
transform 1 0 1350 0 -1 845
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_7
timestamp 1704896540
transform 1 0 5132 0 1 679
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_8
timestamp 1704896540
transform 1 0 5132 0 1 1524
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_9
timestamp 1704896540
transform 1 0 4976 0 1 1355
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_10
timestamp 1704896540
transform 1 0 1163 0 1 1604
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_11
timestamp 1704896540
transform 1 0 2414 0 1 1604
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_12
timestamp 1704896540
transform 1 0 2414 0 1 447
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_0
timestamp 1704896540
transform 0 -1 1215 -1 0 1157
box 0 0 1 1
use M1M2_CDNS_524688791851031  M1M2_CDNS_524688791851031_0
timestamp 1704896540
transform -1 0 9 0 -1 834
box 0 0 128 372
use nfet_CDNS_52468879185310  nfet_CDNS_52468879185310_0
timestamp 1704896540
transform -1 0 811 0 1 279
box -79 -26 199 626
use nfet_CDNS_52468879185319  nfet_CDNS_52468879185319_0
timestamp 1704896540
transform 1 0 4959 0 1 279
box -79 -26 375 626
use nfet_CDNS_52468879185319  nfet_CDNS_52468879185319_1
timestamp 1704896540
transform 1 0 5311 0 1 279
box -79 -26 375 626
use nfet_CDNS_52468879185319  nfet_CDNS_52468879185319_2
timestamp 1704896540
transform 1 0 4607 0 1 279
box -79 -26 375 626
use nfet_CDNS_52468879185365  nfet_CDNS_52468879185365_0
timestamp 1704896540
transform 1 0 1681 0 1 279
box -79 -26 375 626
use nfet_CDNS_52468879185365  nfet_CDNS_52468879185365_1
timestamp 1704896540
transform 1 0 2033 0 1 279
box -79 -26 375 626
use nfet_CDNS_52468879185417  nfet_CDNS_52468879185417_0
timestamp 1704896540
transform -1 0 349 0 1 279
box -79 -26 199 626
use nfet_CDNS_52468879185450  nfet_CDNS_52468879185450_0
timestamp 1704896540
transform -1 0 1515 0 1 279
box -79 -26 727 626
use nfet_CDNS_52468879185451  nfet_CDNS_52468879185451_0
timestamp 1704896540
transform -1 0 3495 0 1 279
box -79 -26 1079 626
use nfet_CDNS_52468879185451  nfet_CDNS_52468879185451_1
timestamp 1704896540
transform 1 0 3551 0 1 279
box -79 -26 1079 626
use nfet_CDNS_52468879185452  nfet_CDNS_52468879185452_0
timestamp 1704896540
transform 1 0 405 0 1 279
box -82 -26 199 626
use pfet_CDNS_52468879185355  pfet_CDNS_52468879185355_0
timestamp 1704896540
transform -1 0 6007 0 -1 2193
box -119 -66 687 1066
use pfet_CDNS_52468879185355  pfet_CDNS_52468879185355_1
timestamp 1704896540
transform 1 0 4815 0 -1 2193
box -119 -66 687 1066
use pfet_CDNS_52468879185453  pfet_CDNS_52468879185453_0
timestamp 1704896540
transform -1 0 3241 0 -1 2193
box -119 -66 999 1066
use pfet_CDNS_52468879185454  pfet_CDNS_52468879185454_0
timestamp 1704896540
transform 1 0 3297 0 -1 2193
box -119 -66 1471 1066
use pfet_CDNS_52468879185455  pfet_CDNS_52468879185455_0
timestamp 1704896540
transform -1 0 1103 0 -1 2193
box -119 -66 219 1066
use pfet_CDNS_52468879185455  pfet_CDNS_52468879185455_1
timestamp 1704896540
transform -1 0 349 0 -1 2193
box -119 -66 219 1066
use pfet_CDNS_52468879185455  pfet_CDNS_52468879185455_2
timestamp 1704896540
transform -1 0 947 0 -1 2193
box -119 -66 219 1066
use pfet_CDNS_52468879185455  pfet_CDNS_52468879185455_3
timestamp 1704896540
transform 1 0 405 0 -1 2193
box -119 -66 219 1066
use pfet_CDNS_52468879185455  pfet_CDNS_52468879185455_4
timestamp 1704896540
transform 1 0 1159 0 -1 2193
box -119 -66 219 1066
use pfet_CDNS_52468879185455  pfet_CDNS_52468879185455_5
timestamp 1704896540
transform 1 0 691 0 -1 2193
box -119 -66 219 1066
use pfet_CDNS_52468879185456  pfet_CDNS_52468879185456_0
timestamp 1704896540
transform -1 0 2305 0 -1 2193
box -119 -66 999 1066
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_0
timestamp 1704896540
transform -1 0 346 0 1 1027
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_1
timestamp 1704896540
transform 1 0 704 0 -1 1145
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_2
timestamp 1704896540
transform 1 0 1159 0 -1 1161
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_3
timestamp 1704896540
transform 1 0 874 0 -1 1145
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_4
timestamp 1704896540
transform 1 0 1020 0 1 1027
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_0
timestamp 1704896540
transform -1 0 486 0 -1 1158
box 0 0 1 1
use PYL1_CDNS_52468879185309  PYL1_CDNS_52468879185309_0
timestamp 1704896540
transform 0 -1 1971 -1 0 977
box 0 0 1 1
use PYL1_CDNS_52468879185309  PYL1_CDNS_52468879185309_1
timestamp 1704896540
transform 0 -1 2318 -1 0 977
box 0 0 1 1
use PYL1_CDNS_52468879185309  PYL1_CDNS_52468879185309_2
timestamp 1704896540
transform 0 1 5322 1 0 911
box 0 0 1 1
use PYL1_CDNS_52468879185318  PYL1_CDNS_52468879185318_0
timestamp 1704896540
transform 0 1 4819 -1 0 1161
box 0 0 66 542
use PYL1_CDNS_52468879185318  PYL1_CDNS_52468879185318_1
timestamp 1704896540
transform 0 1 5455 -1 0 1161
box 0 0 66 542
use PYL1_CDNS_52468879185332  PYL1_CDNS_52468879185332_0
timestamp 1704896540
transform 0 -1 3217 -1 0 1161
box 0 0 66 814
use PYL1_CDNS_52468879185332  PYL1_CDNS_52468879185332_1
timestamp 1704896540
transform 0 -1 2281 -1 0 1161
box 0 0 66 814
use PYL1_CDNS_52468879185383  PYL1_CDNS_52468879185383_0
timestamp 1704896540
transform 0 1 884 -1 0 985
box 0 0 66 610
use PYL1_CDNS_52468879185407  PYL1_CDNS_52468879185407_0
timestamp 1704896540
transform 0 -1 3479 -1 0 977
box 0 0 66 950
use PYL1_CDNS_52468879185407  PYL1_CDNS_52468879185407_1
timestamp 1704896540
transform 0 -1 4529 -1 0 977
box 0 0 66 950
use PYL1_CDNS_52468879185444  PYL1_CDNS_52468879185444_0
timestamp 1704896540
transform 1 0 5439 0 1 1027
box 0 0 1 1
use PYL1_CDNS_52468879185445  PYL1_CDNS_52468879185445_0
timestamp 1704896540
transform 0 1 4618 1 0 911
box 0 0 134 270
use PYL1_CDNS_52468879185445  PYL1_CDNS_52468879185445_1
timestamp 1704896540
transform 0 1 4970 1 0 911
box 0 0 134 270
use PYL1_CDNS_52468879185446  PYL1_CDNS_52468879185446_0
timestamp 1704896540
transform 0 1 3319 -1 0 1161
box 0 0 66 1426
use PYL1_CDNS_52468879185447  PYL1_CDNS_52468879185447_0
timestamp 1704896540
transform -1 0 3241 0 1 1007
box 0 0 1 1
<< labels >>
flabel comment s 5733 1093 5733 1093 0 FreeSans 300 180 0 0 pd_dis_h
flabel comment s 449 898 449 898 0 FreeSans 300 90 0 0 oe_i_h
flabel comment s 892 920 892 920 0 FreeSans 300 90 0 0 oe_i_h
flabel comment s 1165 1134 1165 1134 0 FreeSans 300 90 0 0 drvlo_h_n
flabel comment s 1851 1155 1851 1155 0 FreeSans 300 180 0 0 n0
flabel comment s 1024 1139 1024 1139 0 FreeSans 300 90 0 0 pu_dis_h_n
flabel comment s 2803 1098 2803 1098 0 FreeSans 300 180 0 0 n1
flabel comment s 4863 1097 4863 1097 0 FreeSans 300 180 0 0 drvhi_h
flabel comment s 4016 1098 4016 1098 0 FreeSans 300 180 0 0 oe_i_h_n
flabel comment s 536 1006 536 1006 0 FreeSans 300 90 0 0 oe_i_h_n
flabel comment s 2214 986 2214 986 0 FreeSans 300 0 0 0 pu_dis_h_n
flabel comment s 203 1006 203 1006 0 FreeSans 300 90 0 0 oe_i_h
flabel comment s 1808 1477 1808 1477 0 FreeSans 300 0 0 0 drvhi_h
flabel comment s 5446 975 5446 975 0 FreeSans 300 180 0 0 pd_dis_h
flabel comment s 3804 977 3804 977 0 FreeSans 300 180 0 0 n0
flabel comment s 1161 984 1161 984 0 FreeSans 300 0 0 0 oe_i_h
flabel comment s 1823 984 1823 984 0 FreeSans 300 0 0 0 drvlo_h_n
flabel comment s 740 904 740 904 0 FreeSans 300 270 0 0 pu_dis_h
flabel comment s 2946 986 2946 986 0 FreeSans 300 180 0 0 n1
flabel comment s 3833 786 3833 786 0 FreeSans 300 0 0 0 drvhi_h
flabel comment s 2777 474 2777 474 0 FreeSans 300 0 0 0 drvlo_h_n
flabel comment s 5673 1564 5673 1564 0 FreeSans 300 180 0 0 n1
flabel comment s 3108 1649 3108 1649 0 FreeSans 300 0 0 0 drvlo_h_n
flabel comment s 1069 552 1069 552 0 FreeSans 300 0 0 0 int_nand_n0
flabel comment s 1712 560 1712 560 0 FreeSans 300 0 0 0 int_nand_n1
flabel comment s 2238 560 2238 560 0 FreeSans 300 0 0 0 n0
flabel comment s 1233 1380 1233 1380 0 FreeSans 300 180 0 0 n0
flabel comment s 4906 1474 4906 1474 0 FreeSans 300 180 0 0 int_nor_n<1>
flabel comment s 311 872 311 872 0 FreeSans 300 270 0 0 oe_h_n
flabel comment s 4157 1645 4157 1645 0 FreeSans 300 180 0 0 int_nor_n<0>
flabel comment s 4722 1065 4722 1065 0 FreeSans 300 180 0 0 oe_i_h_n
flabel comment s 3050 1483 3050 1483 0 FreeSans 300 0 0 0 drvhi_h
flabel comment s 2486 1647 2486 1647 0 FreeSans 300 0 0 0 drvlo_h_n
flabel comment s 1696 1637 1696 1637 0 FreeSans 300 0 0 0 drvlo_h_n
flabel comment s 4861 709 4861 709 0 FreeSans 300 180 0 0 n1
flabel comment s 5095 971 5095 971 0 FreeSans 300 0 0 0 drvhi_h
flabel metal1 s 1163 1604 1215 1656 3 FreeSans 300 0 0 0 drvlo_h_n
port 2 nsew
flabel metal1 s 82 1684 122 1886 3 FreeSans 300 0 0 0 vcc_io
port 4 nsew
flabel metal1 s -22 217 18 419 3 FreeSans 300 0 0 0 vgnd
port 3 nsew
flabel metal1 s 6194 1684 6234 1886 3 FreeSans 300 180 0 0 vcc_io
port 4 nsew
flabel metal1 s 5754 217 5794 419 3 FreeSans 300 180 0 0 vgnd
port 3 nsew
flabel metal1 s 1486 1444 1536 1496 3 FreeSans 300 0 0 0 drvhi_h
port 5 nsew
flabel metal1 s 1189 1630 1189 1630 3 FreeSans 300 0 0 0 drvlo_h_n
flabel locali s 5947 1111 5997 1145 3 FreeSans 300 0 0 0 pd_dis_h
port 6 nsew
flabel locali s 720 1111 754 1145 3 FreeSans 300 0 0 0 pu_dis_h
port 7 nsew
flabel locali s 296 1077 330 1111 0 FreeSans 200 0 0 0 oe_h_n
port 8 nsew
flabel metal2 s -72 503 -38 537 0 FreeSans 200 0 0 0 vgnd
port 3 nsew
<< properties >>
string GDS_END 87629248
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 87590090
string path 2.625 56.025 2.625 29.175 
<< end >>
