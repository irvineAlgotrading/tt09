magic
tech sky130A
timestamp 1704896540
<< metal1 >>
rect 0 0 3 90
rect 189 0 192 90
<< via1 >>
rect 3 0 189 90
<< metal2 >>
rect 0 0 3 90
rect 189 0 192 90
<< properties >>
string GDS_END 79749016
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 79747732
<< end >>
