magic
tech sky130B
timestamp 1704896540
<< viali >>
rect 0 0 125 53
<< metal1 >>
rect -6 53 131 56
rect -6 0 0 53
rect 125 0 131 53
rect -6 -3 131 0
<< properties >>
string GDS_END 94937330
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 94936686
<< end >>
