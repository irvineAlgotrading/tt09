magic
tech sky130B
timestamp 1704896540
<< metal1 >>
rect 0 0 3 474
rect 61 0 64 474
<< via1 >>
rect 3 0 61 474
<< metal2 >>
rect 0 0 3 474
rect 61 0 64 474
<< properties >>
string GDS_END 85847216
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85845164
<< end >>
