magic
tech sky130A
timestamp 1704896540
<< viali >>
rect 0 0 53 1817
<< metal1 >>
rect -6 1817 59 1820
rect -6 0 0 1817
rect 53 0 59 1817
rect -6 -3 59 0
<< properties >>
string GDS_END 34469872
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 34463212
<< end >>
