magic
tech sky130B
timestamp 1704896540
<< metal1 >>
rect 0 0 3 762
rect 93 0 96 762
<< via1 >>
rect 3 0 93 762
<< metal2 >>
rect 0 0 3 762
rect 93 0 96 762
<< properties >>
string GDS_END 91738872
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 91734132
<< end >>
