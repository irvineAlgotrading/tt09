magic
tech sky130B
magscale 1 2
timestamp 1704896540
use hvnTran_CDNS_5246887918586  hvnTran_CDNS_5246887918586_0
timestamp 1704896540
transform 1 0 119 0 -1 -26
box -79 -26 199 166
use hvpTran_CDNS_5246887918588  hvpTran_CDNS_5246887918588_0
timestamp 1704896540
transform 1 0 119 0 -1 682
box -119 -66 239 266
use hvpTran_CDNS_5246887918588  hvpTran_CDNS_5246887918588_1
timestamp 1704896540
transform 1 0 119 0 1 750
box -119 -66 239 266
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1704896540
transform 0 -1 108 -1 0 -84
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1704896540
transform 0 -1 108 1 0 872
box 0 0 1 1
<< properties >>
string GDS_END 85589900
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85587840
string path 4.425 0.725 4.425 10.975 
<< end >>
