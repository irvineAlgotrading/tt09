magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< pwell >>
rect 79 639 89 658
<< obsli1 >>
rect 137 717 679 733
rect 137 683 139 717
rect 173 683 211 717
rect 245 683 283 717
rect 317 683 355 717
rect 389 683 427 717
rect 461 683 499 717
rect 533 683 571 717
rect 605 683 643 717
rect 677 683 679 717
rect 137 667 679 683
rect 47 605 81 621
rect 47 533 81 571
rect 47 461 81 499
rect 47 389 81 427
rect 47 317 81 355
rect 47 245 81 283
rect 47 173 81 211
rect 47 101 81 139
rect 47 51 81 67
rect 133 51 167 621
rect 219 605 253 621
rect 219 533 253 571
rect 219 461 253 499
rect 219 389 253 427
rect 219 317 253 355
rect 219 245 253 283
rect 219 173 253 211
rect 219 101 253 139
rect 219 51 253 67
rect 305 51 339 621
rect 391 605 425 621
rect 391 533 425 571
rect 391 461 425 499
rect 391 389 425 427
rect 391 317 425 355
rect 391 245 425 283
rect 391 173 425 211
rect 391 101 425 139
rect 391 51 425 67
rect 477 51 511 621
rect 563 605 597 621
rect 563 533 597 571
rect 563 461 597 499
rect 563 389 597 427
rect 563 317 597 355
rect 563 245 597 283
rect 563 173 597 211
rect 563 101 597 139
rect 563 51 597 67
rect 649 51 683 621
rect 735 605 769 621
rect 735 533 769 571
rect 735 461 769 499
rect 735 389 769 427
rect 735 317 769 355
rect 735 245 769 283
rect 735 173 769 211
rect 735 101 769 139
rect 735 51 769 67
<< obsli1c >>
rect 139 683 173 717
rect 211 683 245 717
rect 283 683 317 717
rect 355 683 389 717
rect 427 683 461 717
rect 499 683 533 717
rect 571 683 605 717
rect 643 683 677 717
rect 47 571 81 605
rect 47 499 81 533
rect 47 427 81 461
rect 47 355 81 389
rect 47 283 81 317
rect 47 211 81 245
rect 47 139 81 173
rect 47 67 81 101
rect 219 571 253 605
rect 219 499 253 533
rect 219 427 253 461
rect 219 355 253 389
rect 219 283 253 317
rect 219 211 253 245
rect 219 139 253 173
rect 219 67 253 101
rect 391 571 425 605
rect 391 499 425 533
rect 391 427 425 461
rect 391 355 425 389
rect 391 283 425 317
rect 391 211 425 245
rect 391 139 425 173
rect 391 67 425 101
rect 563 571 597 605
rect 563 499 597 533
rect 563 427 597 461
rect 563 355 597 389
rect 563 283 597 317
rect 563 211 597 245
rect 563 139 597 173
rect 563 67 597 101
rect 735 571 769 605
rect 735 499 769 533
rect 735 427 769 461
rect 735 355 769 389
rect 735 283 769 317
rect 735 211 769 245
rect 735 139 769 173
rect 735 67 769 101
<< metal1 >>
rect 127 717 689 729
rect 127 683 139 717
rect 173 683 211 717
rect 245 683 283 717
rect 317 683 355 717
rect 389 683 427 717
rect 461 683 499 717
rect 533 683 571 717
rect 605 683 643 717
rect 677 683 689 717
rect 127 671 689 683
rect 41 605 87 621
rect 41 571 47 605
rect 81 571 87 605
rect 41 533 87 571
rect 41 499 47 533
rect 81 499 87 533
rect 41 461 87 499
rect 41 427 47 461
rect 81 427 87 461
rect 41 389 87 427
rect 41 355 47 389
rect 81 355 87 389
rect 41 317 87 355
rect 41 283 47 317
rect 81 283 87 317
rect 41 245 87 283
rect 41 211 47 245
rect 81 211 87 245
rect 41 173 87 211
rect 41 139 47 173
rect 81 139 87 173
rect 41 101 87 139
rect 41 67 47 101
rect 81 67 87 101
rect 41 -29 87 67
rect 213 605 259 621
rect 213 571 219 605
rect 253 571 259 605
rect 213 533 259 571
rect 213 499 219 533
rect 253 499 259 533
rect 213 461 259 499
rect 213 427 219 461
rect 253 427 259 461
rect 213 389 259 427
rect 213 355 219 389
rect 253 355 259 389
rect 213 317 259 355
rect 213 283 219 317
rect 253 283 259 317
rect 213 245 259 283
rect 213 211 219 245
rect 253 211 259 245
rect 213 173 259 211
rect 213 139 219 173
rect 253 139 259 173
rect 213 101 259 139
rect 213 67 219 101
rect 253 67 259 101
rect 213 -29 259 67
rect 385 605 431 621
rect 385 571 391 605
rect 425 571 431 605
rect 385 533 431 571
rect 385 499 391 533
rect 425 499 431 533
rect 385 461 431 499
rect 385 427 391 461
rect 425 427 431 461
rect 385 389 431 427
rect 385 355 391 389
rect 425 355 431 389
rect 385 317 431 355
rect 385 283 391 317
rect 425 283 431 317
rect 385 245 431 283
rect 385 211 391 245
rect 425 211 431 245
rect 385 173 431 211
rect 385 139 391 173
rect 425 139 431 173
rect 385 101 431 139
rect 385 67 391 101
rect 425 67 431 101
rect 385 -29 431 67
rect 557 605 603 621
rect 557 571 563 605
rect 597 571 603 605
rect 557 533 603 571
rect 557 499 563 533
rect 597 499 603 533
rect 557 461 603 499
rect 557 427 563 461
rect 597 427 603 461
rect 557 389 603 427
rect 557 355 563 389
rect 597 355 603 389
rect 557 317 603 355
rect 557 283 563 317
rect 597 283 603 317
rect 557 245 603 283
rect 557 211 563 245
rect 597 211 603 245
rect 557 173 603 211
rect 557 139 563 173
rect 597 139 603 173
rect 557 101 603 139
rect 557 67 563 101
rect 597 67 603 101
rect 557 -29 603 67
rect 729 605 775 621
rect 729 571 735 605
rect 769 571 775 605
rect 729 533 775 571
rect 729 499 735 533
rect 769 499 775 533
rect 729 461 775 499
rect 729 427 735 461
rect 769 427 775 461
rect 729 389 775 427
rect 729 355 735 389
rect 769 355 775 389
rect 729 317 775 355
rect 729 283 735 317
rect 769 283 775 317
rect 729 245 775 283
rect 729 211 735 245
rect 769 211 775 245
rect 729 173 775 211
rect 729 139 735 173
rect 769 139 775 173
rect 729 101 775 139
rect 729 67 735 101
rect 769 67 775 101
rect 729 -29 775 67
rect 41 -89 775 -29
<< obsm1 >>
rect 124 51 176 621
rect 296 51 348 621
rect 468 51 520 621
rect 640 51 692 621
<< obsm2 >>
rect 117 473 183 627
rect 289 473 355 627
rect 461 473 527 627
rect 633 473 699 627
<< metal3 >>
rect 117 561 699 627
rect 117 473 183 561
rect 289 473 355 561
rect 461 473 527 561
rect 633 473 699 561
<< labels >>
rlabel metal3 s 633 473 699 561 6 DRAIN
port 1 nsew
rlabel metal3 s 461 473 527 561 6 DRAIN
port 1 nsew
rlabel metal3 s 289 473 355 561 6 DRAIN
port 1 nsew
rlabel metal3 s 117 561 699 627 6 DRAIN
port 1 nsew
rlabel metal3 s 117 473 183 561 6 DRAIN
port 1 nsew
rlabel metal1 s 127 671 689 729 6 GATE
port 2 nsew
rlabel metal1 s 729 -29 775 621 6 SOURCE
port 3 nsew
rlabel metal1 s 557 -29 603 621 6 SOURCE
port 3 nsew
rlabel metal1 s 385 -29 431 621 6 SOURCE
port 3 nsew
rlabel metal1 s 213 -29 259 621 6 SOURCE
port 3 nsew
rlabel metal1 s 41 -29 87 621 6 SOURCE
port 3 nsew
rlabel metal1 s 41 -89 775 -29 8 SOURCE
port 3 nsew
rlabel pwell s 79 639 89 658 6 SUBSTRATE
port 4 nsew
<< properties >>
string FIXED_BBOX 36 -89 780 733
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 10440928
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 10421650
string device primitive
<< end >>
