magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -38 261 1970 582
<< pwell >>
rect 273 157 457 201
rect 1576 181 1930 203
rect 1390 157 1930 181
rect 1 21 1930 157
rect 29 -17 63 21
<< locali >>
rect 17 195 87 325
rect 354 201 436 325
rect 1762 323 1828 492
rect 1762 299 1915 323
rect 1795 289 1915 299
rect 1804 179 1915 289
rect 1798 171 1915 179
rect 1795 165 1915 171
rect 1778 153 1915 165
rect 1778 53 1827 153
<< obsli1 >>
rect 0 527 1932 561
rect 17 393 69 493
rect 103 427 169 527
rect 203 409 247 493
rect 291 427 357 527
rect 17 359 167 393
rect 121 161 167 359
rect 17 127 167 161
rect 17 69 69 127
rect 201 113 247 409
rect 391 393 425 493
rect 472 450 638 484
rect 686 451 762 527
rect 286 359 425 393
rect 286 165 320 359
rect 470 315 570 391
rect 286 127 425 165
rect 470 141 514 315
rect 604 281 638 450
rect 798 417 832 475
rect 866 451 932 527
rect 1022 433 1148 483
rect 1184 451 1268 527
rect 1114 417 1148 433
rect 1308 417 1356 475
rect 672 367 942 417
rect 672 315 722 367
rect 824 281 874 313
rect 604 247 874 281
rect 604 239 688 247
rect 550 129 620 203
rect 103 17 169 93
rect 203 69 247 113
rect 291 17 357 93
rect 391 61 425 127
rect 654 93 688 239
rect 908 213 942 367
rect 722 147 804 213
rect 862 145 942 213
rect 976 331 1080 393
rect 1114 383 1356 417
rect 1402 389 1468 527
rect 976 179 1010 331
rect 1044 213 1080 295
rect 1114 281 1148 383
rect 1502 353 1536 475
rect 1594 383 1660 485
rect 1502 349 1576 353
rect 1182 315 1576 349
rect 1114 247 1498 281
rect 1160 179 1230 203
rect 976 145 1230 179
rect 485 53 688 93
rect 722 17 804 105
rect 862 59 912 145
rect 952 17 1016 109
rect 1264 95 1298 247
rect 1428 235 1498 247
rect 1332 201 1402 213
rect 1332 147 1468 201
rect 1538 136 1576 315
rect 1128 61 1298 95
rect 1338 17 1466 113
rect 1506 70 1576 136
rect 1610 265 1660 383
rect 1694 299 1728 527
rect 1862 357 1915 527
rect 1610 199 1770 265
rect 1610 69 1644 199
rect 1678 17 1744 165
rect 1861 17 1915 119
rect 0 -17 1932 17
<< metal1 >>
rect 0 496 1932 592
rect 753 184 811 193
rect 1397 184 1455 193
rect 753 156 1455 184
rect 753 147 811 156
rect 1397 147 1455 156
rect 0 -48 1932 48
<< obsm1 >>
rect 109 388 167 397
rect 477 388 535 397
rect 1029 388 1087 397
rect 109 360 1087 388
rect 109 351 167 360
rect 477 351 535 360
rect 1029 351 1087 360
rect 1033 252 1091 261
rect 584 224 1091 252
rect 584 193 627 224
rect 1033 215 1091 224
rect 201 184 259 193
rect 569 184 627 193
rect 201 156 627 184
rect 201 147 259 156
rect 569 147 627 156
<< labels >>
rlabel locali s 17 195 87 325 6 CLK
port 1 nsew clock input
rlabel locali s 354 201 436 325 6 D
port 2 nsew signal input
rlabel metal1 s 1397 147 1455 156 6 SET_B
port 3 nsew signal input
rlabel metal1 s 753 147 811 156 6 SET_B
port 3 nsew signal input
rlabel metal1 s 753 156 1455 184 6 SET_B
port 3 nsew signal input
rlabel metal1 s 1397 184 1455 193 6 SET_B
port 3 nsew signal input
rlabel metal1 s 753 184 811 193 6 SET_B
port 3 nsew signal input
rlabel metal1 s 0 -48 1932 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 21 1930 157 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1390 157 1930 181 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1576 181 1930 203 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 273 157 457 201 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 1970 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 1932 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1778 53 1827 153 6 Q
port 8 nsew signal output
rlabel locali s 1778 153 1915 165 6 Q
port 8 nsew signal output
rlabel locali s 1795 165 1915 171 6 Q
port 8 nsew signal output
rlabel locali s 1798 171 1915 179 6 Q
port 8 nsew signal output
rlabel locali s 1804 179 1915 289 6 Q
port 8 nsew signal output
rlabel locali s 1795 289 1915 299 6 Q
port 8 nsew signal output
rlabel locali s 1762 299 1915 323 6 Q
port 8 nsew signal output
rlabel locali s 1762 323 1828 492 6 Q
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1932 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2547008
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2530896
<< end >>
