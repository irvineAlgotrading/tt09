magic
tech sky130A
timestamp 1704896540
<< metal1 >>
rect 0 0 3 186
rect 253 0 256 186
<< via1 >>
rect 3 0 253 186
<< metal2 >>
rect 0 0 3 186
rect 253 0 256 186
<< properties >>
string GDS_END 88434074
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 88430870
<< end >>
