magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -38 261 1602 582
<< pwell >>
rect 1 21 1513 203
rect 30 -17 64 21
<< locali >>
rect 361 405 694 421
rect 809 405 1536 421
rect 361 371 1536 405
rect 193 303 726 337
rect 193 266 282 303
rect 80 215 282 266
rect 341 215 636 269
rect 670 199 726 303
rect 852 303 1400 337
rect 852 282 995 303
rect 760 199 995 282
rect 1074 215 1288 269
rect 1366 199 1400 303
rect 1434 268 1536 371
rect 1434 165 1470 268
rect 1313 131 1470 165
rect 1313 90 1347 131
rect 1056 54 1347 90
<< obsli1 >>
rect 0 527 1564 561
rect 18 333 77 527
rect 191 455 257 527
rect 291 455 687 493
rect 111 421 155 438
rect 291 421 327 455
rect 723 439 777 527
rect 887 455 953 527
rect 1056 455 1122 527
rect 1224 455 1291 527
rect 1471 455 1537 527
rect 111 387 327 421
rect 111 372 155 387
rect 31 173 359 181
rect 31 159 626 173
rect 31 139 767 159
rect 31 125 248 139
rect 355 125 767 139
rect 801 127 1234 163
rect 31 107 71 125
rect 105 17 171 89
rect 205 85 248 125
rect 293 17 327 105
rect 721 91 767 125
rect 449 17 515 89
rect 621 17 687 89
rect 721 51 984 91
rect 1502 96 1536 119
rect 1396 62 1536 96
rect 0 -17 1564 17
<< metal1 >>
rect 0 496 1564 592
rect 0 -48 1564 48
<< obsm1 >>
rect 202 116 260 125
rect 1490 116 1548 125
rect 202 88 1548 116
rect 202 79 260 88
rect 1490 79 1548 88
<< labels >>
rlabel locali s 670 199 726 303 6 A1
port 1 nsew signal input
rlabel locali s 80 215 282 266 6 A1
port 1 nsew signal input
rlabel locali s 193 266 282 303 6 A1
port 1 nsew signal input
rlabel locali s 193 303 726 337 6 A1
port 1 nsew signal input
rlabel locali s 341 215 636 269 6 A2
port 2 nsew signal input
rlabel locali s 1366 199 1400 303 6 B1
port 3 nsew signal input
rlabel locali s 760 199 995 282 6 B1
port 3 nsew signal input
rlabel locali s 852 282 995 303 6 B1
port 3 nsew signal input
rlabel locali s 852 303 1400 337 6 B1
port 3 nsew signal input
rlabel locali s 1074 215 1288 269 6 C1
port 4 nsew signal input
rlabel metal1 s 0 -48 1564 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1 21 1513 203 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 1602 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 1564 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1056 54 1347 90 6 Y
port 9 nsew signal output
rlabel locali s 1313 90 1347 131 6 Y
port 9 nsew signal output
rlabel locali s 1313 131 1470 165 6 Y
port 9 nsew signal output
rlabel locali s 1434 165 1470 268 6 Y
port 9 nsew signal output
rlabel locali s 1434 268 1536 371 6 Y
port 9 nsew signal output
rlabel locali s 361 371 1536 405 6 Y
port 9 nsew signal output
rlabel locali s 809 405 1536 421 6 Y
port 9 nsew signal output
rlabel locali s 361 405 694 421 6 Y
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1564 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 793882
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 783862
<< end >>
