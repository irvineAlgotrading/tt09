magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< pwell >>
rect -79 -26 879 110
<< mvnmos >>
rect 0 0 800 84
<< mvndiff >>
rect -53 46 0 84
rect -53 12 -45 46
rect -11 12 0 46
rect -53 0 0 12
rect 800 46 853 84
rect 800 12 811 46
rect 845 12 853 46
rect 800 0 853 12
<< mvndiffc >>
rect -45 12 -11 46
rect 811 12 845 46
<< poly >>
rect 0 84 800 110
rect 0 -26 800 0
<< locali >>
rect -45 46 -11 62
rect -45 -4 -11 12
rect 811 46 845 62
rect 811 -4 845 12
use hvDFL1sd_CDNS_52468879185349  hvDFL1sd_CDNS_52468879185349_0
timestamp 1704896540
transform -1 0 0 0 1 0
box 0 0 1 1
use hvDFL1sd_CDNS_52468879185349  hvDFL1sd_CDNS_52468879185349_1
timestamp 1704896540
transform 1 0 800 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s -28 29 -28 29 0 FreeSans 300 0 0 0 S
flabel comment s 828 29 828 29 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 87731162
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 87730272
<< end >>
