magic
tech sky130B
timestamp 1704896540
<< metal1 >>
rect 0 0 3 58
rect 573 0 576 58
<< via1 >>
rect 3 0 573 58
<< metal2 >>
rect 0 0 3 58
rect 573 0 576 58
<< properties >>
string GDS_END 78967556
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 78965120
<< end >>
