magic
tech sky130B
timestamp 1704896540
<< metal1 >>
rect 0 0 3 58
rect 765 0 768 58
<< via1 >>
rect 3 0 765 58
<< metal2 >>
rect 0 0 3 58
rect 765 0 768 58
<< properties >>
string GDS_END 88497828
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 88494624
<< end >>
