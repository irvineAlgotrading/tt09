magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< pwell >>
rect -76 -26 199 166
<< mvnmos >>
rect 0 0 120 140
<< mvndiff >>
rect -50 0 0 140
rect 120 114 173 140
rect 120 80 131 114
rect 165 80 173 114
rect 120 46 173 80
rect 120 12 131 46
rect 165 12 173 46
rect 120 0 173 12
<< mvndiffc >>
rect 131 80 165 114
rect 131 12 165 46
<< poly >>
rect 0 140 120 166
rect 0 -26 120 0
<< locali >>
rect 131 114 165 130
rect 131 46 165 80
rect 131 -4 165 12
use DFL1sd_CDNS_5246887918531  DFL1sd_CDNS_5246887918531_0
timestamp 1704896540
transform 1 0 120 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s -25 70 -25 70 0 FreeSans 300 0 0 0 S
flabel comment s 148 63 148 63 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 3492
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 2738
<< end >>
