magic
tech sky130B
magscale 1 2
timestamp 1704896540
use sky130_fd_pr__nfet_01v8__example_55959141808637  sky130_fd_pr__nfet_01v8__example_55959141808637_0
timestamp 1704896540
transform 1 0 1401 0 1 -1273
box -1 0 297 1
use sky130_fd_pr__nfet_01v8__example_55959141808638  sky130_fd_pr__nfet_01v8__example_55959141808638_0
timestamp 1704896540
transform 1 0 1753 0 1 -1273
box -1 0 825 1
use sky130_fd_pr__pfet_01v8__example_55959141808481  sky130_fd_pr__pfet_01v8__example_55959141808481_0
timestamp 1704896540
transform 1 0 2377 0 1 -356
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808481  sky130_fd_pr__pfet_01v8__example_55959141808481_1
timestamp 1704896540
transform 1 0 2533 0 1 -356
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808481  sky130_fd_pr__pfet_01v8__example_55959141808481_2
timestamp 1704896540
transform -1 0 2789 0 1 -356
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808481  sky130_fd_pr__pfet_01v8__example_55959141808481_3
timestamp 1704896540
transform -1 0 2321 0 1 -356
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808630  sky130_fd_pr__pfet_01v8__example_55959141808630_0
timestamp 1704896540
transform 1 0 1192 0 1 -250
box -1 0 801 1
use sky130_fd_pr__pfet_01v8__example_55959141808632  sky130_fd_pr__pfet_01v8__example_55959141808632_0
timestamp 1704896540
transform -1 0 2017 0 1 456
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_55959141808634  sky130_fd_pr__pfet_01v8__example_55959141808634_0
timestamp 1704896540
transform 1 0 2197 0 1 456
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808634  sky130_fd_pr__pfet_01v8__example_55959141808634_1
timestamp 1704896540
transform -1 0 2453 0 1 456
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808635  sky130_fd_pr__pfet_01v8__example_55959141808635_0
timestamp 1704896540
transform 1 0 2699 0 1 456
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_55959141808636  sky130_fd_pr__pfet_01v8__example_55959141808636_0
timestamp 1704896540
transform 1 0 1192 0 1 172
box -1 0 401 1
use sky130_fd_pr__pfet_01v8__example_55959141808636  sky130_fd_pr__pfet_01v8__example_55959141808636_1
timestamp 1704896540
transform -1 0 2504 0 1 172
box -1 0 401 1
use sky130_fd_pr__pfet_01v8__example_55959141808636  sky130_fd_pr__pfet_01v8__example_55959141808636_2
timestamp 1704896540
transform 1 0 1648 0 1 172
box -1 0 401 1
<< properties >>
string GDS_END 21024262
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 20996144
<< end >>
