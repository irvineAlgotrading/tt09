magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -36 679 5808 1471
<< locali >>
rect 0 1397 5772 1431
rect 64 636 98 702
rect 196 652 449 686
rect 547 664 817 698
rect 919 690 1293 724
rect 1518 690 1877 724
rect 2320 690 3001 724
rect 4291 690 4325 724
rect 919 681 953 690
rect 0 -17 5772 17
use sky130_sram_1kbyte_1rw1r_32x256_8_pinv_6  sky130_sram_1kbyte_1rw1r_32x256_8_pinv_6_0
timestamp 1704896540
transform 1 0 368 0 1 0
box -36 -17 404 1471
use sky130_sram_1kbyte_1rw1r_32x256_8_pinv_6  sky130_sram_1kbyte_1rw1r_32x256_8_pinv_6_1
timestamp 1704896540
transform 1 0 0 0 1 0
box -36 -17 404 1471
use sky130_sram_1kbyte_1rw1r_32x256_8_pinv_11  sky130_sram_1kbyte_1rw1r_32x256_8_pinv_11_0
timestamp 1704896540
transform 1 0 736 0 1 0
box -36 -17 512 1471
use sky130_sram_1kbyte_1rw1r_32x256_8_pinv_12  sky130_sram_1kbyte_1rw1r_32x256_8_pinv_12_0
timestamp 1704896540
transform 1 0 1212 0 1 0
box -36 -17 620 1471
use sky130_sram_1kbyte_1rw1r_32x256_8_pinv_13  sky130_sram_1kbyte_1rw1r_32x256_8_pinv_13_0
timestamp 1704896540
transform 1 0 1796 0 1 0
box -36 -17 1160 1471
use sky130_sram_1kbyte_1rw1r_32x256_8_pinv_14  sky130_sram_1kbyte_1rw1r_32x256_8_pinv_14_0
timestamp 1704896540
transform 1 0 2920 0 1 0
box -36 -17 2888 1471
<< labels >>
rlabel locali s 4308 707 4308 707 4 Z
rlabel locali s 81 669 81 669 4 A
rlabel locali s 2886 0 2886 0 4 gnd
rlabel locali s 2886 1414 2886 1414 4 vdd
<< properties >>
string FIXED_BBOX 0 0 5772 1414
string GDS_END 6272022
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_32x256_8.gds
string GDS_START 6270258
<< end >>
