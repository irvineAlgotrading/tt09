magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -66 377 1122 897
<< pwell >>
rect 4 43 998 283
rect -26 -43 1082 43
<< locali >>
rect 112 355 302 411
rect 409 355 647 430
rect 268 319 302 355
rect 683 319 743 367
rect 268 301 743 319
rect 268 285 717 301
rect 793 265 874 485
rect 770 99 874 265
<< obsli1 >>
rect 0 797 1056 831
rect 26 521 76 751
rect 112 557 506 751
rect 542 625 576 751
rect 612 661 944 751
rect 980 625 1030 751
rect 542 591 1030 625
rect 542 557 576 591
rect 612 521 944 555
rect 26 487 646 521
rect 26 319 76 487
rect 26 285 232 319
rect 18 73 136 249
rect 182 99 232 285
rect 910 399 944 521
rect 980 435 1030 591
rect 910 333 976 399
rect 268 73 734 249
rect 910 73 1028 265
rect 0 -17 1056 17
<< metal1 >>
rect 0 791 1056 837
rect 0 689 1056 763
rect 0 51 1056 125
rect 0 -23 1056 23
<< labels >>
rlabel locali s 409 355 647 430 6 A
port 1 nsew signal input
rlabel locali s 268 285 717 301 6 B
port 2 nsew signal input
rlabel locali s 268 301 743 319 6 B
port 2 nsew signal input
rlabel locali s 683 319 743 367 6 B
port 2 nsew signal input
rlabel locali s 268 319 302 355 6 B
port 2 nsew signal input
rlabel locali s 112 355 302 411 6 B
port 2 nsew signal input
rlabel metal1 s 0 51 1056 125 6 VGND
port 3 nsew ground bidirectional
rlabel metal1 s 0 -23 1056 23 8 VNB
port 4 nsew ground bidirectional
rlabel pwell s -26 -43 1082 43 8 VNB
port 4 nsew ground bidirectional
rlabel pwell s 4 43 998 283 6 VNB
port 4 nsew ground bidirectional
rlabel metal1 s 0 791 1056 837 6 VPB
port 5 nsew power bidirectional
rlabel nwell s -66 377 1122 897 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 689 1056 763 6 VPWR
port 6 nsew power bidirectional
rlabel locali s 770 99 874 265 6 X
port 7 nsew signal output
rlabel locali s 793 265 874 485 6 X
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1056 814
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 743414
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 731354
<< end >>
