magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -36 679 1052 1471
<< pwell >>
rect 880 25 982 159
<< psubdiff >>
rect 906 109 956 133
rect 906 75 914 109
rect 948 75 956 109
rect 906 51 956 75
<< nsubdiff >>
rect 906 1339 956 1363
rect 906 1305 914 1339
rect 948 1305 956 1339
rect 906 1281 956 1305
<< psubdiffcont >>
rect 914 75 948 109
<< nsubdiffcont >>
rect 914 1305 948 1339
<< poly >>
rect 114 724 144 907
rect 48 708 144 724
rect 48 674 64 708
rect 98 674 144 708
rect 48 658 144 674
rect 114 443 144 658
<< polycont >>
rect 64 674 98 708
<< locali >>
rect 0 1397 1016 1431
rect 62 1130 96 1397
rect 274 1130 308 1397
rect 490 1130 524 1397
rect 706 1130 740 1397
rect 914 1339 948 1397
rect 914 1289 948 1305
rect 64 708 98 724
rect 64 658 98 674
rect 488 708 522 1096
rect 488 674 539 708
rect 488 286 522 674
rect 62 17 96 186
rect 274 17 308 186
rect 490 17 524 186
rect 706 17 740 186
rect 914 109 948 125
rect 914 17 948 75
rect 0 -17 1016 17
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_16  sky130_sram_2kbyte_1rw1r_32x512_8_contact_16_0
timestamp 1704896540
transform 1 0 48 0 1 658
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_28  sky130_sram_2kbyte_1rw1r_32x512_8_contact_28_0
timestamp 1704896540
transform 1 0 906 0 1 1281
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_29  sky130_sram_2kbyte_1rw1r_32x512_8_contact_29_0
timestamp 1704896540
transform 1 0 906 0 1 51
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_nmos_m7_w1_680_sli_dli_da_p  sky130_sram_2kbyte_1rw1r_32x512_8_nmos_m7_w1_680_sli_dli_da_p_0
timestamp 1704896540
transform 1 0 54 0 1 51
box -26 -26 824 392
use sky130_sram_2kbyte_1rw1r_32x512_8_pmos_m7_w2_000_sli_dli_da_p  sky130_sram_2kbyte_1rw1r_32x512_8_pmos_m7_w2_000_sli_dli_da_p_0
timestamp 1704896540
transform 1 0 54 0 1 963
box -59 -56 857 454
<< labels >>
rlabel locali s 81 691 81 691 4 A
rlabel locali s 522 691 522 691 4 Z
rlabel locali s 508 0 508 0 4 gnd
rlabel locali s 508 1414 508 1414 4 vdd
<< properties >>
string FIXED_BBOX 0 0 1016 1414
string GDS_END 129572
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_2kbyte_1rw1r_32x512_8.gds
string GDS_START 127318
<< end >>
