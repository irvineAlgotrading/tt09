magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< pwell >>
rect -76 -26 964 226
<< mvnnmos >>
rect 0 0 180 200
rect 236 0 416 200
rect 472 0 652 200
rect 708 0 888 200
<< mvndiff >>
rect -50 0 0 200
rect 888 0 938 200
<< poly >>
rect 0 200 180 226
rect 0 -26 180 0
rect 236 200 416 226
rect 236 -26 416 0
rect 472 200 652 226
rect 472 -26 652 0
rect 708 200 888 226
rect 708 -26 888 0
<< metal1 >>
rect -51 -16 -5 186
rect 185 -16 231 186
rect 421 -16 467 186
rect 657 -16 703 186
rect 893 -16 939 186
use hvDFM1sd2_CDNS_52468879185104  hvDFM1sd2_CDNS_52468879185104_0
timestamp 1704896540
transform 1 0 652 0 1 0
box -26 -26 82 226
use hvDFM1sd2_CDNS_52468879185104  hvDFM1sd2_CDNS_52468879185104_1
timestamp 1704896540
transform 1 0 416 0 1 0
box -26 -26 82 226
use hvDFM1sd2_CDNS_52468879185104  hvDFM1sd2_CDNS_52468879185104_2
timestamp 1704896540
transform 1 0 180 0 1 0
box -26 -26 82 226
use hvDFM1sd_CDNS_52468879185147  hvDFM1sd_CDNS_52468879185147_0
timestamp 1704896540
transform -1 0 0 0 1 0
box -26 -26 79 226
use hvDFM1sd_CDNS_52468879185147  hvDFM1sd_CDNS_52468879185147_1
timestamp 1704896540
transform 1 0 888 0 1 0
box -26 -26 79 226
<< labels >>
flabel comment s -28 85 -28 85 0 FreeSans 300 0 0 0 S
flabel comment s 208 85 208 85 0 FreeSans 300 0 0 0 D
flabel comment s 444 85 444 85 0 FreeSans 300 0 0 0 S
flabel comment s 680 85 680 85 0 FreeSans 300 0 0 0 D
flabel comment s 916 85 916 85 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 86862302
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86859848
<< end >>
