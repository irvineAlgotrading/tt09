magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect 21 1931 731 1967
<< poly >>
rect 316 1947 612 1967
rect 316 1913 345 1947
rect 379 1913 413 1947
rect 447 1913 481 1947
rect 515 1913 549 1947
rect 583 1913 612 1947
rect 316 1891 612 1913
rect 115 803 260 839
rect 115 769 135 803
rect 169 769 203 803
rect 237 769 260 803
rect 115 728 260 769
rect 336 807 673 839
rect 336 773 551 807
rect 585 773 619 807
rect 653 773 673 807
rect 336 728 673 773
rect 138 57 280 76
rect 138 23 158 57
rect 192 23 226 57
rect 260 23 280 57
rect 138 7 280 23
rect 336 57 480 76
rect 336 23 358 57
rect 392 23 426 57
rect 460 23 480 57
rect 336 7 480 23
<< polycont >>
rect 345 1913 379 1947
rect 413 1913 447 1947
rect 481 1913 515 1947
rect 549 1913 583 1947
rect 135 769 169 803
rect 203 769 237 803
rect 551 773 585 807
rect 619 773 653 807
rect 158 23 192 57
rect 226 23 260 57
rect 358 23 392 57
rect 426 23 460 57
<< locali >>
rect 329 1913 345 1947
rect 379 1913 413 1947
rect 447 1913 481 1947
rect 515 1913 549 1947
rect 583 1913 599 1947
rect 129 1221 167 1255
rect 443 1221 481 1255
rect 271 1029 305 1067
rect 271 957 305 995
rect 623 1029 657 1067
rect 623 957 657 995
rect 447 803 481 919
rect 119 769 135 803
rect 169 769 203 803
rect 237 769 253 803
rect 447 769 501 803
rect 535 773 551 807
rect 585 773 619 807
rect 653 773 669 807
rect 467 638 501 769
rect 115 496 149 534
rect 115 424 149 462
rect 142 23 158 57
rect 192 23 226 57
rect 260 23 276 57
rect 342 23 358 57
rect 392 23 426 57
rect 460 23 476 57
<< viali >>
rect 95 1221 129 1255
rect 167 1221 201 1255
rect 409 1221 443 1255
rect 481 1221 515 1255
rect 271 1067 305 1101
rect 271 995 305 1029
rect 271 923 305 957
rect 623 1067 657 1101
rect 623 995 657 1029
rect 623 923 657 957
rect 115 534 149 568
rect 115 462 149 496
rect 115 390 149 424
<< metal1 >>
rect 83 1255 527 1261
rect 83 1221 95 1255
rect 129 1221 167 1255
rect 201 1221 409 1255
rect 443 1221 481 1255
rect 515 1221 527 1255
rect 83 1215 527 1221
rect 21 1101 731 1107
rect 21 1067 271 1101
rect 305 1067 623 1101
rect 657 1067 731 1101
rect 21 1029 731 1067
rect 21 995 271 1029
rect 305 995 623 1029
rect 657 995 731 1029
rect 21 957 731 995
rect 21 923 271 957
rect 305 923 623 957
rect 657 923 731 957
rect 21 905 731 923
rect 21 568 731 581
rect 21 534 115 568
rect 149 534 731 568
rect 21 496 731 534
rect 21 462 115 496
rect 149 462 731 496
rect 21 424 731 462
rect 21 390 115 424
rect 149 390 731 424
rect 21 379 731 390
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1704896540
transform -1 0 515 0 -1 1255
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1704896540
transform -1 0 201 0 -1 1255
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_0
timestamp 1704896540
transform 1 0 623 0 -1 1101
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_1
timestamp 1704896540
transform 1 0 271 0 -1 1101
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_2
timestamp 1704896540
transform 1 0 115 0 1 390
box 0 0 1 1
use nfet_CDNS_52468879185310  nfet_CDNS_52468879185310_0
timestamp 1704896540
transform 1 0 160 0 1 102
box -79 -26 199 626
use nfet_CDNS_52468879185310  nfet_CDNS_52468879185310_1
timestamp 1704896540
transform 1 0 336 0 1 102
box -79 -26 199 626
use pfet_CDNS_52468879185312  pfet_CDNS_52468879185312_0
timestamp 1704896540
transform -1 0 612 0 -1 1865
box -119 -66 415 1066
use pfet_CDNS_52468879185313  pfet_CDNS_52468879185313_0
timestamp 1704896540
transform -1 0 260 0 -1 1865
box -119 -66 239 1066
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_0
timestamp 1704896540
transform 0 1 535 1 0 757
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_1
timestamp 1704896540
transform 0 -1 276 1 0 7
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_2
timestamp 1704896540
transform 0 -1 476 1 0 7
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_3
timestamp 1704896540
transform 0 -1 253 1 0 753
box 0 0 1 1
use PYL1_CDNS_52468879185309  PYL1_CDNS_52468879185309_0
timestamp 1704896540
transform 0 1 329 1 0 1897
box 0 0 1 1
<< labels >>
flabel metal1 s 487 1215 527 1261 3 FreeSans 300 0 0 0 pu_h_n
port 1 nsew
flabel metal1 s 694 905 731 1107 6 FreeSans 300 180 0 0 vcc_io
port 2 nsew
flabel metal1 s 21 905 58 1107 7 FreeSans 300 0 0 0 vcc_io
port 2 nsew
flabel metal1 s 689 379 731 581 7 FreeSans 300 180 0 0 vgnd_io
port 3 nsew
flabel metal1 s 21 379 63 581 7 FreeSans 300 0 0 0 vgnd_io
port 3 nsew
flabel metal1 s 83 1215 123 1261 3 FreeSans 300 180 0 0 pu_h_n
port 1 nsew
flabel locali s 147 769 188 803 8 FreeSans 300 0 0 0 puen_h
port 5 nsew
flabel locali s 541 773 575 807 2 FreeSans 300 0 0 0 drvhi_h
port 6 nsew
<< properties >>
string GDS_END 87978790
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 87975866
<< end >>
