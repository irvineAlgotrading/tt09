magic
tech sky130B
magscale 1 2
timestamp 1704896540
use sky130_fd_pr__hvdfm1sd__example_55959141808237  sky130_fd_pr__hvdfm1sd__example_55959141808237_0
timestamp 1704896540
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd__example_55959141808237  sky130_fd_pr__hvdfm1sd__example_55959141808237_1
timestamp 1704896540
transform 1 0 180 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 68114782
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 68113792
<< end >>
