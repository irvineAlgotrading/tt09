magic
tech sky130B
magscale 1 2
timestamp 1704896540
use sky130_fd_io__refgen_compl_switch  sky130_fd_io__refgen_compl_switch_0
timestamp 1704896540
transform -1 0 10851 0 1 11
box 43 4 1501 2827
use sky130_fd_io__refgen_compl_switch  sky130_fd_io__refgen_compl_switch_1
timestamp 1704896540
transform -1 0 5447 0 1 11
box 43 4 1501 2827
use sky130_fd_io__refgen_compl_switch  sky130_fd_io__refgen_compl_switch_2
timestamp 1704896540
transform -1 0 8149 0 1 11
box 43 4 1501 2827
use sky130_fd_io__refgen_compl_switch  sky130_fd_io__refgen_compl_switch_3
timestamp 1704896540
transform -1 0 2745 0 1 11
box 43 4 1501 2827
use sky130_fd_io__refgen_compl_switch  sky130_fd_io__refgen_compl_switch_4
timestamp 1704896540
transform 1 0 5361 0 1 11
box 43 4 1501 2827
use sky130_fd_io__refgen_compl_switch  sky130_fd_io__refgen_compl_switch_5
timestamp 1704896540
transform 1 0 8063 0 1 11
box 43 4 1501 2827
use sky130_fd_io__refgen_compl_switch  sky130_fd_io__refgen_compl_switch_6
timestamp 1704896540
transform 1 0 2659 0 1 11
box 43 4 1501 2827
use sky130_fd_io__refgen_compl_switch  sky130_fd_io__refgen_compl_switch_7
timestamp 1704896540
transform 1 0 -43 0 1 11
box 43 4 1501 2827
<< properties >>
string GDS_END 80607104
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 80606564
<< end >>
