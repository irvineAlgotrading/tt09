magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< locali >>
rect 248 961 394 980
rect 248 927 262 961
rect 296 927 346 961
rect 380 927 394 961
rect 248 889 394 927
rect 248 855 262 889
rect 296 855 346 889
rect 380 855 394 889
rect 248 841 394 855
rect 248 125 394 139
rect 248 91 262 125
rect 296 91 346 125
rect 380 91 394 125
rect 248 53 394 91
rect 248 19 262 53
rect 296 19 346 53
rect 380 19 394 53
rect 248 0 394 19
<< viali >>
rect 262 927 296 961
rect 346 927 380 961
rect 262 855 296 889
rect 346 855 380 889
rect 262 91 296 125
rect 346 91 380 125
rect 262 19 296 53
rect 346 19 380 53
<< obsli1 >>
rect 120 817 186 883
rect 456 817 522 883
rect 120 795 160 817
rect 482 795 522 817
rect 41 759 160 795
rect 41 725 60 759
rect 94 725 160 759
rect 41 687 160 725
rect 41 653 60 687
rect 94 653 160 687
rect 41 615 160 653
rect 41 581 60 615
rect 94 581 160 615
rect 41 543 160 581
rect 41 509 60 543
rect 94 509 160 543
rect 41 471 160 509
rect 41 437 60 471
rect 94 437 160 471
rect 41 399 160 437
rect 41 365 60 399
rect 94 365 160 399
rect 41 327 160 365
rect 41 293 60 327
rect 94 293 160 327
rect 41 255 160 293
rect 41 221 60 255
rect 94 221 160 255
rect 41 185 160 221
rect 212 185 246 795
rect 304 185 338 795
rect 396 185 430 795
rect 482 759 601 795
rect 482 725 548 759
rect 582 725 601 759
rect 482 687 601 725
rect 482 653 548 687
rect 582 653 601 687
rect 482 615 601 653
rect 482 581 548 615
rect 582 581 601 615
rect 482 543 601 581
rect 482 509 548 543
rect 582 509 601 543
rect 482 471 601 509
rect 482 437 548 471
rect 582 437 601 471
rect 482 399 601 437
rect 482 365 548 399
rect 582 365 601 399
rect 482 327 601 365
rect 482 293 548 327
rect 582 293 601 327
rect 482 255 601 293
rect 482 221 548 255
rect 582 221 601 255
rect 482 185 601 221
rect 120 163 160 185
rect 482 163 522 185
rect 120 97 186 163
rect 456 97 522 163
<< obsli1c >>
rect 60 725 94 759
rect 60 653 94 687
rect 60 581 94 615
rect 60 509 94 543
rect 60 437 94 471
rect 60 365 94 399
rect 60 293 94 327
rect 60 221 94 255
rect 548 725 582 759
rect 548 653 582 687
rect 548 581 582 615
rect 548 509 582 543
rect 548 437 582 471
rect 548 365 582 399
rect 548 293 582 327
rect 548 221 582 255
<< metal1 >>
rect 250 961 392 980
rect 250 927 262 961
rect 296 927 346 961
rect 380 927 392 961
rect 250 889 392 927
rect 250 855 262 889
rect 296 855 346 889
rect 380 855 392 889
rect 250 843 392 855
rect 41 759 100 771
rect 41 725 60 759
rect 94 725 100 759
rect 41 687 100 725
rect 41 653 60 687
rect 94 653 100 687
rect 41 615 100 653
rect 41 581 60 615
rect 94 581 100 615
rect 41 543 100 581
rect 41 509 60 543
rect 94 509 100 543
rect 41 471 100 509
rect 41 437 60 471
rect 94 437 100 471
rect 41 399 100 437
rect 41 365 60 399
rect 94 365 100 399
rect 41 327 100 365
rect 41 293 60 327
rect 94 293 100 327
rect 41 255 100 293
rect 41 221 60 255
rect 94 221 100 255
rect 41 209 100 221
rect 542 759 601 771
rect 542 725 548 759
rect 582 725 601 759
rect 542 687 601 725
rect 542 653 548 687
rect 582 653 601 687
rect 542 615 601 653
rect 542 581 548 615
rect 582 581 601 615
rect 542 543 601 581
rect 542 509 548 543
rect 582 509 601 543
rect 542 471 601 509
rect 542 437 548 471
rect 582 437 601 471
rect 542 399 601 437
rect 542 365 548 399
rect 582 365 601 399
rect 542 327 601 365
rect 542 293 548 327
rect 582 293 601 327
rect 542 255 601 293
rect 542 221 548 255
rect 582 221 601 255
rect 542 209 601 221
rect 250 125 392 137
rect 250 91 262 125
rect 296 91 346 125
rect 380 91 392 125
rect 250 53 392 91
rect 250 19 262 53
rect 296 19 346 53
rect 380 19 392 53
rect 250 0 392 19
<< obsm1 >>
rect 203 209 255 771
rect 295 209 347 771
rect 387 209 439 771
<< metal2 >>
rect 14 515 628 771
rect 14 209 628 465
<< labels >>
rlabel metal2 s 14 515 628 771 6 DRAIN
port 1 nsew
rlabel viali s 346 927 380 961 6 GATE
port 2 nsew
rlabel viali s 346 855 380 889 6 GATE
port 2 nsew
rlabel viali s 346 91 380 125 6 GATE
port 2 nsew
rlabel viali s 346 19 380 53 6 GATE
port 2 nsew
rlabel viali s 262 927 296 961 6 GATE
port 2 nsew
rlabel viali s 262 855 296 889 6 GATE
port 2 nsew
rlabel viali s 262 91 296 125 6 GATE
port 2 nsew
rlabel viali s 262 19 296 53 6 GATE
port 2 nsew
rlabel locali s 248 841 394 980 6 GATE
port 2 nsew
rlabel locali s 248 0 394 139 6 GATE
port 2 nsew
rlabel metal1 s 250 843 392 980 6 GATE
port 2 nsew
rlabel metal1 s 250 0 392 137 6 GATE
port 2 nsew
rlabel metal2 s 14 209 628 465 6 SOURCE
port 3 nsew
rlabel metal1 s 41 209 100 771 6 SUBSTRATE
port 4 nsew
rlabel metal1 s 542 209 601 771 6 SUBSTRATE
port 4 nsew
<< properties >>
string FIXED_BBOX 14 0 628 980
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 6210800
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 6196208
<< end >>
