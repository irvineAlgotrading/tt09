magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< pwell >>
rect -161 398 -75 434
rect -161 -26 91 398
rect 1748 -26 1818 398
rect 3475 -26 3595 398
rect -161 -62 -75 -26
<< mvndiff >>
rect -3 334 65 372
rect -3 300 5 334
rect 39 300 65 334
rect -3 288 65 300
rect 1774 288 1792 372
rect 3501 334 3569 372
rect 3501 300 3527 334
rect 3561 300 3569 334
rect 3501 288 3569 300
rect -3 190 65 228
rect -3 156 5 190
rect 39 156 65 190
rect -3 144 65 156
rect 1774 144 1792 228
rect 3501 190 3569 228
rect 3501 156 3527 190
rect 3561 156 3569 190
rect 3501 144 3569 156
rect -3 46 65 84
rect -3 12 5 46
rect 39 12 65 46
rect -3 0 65 12
rect 1774 0 1792 84
rect 3501 46 3569 84
rect 3501 12 3527 46
rect 3561 12 3569 46
rect 3501 0 3569 12
<< mvndiffc >>
rect 5 300 39 334
rect 3527 300 3561 334
rect 5 156 39 190
rect 3527 156 3561 190
rect 5 12 39 46
rect 3527 12 3561 46
<< mvpsubdiff >>
rect -135 342 -101 408
rect -135 272 -101 308
rect -135 204 -101 238
rect -135 136 -101 170
rect -135 68 -101 102
rect -135 -36 -101 34
<< mvpsubdiffcont >>
rect -135 308 -101 342
rect -135 238 -101 272
rect -135 170 -101 204
rect -135 102 -101 136
rect -135 34 -101 68
<< poly >>
rect 121 372 1721 398
rect 1845 372 3444 398
rect 121 254 1721 262
rect 1845 254 3445 262
rect 121 110 1721 118
rect 1845 110 3445 118
<< locali >>
rect -135 342 -101 408
rect -135 272 -101 308
rect 5 334 781 350
rect 39 316 781 334
rect 815 316 853 350
rect 887 316 896 350
rect 39 300 896 316
rect 5 284 896 300
rect 946 316 952 350
rect 986 316 1024 350
rect 1058 316 1732 350
rect 946 284 1732 316
rect 1766 284 1800 350
rect 1834 338 2620 350
rect 1834 304 2514 338
rect 2548 304 2586 338
rect 1834 284 2620 304
rect 2670 338 3456 350
rect 2704 304 2742 338
rect 2776 304 3456 338
rect 2670 284 3456 304
rect 3490 334 3561 350
rect 3490 300 3527 334
rect 3490 284 3561 300
rect -135 204 -101 238
rect 3445 206 3561 284
rect -135 136 -101 170
rect -135 68 -101 102
rect -135 -36 -101 34
rect 5 190 781 206
rect 39 172 781 190
rect 815 172 853 206
rect 887 172 896 206
rect 39 156 896 172
rect 5 140 896 156
rect 946 172 952 206
rect 986 172 1024 206
rect 1058 172 1732 206
rect 946 140 1732 172
rect 1766 140 1800 206
rect 1834 194 2620 206
rect 1834 160 2514 194
rect 2548 160 2586 194
rect 1834 140 2620 160
rect 2670 194 3456 206
rect 2704 160 2742 194
rect 2776 160 3456 194
rect 2670 140 3456 160
rect 3490 190 3561 206
rect 3490 156 3527 190
rect 3490 140 3561 156
rect 5 62 121 140
rect 5 46 781 62
rect 39 28 781 46
rect 815 28 853 62
rect 887 28 896 62
rect 39 12 896 28
rect 5 -4 896 12
rect 946 28 952 62
rect 986 28 1024 62
rect 1058 28 1732 62
rect 946 -4 1732 28
rect 1766 -4 1800 62
rect 1834 50 2620 62
rect 1834 16 2514 50
rect 2548 16 2586 50
rect 1834 -4 2620 16
rect 2670 50 3561 62
rect 2704 16 2742 50
rect 2776 46 3561 50
rect 2776 16 3527 46
rect 2670 12 3527 16
rect 2670 -4 3561 12
<< viali >>
rect 781 316 815 350
rect 853 316 887 350
rect 952 316 986 350
rect 1024 316 1058 350
rect 2514 304 2548 338
rect 2586 304 2620 338
rect 2670 304 2704 338
rect 2742 304 2776 338
rect 781 172 815 206
rect 853 172 887 206
rect 952 172 986 206
rect 1024 172 1058 206
rect 2514 160 2548 194
rect 2586 160 2620 194
rect 2670 160 2704 194
rect 2742 160 2776 194
rect 781 28 815 62
rect 853 28 887 62
rect 952 28 986 62
rect 1024 28 1058 62
rect 2514 16 2548 50
rect 2586 16 2620 50
rect 2670 16 2704 50
rect 2742 16 2776 50
<< metal1 >>
rect 769 350 902 356
rect 769 316 781 350
rect 815 316 853 350
rect 887 316 902 350
rect 769 310 902 316
rect 903 311 904 355
rect 932 311 933 355
rect 934 350 1070 356
rect 934 316 952 350
rect 986 316 1024 350
rect 1058 316 1070 350
rect 934 310 1070 316
rect 2508 338 2625 350
rect 2508 304 2514 338
rect 2548 304 2586 338
rect 2620 304 2625 338
rect 2508 292 2625 304
rect 2626 293 2627 349
rect 2663 293 2664 349
rect 2665 338 2782 350
rect 2665 304 2670 338
rect 2704 304 2742 338
rect 2776 304 2782 338
rect 2665 292 2782 304
rect 769 206 902 212
rect 769 172 781 206
rect 815 172 853 206
rect 887 172 902 206
rect 769 166 902 172
rect 903 167 904 211
rect 932 167 933 211
rect 934 206 1070 212
rect 934 172 952 206
rect 986 172 1024 206
rect 1058 172 1070 206
rect 934 166 1070 172
rect 2508 194 2627 206
rect 2508 160 2514 194
rect 2548 160 2586 194
rect 2620 160 2627 194
rect 2508 148 2627 160
rect 2628 149 2629 205
rect 2664 205 2665 206
rect 2664 149 2666 205
rect 2667 194 2782 206
rect 2667 160 2670 194
rect 2704 160 2742 194
rect 2776 160 2782 194
rect 2664 148 2665 149
rect 2667 148 2782 160
rect 769 62 902 68
rect 769 28 781 62
rect 815 28 853 62
rect 887 28 902 62
rect 769 22 902 28
rect 903 23 904 67
rect 932 23 933 67
rect 934 62 1070 68
rect 934 28 952 62
rect 986 28 1024 62
rect 1058 28 1070 62
rect 934 22 1070 28
rect 2508 50 2627 62
rect 2508 16 2514 50
rect 2548 16 2586 50
rect 2620 16 2627 50
rect 2508 4 2627 16
rect 2628 5 2629 61
rect 2664 61 2665 62
rect 2664 5 2666 61
rect 2667 50 2782 62
rect 2667 16 2670 50
rect 2704 16 2742 50
rect 2776 16 2782 50
rect 2664 4 2665 5
rect 2667 4 2782 16
<< rmetal1 >>
rect 902 355 904 356
rect 902 311 903 355
rect 902 310 904 311
rect 932 355 934 356
rect 933 311 934 355
rect 932 310 934 311
rect 2625 349 2627 350
rect 2625 293 2626 349
rect 2625 292 2627 293
rect 2663 349 2665 350
rect 2664 293 2665 349
rect 2663 292 2665 293
rect 902 211 904 212
rect 902 167 903 211
rect 902 166 904 167
rect 932 211 934 212
rect 933 167 934 211
rect 932 166 934 167
rect 2627 205 2629 206
rect 2627 149 2628 205
rect 2627 148 2629 149
rect 2665 205 2667 206
rect 2666 149 2667 205
rect 2665 148 2667 149
rect 902 67 904 68
rect 902 23 903 67
rect 902 22 904 23
rect 932 67 934 68
rect 933 23 934 67
rect 932 22 934 23
rect 2627 61 2629 62
rect 2627 5 2628 61
rect 2627 4 2629 5
rect 2665 61 2667 62
rect 2666 5 2667 61
rect 2665 4 2667 5
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_0
timestamp 1704896540
transform -1 0 47 0 -1 346
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_1
timestamp 1704896540
transform -1 0 47 0 -1 202
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_2
timestamp 1704896540
transform -1 0 47 0 -1 58
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_3
timestamp 1704896540
transform 1 0 3519 0 -1 58
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_4
timestamp 1704896540
transform 1 0 3519 0 -1 202
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_5
timestamp 1704896540
transform 1 0 3519 0 -1 346
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_0
timestamp 1704896540
transform 0 1 2514 -1 0 194
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_1
timestamp 1704896540
transform 0 1 2670 -1 0 194
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_2
timestamp 1704896540
transform 0 1 2514 -1 0 50
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_3
timestamp 1704896540
transform 0 1 2670 -1 0 50
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_4
timestamp 1704896540
transform 0 1 2514 -1 0 338
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_5
timestamp 1704896540
transform 0 1 2670 -1 0 338
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1704896540
transform 1 0 781 0 1 316
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1704896540
transform 1 0 952 0 1 172
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1704896540
transform 1 0 781 0 1 172
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1704896540
transform 1 0 781 0 1 28
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_4
timestamp 1704896540
transform 1 0 952 0 1 28
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_5
timestamp 1704896540
transform 1 0 952 0 1 316
box 0 0 1 1
use nfet_CDNS_524688791851480  nfet_CDNS_524688791851480_0
timestamp 1704896540
transform -1 0 3445 0 1 288
box -82 -26 1679 110
use nfet_CDNS_524688791851480  nfet_CDNS_524688791851480_1
timestamp 1704896540
transform -1 0 3445 0 1 144
box -82 -26 1679 110
use nfet_CDNS_524688791851480  nfet_CDNS_524688791851480_2
timestamp 1704896540
transform -1 0 3445 0 1 0
box -82 -26 1679 110
use nfet_CDNS_524688791851480  nfet_CDNS_524688791851480_3
timestamp 1704896540
transform 1 0 121 0 1 288
box -82 -26 1679 110
use nfet_CDNS_524688791851480  nfet_CDNS_524688791851480_4
timestamp 1704896540
transform 1 0 121 0 1 144
box -82 -26 1679 110
use nfet_CDNS_524688791851480  nfet_CDNS_524688791851480_5
timestamp 1704896540
transform 1 0 121 0 1 0
box -82 -26 1679 110
use sky130_fd_io__tk_em1o_b_CDNS_524688791851479  sky130_fd_io__tk_em1o_b_CDNS_524688791851479_0
timestamp 1704896540
transform 1 0 850 0 1 310
box 0 0 1 1
use sky130_fd_io__tk_em1o_b_CDNS_524688791851479  sky130_fd_io__tk_em1o_b_CDNS_524688791851479_1
timestamp 1704896540
transform 1 0 850 0 1 166
box 0 0 1 1
use sky130_fd_io__tk_em1o_b_CDNS_524688791851479  sky130_fd_io__tk_em1o_b_CDNS_524688791851479_2
timestamp 1704896540
transform 1 0 850 0 1 22
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_0
timestamp 1704896540
transform -1 0 2719 0 1 148
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_1
timestamp 1704896540
transform -1 0 2719 0 1 4
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_2
timestamp 1704896540
transform 1 0 2573 0 1 292
box 0 0 1 1
<< labels >>
flabel locali s -135 340 -101 356 0 FreeSans 200 0 0 0 vgnd
port 2 nsew
flabel locali s 3445 -4 3490 62 0 FreeSans 200 0 0 0 out
port 3 nsew
flabel locali s 58 284 121 350 0 FreeSans 200 0 0 0 vgnd
port 2 nsew
flabel poly s 121 372 1721 398 0 FreeSans 200 0 0 0 en
port 5 nsew
flabel poly s 1845 372 3444 398 0 FreeSans 200 0 0 0 en
port 5 nsew
<< properties >>
string GDS_END 88567270
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 88561466
<< end >>
