magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -77 660 1861 1066
<< pwell >>
rect -67 0 1851 86
<< psubdiff >>
rect -41 26 -17 60
rect 17 26 63 60
rect 97 26 134 60
rect 168 26 205 60
rect 239 26 276 60
rect 310 26 347 60
rect 381 26 418 60
rect 452 26 489 60
rect 523 26 560 60
rect 594 26 631 60
rect 665 26 702 60
rect 736 26 773 60
rect 807 26 844 60
rect 878 26 915 60
rect 949 26 985 60
rect 1019 26 1055 60
rect 1089 26 1125 60
rect 1159 26 1195 60
rect 1229 26 1265 60
rect 1299 26 1335 60
rect 1369 26 1405 60
rect 1439 26 1475 60
rect 1509 26 1545 60
rect 1579 26 1615 60
rect 1649 26 1685 60
rect 1719 26 1767 60
rect 1801 26 1825 60
<< nsubdiff >>
rect -41 996 -17 1030
rect 17 996 75 1030
rect 109 996 145 1030
rect 179 996 215 1030
rect 249 996 285 1030
rect 319 996 355 1030
rect 389 996 425 1030
rect 459 996 495 1030
rect 529 996 565 1030
rect 599 996 635 1030
rect 669 996 705 1030
rect 739 996 775 1030
rect 809 996 845 1030
rect 879 996 915 1030
rect 949 996 985 1030
rect 1019 996 1055 1030
rect 1089 996 1125 1030
rect 1159 996 1194 1030
rect 1228 996 1263 1030
rect 1297 996 1332 1030
rect 1366 996 1401 1030
rect 1435 996 1470 1030
rect 1504 996 1539 1030
rect 1573 996 1608 1030
rect 1642 996 1677 1030
rect 1711 996 1767 1030
rect 1801 996 1825 1030
rect 879 948 913 996
rect 879 851 913 914
rect 879 754 913 817
rect 879 696 913 720
<< psubdiffcont >>
rect -17 26 17 60
rect 63 26 97 60
rect 134 26 168 60
rect 205 26 239 60
rect 276 26 310 60
rect 347 26 381 60
rect 418 26 452 60
rect 489 26 523 60
rect 560 26 594 60
rect 631 26 665 60
rect 702 26 736 60
rect 773 26 807 60
rect 844 26 878 60
rect 915 26 949 60
rect 985 26 1019 60
rect 1055 26 1089 60
rect 1125 26 1159 60
rect 1195 26 1229 60
rect 1265 26 1299 60
rect 1335 26 1369 60
rect 1405 26 1439 60
rect 1475 26 1509 60
rect 1545 26 1579 60
rect 1615 26 1649 60
rect 1685 26 1719 60
rect 1767 26 1801 60
<< nsubdiffcont >>
rect -17 996 17 1030
rect 75 996 109 1030
rect 145 996 179 1030
rect 215 996 249 1030
rect 285 996 319 1030
rect 355 996 389 1030
rect 425 996 459 1030
rect 495 996 529 1030
rect 565 996 599 1030
rect 635 996 669 1030
rect 705 996 739 1030
rect 775 996 809 1030
rect 845 996 879 1030
rect 915 996 949 1030
rect 985 996 1019 1030
rect 1055 996 1089 1030
rect 1125 996 1159 1030
rect 1194 996 1228 1030
rect 1263 996 1297 1030
rect 1332 996 1366 1030
rect 1401 996 1435 1030
rect 1470 996 1504 1030
rect 1539 996 1573 1030
rect 1608 996 1642 1030
rect 1677 996 1711 1030
rect 1767 996 1801 1030
rect 879 914 913 948
rect 879 817 913 851
rect 879 720 913 754
<< poly >>
rect 28 664 228 671
rect 284 664 484 671
rect 540 664 740 670
rect 1044 664 1244 671
rect 1556 670 1756 671
rect 1300 664 1756 670
rect 28 648 953 664
rect 28 614 323 648
rect 357 614 391 648
rect 425 614 459 648
rect 493 614 527 648
rect 561 614 595 648
rect 629 614 663 648
rect 697 614 835 648
rect 869 614 903 648
rect 937 614 953 648
rect 28 598 953 614
rect 1044 648 1756 664
rect 1044 614 1087 648
rect 1121 614 1155 648
rect 1189 614 1223 648
rect 1257 614 1291 648
rect 1325 614 1359 648
rect 1393 614 1427 648
rect 1461 614 1756 648
rect 1044 598 1756 614
rect 28 510 228 598
rect 1556 510 1756 598
rect 408 142 864 158
rect 408 108 449 142
rect 483 108 517 142
rect 551 108 585 142
rect 619 108 653 142
rect 687 108 721 142
rect 755 108 789 142
rect 823 108 864 142
rect 408 92 864 108
rect 920 142 1376 158
rect 920 108 961 142
rect 995 108 1029 142
rect 1063 108 1097 142
rect 1131 108 1165 142
rect 1199 108 1233 142
rect 1267 108 1301 142
rect 1335 108 1376 142
rect 920 92 1376 108
<< polycont >>
rect 323 614 357 648
rect 391 614 425 648
rect 459 614 493 648
rect 527 614 561 648
rect 595 614 629 648
rect 663 614 697 648
rect 835 614 869 648
rect 903 614 937 648
rect 1087 614 1121 648
rect 1155 614 1189 648
rect 1223 614 1257 648
rect 1291 614 1325 648
rect 1359 614 1393 648
rect 1427 614 1461 648
rect 449 108 483 142
rect 517 108 551 142
rect 585 108 619 142
rect 653 108 687 142
rect 721 108 755 142
rect 789 108 823 142
rect 961 108 995 142
rect 1029 108 1063 142
rect 1097 108 1131 142
rect 1165 108 1199 142
rect 1233 108 1267 142
rect 1301 108 1335 142
<< locali >>
rect -33 996 -17 1030
rect 17 996 75 1030
rect 109 996 145 1030
rect 179 996 215 1030
rect 249 996 285 1030
rect 319 996 355 1030
rect 389 996 425 1030
rect 459 996 495 1030
rect 529 996 565 1030
rect 599 996 635 1030
rect 669 996 705 1030
rect 739 996 775 1030
rect 809 996 845 1030
rect 879 996 915 1030
rect 949 996 985 1030
rect 1019 996 1055 1030
rect 1089 996 1125 1030
rect 1159 996 1194 1030
rect 1228 996 1263 1030
rect 1297 996 1332 1030
rect 1366 996 1401 1030
rect 1435 996 1470 1030
rect 1504 996 1539 1030
rect 1573 996 1608 1030
rect 1642 996 1677 1030
rect 1711 996 1767 1030
rect 1801 996 1817 1030
rect 879 948 913 996
rect -17 790 17 824
rect 495 790 529 824
rect 751 788 785 900
rect 879 851 913 914
rect 751 754 811 788
rect 239 482 273 743
rect 751 716 845 754
rect 751 682 811 716
rect 879 754 913 817
rect 1255 790 1289 824
rect 1767 790 1801 824
rect 879 696 913 720
rect 1067 716 1101 754
rect 307 614 323 648
rect 357 614 391 648
rect 425 614 459 648
rect 493 614 527 648
rect 561 614 595 648
rect 629 614 663 648
rect 697 614 713 648
rect 751 488 785 682
rect 999 648 1033 698
rect 819 614 835 648
rect 869 614 903 648
rect 937 614 1033 648
rect 1067 648 1101 682
rect 1067 614 1087 648
rect 1121 614 1155 648
rect 1189 614 1223 648
rect 1257 614 1291 648
rect 1325 614 1359 648
rect 1393 614 1427 648
rect 1461 614 1477 648
rect 639 454 785 488
rect 999 488 1033 614
rect 999 454 1145 488
rect 1511 482 1545 698
rect -17 370 17 404
rect 363 370 397 404
rect 875 370 909 404
rect 1387 370 1421 404
rect 1767 370 1801 404
rect 433 108 449 142
rect 483 108 517 142
rect 551 108 585 142
rect 619 108 653 142
rect 687 108 721 142
rect 755 108 789 142
rect 823 108 839 142
rect 945 108 961 142
rect 995 108 1029 142
rect 1063 108 1097 142
rect 1131 108 1165 142
rect 1199 108 1233 142
rect 1267 108 1301 142
rect 1335 108 1351 142
rect -33 26 -17 60
rect 17 26 63 60
rect 97 26 134 60
rect 168 26 205 60
rect 239 26 276 60
rect 310 26 347 60
rect 381 26 418 60
rect 452 26 489 60
rect 523 26 560 60
rect 594 26 631 60
rect 665 26 702 60
rect 736 26 773 60
rect 807 26 844 60
rect 878 26 915 60
rect 949 26 985 60
rect 1019 26 1055 60
rect 1089 26 1125 60
rect 1159 26 1195 60
rect 1229 26 1265 60
rect 1299 26 1335 60
rect 1369 26 1405 60
rect 1439 26 1475 60
rect 1509 26 1545 60
rect 1579 26 1615 60
rect 1649 26 1685 60
rect 1719 26 1767 60
rect 1801 26 1817 60
<< viali >>
rect 811 754 845 788
rect 811 682 845 716
rect 1067 754 1101 788
rect 1067 682 1101 716
<< metal1 >>
rect 805 788 1107 800
rect 805 754 811 788
rect 845 754 1067 788
rect 1101 754 1107 788
rect 805 716 1107 754
rect 805 682 811 716
rect 845 682 1067 716
rect 1101 682 1107 716
rect 805 670 1107 682
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1704896540
transform 0 -1 1101 1 0 682
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1704896540
transform 0 -1 845 1 0 682
box 0 0 1 1
use nfet_CDNS_524688791851172  nfet_CDNS_524688791851172_0
timestamp 1704896540
transform -1 0 1756 0 1 284
box -79 -26 279 226
use nfet_CDNS_524688791851172  nfet_CDNS_524688791851172_1
timestamp 1704896540
transform 1 0 28 0 1 284
box -79 -26 279 226
use nfet_CDNS_524688791851605  nfet_CDNS_524688791851605_0
timestamp 1704896540
transform 1 0 408 0 -1 484
box -79 -26 1047 326
use pfet_CDNS_524688791851170  pfet_CDNS_524688791851170_0
timestamp 1704896540
transform -1 0 1244 0 1 696
box -89 -36 289 236
use pfet_CDNS_524688791851170  pfet_CDNS_524688791851170_1
timestamp 1704896540
transform 1 0 540 0 1 696
box -89 -36 289 236
use pfet_CDNS_524688791851171  pfet_CDNS_524688791851171_0
timestamp 1704896540
transform 1 0 28 0 1 696
box -89 -36 545 236
use pfet_CDNS_524688791851171  pfet_CDNS_524688791851171_1
timestamp 1704896540
transform 1 0 1300 0 1 696
box -89 -36 545 236
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_0
timestamp 1704896540
transform 0 1 819 1 0 598
box 0 0 1 1
use PYL1_CDNS_52468879185327  PYL1_CDNS_52468879185327_0
timestamp 1704896540
transform 0 -1 1477 -1 0 664
box 0 0 1 1
use PYL1_CDNS_52468879185327  PYL1_CDNS_52468879185327_1
timestamp 1704896540
transform 0 1 433 1 0 92
box 0 0 1 1
use PYL1_CDNS_52468879185327  PYL1_CDNS_52468879185327_2
timestamp 1704896540
transform 0 1 945 1 0 92
box 0 0 1 1
use PYL1_CDNS_52468879185327  PYL1_CDNS_52468879185327_3
timestamp 1704896540
transform 0 -1 713 1 0 598
box 0 0 1 1
<< labels >>
flabel comment s 252 593 252 593 0 FreeSans 200 0 0 0 out_c
flabel comment s 1150 89 1150 89 0 FreeSans 200 0 0 0 in_c
flabel comment s 1531 593 1531 593 0 FreeSans 200 0 0 0 out_t
flabel comment s 640 89 640 89 0 FreeSans 200 0 0 0 in_t
flabel locali s 1387 370 1421 404 0 FreeSans 200 0 0 0 vgnd
port 2 nsew
flabel locali s 875 370 909 404 0 FreeSans 200 0 0 0 vgnd
port 2 nsew
flabel locali s -17 790 17 824 0 FreeSans 200 0 0 0 vpwr
port 3 nsew
flabel locali s 495 790 529 824 0 FreeSans 200 0 0 0 vpwr
port 3 nsew
flabel locali s 1255 790 1289 824 0 FreeSans 200 0 0 0 vpwr
port 3 nsew
flabel locali s 1767 790 1801 824 0 FreeSans 200 0 0 0 vpwr
port 3 nsew
flabel locali s 1767 370 1801 404 0 FreeSans 200 0 0 0 vgnd
port 2 nsew
flabel locali s 619 108 653 142 0 FreeSans 200 0 0 0 in_t
port 4 nsew
flabel locali s 1511 615 1545 648 0 FreeSans 200 0 0 0 out_t
port 5 nsew
flabel locali s -17 370 17 404 0 FreeSans 200 0 0 0 vgnd
port 2 nsew
flabel locali s 239 611 273 641 0 FreeSans 200 0 0 0 out_c
port 6 nsew
flabel locali s 1131 108 1165 142 0 FreeSans 200 0 0 0 in_c
port 7 nsew
flabel locali s 363 370 397 404 0 FreeSans 200 0 0 0 vgnd
port 2 nsew
<< properties >>
string GDS_END 98002872
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 97993380
string path 0.375 25.325 44.275 25.325 
<< end >>
