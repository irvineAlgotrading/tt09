magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect 7676 2269 8992 2779
<< pwell >>
rect 3510 2033 9190 2119
rect 3510 1481 3871 2033
rect 4590 1733 4660 1851
rect 5492 1733 5562 1851
rect 5135 1481 5205 1725
rect 6394 1481 6464 1851
rect 7653 1481 7723 1851
rect 8858 1574 9190 2033
rect 8858 1488 10905 1574
rect 8858 1481 9036 1488
rect 3510 1448 3596 1481
rect -71 1362 3596 1448
rect -71 66 215 1362
rect 5202 1340 5205 1481
rect 5449 1340 5627 1466
rect 5202 693 5627 1340
rect 10614 693 10905 1488
rect 5202 607 10905 693
rect 5202 66 5488 607
rect -71 -20 5488 66
<< mvndiff >>
rect 3719 1935 3845 1951
rect 3719 1901 3731 1935
rect 3765 1901 3799 1935
rect 3833 1901 3845 1935
rect 3719 1885 3845 1901
rect 8884 1935 9010 1951
rect 8884 1901 8896 1935
rect 8930 1901 8964 1935
rect 8998 1901 9010 1935
rect 8884 1885 9010 1901
rect 3719 1809 3845 1825
rect 3719 1775 3731 1809
rect 3765 1775 3799 1809
rect 3833 1775 3845 1809
rect 3719 1759 3845 1775
rect 4616 1759 4634 1825
rect 5518 1759 5536 1825
rect 6420 1759 6438 1825
rect 7679 1759 7697 1825
rect 8884 1809 9010 1825
rect 8884 1775 8896 1809
rect 8930 1775 8964 1809
rect 8998 1775 9010 1809
rect 8884 1759 9010 1775
rect 3719 1683 3845 1699
rect 3719 1649 3731 1683
rect 3765 1649 3799 1683
rect 3833 1649 3845 1683
rect 3719 1633 3845 1649
rect 5161 1633 5179 1699
rect 6420 1633 6438 1699
rect 7679 1633 7697 1699
rect 8884 1683 9010 1699
rect 8884 1649 8896 1683
rect 8930 1649 8964 1683
rect 8998 1649 9010 1683
rect 8884 1633 9010 1649
rect 3719 1557 3845 1573
rect 3719 1523 3731 1557
rect 3765 1523 3799 1557
rect 3833 1523 3845 1557
rect 3719 1507 3845 1523
rect 5161 1507 5179 1573
rect 6420 1507 6438 1573
rect 7679 1507 7697 1573
rect 8884 1557 9010 1573
rect 8884 1523 8896 1557
rect 8930 1523 8964 1557
rect 8998 1523 9010 1557
rect 8884 1507 9010 1523
rect 5475 1424 5601 1440
rect 5475 1390 5487 1424
rect 5521 1390 5555 1424
rect 5589 1390 5601 1424
rect 5475 1374 5601 1390
rect 10640 1424 10766 1440
rect 10640 1390 10652 1424
rect 10686 1390 10720 1424
rect 10754 1390 10766 1424
rect 10640 1374 10766 1390
rect 63 1298 189 1314
rect 63 1264 75 1298
rect 109 1264 143 1298
rect 177 1264 189 1298
rect 63 1248 189 1264
rect 5228 1298 5354 1314
rect 5228 1264 5240 1298
rect 5274 1264 5308 1298
rect 5342 1264 5354 1298
rect 5228 1248 5354 1264
rect 5475 1298 5601 1314
rect 5475 1264 5487 1298
rect 5521 1264 5555 1298
rect 5589 1264 5601 1298
rect 5475 1248 5601 1264
rect 10640 1298 10766 1314
rect 10640 1264 10652 1298
rect 10686 1264 10720 1298
rect 10754 1264 10766 1298
rect 10640 1248 10766 1264
rect 63 1172 189 1188
rect 63 1138 75 1172
rect 109 1138 143 1172
rect 177 1138 189 1172
rect 63 1122 189 1138
rect 5228 1172 5354 1188
rect 5228 1138 5240 1172
rect 5274 1138 5308 1172
rect 5342 1138 5354 1172
rect 5228 1122 5354 1138
rect 5475 1172 5601 1188
rect 5475 1138 5487 1172
rect 5521 1138 5555 1172
rect 5589 1138 5601 1172
rect 5475 1122 5601 1138
rect 10640 1172 10766 1188
rect 10640 1138 10652 1172
rect 10686 1138 10720 1172
rect 10754 1138 10766 1172
rect 10640 1122 10766 1138
rect 63 1046 189 1062
rect 63 1012 75 1046
rect 109 1012 143 1046
rect 177 1012 189 1046
rect 63 996 189 1012
rect 5228 1046 5354 1062
rect 5228 1012 5240 1046
rect 5274 1012 5308 1046
rect 5342 1012 5354 1046
rect 5228 996 5354 1012
rect 5475 1046 5601 1062
rect 5475 1012 5487 1046
rect 5521 1012 5555 1046
rect 5589 1012 5601 1046
rect 5475 996 5601 1012
rect 10640 1046 10766 1062
rect 10640 1012 10652 1046
rect 10686 1012 10720 1046
rect 10754 1012 10766 1046
rect 10640 996 10766 1012
rect 63 920 189 936
rect 63 886 75 920
rect 109 886 143 920
rect 177 886 189 920
rect 63 870 189 886
rect 5228 920 5354 936
rect 5228 886 5240 920
rect 5274 886 5308 920
rect 5342 886 5354 920
rect 5228 870 5354 886
rect 5475 920 5601 936
rect 5475 886 5487 920
rect 5521 886 5555 920
rect 5589 886 5601 920
rect 5475 870 5601 886
rect 10640 920 10766 936
rect 10640 886 10652 920
rect 10686 886 10720 920
rect 10754 886 10766 920
rect 10640 870 10766 886
rect 63 794 189 810
rect 63 760 75 794
rect 109 760 143 794
rect 177 760 189 794
rect 63 744 189 760
rect 5228 794 5354 810
rect 5228 760 5240 794
rect 5274 760 5308 794
rect 5342 760 5354 794
rect 5228 744 5354 760
rect 5475 794 5601 810
rect 5475 760 5487 794
rect 5521 760 5555 794
rect 5589 760 5601 794
rect 5475 744 5601 760
rect 10640 794 10766 810
rect 10640 760 10652 794
rect 10686 760 10720 794
rect 10754 760 10766 794
rect 10640 744 10766 760
rect 63 668 189 684
rect 63 634 75 668
rect 109 634 143 668
rect 177 634 189 668
rect 63 618 189 634
rect 5228 668 5354 684
rect 5228 634 5240 668
rect 5274 634 5308 668
rect 5342 634 5354 668
rect 5228 618 5354 634
rect 63 542 189 558
rect 63 508 75 542
rect 109 508 143 542
rect 177 508 189 542
rect 63 492 189 508
rect 5228 542 5354 558
rect 5228 508 5240 542
rect 5274 508 5308 542
rect 5342 508 5354 542
rect 5228 492 5354 508
rect 63 416 189 432
rect 63 382 75 416
rect 109 382 143 416
rect 177 382 189 416
rect 63 366 189 382
rect 5228 416 5354 432
rect 5228 382 5240 416
rect 5274 382 5308 416
rect 5342 382 5354 416
rect 5228 366 5354 382
rect 63 290 189 306
rect 63 256 75 290
rect 109 256 143 290
rect 177 256 189 290
rect 63 240 189 256
rect 5228 290 5354 306
rect 5228 256 5240 290
rect 5274 256 5308 290
rect 5342 256 5354 290
rect 5228 240 5354 256
rect 63 164 189 180
rect 63 130 75 164
rect 109 130 143 164
rect 177 130 189 164
rect 63 114 189 130
rect 5228 164 5354 180
rect 5228 130 5240 164
rect 5274 130 5308 164
rect 5342 130 5354 164
rect 5228 114 5354 130
<< ndiffc >>
rect 3799 1901 3833 1935
rect 8896 1901 8930 1935
rect 3799 1775 3833 1809
rect 8896 1775 8930 1809
rect 3799 1649 3833 1683
rect 8896 1649 8930 1683
rect 3799 1523 3833 1557
rect 8896 1523 8930 1557
rect 5555 1390 5589 1424
rect 10652 1390 10686 1424
rect 143 1264 177 1298
rect 5240 1264 5274 1298
rect 5555 1264 5589 1298
rect 10652 1264 10686 1298
rect 143 1138 177 1172
rect 5240 1138 5274 1172
rect 5555 1138 5589 1172
rect 10652 1138 10686 1172
rect 143 1012 177 1046
rect 5240 1012 5274 1046
rect 5555 1012 5589 1046
rect 10652 1012 10686 1046
rect 143 886 177 920
rect 5240 886 5274 920
rect 5555 886 5589 920
rect 10652 886 10686 920
rect 143 760 177 794
rect 5240 760 5274 794
rect 5555 760 5589 794
rect 10652 760 10686 794
rect 143 634 177 668
rect 5240 634 5274 668
rect 143 508 177 542
rect 5240 508 5274 542
rect 143 382 177 416
rect 5240 382 5274 416
rect 143 256 177 290
rect 5240 256 5274 290
rect 143 130 177 164
rect 5240 130 5274 164
<< mvndiffc >>
rect 3731 1901 3765 1935
rect 8964 1901 8998 1935
rect 3731 1775 3765 1809
rect 8964 1775 8998 1809
rect 3731 1649 3765 1683
rect 8964 1649 8998 1683
rect 3731 1523 3765 1557
rect 8964 1523 8998 1557
rect 5487 1390 5521 1424
rect 10720 1390 10754 1424
rect 75 1264 109 1298
rect 5308 1264 5342 1298
rect 5487 1264 5521 1298
rect 10720 1264 10754 1298
rect 75 1138 109 1172
rect 5308 1138 5342 1172
rect 5487 1138 5521 1172
rect 10720 1138 10754 1172
rect 75 1012 109 1046
rect 5308 1012 5342 1046
rect 5487 1012 5521 1046
rect 10720 1012 10754 1046
rect 75 886 109 920
rect 5308 886 5342 920
rect 5487 886 5521 920
rect 10720 886 10754 920
rect 75 760 109 794
rect 5308 760 5342 794
rect 5487 760 5521 794
rect 10720 760 10754 794
rect 75 634 109 668
rect 5308 634 5342 668
rect 75 508 109 542
rect 5308 508 5342 542
rect 75 382 109 416
rect 5308 382 5342 416
rect 75 256 109 290
rect 5308 256 5342 290
rect 75 130 109 164
rect 5308 130 5342 164
<< nsubdiff >>
rect 7712 2709 7820 2743
rect 7854 2709 7891 2743
rect 7925 2709 7962 2743
rect 7996 2709 8033 2743
rect 8067 2709 8104 2743
rect 8138 2709 8175 2743
rect 8209 2709 8246 2743
rect 8280 2709 8317 2743
rect 8351 2709 8388 2743
rect 8422 2709 8459 2743
rect 8493 2709 8530 2743
rect 8564 2709 8601 2743
rect 8635 2709 8672 2743
rect 8706 2709 8744 2743
rect 8778 2709 8816 2743
rect 8850 2709 8888 2743
rect 7712 2613 7746 2675
rect 8922 2616 8956 2743
rect 7712 2459 7746 2579
rect 8922 2535 8956 2582
rect 8922 2454 8956 2501
rect 7712 2305 7746 2425
rect 8922 2373 8956 2420
rect 7780 2305 7818 2339
rect 7852 2305 7890 2339
rect 7924 2305 7962 2339
rect 7996 2305 8033 2339
rect 8067 2305 8104 2339
rect 8138 2305 8175 2339
rect 8209 2305 8246 2339
rect 8280 2305 8317 2339
rect 8351 2305 8388 2339
rect 8422 2305 8459 2339
rect 8493 2305 8530 2339
rect 8564 2305 8601 2339
rect 8635 2305 8672 2339
rect 8706 2305 8743 2339
rect 8777 2305 8814 2339
rect 8848 2305 8956 2339
<< mvpsubdiff >>
rect 3536 2059 3604 2093
rect 3638 2059 3672 2093
rect 3706 2059 3740 2093
rect 3774 2059 3808 2093
rect 3842 2059 3876 2093
rect 3910 2059 3944 2093
rect 3978 2059 4012 2093
rect 4046 2059 4080 2093
rect 4114 2059 4148 2093
rect 4182 2059 4216 2093
rect 4250 2059 4284 2093
rect 4318 2059 4352 2093
rect 4386 2059 4420 2093
rect 4454 2059 4488 2093
rect 4522 2059 4556 2093
rect 4590 2059 4624 2093
rect 4658 2059 4692 2093
rect 4726 2059 4760 2093
rect 4794 2059 4828 2093
rect 4862 2059 4896 2093
rect 4930 2059 4964 2093
rect 4998 2059 5032 2093
rect 5066 2059 5100 2093
rect 5134 2059 5168 2093
rect 5202 2059 5236 2093
rect 5270 2059 5304 2093
rect 5338 2059 5372 2093
rect 5406 2059 5440 2093
rect 5474 2059 5508 2093
rect 5542 2059 5576 2093
rect 5610 2059 5644 2093
rect 5678 2059 5712 2093
rect 5746 2059 5780 2093
rect 5814 2059 5848 2093
rect 5882 2059 5916 2093
rect 5950 2059 5984 2093
rect 6018 2059 6052 2093
rect 6086 2059 6120 2093
rect 6154 2059 6188 2093
rect 6222 2059 6256 2093
rect 6290 2059 6324 2093
rect 6358 2059 6392 2093
rect 6426 2059 6460 2093
rect 6494 2059 6528 2093
rect 6562 2059 6596 2093
rect 6630 2059 6664 2093
rect 6698 2059 6732 2093
rect 6766 2059 6800 2093
rect 6834 2059 6868 2093
rect 6902 2059 6936 2093
rect 6970 2059 7004 2093
rect 7038 2059 7072 2093
rect 7106 2059 7140 2093
rect 7174 2059 7208 2093
rect 7242 2059 7276 2093
rect 7310 2059 7344 2093
rect 7378 2059 7412 2093
rect 7446 2059 7480 2093
rect 7514 2059 7548 2093
rect 7582 2059 7616 2093
rect 7650 2059 7684 2093
rect 7718 2059 7752 2093
rect 7786 2059 7820 2093
rect 7854 2059 7888 2093
rect 7922 2059 7956 2093
rect 7990 2059 8024 2093
rect 8058 2059 8092 2093
rect 8126 2059 8160 2093
rect 8194 2059 8228 2093
rect 8262 2059 8296 2093
rect 8330 2059 8364 2093
rect 8398 2059 8432 2093
rect 8466 2059 8500 2093
rect 8534 2059 8568 2093
rect 8602 2059 8636 2093
rect 8670 2059 8704 2093
rect 8738 2059 8772 2093
rect 8806 2059 8840 2093
rect 8874 2059 8908 2093
rect 8942 2059 8976 2093
rect 9010 2059 9044 2093
rect 9078 2059 9164 2093
rect 3536 1966 3570 2059
rect 9130 2025 9164 2059
rect 9130 1957 9164 1991
rect 3536 1898 3570 1932
rect 9130 1889 9164 1923
rect 3536 1830 3570 1864
rect 3536 1762 3570 1796
rect 9130 1821 9164 1855
rect 3536 1694 3570 1728
rect 9130 1753 9164 1787
rect 3536 1626 3570 1660
rect 9130 1685 9164 1719
rect 3536 1558 3570 1592
rect 9130 1617 9164 1651
rect 3536 1490 3570 1524
rect 9130 1548 9164 1583
rect 9130 1514 9198 1548
rect 9232 1514 9266 1548
rect 9300 1514 9334 1548
rect 9368 1514 9402 1548
rect 9436 1514 9470 1548
rect 9504 1514 9538 1548
rect 9572 1514 9606 1548
rect 9640 1514 9674 1548
rect 9708 1514 9742 1548
rect 9776 1514 9810 1548
rect 9844 1514 9878 1548
rect 9912 1514 9946 1548
rect 9980 1514 10014 1548
rect 10048 1514 10082 1548
rect 10116 1514 10150 1548
rect 10184 1514 10218 1548
rect 10252 1514 10286 1548
rect 10320 1514 10354 1548
rect 10388 1514 10422 1548
rect 10456 1514 10490 1548
rect 10524 1514 10558 1548
rect 10592 1514 10626 1548
rect 10660 1514 10694 1548
rect 10728 1514 10762 1548
rect 10796 1514 10879 1548
rect 3536 1422 3570 1456
rect 10845 1480 10879 1514
rect -45 1388 23 1422
rect 57 1388 91 1422
rect 125 1388 159 1422
rect 193 1388 227 1422
rect 261 1388 295 1422
rect 329 1388 363 1422
rect 397 1388 431 1422
rect 465 1388 499 1422
rect 533 1388 567 1422
rect 601 1388 635 1422
rect 669 1388 703 1422
rect 737 1388 771 1422
rect 805 1388 839 1422
rect 873 1388 907 1422
rect 941 1388 975 1422
rect 1009 1388 1043 1422
rect 1077 1388 1111 1422
rect 1145 1388 1179 1422
rect 1213 1388 1247 1422
rect 1281 1388 1315 1422
rect 1349 1388 1383 1422
rect 1417 1388 1451 1422
rect 1485 1388 1519 1422
rect 1553 1388 1587 1422
rect 1621 1388 1655 1422
rect 1689 1388 1723 1422
rect 1757 1388 1791 1422
rect 1825 1388 1859 1422
rect 1893 1388 1927 1422
rect 1961 1388 1995 1422
rect 2029 1388 2063 1422
rect 2097 1388 2131 1422
rect 2165 1388 2199 1422
rect 2233 1388 2267 1422
rect 2301 1388 2335 1422
rect 2369 1388 2403 1422
rect 2437 1388 2471 1422
rect 2505 1388 2539 1422
rect 2573 1388 2607 1422
rect 2641 1388 2675 1422
rect 2709 1388 2743 1422
rect 2777 1388 2811 1422
rect 2845 1388 2879 1422
rect 2913 1388 2947 1422
rect 2981 1388 3015 1422
rect 3049 1388 3083 1422
rect 3117 1388 3151 1422
rect 3185 1388 3219 1422
rect 3253 1388 3287 1422
rect 3321 1388 3355 1422
rect 3389 1388 3423 1422
rect 3457 1388 3570 1422
rect -45 1196 -11 1388
rect 10845 1412 10879 1446
rect 10845 1344 10879 1378
rect 10845 1276 10879 1310
rect 10845 1208 10879 1242
rect -45 1128 -11 1162
rect 10845 1140 10879 1174
rect -45 1060 -11 1094
rect 10845 1072 10879 1106
rect -45 992 -11 1026
rect 10845 1004 10879 1038
rect -45 924 -11 958
rect 10845 936 10879 970
rect -45 856 -11 890
rect -45 788 -11 822
rect 10845 868 10879 902
rect -45 720 -11 754
rect 10845 800 10879 834
rect -45 652 -11 686
rect 10845 667 10879 766
rect 5428 633 5541 667
rect 5575 633 5609 667
rect 5643 633 5677 667
rect 5711 633 5745 667
rect 5779 633 5813 667
rect 5847 633 5881 667
rect 5915 633 5949 667
rect 5983 633 6017 667
rect 6051 633 6085 667
rect 6119 633 6153 667
rect 6187 633 6221 667
rect 6255 633 6289 667
rect 6323 633 6357 667
rect 6391 633 6425 667
rect 6459 633 6493 667
rect 6527 633 6561 667
rect 6595 633 6629 667
rect 6663 633 6697 667
rect 6731 633 6765 667
rect 6799 633 6833 667
rect 6867 633 6901 667
rect 6935 633 6969 667
rect 7003 633 7037 667
rect 7071 633 7105 667
rect 7139 633 7173 667
rect 7207 633 7241 667
rect 7275 633 7309 667
rect 7343 633 7377 667
rect 7411 633 7445 667
rect 7479 633 7513 667
rect 7547 633 7581 667
rect 7615 633 7649 667
rect 7683 633 7717 667
rect 7751 633 7785 667
rect 7819 633 7853 667
rect 7887 633 7921 667
rect 7955 633 7989 667
rect 8023 633 8057 667
rect 8091 633 8125 667
rect 8159 633 8193 667
rect 8227 633 8261 667
rect 8295 633 8329 667
rect 8363 633 8397 667
rect 8431 633 8465 667
rect 8499 633 8533 667
rect 8567 633 8601 667
rect 8635 633 8669 667
rect 8703 633 8737 667
rect 8771 633 8805 667
rect 8839 633 8873 667
rect 8907 633 8941 667
rect 8975 633 9009 667
rect 9043 633 9077 667
rect 9111 633 9145 667
rect 9179 633 9213 667
rect 9247 633 9281 667
rect 9315 633 9349 667
rect 9383 633 9417 667
rect 9451 633 9485 667
rect 9519 633 9553 667
rect 9587 633 9621 667
rect 9655 633 9689 667
rect 9723 633 9757 667
rect 9791 633 9825 667
rect 9859 633 9893 667
rect 9927 633 9961 667
rect 9995 633 10029 667
rect 10063 633 10097 667
rect 10131 633 10165 667
rect 10199 633 10233 667
rect 10267 633 10301 667
rect 10335 633 10369 667
rect 10403 633 10437 667
rect 10471 633 10505 667
rect 10539 633 10573 667
rect 10607 633 10641 667
rect 10675 633 10709 667
rect 10743 633 10777 667
rect 10811 633 10879 667
rect -45 584 -11 618
rect 5428 599 5462 633
rect -45 516 -11 550
rect 5428 531 5462 565
rect -45 448 -11 482
rect 5428 463 5462 497
rect -45 380 -11 414
rect 5428 395 5462 429
rect -45 312 -11 346
rect 5428 327 5462 361
rect -45 244 -11 278
rect 5428 259 5462 293
rect -45 176 -11 210
rect 5428 191 5462 225
rect -45 108 -11 142
rect 5428 123 5462 157
rect -45 40 -11 74
rect 5428 40 5462 89
rect -45 6 56 40
rect 90 6 124 40
rect 158 6 192 40
rect 226 6 260 40
rect 294 6 328 40
rect 362 6 396 40
rect 430 6 464 40
rect 498 6 532 40
rect 566 6 600 40
rect 634 6 668 40
rect 702 6 736 40
rect 770 6 804 40
rect 838 6 872 40
rect 906 6 940 40
rect 974 6 1008 40
rect 1042 6 1076 40
rect 1110 6 1144 40
rect 1178 6 1212 40
rect 1246 6 1280 40
rect 1314 6 1348 40
rect 1382 6 1416 40
rect 1450 6 1484 40
rect 1518 6 1552 40
rect 1586 6 1620 40
rect 1654 6 1688 40
rect 1722 6 1756 40
rect 1790 6 1824 40
rect 1858 6 1892 40
rect 1926 6 1960 40
rect 1994 6 2028 40
rect 2062 6 2096 40
rect 2130 6 2164 40
rect 2198 6 2232 40
rect 2266 6 2300 40
rect 2334 6 2368 40
rect 2402 6 2436 40
rect 2470 6 2504 40
rect 2538 6 2572 40
rect 2606 6 2640 40
rect 2674 6 2708 40
rect 2742 6 2776 40
rect 2810 6 2844 40
rect 2878 6 2912 40
rect 2946 6 2980 40
rect 3014 6 3048 40
rect 3082 6 3116 40
rect 3150 6 3184 40
rect 3218 6 3252 40
rect 3286 6 3320 40
rect 3354 6 3388 40
rect 3422 6 3456 40
rect 3490 6 3524 40
rect 3558 6 3592 40
rect 3626 6 3660 40
rect 3694 6 3728 40
rect 3762 6 3796 40
rect 3830 6 3864 40
rect 3898 6 3932 40
rect 3966 6 4000 40
rect 4034 6 4068 40
rect 4102 6 4136 40
rect 4170 6 4204 40
rect 4238 6 4272 40
rect 4306 6 4340 40
rect 4374 6 4408 40
rect 4442 6 4476 40
rect 4510 6 4544 40
rect 4578 6 4612 40
rect 4646 6 4680 40
rect 4714 6 4748 40
rect 4782 6 4816 40
rect 4850 6 4884 40
rect 4918 6 4952 40
rect 4986 6 5020 40
rect 5054 6 5088 40
rect 5122 6 5156 40
rect 5190 6 5224 40
rect 5258 6 5292 40
rect 5326 6 5360 40
rect 5394 6 5462 40
<< nsubdiffcont >>
rect 7820 2709 7854 2743
rect 7891 2709 7925 2743
rect 7962 2709 7996 2743
rect 8033 2709 8067 2743
rect 8104 2709 8138 2743
rect 8175 2709 8209 2743
rect 8246 2709 8280 2743
rect 8317 2709 8351 2743
rect 8388 2709 8422 2743
rect 8459 2709 8493 2743
rect 8530 2709 8564 2743
rect 8601 2709 8635 2743
rect 8672 2709 8706 2743
rect 8744 2709 8778 2743
rect 8816 2709 8850 2743
rect 8888 2709 8922 2743
rect 7712 2675 7746 2709
rect 7712 2579 7746 2613
rect 7712 2425 7746 2459
rect 8922 2582 8956 2616
rect 8922 2501 8956 2535
rect 8922 2420 8956 2454
rect 8922 2339 8956 2373
rect 7746 2305 7780 2339
rect 7818 2305 7852 2339
rect 7890 2305 7924 2339
rect 7962 2305 7996 2339
rect 8033 2305 8067 2339
rect 8104 2305 8138 2339
rect 8175 2305 8209 2339
rect 8246 2305 8280 2339
rect 8317 2305 8351 2339
rect 8388 2305 8422 2339
rect 8459 2305 8493 2339
rect 8530 2305 8564 2339
rect 8601 2305 8635 2339
rect 8672 2305 8706 2339
rect 8743 2305 8777 2339
rect 8814 2305 8848 2339
<< mvpsubdiffcont >>
rect 3604 2059 3638 2093
rect 3672 2059 3706 2093
rect 3740 2059 3774 2093
rect 3808 2059 3842 2093
rect 3876 2059 3910 2093
rect 3944 2059 3978 2093
rect 4012 2059 4046 2093
rect 4080 2059 4114 2093
rect 4148 2059 4182 2093
rect 4216 2059 4250 2093
rect 4284 2059 4318 2093
rect 4352 2059 4386 2093
rect 4420 2059 4454 2093
rect 4488 2059 4522 2093
rect 4556 2059 4590 2093
rect 4624 2059 4658 2093
rect 4692 2059 4726 2093
rect 4760 2059 4794 2093
rect 4828 2059 4862 2093
rect 4896 2059 4930 2093
rect 4964 2059 4998 2093
rect 5032 2059 5066 2093
rect 5100 2059 5134 2093
rect 5168 2059 5202 2093
rect 5236 2059 5270 2093
rect 5304 2059 5338 2093
rect 5372 2059 5406 2093
rect 5440 2059 5474 2093
rect 5508 2059 5542 2093
rect 5576 2059 5610 2093
rect 5644 2059 5678 2093
rect 5712 2059 5746 2093
rect 5780 2059 5814 2093
rect 5848 2059 5882 2093
rect 5916 2059 5950 2093
rect 5984 2059 6018 2093
rect 6052 2059 6086 2093
rect 6120 2059 6154 2093
rect 6188 2059 6222 2093
rect 6256 2059 6290 2093
rect 6324 2059 6358 2093
rect 6392 2059 6426 2093
rect 6460 2059 6494 2093
rect 6528 2059 6562 2093
rect 6596 2059 6630 2093
rect 6664 2059 6698 2093
rect 6732 2059 6766 2093
rect 6800 2059 6834 2093
rect 6868 2059 6902 2093
rect 6936 2059 6970 2093
rect 7004 2059 7038 2093
rect 7072 2059 7106 2093
rect 7140 2059 7174 2093
rect 7208 2059 7242 2093
rect 7276 2059 7310 2093
rect 7344 2059 7378 2093
rect 7412 2059 7446 2093
rect 7480 2059 7514 2093
rect 7548 2059 7582 2093
rect 7616 2059 7650 2093
rect 7684 2059 7718 2093
rect 7752 2059 7786 2093
rect 7820 2059 7854 2093
rect 7888 2059 7922 2093
rect 7956 2059 7990 2093
rect 8024 2059 8058 2093
rect 8092 2059 8126 2093
rect 8160 2059 8194 2093
rect 8228 2059 8262 2093
rect 8296 2059 8330 2093
rect 8364 2059 8398 2093
rect 8432 2059 8466 2093
rect 8500 2059 8534 2093
rect 8568 2059 8602 2093
rect 8636 2059 8670 2093
rect 8704 2059 8738 2093
rect 8772 2059 8806 2093
rect 8840 2059 8874 2093
rect 8908 2059 8942 2093
rect 8976 2059 9010 2093
rect 9044 2059 9078 2093
rect 3536 1932 3570 1966
rect 9130 1991 9164 2025
rect 3536 1864 3570 1898
rect 9130 1923 9164 1957
rect 3536 1796 3570 1830
rect 9130 1855 9164 1889
rect 3536 1728 3570 1762
rect 9130 1787 9164 1821
rect 9130 1719 9164 1753
rect 3536 1660 3570 1694
rect 9130 1651 9164 1685
rect 3536 1592 3570 1626
rect 9130 1583 9164 1617
rect 3536 1524 3570 1558
rect 9198 1514 9232 1548
rect 9266 1514 9300 1548
rect 9334 1514 9368 1548
rect 9402 1514 9436 1548
rect 9470 1514 9504 1548
rect 9538 1514 9572 1548
rect 9606 1514 9640 1548
rect 9674 1514 9708 1548
rect 9742 1514 9776 1548
rect 9810 1514 9844 1548
rect 9878 1514 9912 1548
rect 9946 1514 9980 1548
rect 10014 1514 10048 1548
rect 10082 1514 10116 1548
rect 10150 1514 10184 1548
rect 10218 1514 10252 1548
rect 10286 1514 10320 1548
rect 10354 1514 10388 1548
rect 10422 1514 10456 1548
rect 10490 1514 10524 1548
rect 10558 1514 10592 1548
rect 10626 1514 10660 1548
rect 10694 1514 10728 1548
rect 10762 1514 10796 1548
rect 3536 1456 3570 1490
rect 10845 1446 10879 1480
rect 23 1388 57 1422
rect 91 1388 125 1422
rect 159 1388 193 1422
rect 227 1388 261 1422
rect 295 1388 329 1422
rect 363 1388 397 1422
rect 431 1388 465 1422
rect 499 1388 533 1422
rect 567 1388 601 1422
rect 635 1388 669 1422
rect 703 1388 737 1422
rect 771 1388 805 1422
rect 839 1388 873 1422
rect 907 1388 941 1422
rect 975 1388 1009 1422
rect 1043 1388 1077 1422
rect 1111 1388 1145 1422
rect 1179 1388 1213 1422
rect 1247 1388 1281 1422
rect 1315 1388 1349 1422
rect 1383 1388 1417 1422
rect 1451 1388 1485 1422
rect 1519 1388 1553 1422
rect 1587 1388 1621 1422
rect 1655 1388 1689 1422
rect 1723 1388 1757 1422
rect 1791 1388 1825 1422
rect 1859 1388 1893 1422
rect 1927 1388 1961 1422
rect 1995 1388 2029 1422
rect 2063 1388 2097 1422
rect 2131 1388 2165 1422
rect 2199 1388 2233 1422
rect 2267 1388 2301 1422
rect 2335 1388 2369 1422
rect 2403 1388 2437 1422
rect 2471 1388 2505 1422
rect 2539 1388 2573 1422
rect 2607 1388 2641 1422
rect 2675 1388 2709 1422
rect 2743 1388 2777 1422
rect 2811 1388 2845 1422
rect 2879 1388 2913 1422
rect 2947 1388 2981 1422
rect 3015 1388 3049 1422
rect 3083 1388 3117 1422
rect 3151 1388 3185 1422
rect 3219 1388 3253 1422
rect 3287 1388 3321 1422
rect 3355 1388 3389 1422
rect 3423 1388 3457 1422
rect 10845 1378 10879 1412
rect 10845 1310 10879 1344
rect -45 1162 -11 1196
rect 10845 1242 10879 1276
rect -45 1094 -11 1128
rect 10845 1174 10879 1208
rect 10845 1106 10879 1140
rect -45 1026 -11 1060
rect 10845 1038 10879 1072
rect -45 958 -11 992
rect 10845 970 10879 1004
rect -45 890 -11 924
rect 10845 902 10879 936
rect -45 822 -11 856
rect 10845 834 10879 868
rect -45 754 -11 788
rect 10845 766 10879 800
rect -45 686 -11 720
rect -45 618 -11 652
rect 5541 633 5575 667
rect 5609 633 5643 667
rect 5677 633 5711 667
rect 5745 633 5779 667
rect 5813 633 5847 667
rect 5881 633 5915 667
rect 5949 633 5983 667
rect 6017 633 6051 667
rect 6085 633 6119 667
rect 6153 633 6187 667
rect 6221 633 6255 667
rect 6289 633 6323 667
rect 6357 633 6391 667
rect 6425 633 6459 667
rect 6493 633 6527 667
rect 6561 633 6595 667
rect 6629 633 6663 667
rect 6697 633 6731 667
rect 6765 633 6799 667
rect 6833 633 6867 667
rect 6901 633 6935 667
rect 6969 633 7003 667
rect 7037 633 7071 667
rect 7105 633 7139 667
rect 7173 633 7207 667
rect 7241 633 7275 667
rect 7309 633 7343 667
rect 7377 633 7411 667
rect 7445 633 7479 667
rect 7513 633 7547 667
rect 7581 633 7615 667
rect 7649 633 7683 667
rect 7717 633 7751 667
rect 7785 633 7819 667
rect 7853 633 7887 667
rect 7921 633 7955 667
rect 7989 633 8023 667
rect 8057 633 8091 667
rect 8125 633 8159 667
rect 8193 633 8227 667
rect 8261 633 8295 667
rect 8329 633 8363 667
rect 8397 633 8431 667
rect 8465 633 8499 667
rect 8533 633 8567 667
rect 8601 633 8635 667
rect 8669 633 8703 667
rect 8737 633 8771 667
rect 8805 633 8839 667
rect 8873 633 8907 667
rect 8941 633 8975 667
rect 9009 633 9043 667
rect 9077 633 9111 667
rect 9145 633 9179 667
rect 9213 633 9247 667
rect 9281 633 9315 667
rect 9349 633 9383 667
rect 9417 633 9451 667
rect 9485 633 9519 667
rect 9553 633 9587 667
rect 9621 633 9655 667
rect 9689 633 9723 667
rect 9757 633 9791 667
rect 9825 633 9859 667
rect 9893 633 9927 667
rect 9961 633 9995 667
rect 10029 633 10063 667
rect 10097 633 10131 667
rect 10165 633 10199 667
rect 10233 633 10267 667
rect 10301 633 10335 667
rect 10369 633 10403 667
rect 10437 633 10471 667
rect 10505 633 10539 667
rect 10573 633 10607 667
rect 10641 633 10675 667
rect 10709 633 10743 667
rect 10777 633 10811 667
rect -45 550 -11 584
rect 5428 565 5462 599
rect -45 482 -11 516
rect 5428 497 5462 531
rect -45 414 -11 448
rect -45 346 -11 380
rect 5428 429 5462 463
rect -45 278 -11 312
rect 5428 361 5462 395
rect -45 210 -11 244
rect 5428 293 5462 327
rect 5428 225 5462 259
rect -45 142 -11 176
rect 5428 157 5462 191
rect -45 74 -11 108
rect 5428 89 5462 123
rect 56 6 90 40
rect 124 6 158 40
rect 192 6 226 40
rect 260 6 294 40
rect 328 6 362 40
rect 396 6 430 40
rect 464 6 498 40
rect 532 6 566 40
rect 600 6 634 40
rect 668 6 702 40
rect 736 6 770 40
rect 804 6 838 40
rect 872 6 906 40
rect 940 6 974 40
rect 1008 6 1042 40
rect 1076 6 1110 40
rect 1144 6 1178 40
rect 1212 6 1246 40
rect 1280 6 1314 40
rect 1348 6 1382 40
rect 1416 6 1450 40
rect 1484 6 1518 40
rect 1552 6 1586 40
rect 1620 6 1654 40
rect 1688 6 1722 40
rect 1756 6 1790 40
rect 1824 6 1858 40
rect 1892 6 1926 40
rect 1960 6 1994 40
rect 2028 6 2062 40
rect 2096 6 2130 40
rect 2164 6 2198 40
rect 2232 6 2266 40
rect 2300 6 2334 40
rect 2368 6 2402 40
rect 2436 6 2470 40
rect 2504 6 2538 40
rect 2572 6 2606 40
rect 2640 6 2674 40
rect 2708 6 2742 40
rect 2776 6 2810 40
rect 2844 6 2878 40
rect 2912 6 2946 40
rect 2980 6 3014 40
rect 3048 6 3082 40
rect 3116 6 3150 40
rect 3184 6 3218 40
rect 3252 6 3286 40
rect 3320 6 3354 40
rect 3388 6 3422 40
rect 3456 6 3490 40
rect 3524 6 3558 40
rect 3592 6 3626 40
rect 3660 6 3694 40
rect 3728 6 3762 40
rect 3796 6 3830 40
rect 3864 6 3898 40
rect 3932 6 3966 40
rect 4000 6 4034 40
rect 4068 6 4102 40
rect 4136 6 4170 40
rect 4204 6 4238 40
rect 4272 6 4306 40
rect 4340 6 4374 40
rect 4408 6 4442 40
rect 4476 6 4510 40
rect 4544 6 4578 40
rect 4612 6 4646 40
rect 4680 6 4714 40
rect 4748 6 4782 40
rect 4816 6 4850 40
rect 4884 6 4918 40
rect 4952 6 4986 40
rect 5020 6 5054 40
rect 5088 6 5122 40
rect 5156 6 5190 40
rect 5224 6 5258 40
rect 5292 6 5326 40
rect 5360 6 5394 40
<< poly >>
rect 8826 2586 8898 2602
rect 8826 2552 8848 2586
rect 8882 2552 8898 2586
rect 8832 2496 8898 2552
rect 8826 2462 8848 2496
rect 8882 2462 8898 2496
rect 8826 2446 8898 2462
<< polycont >>
rect 8848 2552 8882 2586
rect 8848 2462 8882 2496
<< locali >>
rect 7712 2711 7735 2743
rect 7769 2711 7810 2745
rect 7844 2743 7885 2745
rect 7919 2743 7960 2745
rect 7994 2743 8035 2745
rect 8069 2743 8109 2745
rect 8143 2743 8183 2745
rect 8217 2743 8257 2745
rect 8291 2743 8331 2745
rect 8365 2743 8405 2745
rect 8439 2743 8479 2745
rect 8513 2743 8553 2745
rect 8587 2743 8627 2745
rect 8661 2743 8701 2745
rect 8735 2743 8775 2745
rect 8809 2743 8849 2745
rect 8883 2743 8957 2745
rect 7854 2711 7885 2743
rect 7925 2711 7960 2743
rect 7712 2709 7820 2711
rect 7854 2709 7891 2711
rect 7925 2709 7962 2711
rect 7996 2709 8033 2743
rect 8069 2711 8104 2743
rect 8143 2711 8175 2743
rect 8217 2711 8246 2743
rect 8291 2711 8317 2743
rect 8365 2711 8388 2743
rect 8439 2711 8459 2743
rect 8513 2711 8530 2743
rect 8587 2711 8601 2743
rect 8661 2711 8672 2743
rect 8735 2711 8744 2743
rect 8809 2711 8816 2743
rect 8883 2711 8888 2743
rect 8067 2709 8104 2711
rect 8138 2709 8175 2711
rect 8209 2709 8246 2711
rect 8280 2709 8317 2711
rect 8351 2709 8388 2711
rect 8422 2709 8459 2711
rect 8493 2709 8530 2711
rect 8564 2709 8601 2711
rect 8635 2709 8672 2711
rect 8706 2709 8744 2711
rect 8778 2709 8816 2711
rect 8850 2709 8888 2711
rect 7712 2613 7746 2675
rect 8922 2673 8957 2743
rect 7888 2611 7930 2645
rect 7964 2611 8006 2645
rect 8040 2611 8082 2645
rect 8116 2611 8158 2645
rect 8192 2611 8234 2645
rect 8268 2611 8310 2645
rect 8344 2611 8386 2645
rect 8420 2611 8461 2645
rect 8495 2611 8536 2645
rect 8570 2611 8611 2645
rect 8645 2611 8686 2645
rect 8720 2611 8761 2645
rect 8922 2639 8923 2673
rect 8922 2616 8957 2639
rect 7712 2555 7746 2579
rect 8848 2586 8882 2602
rect 7888 2507 7930 2541
rect 7964 2507 8006 2541
rect 8040 2507 8082 2541
rect 8116 2507 8158 2541
rect 8192 2507 8234 2541
rect 8268 2507 8310 2541
rect 8344 2507 8386 2541
rect 8420 2507 8461 2541
rect 8495 2507 8536 2541
rect 8570 2507 8611 2541
rect 8645 2507 8686 2541
rect 8720 2507 8761 2541
rect 8848 2509 8882 2547
rect 7712 2459 7746 2483
rect 8848 2446 8882 2462
rect 8956 2588 8957 2616
rect 8922 2554 8923 2582
rect 8922 2535 8957 2554
rect 8956 2503 8957 2535
rect 8922 2469 8923 2501
rect 8922 2454 8957 2469
rect 7712 2305 7746 2425
rect 7888 2401 7930 2435
rect 7964 2401 8006 2435
rect 8040 2401 8082 2435
rect 8116 2401 8158 2435
rect 8192 2401 8234 2435
rect 8268 2401 8310 2435
rect 8344 2401 8386 2435
rect 8420 2401 8461 2435
rect 8495 2401 8536 2435
rect 8570 2401 8611 2435
rect 8645 2401 8686 2435
rect 8720 2401 8761 2435
rect 8956 2420 8957 2454
rect 8922 2418 8957 2420
rect 8922 2384 8923 2418
rect 8922 2373 8957 2384
rect 8956 2339 8957 2373
rect 7780 2305 7818 2339
rect 7852 2333 7890 2339
rect 7852 2305 7854 2333
rect 7888 2305 7890 2333
rect 7924 2333 7962 2339
rect 7996 2333 8033 2339
rect 8067 2333 8104 2339
rect 8138 2333 8175 2339
rect 8209 2333 8246 2339
rect 8280 2333 8317 2339
rect 7924 2305 7930 2333
rect 7996 2305 8006 2333
rect 8067 2305 8082 2333
rect 8138 2305 8158 2333
rect 8209 2305 8235 2333
rect 8280 2305 8312 2333
rect 8351 2305 8388 2339
rect 8422 2333 8459 2339
rect 8493 2333 8530 2339
rect 8564 2333 8601 2339
rect 8635 2333 8672 2339
rect 8706 2333 8743 2339
rect 8777 2333 8814 2339
rect 8423 2305 8459 2333
rect 8500 2305 8530 2333
rect 8577 2305 8601 2333
rect 8654 2305 8672 2333
rect 8731 2305 8743 2333
rect 8808 2305 8814 2333
rect 8848 2333 8957 2339
rect 8848 2305 8851 2333
rect 7888 2299 7930 2305
rect 7964 2299 8006 2305
rect 8040 2299 8082 2305
rect 8116 2299 8158 2305
rect 8192 2299 8235 2305
rect 8269 2299 8312 2305
rect 8346 2299 8389 2305
rect 8423 2299 8466 2305
rect 8500 2299 8543 2305
rect 8577 2299 8620 2305
rect 8654 2299 8697 2305
rect 8731 2299 8774 2305
rect 8808 2299 8851 2305
rect 8885 2299 8957 2333
rect 3536 2059 3604 2093
rect 3638 2059 3648 2093
rect 3706 2059 3721 2093
rect 3774 2059 3794 2093
rect 3842 2059 3867 2093
rect 3910 2059 3940 2093
rect 3978 2059 4012 2093
rect 4047 2059 4080 2093
rect 4120 2059 4148 2093
rect 4193 2059 4216 2093
rect 4266 2059 4284 2093
rect 4339 2059 4352 2093
rect 4412 2059 4420 2093
rect 4485 2059 4488 2093
rect 4522 2059 4524 2093
rect 4590 2059 4597 2093
rect 4658 2059 4670 2093
rect 4726 2059 4743 2093
rect 4794 2059 4816 2093
rect 4862 2059 4889 2093
rect 4930 2059 4962 2093
rect 4998 2059 5032 2093
rect 5069 2059 5100 2093
rect 5142 2059 5168 2093
rect 5215 2059 5236 2093
rect 5288 2059 5304 2093
rect 5361 2059 5372 2093
rect 5434 2059 5440 2093
rect 5507 2059 5508 2093
rect 5542 2059 5546 2093
rect 5610 2059 5619 2093
rect 5678 2059 5692 2093
rect 5746 2059 5765 2093
rect 5814 2059 5838 2093
rect 5882 2059 5911 2093
rect 5950 2059 5984 2093
rect 6018 2059 6052 2093
rect 6091 2059 6120 2093
rect 6164 2059 6188 2093
rect 6237 2059 6256 2093
rect 6310 2059 6324 2093
rect 6383 2059 6392 2093
rect 6456 2059 6460 2093
rect 6494 2059 6495 2093
rect 6562 2059 6568 2093
rect 6630 2059 6641 2093
rect 6698 2059 6714 2093
rect 6766 2059 6787 2093
rect 6834 2059 6861 2093
rect 6902 2059 6935 2093
rect 6970 2059 7004 2093
rect 7043 2059 7072 2093
rect 7117 2059 7140 2093
rect 7191 2059 7208 2093
rect 7265 2059 7276 2093
rect 7339 2059 7344 2093
rect 7378 2059 7379 2093
rect 7446 2059 7480 2093
rect 7514 2059 7548 2093
rect 7582 2059 7616 2093
rect 7650 2059 7684 2093
rect 7718 2059 7752 2093
rect 7786 2059 7820 2093
rect 7854 2059 7888 2093
rect 7922 2059 7956 2093
rect 7990 2059 8024 2093
rect 8058 2059 8092 2093
rect 8126 2059 8160 2093
rect 8194 2059 8228 2093
rect 8262 2059 8296 2093
rect 8330 2059 8364 2093
rect 8398 2059 8432 2093
rect 8466 2059 8500 2093
rect 8534 2059 8568 2093
rect 8602 2059 8636 2093
rect 8670 2059 8698 2093
rect 8738 2059 8770 2093
rect 8806 2059 8840 2093
rect 8876 2059 8908 2093
rect 8948 2059 8976 2093
rect 9021 2059 9044 2093
rect 9094 2059 9164 2093
rect 3536 2055 3570 2059
rect 3536 1966 3570 2021
rect 9130 2025 9164 2059
rect 9130 1957 9164 1991
rect 3570 1935 7708 1951
rect 3570 1931 3731 1935
rect 3536 1901 3731 1931
rect 3765 1932 7708 1935
rect 3765 1901 7602 1932
rect 3536 1898 7602 1901
rect 7636 1898 7674 1932
rect 3570 1885 7708 1898
rect 8856 1935 9106 1951
rect 8856 1901 8964 1935
rect 8998 1901 9106 1935
rect 8856 1885 9106 1901
rect 9130 1889 9164 1923
rect 3536 1830 3570 1841
rect 3795 1817 3873 1825
rect 3536 1785 3570 1796
rect 3715 1809 3873 1817
rect 3715 1806 3731 1809
rect 3765 1806 3873 1809
rect 4608 1806 4642 1825
rect 5510 1806 5544 1825
rect 6412 1806 6446 1825
rect 7671 1806 7705 1825
rect 8880 1809 9014 1825
rect 8880 1806 8964 1809
rect 8998 1806 9014 1809
rect 3715 1772 3729 1806
rect 3765 1775 3801 1806
rect 3763 1772 3801 1775
rect 3835 1772 3873 1806
rect 4606 1772 4644 1806
rect 5508 1772 5546 1806
rect 6410 1772 6448 1806
rect 7669 1772 7707 1806
rect 8880 1772 8894 1806
rect 8928 1775 8964 1806
rect 8928 1772 8966 1775
rect 9000 1772 9014 1806
rect 3715 1767 3873 1772
rect 3795 1759 3873 1767
rect 4608 1759 4642 1772
rect 5510 1759 5544 1772
rect 6412 1759 6446 1772
rect 7671 1759 7705 1772
rect 3536 1694 3570 1728
rect 3536 1626 3570 1660
rect 3536 1558 3570 1592
rect 3536 1490 3570 1513
rect 3715 1683 4778 1699
rect 3715 1649 3731 1683
rect 3765 1680 4778 1683
rect 5153 1680 5187 1699
rect 6412 1680 6446 1699
rect 7671 1680 7705 1699
rect 8880 1684 9014 1772
rect 3765 1649 4672 1680
rect 3715 1646 4672 1649
rect 4706 1646 4744 1680
rect 5151 1646 5189 1680
rect 6410 1646 6448 1680
rect 7669 1646 7707 1680
rect 8880 1650 8894 1684
rect 8928 1683 8966 1684
rect 8928 1650 8964 1683
rect 9000 1650 9014 1684
rect 8880 1649 8964 1650
rect 8998 1649 9014 1650
rect 3715 1633 4778 1646
rect 5153 1633 5187 1646
rect 6412 1633 6446 1646
rect 7671 1633 7705 1646
rect 8880 1633 9014 1649
rect 9130 1821 9164 1855
rect 9130 1753 9164 1787
rect 9130 1685 9164 1719
rect 3715 1573 3849 1633
rect 9130 1617 9164 1651
rect 3715 1557 4778 1573
rect 3715 1523 3731 1557
rect 3765 1523 4672 1557
rect 4706 1523 4744 1557
rect 5153 1556 5187 1573
rect 6412 1557 6446 1573
rect 3715 1507 4778 1523
rect 5151 1522 5189 1556
rect 6410 1523 6448 1557
rect 7671 1555 7705 1573
rect 8878 1557 9014 1573
rect 8878 1556 8964 1557
rect 8998 1556 9014 1557
rect 5153 1507 5187 1522
rect 6412 1507 6446 1523
rect 7669 1521 7707 1555
rect 8878 1522 8894 1556
rect 8928 1523 8964 1556
rect 8928 1522 8966 1523
rect 9000 1522 9014 1556
rect 7671 1507 7705 1521
rect 3536 1422 3570 1456
rect 8878 1440 9014 1522
rect 9130 1548 9164 1583
rect 9130 1514 9198 1548
rect 9232 1514 9266 1548
rect 9300 1514 9334 1548
rect 9368 1514 9402 1548
rect 9436 1514 9470 1548
rect 9504 1514 9538 1548
rect 9572 1514 9606 1548
rect 9640 1514 9674 1548
rect 9708 1514 9742 1548
rect 9776 1514 9810 1548
rect 9844 1514 9878 1548
rect 9912 1514 9946 1548
rect 9980 1514 10014 1548
rect 10048 1514 10082 1548
rect 10116 1514 10150 1548
rect 10184 1514 10218 1548
rect 10252 1514 10286 1548
rect 10320 1514 10354 1548
rect 10388 1514 10422 1548
rect 10456 1514 10490 1548
rect 10524 1514 10558 1548
rect 10592 1514 10626 1548
rect 10660 1514 10694 1548
rect 10728 1514 10762 1548
rect 10796 1514 10879 1548
rect 10845 1480 10879 1514
rect -45 1388 23 1422
rect 57 1388 91 1422
rect 125 1388 159 1422
rect 193 1388 227 1422
rect 261 1388 295 1422
rect 329 1388 363 1422
rect 397 1388 431 1422
rect 465 1388 499 1422
rect 533 1388 567 1422
rect 601 1388 635 1422
rect 669 1388 703 1422
rect 737 1388 771 1422
rect 805 1388 839 1422
rect 873 1388 907 1422
rect 941 1388 975 1422
rect 1009 1388 1043 1422
rect 1077 1388 1111 1422
rect 1145 1388 1179 1422
rect 1213 1388 1247 1422
rect 1281 1388 1315 1422
rect 1349 1388 1383 1422
rect 1417 1388 1451 1422
rect 1485 1388 1519 1422
rect 1553 1388 1587 1422
rect 1621 1388 1655 1422
rect 1689 1388 1723 1422
rect 1757 1388 1791 1422
rect 1825 1388 1859 1422
rect 1893 1388 1927 1422
rect 1961 1388 1995 1422
rect 2029 1388 2063 1422
rect 2097 1388 2131 1422
rect 2165 1388 2199 1422
rect 2233 1388 2267 1422
rect 2301 1388 2335 1422
rect 2369 1388 2403 1422
rect 2437 1388 2471 1422
rect 2505 1388 2539 1422
rect 2573 1388 2607 1422
rect 2641 1388 2675 1422
rect 2709 1388 2743 1422
rect 2777 1388 2811 1422
rect 2845 1388 2879 1422
rect 2913 1388 2947 1422
rect 2981 1388 3015 1422
rect 3049 1388 3083 1422
rect 3117 1388 3151 1422
rect 3185 1388 3219 1422
rect 3253 1388 3287 1422
rect 3321 1388 3355 1422
rect 3389 1388 3422 1422
rect 3457 1388 3498 1422
rect 3532 1388 3570 1422
rect 5471 1424 5605 1440
rect 5471 1421 5487 1424
rect 5521 1421 5605 1424
rect -45 1196 -11 1388
rect 5471 1387 5485 1421
rect 5521 1390 5557 1421
rect 5519 1387 5557 1390
rect 5591 1387 5605 1421
rect 59 1303 3661 1314
rect 5199 1303 5358 1314
rect 59 1298 3528 1303
rect 59 1264 75 1298
rect 109 1269 3528 1298
rect 3562 1269 3600 1303
rect 3634 1269 3661 1303
rect 4269 1269 4307 1303
rect 5199 1269 5221 1303
rect 5255 1269 5293 1303
rect 5327 1298 5358 1303
rect 109 1264 3661 1269
rect 59 1248 3661 1264
rect 5199 1264 5308 1269
rect 5342 1264 5358 1298
rect 5199 1248 5358 1264
rect 5471 1298 5605 1387
rect 8878 1432 10652 1440
rect 10686 1432 10770 1440
rect 8878 1424 10770 1432
rect 8878 1421 10720 1424
rect 10754 1421 10770 1424
rect 8878 1387 10650 1421
rect 10684 1390 10720 1421
rect 10684 1387 10722 1390
rect 10756 1387 10770 1421
rect 8878 1382 10770 1387
rect 8878 1374 10652 1382
rect 10686 1374 10770 1382
rect 10845 1412 10879 1446
rect 10845 1344 10879 1378
rect 5471 1296 5487 1298
rect 5521 1296 5605 1298
rect 5471 1262 5485 1296
rect 5521 1264 5557 1296
rect 5519 1262 5557 1264
rect 5591 1262 5605 1296
rect 5471 1248 5605 1262
rect 10636 1299 10770 1314
rect 10636 1265 10650 1299
rect 10684 1298 10722 1299
rect 10684 1265 10720 1298
rect 10756 1265 10770 1299
rect 10636 1264 10720 1265
rect 10754 1264 10770 1265
rect -45 1128 -11 1162
rect -45 1060 -11 1094
rect -45 992 -11 1026
rect 59 1172 4482 1188
rect 59 1138 75 1172
rect 109 1138 4376 1172
rect 4410 1138 4448 1172
rect 59 1122 4482 1138
rect 5200 1172 5605 1188
rect 5200 1138 5238 1172
rect 5272 1138 5308 1172
rect 5344 1169 5487 1172
rect 5521 1169 5605 1172
rect 5344 1138 5485 1169
rect 5521 1138 5557 1169
rect 5200 1135 5485 1138
rect 5519 1135 5557 1138
rect 5591 1135 5605 1169
rect 5200 1122 5605 1135
rect 10636 1172 10770 1264
rect 10636 1169 10720 1172
rect 10754 1169 10770 1172
rect 10636 1135 10650 1169
rect 10684 1138 10720 1169
rect 10684 1135 10722 1138
rect 10756 1135 10770 1169
rect 10636 1122 10770 1135
rect 10845 1276 10879 1310
rect 10845 1208 10879 1242
rect 10845 1140 10879 1174
rect 59 1062 193 1122
rect 10845 1072 10879 1106
rect 59 1046 4482 1062
rect 59 1012 75 1046
rect 109 1012 4376 1046
rect 4410 1012 4448 1046
rect 59 996 4482 1012
rect 5200 1046 5605 1062
rect 5200 1012 5238 1046
rect 5272 1012 5308 1046
rect 5344 1043 5487 1046
rect 5521 1043 5605 1046
rect 5344 1012 5485 1043
rect 5521 1012 5557 1043
rect 5200 1009 5485 1012
rect 5519 1009 5557 1012
rect 5591 1009 5605 1043
rect 5200 996 5605 1009
rect 10636 1046 10770 1062
rect 10636 1043 10720 1046
rect 10754 1043 10770 1046
rect 10636 1009 10650 1043
rect 10684 1012 10720 1043
rect 10684 1009 10722 1012
rect 10756 1009 10770 1043
rect -45 924 -11 958
rect -45 856 -11 890
rect -45 788 -11 822
rect -45 720 -11 754
rect 59 920 4482 936
rect 59 886 75 920
rect 109 886 4376 920
rect 4410 886 4448 920
rect 59 870 4482 886
rect 5200 920 5605 936
rect 5200 886 5238 920
rect 5272 886 5308 920
rect 5344 917 5487 920
rect 5521 917 5605 920
rect 5344 886 5485 917
rect 5521 886 5557 917
rect 5200 883 5485 886
rect 5519 883 5557 886
rect 5591 883 5605 917
rect 5200 870 5605 883
rect 10636 920 10770 1009
rect 10636 917 10720 920
rect 10754 917 10770 920
rect 10636 883 10650 917
rect 10684 886 10720 917
rect 10684 883 10722 886
rect 10756 883 10770 917
rect 10636 870 10770 883
rect 10845 1004 10879 1038
rect 10845 936 10879 970
rect 59 810 193 870
rect 10845 868 10879 902
rect 59 794 4482 810
rect 59 760 75 794
rect 109 760 4376 794
rect 4410 760 4448 794
rect 59 744 4482 760
rect 5200 794 5358 810
rect 5200 760 5238 794
rect 5272 760 5308 794
rect 5344 760 5358 794
rect -45 652 -11 686
rect -45 584 -11 618
rect -45 516 -11 550
rect 59 668 4482 684
rect 59 634 75 668
rect 109 634 4376 668
rect 4410 634 4448 668
rect 59 618 4482 634
rect 5200 668 5358 760
rect 5471 794 10770 810
rect 5471 791 5487 794
rect 5521 791 10720 794
rect 10754 791 10770 794
rect 5471 757 5485 791
rect 5521 760 5557 791
rect 5519 757 5557 760
rect 5591 757 10650 791
rect 10684 760 10720 791
rect 10684 757 10722 760
rect 10756 757 10770 791
rect 5471 744 10770 757
rect 10845 800 10879 834
rect 5200 634 5238 668
rect 5272 634 5308 668
rect 5344 634 5358 668
rect 10845 667 10879 766
rect 5200 618 5358 634
rect 5428 633 5483 667
rect 5517 633 5541 667
rect 5590 633 5609 667
rect 5663 633 5677 667
rect 5736 633 5745 667
rect 5809 633 5813 667
rect 5847 633 5848 667
rect 5915 633 5920 667
rect 5983 633 5992 667
rect 6051 633 6064 667
rect 6119 633 6136 667
rect 6187 633 6208 667
rect 6255 633 6280 667
rect 6323 633 6352 667
rect 6391 633 6424 667
rect 6459 633 6493 667
rect 6530 633 6561 667
rect 6602 633 6629 667
rect 6674 633 6697 667
rect 6746 633 6765 667
rect 6818 633 6833 667
rect 6890 633 6901 667
rect 6962 633 6969 667
rect 7034 633 7037 667
rect 7071 633 7072 667
rect 7139 633 7144 667
rect 7207 633 7216 667
rect 7275 633 7288 667
rect 7343 633 7360 667
rect 7411 633 7432 667
rect 7479 633 7504 667
rect 7547 633 7576 667
rect 7615 633 7648 667
rect 7683 633 7717 667
rect 7754 633 7785 667
rect 7826 633 7853 667
rect 7898 633 7921 667
rect 7970 633 7989 667
rect 8042 633 8057 667
rect 8114 633 8125 667
rect 8186 633 8193 667
rect 8258 633 8261 667
rect 8295 633 8296 667
rect 8363 633 8368 667
rect 8431 633 8440 667
rect 8499 633 8512 667
rect 8567 633 8584 667
rect 8635 633 8656 667
rect 8703 633 8728 667
rect 8771 633 8800 667
rect 8839 633 8872 667
rect 8907 633 8941 667
rect 8978 633 9009 667
rect 9050 633 9077 667
rect 9122 633 9145 667
rect 9194 633 9213 667
rect 9266 633 9281 667
rect 9338 633 9349 667
rect 9410 633 9417 667
rect 9482 633 9485 667
rect 9519 633 9520 667
rect 9587 633 9592 667
rect 9655 633 9664 667
rect 9723 633 9736 667
rect 9791 633 9808 667
rect 9859 633 9880 667
rect 9927 633 9952 667
rect 9995 633 10024 667
rect 10063 633 10096 667
rect 10131 633 10165 667
rect 10202 633 10233 667
rect 10274 633 10301 667
rect 10346 633 10369 667
rect 10418 633 10437 667
rect 10490 633 10505 667
rect 10562 633 10573 667
rect 10634 633 10641 667
rect 10706 633 10709 667
rect 10743 633 10744 667
rect 10811 633 10816 667
rect 10850 633 10879 667
rect 59 558 193 618
rect 5428 599 5462 633
rect 59 542 4482 558
rect 59 508 75 542
rect 109 508 4376 542
rect 4410 508 4448 542
rect 59 492 4482 508
rect 5200 542 5358 558
rect 5200 508 5238 542
rect 5272 508 5308 542
rect 5344 508 5358 542
rect -45 448 -11 482
rect -45 380 -11 414
rect -45 312 -11 346
rect -45 244 -11 278
rect 59 416 4482 432
rect 59 382 75 416
rect 109 382 4376 416
rect 4410 382 4448 416
rect 59 366 4482 382
rect 5200 416 5358 508
rect 5200 382 5238 416
rect 5272 382 5308 416
rect 5344 382 5358 416
rect 5200 366 5358 382
rect 5428 531 5462 565
rect 5428 463 5462 497
rect 5428 395 5462 429
rect 59 306 193 366
rect 5428 327 5462 361
rect 59 290 4482 306
rect 59 256 75 290
rect 109 256 4376 290
rect 4410 256 4448 290
rect 59 240 4482 256
rect 5200 290 5358 306
rect 5200 256 5238 290
rect 5272 256 5308 290
rect 5344 256 5358 290
rect 5200 240 5358 256
rect 5428 259 5462 293
rect -45 176 -11 210
rect 5428 191 5462 225
rect -45 108 -11 142
rect 59 164 3648 180
rect 59 130 75 164
rect 109 163 3648 164
rect 5196 164 5358 180
rect 5196 163 5308 164
rect 109 130 3528 163
rect 59 129 3528 130
rect 3562 129 3600 163
rect 3634 129 3648 163
rect 4269 129 4307 163
rect 5196 129 5226 163
rect 5260 129 5298 163
rect 5342 130 5358 164
rect 5332 129 5358 130
rect 59 114 3648 129
rect 5196 114 5358 129
rect 5428 123 5462 157
rect -45 40 -11 74
rect 5428 40 5462 89
rect -45 6 56 40
rect 90 6 124 40
rect 158 6 192 40
rect 226 6 260 40
rect 294 6 328 40
rect 362 6 396 40
rect 430 6 464 40
rect 498 6 532 40
rect 566 6 600 40
rect 634 6 668 40
rect 702 6 736 40
rect 770 6 804 40
rect 838 6 872 40
rect 906 6 940 40
rect 974 6 1008 40
rect 1042 6 1076 40
rect 1110 6 1144 40
rect 1178 6 1212 40
rect 1246 6 1280 40
rect 1314 6 1348 40
rect 1382 6 1416 40
rect 1450 6 1484 40
rect 1518 6 1552 40
rect 1586 6 1620 40
rect 1654 6 1688 40
rect 1722 6 1756 40
rect 1790 6 1824 40
rect 1858 6 1892 40
rect 1926 6 1960 40
rect 1994 6 2028 40
rect 2062 6 2096 40
rect 2130 6 2164 40
rect 2198 6 2232 40
rect 2266 6 2300 40
rect 2334 6 2368 40
rect 2402 6 2436 40
rect 2470 6 2504 40
rect 2538 6 2572 40
rect 2606 6 2640 40
rect 2674 6 2708 40
rect 2742 6 2776 40
rect 2810 6 2844 40
rect 2878 6 2912 40
rect 2946 6 2980 40
rect 3014 6 3048 40
rect 3082 6 3116 40
rect 3150 6 3184 40
rect 3218 6 3252 40
rect 3286 6 3320 40
rect 3354 6 3388 40
rect 3490 6 3496 40
rect 3558 6 3570 40
rect 3626 6 3644 40
rect 3694 6 3718 40
rect 3762 6 3792 40
rect 3830 6 3864 40
rect 3900 6 3932 40
rect 3974 6 4000 40
rect 4048 6 4068 40
rect 4122 6 4136 40
rect 4196 6 4204 40
rect 4270 6 4272 40
rect 4306 6 4310 40
rect 4374 6 4384 40
rect 4442 6 4458 40
rect 4510 6 4532 40
rect 4578 6 4606 40
rect 4646 6 4680 40
rect 4714 6 4748 40
rect 4788 6 4816 40
rect 4862 6 4884 40
rect 4936 6 4952 40
rect 5010 6 5020 40
rect 5084 6 5088 40
rect 5122 6 5124 40
rect 5190 6 5198 40
rect 5258 6 5272 40
rect 5326 6 5347 40
rect 5394 6 5422 40
rect 5456 6 5462 40
<< viali >>
rect 7735 2711 7769 2745
rect 7810 2743 7844 2745
rect 7885 2743 7919 2745
rect 7960 2743 7994 2745
rect 8035 2743 8069 2745
rect 8109 2743 8143 2745
rect 8183 2743 8217 2745
rect 8257 2743 8291 2745
rect 8331 2743 8365 2745
rect 8405 2743 8439 2745
rect 8479 2743 8513 2745
rect 8553 2743 8587 2745
rect 8627 2743 8661 2745
rect 8701 2743 8735 2745
rect 8775 2743 8809 2745
rect 8849 2743 8883 2745
rect 7810 2711 7820 2743
rect 7820 2711 7844 2743
rect 7885 2711 7891 2743
rect 7891 2711 7919 2743
rect 7960 2711 7962 2743
rect 7962 2711 7994 2743
rect 8035 2711 8067 2743
rect 8067 2711 8069 2743
rect 8109 2711 8138 2743
rect 8138 2711 8143 2743
rect 8183 2711 8209 2743
rect 8209 2711 8217 2743
rect 8257 2711 8280 2743
rect 8280 2711 8291 2743
rect 8331 2711 8351 2743
rect 8351 2711 8365 2743
rect 8405 2711 8422 2743
rect 8422 2711 8439 2743
rect 8479 2711 8493 2743
rect 8493 2711 8513 2743
rect 8553 2711 8564 2743
rect 8564 2711 8587 2743
rect 8627 2711 8635 2743
rect 8635 2711 8661 2743
rect 8701 2711 8706 2743
rect 8706 2711 8735 2743
rect 8775 2711 8778 2743
rect 8778 2711 8809 2743
rect 8849 2711 8850 2743
rect 8850 2711 8883 2743
rect 7854 2611 7888 2645
rect 7930 2611 7964 2645
rect 8006 2611 8040 2645
rect 8082 2611 8116 2645
rect 8158 2611 8192 2645
rect 8234 2611 8268 2645
rect 8310 2611 8344 2645
rect 8386 2611 8420 2645
rect 8461 2611 8495 2645
rect 8536 2611 8570 2645
rect 8611 2611 8645 2645
rect 8686 2611 8720 2645
rect 8761 2611 8795 2645
rect 8923 2639 8957 2673
rect 8848 2552 8882 2581
rect 8848 2547 8882 2552
rect 7854 2507 7888 2541
rect 7930 2507 7964 2541
rect 8006 2507 8040 2541
rect 8082 2507 8116 2541
rect 8158 2507 8192 2541
rect 8234 2507 8268 2541
rect 8310 2507 8344 2541
rect 8386 2507 8420 2541
rect 8461 2507 8495 2541
rect 8536 2507 8570 2541
rect 8611 2507 8645 2541
rect 8686 2507 8720 2541
rect 8761 2507 8795 2541
rect 8848 2496 8882 2509
rect 8848 2475 8882 2496
rect 8923 2582 8956 2588
rect 8956 2582 8957 2588
rect 8923 2554 8957 2582
rect 8923 2501 8956 2503
rect 8956 2501 8957 2503
rect 8923 2469 8957 2501
rect 7854 2401 7888 2435
rect 7930 2401 7964 2435
rect 8006 2401 8040 2435
rect 8082 2401 8116 2435
rect 8158 2401 8192 2435
rect 8234 2401 8268 2435
rect 8310 2401 8344 2435
rect 8386 2401 8420 2435
rect 8461 2401 8495 2435
rect 8536 2401 8570 2435
rect 8611 2401 8645 2435
rect 8686 2401 8720 2435
rect 8761 2401 8795 2435
rect 8923 2384 8957 2418
rect 7854 2299 7888 2333
rect 7930 2305 7962 2333
rect 7962 2305 7964 2333
rect 8006 2305 8033 2333
rect 8033 2305 8040 2333
rect 8082 2305 8104 2333
rect 8104 2305 8116 2333
rect 8158 2305 8175 2333
rect 8175 2305 8192 2333
rect 8235 2305 8246 2333
rect 8246 2305 8269 2333
rect 8312 2305 8317 2333
rect 8317 2305 8346 2333
rect 8389 2305 8422 2333
rect 8422 2305 8423 2333
rect 8466 2305 8493 2333
rect 8493 2305 8500 2333
rect 8543 2305 8564 2333
rect 8564 2305 8577 2333
rect 8620 2305 8635 2333
rect 8635 2305 8654 2333
rect 8697 2305 8706 2333
rect 8706 2305 8731 2333
rect 8774 2305 8777 2333
rect 8777 2305 8808 2333
rect 7930 2299 7964 2305
rect 8006 2299 8040 2305
rect 8082 2299 8116 2305
rect 8158 2299 8192 2305
rect 8235 2299 8269 2305
rect 8312 2299 8346 2305
rect 8389 2299 8423 2305
rect 8466 2299 8500 2305
rect 8543 2299 8577 2305
rect 8620 2299 8654 2305
rect 8697 2299 8731 2305
rect 8774 2299 8808 2305
rect 8851 2299 8885 2333
rect 3648 2059 3672 2093
rect 3672 2059 3682 2093
rect 3721 2059 3740 2093
rect 3740 2059 3755 2093
rect 3794 2059 3808 2093
rect 3808 2059 3828 2093
rect 3867 2059 3876 2093
rect 3876 2059 3901 2093
rect 3940 2059 3944 2093
rect 3944 2059 3974 2093
rect 4013 2059 4046 2093
rect 4046 2059 4047 2093
rect 4086 2059 4114 2093
rect 4114 2059 4120 2093
rect 4159 2059 4182 2093
rect 4182 2059 4193 2093
rect 4232 2059 4250 2093
rect 4250 2059 4266 2093
rect 4305 2059 4318 2093
rect 4318 2059 4339 2093
rect 4378 2059 4386 2093
rect 4386 2059 4412 2093
rect 4451 2059 4454 2093
rect 4454 2059 4485 2093
rect 4524 2059 4556 2093
rect 4556 2059 4558 2093
rect 4597 2059 4624 2093
rect 4624 2059 4631 2093
rect 4670 2059 4692 2093
rect 4692 2059 4704 2093
rect 4743 2059 4760 2093
rect 4760 2059 4777 2093
rect 4816 2059 4828 2093
rect 4828 2059 4850 2093
rect 4889 2059 4896 2093
rect 4896 2059 4923 2093
rect 4962 2059 4964 2093
rect 4964 2059 4996 2093
rect 5035 2059 5066 2093
rect 5066 2059 5069 2093
rect 5108 2059 5134 2093
rect 5134 2059 5142 2093
rect 5181 2059 5202 2093
rect 5202 2059 5215 2093
rect 5254 2059 5270 2093
rect 5270 2059 5288 2093
rect 5327 2059 5338 2093
rect 5338 2059 5361 2093
rect 5400 2059 5406 2093
rect 5406 2059 5434 2093
rect 5473 2059 5474 2093
rect 5474 2059 5507 2093
rect 5546 2059 5576 2093
rect 5576 2059 5580 2093
rect 5619 2059 5644 2093
rect 5644 2059 5653 2093
rect 5692 2059 5712 2093
rect 5712 2059 5726 2093
rect 5765 2059 5780 2093
rect 5780 2059 5799 2093
rect 5838 2059 5848 2093
rect 5848 2059 5872 2093
rect 5911 2059 5916 2093
rect 5916 2059 5945 2093
rect 5984 2059 6018 2093
rect 6057 2059 6086 2093
rect 6086 2059 6091 2093
rect 6130 2059 6154 2093
rect 6154 2059 6164 2093
rect 6203 2059 6222 2093
rect 6222 2059 6237 2093
rect 6276 2059 6290 2093
rect 6290 2059 6310 2093
rect 6349 2059 6358 2093
rect 6358 2059 6383 2093
rect 6422 2059 6426 2093
rect 6426 2059 6456 2093
rect 6495 2059 6528 2093
rect 6528 2059 6529 2093
rect 6568 2059 6596 2093
rect 6596 2059 6602 2093
rect 6641 2059 6664 2093
rect 6664 2059 6675 2093
rect 6714 2059 6732 2093
rect 6732 2059 6748 2093
rect 6787 2059 6800 2093
rect 6800 2059 6821 2093
rect 6861 2059 6868 2093
rect 6868 2059 6895 2093
rect 6935 2059 6936 2093
rect 6936 2059 6969 2093
rect 7009 2059 7038 2093
rect 7038 2059 7043 2093
rect 7083 2059 7106 2093
rect 7106 2059 7117 2093
rect 7157 2059 7174 2093
rect 7174 2059 7191 2093
rect 7231 2059 7242 2093
rect 7242 2059 7265 2093
rect 7305 2059 7310 2093
rect 7310 2059 7339 2093
rect 7379 2059 7412 2093
rect 7412 2059 7413 2093
rect 8698 2059 8704 2093
rect 8704 2059 8732 2093
rect 8770 2059 8772 2093
rect 8772 2059 8804 2093
rect 8842 2059 8874 2093
rect 8874 2059 8876 2093
rect 8914 2059 8942 2093
rect 8942 2059 8948 2093
rect 8987 2059 9010 2093
rect 9010 2059 9021 2093
rect 9060 2059 9078 2093
rect 9078 2059 9094 2093
rect 3536 2021 3570 2055
rect 3536 1932 3570 1965
rect 3536 1931 3570 1932
rect 7602 1898 7636 1932
rect 7674 1898 7708 1932
rect 3536 1864 3570 1875
rect 3536 1841 3570 1864
rect 3536 1762 3570 1785
rect 3729 1775 3731 1806
rect 3731 1775 3763 1806
rect 3729 1772 3763 1775
rect 3801 1772 3835 1806
rect 4572 1772 4606 1806
rect 4644 1772 4678 1806
rect 5474 1772 5508 1806
rect 5546 1772 5580 1806
rect 6376 1772 6410 1806
rect 6448 1772 6482 1806
rect 7635 1772 7669 1806
rect 7707 1772 7741 1806
rect 8894 1772 8928 1806
rect 8966 1775 8998 1806
rect 8998 1775 9000 1806
rect 8966 1772 9000 1775
rect 3536 1751 3570 1762
rect 3536 1524 3570 1547
rect 3536 1513 3570 1524
rect 4672 1646 4706 1680
rect 4744 1646 4778 1680
rect 5117 1646 5151 1680
rect 5189 1646 5223 1680
rect 6376 1646 6410 1680
rect 6448 1646 6482 1680
rect 7635 1646 7669 1680
rect 7707 1646 7741 1680
rect 8894 1650 8928 1684
rect 8966 1683 9000 1684
rect 8966 1650 8998 1683
rect 8998 1650 9000 1683
rect 4672 1523 4706 1557
rect 4744 1523 4778 1557
rect 5117 1522 5151 1556
rect 5189 1522 5223 1556
rect 6376 1523 6410 1557
rect 6448 1523 6482 1557
rect 7635 1521 7669 1555
rect 7707 1521 7741 1555
rect 8894 1522 8928 1556
rect 8966 1523 8998 1556
rect 8998 1523 9000 1556
rect 8966 1522 9000 1523
rect 3422 1388 3423 1422
rect 3423 1388 3456 1422
rect 3498 1388 3532 1422
rect 5485 1390 5487 1421
rect 5487 1390 5519 1421
rect 5485 1387 5519 1390
rect 5557 1387 5591 1421
rect 3528 1269 3562 1303
rect 3600 1269 3634 1303
rect 4235 1269 4269 1303
rect 4307 1269 4341 1303
rect 5221 1269 5255 1303
rect 5293 1298 5327 1303
rect 5293 1269 5308 1298
rect 5308 1269 5327 1298
rect 10650 1387 10684 1421
rect 10722 1390 10754 1421
rect 10754 1390 10756 1421
rect 10722 1387 10756 1390
rect 5485 1264 5487 1296
rect 5487 1264 5519 1296
rect 5485 1262 5519 1264
rect 5557 1262 5591 1296
rect 10650 1265 10684 1299
rect 10722 1298 10756 1299
rect 10722 1265 10754 1298
rect 10754 1265 10756 1298
rect 4376 1138 4410 1172
rect 4448 1138 4482 1172
rect 5238 1138 5272 1172
rect 5310 1138 5342 1172
rect 5342 1138 5344 1172
rect 5485 1138 5487 1169
rect 5487 1138 5519 1169
rect 5485 1135 5519 1138
rect 5557 1135 5591 1169
rect 10650 1135 10684 1169
rect 10722 1138 10754 1169
rect 10754 1138 10756 1169
rect 10722 1135 10756 1138
rect 4376 1012 4410 1046
rect 4448 1012 4482 1046
rect 5238 1012 5272 1046
rect 5310 1012 5342 1046
rect 5342 1012 5344 1046
rect 5485 1012 5487 1043
rect 5487 1012 5519 1043
rect 5485 1009 5519 1012
rect 5557 1009 5591 1043
rect 10650 1009 10684 1043
rect 10722 1012 10754 1043
rect 10754 1012 10756 1043
rect 10722 1009 10756 1012
rect 4376 886 4410 920
rect 4448 886 4482 920
rect 5238 886 5272 920
rect 5310 886 5342 920
rect 5342 886 5344 920
rect 5485 886 5487 917
rect 5487 886 5519 917
rect 5485 883 5519 886
rect 5557 883 5591 917
rect 10650 883 10684 917
rect 10722 886 10754 917
rect 10754 886 10756 917
rect 10722 883 10756 886
rect 4376 760 4410 794
rect 4448 760 4482 794
rect 5238 760 5272 794
rect 5310 760 5342 794
rect 5342 760 5344 794
rect 4376 634 4410 668
rect 4448 634 4482 668
rect 5485 760 5487 791
rect 5487 760 5519 791
rect 5485 757 5519 760
rect 5557 757 5591 791
rect 10650 757 10684 791
rect 10722 760 10754 791
rect 10754 760 10756 791
rect 10722 757 10756 760
rect 5238 634 5272 668
rect 5310 634 5342 668
rect 5342 634 5344 668
rect 5483 633 5517 667
rect 5556 633 5575 667
rect 5575 633 5590 667
rect 5629 633 5643 667
rect 5643 633 5663 667
rect 5702 633 5711 667
rect 5711 633 5736 667
rect 5775 633 5779 667
rect 5779 633 5809 667
rect 5848 633 5881 667
rect 5881 633 5882 667
rect 5920 633 5949 667
rect 5949 633 5954 667
rect 5992 633 6017 667
rect 6017 633 6026 667
rect 6064 633 6085 667
rect 6085 633 6098 667
rect 6136 633 6153 667
rect 6153 633 6170 667
rect 6208 633 6221 667
rect 6221 633 6242 667
rect 6280 633 6289 667
rect 6289 633 6314 667
rect 6352 633 6357 667
rect 6357 633 6386 667
rect 6424 633 6425 667
rect 6425 633 6458 667
rect 6496 633 6527 667
rect 6527 633 6530 667
rect 6568 633 6595 667
rect 6595 633 6602 667
rect 6640 633 6663 667
rect 6663 633 6674 667
rect 6712 633 6731 667
rect 6731 633 6746 667
rect 6784 633 6799 667
rect 6799 633 6818 667
rect 6856 633 6867 667
rect 6867 633 6890 667
rect 6928 633 6935 667
rect 6935 633 6962 667
rect 7000 633 7003 667
rect 7003 633 7034 667
rect 7072 633 7105 667
rect 7105 633 7106 667
rect 7144 633 7173 667
rect 7173 633 7178 667
rect 7216 633 7241 667
rect 7241 633 7250 667
rect 7288 633 7309 667
rect 7309 633 7322 667
rect 7360 633 7377 667
rect 7377 633 7394 667
rect 7432 633 7445 667
rect 7445 633 7466 667
rect 7504 633 7513 667
rect 7513 633 7538 667
rect 7576 633 7581 667
rect 7581 633 7610 667
rect 7648 633 7649 667
rect 7649 633 7682 667
rect 7720 633 7751 667
rect 7751 633 7754 667
rect 7792 633 7819 667
rect 7819 633 7826 667
rect 7864 633 7887 667
rect 7887 633 7898 667
rect 7936 633 7955 667
rect 7955 633 7970 667
rect 8008 633 8023 667
rect 8023 633 8042 667
rect 8080 633 8091 667
rect 8091 633 8114 667
rect 8152 633 8159 667
rect 8159 633 8186 667
rect 8224 633 8227 667
rect 8227 633 8258 667
rect 8296 633 8329 667
rect 8329 633 8330 667
rect 8368 633 8397 667
rect 8397 633 8402 667
rect 8440 633 8465 667
rect 8465 633 8474 667
rect 8512 633 8533 667
rect 8533 633 8546 667
rect 8584 633 8601 667
rect 8601 633 8618 667
rect 8656 633 8669 667
rect 8669 633 8690 667
rect 8728 633 8737 667
rect 8737 633 8762 667
rect 8800 633 8805 667
rect 8805 633 8834 667
rect 8872 633 8873 667
rect 8873 633 8906 667
rect 8944 633 8975 667
rect 8975 633 8978 667
rect 9016 633 9043 667
rect 9043 633 9050 667
rect 9088 633 9111 667
rect 9111 633 9122 667
rect 9160 633 9179 667
rect 9179 633 9194 667
rect 9232 633 9247 667
rect 9247 633 9266 667
rect 9304 633 9315 667
rect 9315 633 9338 667
rect 9376 633 9383 667
rect 9383 633 9410 667
rect 9448 633 9451 667
rect 9451 633 9482 667
rect 9520 633 9553 667
rect 9553 633 9554 667
rect 9592 633 9621 667
rect 9621 633 9626 667
rect 9664 633 9689 667
rect 9689 633 9698 667
rect 9736 633 9757 667
rect 9757 633 9770 667
rect 9808 633 9825 667
rect 9825 633 9842 667
rect 9880 633 9893 667
rect 9893 633 9914 667
rect 9952 633 9961 667
rect 9961 633 9986 667
rect 10024 633 10029 667
rect 10029 633 10058 667
rect 10096 633 10097 667
rect 10097 633 10130 667
rect 10168 633 10199 667
rect 10199 633 10202 667
rect 10240 633 10267 667
rect 10267 633 10274 667
rect 10312 633 10335 667
rect 10335 633 10346 667
rect 10384 633 10403 667
rect 10403 633 10418 667
rect 10456 633 10471 667
rect 10471 633 10490 667
rect 10528 633 10539 667
rect 10539 633 10562 667
rect 10600 633 10607 667
rect 10607 633 10634 667
rect 10672 633 10675 667
rect 10675 633 10706 667
rect 10744 633 10777 667
rect 10777 633 10778 667
rect 10816 633 10850 667
rect 4376 508 4410 542
rect 4448 508 4482 542
rect 5238 508 5272 542
rect 5310 508 5342 542
rect 5342 508 5344 542
rect 4376 382 4410 416
rect 4448 382 4482 416
rect 5238 382 5272 416
rect 5310 382 5342 416
rect 5342 382 5344 416
rect 4376 256 4410 290
rect 4448 256 4482 290
rect 5238 256 5272 290
rect 5310 256 5342 290
rect 5342 256 5344 290
rect 3528 129 3562 163
rect 3600 129 3634 163
rect 4235 129 4269 163
rect 4307 129 4341 163
rect 5226 129 5260 163
rect 5298 130 5308 163
rect 5308 130 5332 163
rect 5298 129 5332 130
rect 3422 6 3456 40
rect 3496 6 3524 40
rect 3524 6 3530 40
rect 3570 6 3592 40
rect 3592 6 3604 40
rect 3644 6 3660 40
rect 3660 6 3678 40
rect 3718 6 3728 40
rect 3728 6 3752 40
rect 3792 6 3796 40
rect 3796 6 3826 40
rect 3866 6 3898 40
rect 3898 6 3900 40
rect 3940 6 3966 40
rect 3966 6 3974 40
rect 4014 6 4034 40
rect 4034 6 4048 40
rect 4088 6 4102 40
rect 4102 6 4122 40
rect 4162 6 4170 40
rect 4170 6 4196 40
rect 4236 6 4238 40
rect 4238 6 4270 40
rect 4310 6 4340 40
rect 4340 6 4344 40
rect 4384 6 4408 40
rect 4408 6 4418 40
rect 4458 6 4476 40
rect 4476 6 4492 40
rect 4532 6 4544 40
rect 4544 6 4566 40
rect 4606 6 4612 40
rect 4612 6 4640 40
rect 4680 6 4714 40
rect 4754 6 4782 40
rect 4782 6 4788 40
rect 4828 6 4850 40
rect 4850 6 4862 40
rect 4902 6 4918 40
rect 4918 6 4936 40
rect 4976 6 4986 40
rect 4986 6 5010 40
rect 5050 6 5054 40
rect 5054 6 5084 40
rect 5124 6 5156 40
rect 5156 6 5158 40
rect 5198 6 5224 40
rect 5224 6 5232 40
rect 5272 6 5292 40
rect 5292 6 5306 40
rect 5347 6 5360 40
rect 5360 6 5381 40
rect 5422 6 5456 40
<< metal1 >>
rect 7723 2745 8963 2751
rect 7723 2711 7735 2745
rect 7769 2711 7810 2745
rect 7844 2711 7885 2745
rect 7919 2711 7960 2745
rect 7994 2711 8035 2745
rect 8069 2711 8109 2745
rect 8143 2711 8183 2745
rect 8217 2711 8257 2745
rect 8291 2711 8331 2745
rect 8365 2711 8405 2745
rect 8439 2711 8479 2745
rect 8513 2711 8553 2745
rect 8587 2711 8627 2745
rect 8661 2711 8701 2745
rect 8735 2711 8775 2745
rect 8809 2711 8849 2745
rect 8883 2711 8963 2745
rect 7723 2705 8963 2711
rect 7723 2645 8807 2705
rect 7723 2611 7854 2645
rect 7888 2611 7930 2645
rect 7964 2611 8006 2645
rect 8040 2611 8082 2645
rect 8116 2611 8158 2645
rect 8192 2611 8234 2645
rect 8268 2611 8310 2645
rect 8344 2611 8386 2645
rect 8420 2611 8461 2645
rect 8495 2611 8536 2645
rect 8570 2611 8611 2645
rect 8645 2611 8686 2645
rect 8720 2611 8761 2645
rect 8795 2611 8807 2645
rect 7723 2605 8807 2611
rect 8917 2673 8963 2705
rect 8917 2639 8923 2673
rect 8957 2639 8963 2673
rect 8842 2581 8888 2593
rect 8842 2547 8848 2581
rect 8882 2547 8888 2581
tri 7676 2541 7682 2547 se
rect 7682 2541 8807 2547
tri 7642 2507 7676 2541 se
rect 7676 2507 7854 2541
rect 7888 2507 7930 2541
rect 7964 2507 8006 2541
rect 8040 2507 8082 2541
rect 8116 2507 8158 2541
rect 8192 2507 8234 2541
rect 8268 2507 8310 2541
rect 8344 2507 8386 2541
rect 8420 2507 8461 2541
rect 8495 2507 8536 2541
rect 8570 2507 8611 2541
rect 8645 2507 8686 2541
rect 8720 2507 8761 2541
rect 8795 2507 8807 2541
tri 7616 2481 7642 2507 se
rect 7642 2501 8807 2507
rect 8842 2509 8888 2547
rect 7642 2481 7682 2501
tri 7682 2481 7702 2501 nw
tri 7610 2475 7616 2481 se
rect 7616 2475 7676 2481
tri 7676 2475 7682 2481 nw
rect 8842 2475 8848 2509
rect 8882 2475 8888 2509
tri 7604 2469 7610 2475 se
rect 7610 2469 7670 2475
tri 7670 2469 7676 2475 nw
tri 7570 2435 7604 2469 se
rect 7604 2435 7636 2469
tri 7636 2435 7670 2469 nw
rect 8842 2463 8888 2475
rect 8917 2588 8963 2639
rect 8917 2554 8923 2588
rect 8957 2554 8963 2588
rect 8917 2503 8963 2554
rect 8917 2469 8923 2503
rect 8957 2469 8963 2503
rect 7842 2435 8807 2441
tri 7550 2415 7570 2435 se
rect 7570 2415 7616 2435
tri 7616 2415 7636 2435 nw
tri 7536 2401 7550 2415 se
rect 7550 2401 7602 2415
tri 7602 2401 7616 2415 nw
rect 7842 2401 7854 2435
rect 7888 2401 7930 2435
rect 7964 2401 8006 2435
rect 8040 2401 8082 2435
rect 8116 2401 8158 2435
rect 8192 2401 8234 2435
rect 8268 2401 8310 2435
rect 8344 2401 8386 2435
rect 8420 2401 8461 2435
rect 8495 2401 8536 2435
rect 8570 2401 8611 2435
rect 8645 2401 8686 2435
rect 8720 2401 8761 2435
rect 8795 2401 8807 2435
tri 7519 2384 7536 2401 se
rect 7536 2384 7585 2401
tri 7585 2384 7602 2401 nw
tri 7504 2369 7519 2384 se
rect 7519 2369 7550 2384
tri 3539 2099 3545 2105 se
rect 3545 2099 3551 2105
rect 3530 2055 3551 2099
rect 3530 2021 3536 2055
rect 3603 2053 3615 2105
rect 3667 2093 3679 2105
rect 3731 2099 3737 2105
tri 3737 2099 3743 2105 sw
tri 4179 2099 4185 2105 se
rect 4185 2099 4191 2105
rect 3731 2093 4191 2099
rect 4243 2093 4256 2105
rect 4308 2093 4321 2105
rect 4373 2093 4386 2105
rect 3755 2059 3794 2093
rect 3828 2059 3867 2093
rect 3901 2059 3940 2093
rect 3974 2059 4013 2093
rect 4047 2059 4086 2093
rect 4120 2059 4159 2093
rect 4373 2059 4378 2093
rect 3667 2053 3679 2059
rect 3731 2053 4191 2059
rect 4243 2053 4256 2059
rect 4308 2053 4321 2059
rect 4373 2053 4386 2059
rect 4438 2053 4450 2105
rect 4502 2053 4514 2105
rect 4566 2053 4578 2105
rect 4630 2099 4636 2105
tri 4636 2099 4642 2105 sw
rect 4630 2093 7425 2099
rect 4631 2059 4670 2093
rect 4704 2059 4743 2093
rect 4777 2059 4816 2093
rect 4850 2059 4889 2093
rect 4923 2059 4962 2093
rect 4996 2059 5035 2093
rect 5069 2059 5108 2093
rect 5142 2059 5181 2093
rect 5215 2059 5254 2093
rect 5288 2059 5327 2093
rect 5361 2059 5400 2093
rect 5434 2059 5473 2093
rect 5507 2059 5546 2093
rect 5580 2059 5619 2093
rect 5653 2059 5692 2093
rect 5726 2059 5765 2093
rect 5799 2059 5838 2093
rect 5872 2059 5911 2093
rect 5945 2059 5984 2093
rect 6018 2059 6057 2093
rect 6091 2059 6130 2093
rect 6164 2059 6203 2093
rect 6237 2059 6276 2093
rect 6310 2059 6349 2093
rect 6383 2059 6422 2093
rect 6456 2059 6495 2093
rect 6529 2059 6568 2093
rect 6602 2059 6641 2093
rect 6675 2059 6714 2093
rect 6748 2059 6787 2093
rect 6821 2059 6861 2093
rect 6895 2059 6935 2093
rect 6969 2059 7009 2093
rect 7043 2059 7083 2093
rect 7117 2059 7157 2093
rect 7191 2059 7231 2093
rect 7265 2059 7305 2093
rect 7339 2059 7379 2093
rect 7413 2059 7425 2093
tri 7472 2059 7504 2091 se
rect 7504 2071 7550 2369
tri 7550 2349 7585 2384 nw
rect 7842 2339 8807 2401
rect 8917 2418 8963 2469
rect 8917 2384 8923 2418
rect 8957 2384 8963 2418
rect 8917 2339 8963 2384
rect 7842 2333 8963 2339
rect 7842 2299 7854 2333
rect 7888 2299 7930 2333
rect 7964 2299 8006 2333
rect 8040 2299 8082 2333
rect 8116 2299 8158 2333
rect 8192 2299 8235 2333
rect 8269 2299 8312 2333
rect 8346 2299 8389 2333
rect 8423 2299 8466 2333
rect 8500 2299 8543 2333
rect 8577 2299 8620 2333
rect 8654 2299 8697 2333
rect 8731 2299 8774 2333
rect 8808 2299 8851 2333
rect 8885 2299 8963 2333
rect 7842 2293 8963 2299
rect 7504 2059 7538 2071
tri 7538 2059 7550 2071 nw
rect 4630 2053 7425 2059
tri 7466 2053 7472 2059 se
rect 7472 2053 7504 2059
rect 3570 2021 3576 2053
tri 7438 2025 7466 2053 se
rect 7466 2025 7504 2053
tri 7504 2025 7538 2059 nw
tri 7436 2023 7438 2025 se
rect 7438 2023 7456 2025
rect 3530 1965 3576 2021
rect 3530 1931 3536 1965
rect 3570 1931 3576 1965
rect 3530 1875 3576 1931
rect 3530 1841 3536 1875
rect 3570 1841 3576 1875
rect 3530 1785 3576 1841
rect 3530 1751 3536 1785
rect 3570 1751 3576 1785
rect 3713 1977 7456 2023
tri 7456 1977 7504 2025 nw
rect 3713 1818 3759 1977
tri 3759 1943 3793 1977 nw
rect 8379 1938 8425 2293
rect 8686 2093 9106 2099
rect 8686 2059 8698 2093
rect 8732 2059 8770 2093
rect 8804 2059 8842 2093
rect 8876 2059 8914 2093
rect 8948 2059 8987 2093
rect 9021 2059 9060 2093
rect 9094 2059 9106 2093
rect 8686 2053 9106 2059
rect 7590 1932 8111 1938
rect 7590 1898 7602 1932
rect 7636 1898 7674 1932
rect 7708 1898 8111 1932
rect 7590 1892 8111 1898
rect 8345 1892 9221 1938
tri 3759 1818 3793 1852 sw
rect 3713 1806 4294 1818
rect 3713 1772 3729 1806
rect 3763 1772 3801 1806
rect 3835 1772 4294 1806
rect 3713 1766 4294 1772
rect 4295 1767 4296 1817
rect 4332 1767 4333 1817
rect 4334 1806 5302 1818
rect 5304 1817 5340 1818
rect 4334 1772 4572 1806
rect 4606 1772 4644 1806
rect 4678 1772 5302 1806
rect 4334 1766 5302 1772
rect 5303 1767 5341 1817
rect 5342 1806 6204 1818
rect 6206 1817 6242 1818
rect 5342 1772 5474 1806
rect 5508 1772 5546 1806
rect 5580 1772 6204 1806
rect 5304 1766 5340 1767
rect 5342 1766 6204 1772
rect 6205 1767 6243 1817
rect 6244 1806 7463 1818
rect 7465 1817 7501 1818
rect 6244 1772 6376 1806
rect 6410 1772 6448 1806
rect 6482 1772 7463 1806
rect 6206 1766 6242 1767
rect 6244 1766 7463 1772
rect 7464 1767 7502 1817
rect 7503 1806 8422 1818
rect 8424 1817 8460 1818
rect 7503 1772 7635 1806
rect 7669 1772 7707 1806
rect 7741 1772 8422 1806
rect 7465 1766 7501 1767
rect 7503 1766 8422 1772
rect 8423 1767 8461 1817
rect 8462 1806 9013 1818
rect 8462 1772 8894 1806
rect 8928 1772 8966 1806
rect 9000 1772 9013 1806
rect 8424 1766 8460 1767
rect 8462 1766 9013 1772
rect 3530 1739 3576 1751
rect 4660 1680 4926 1692
rect 4928 1691 4964 1692
rect 4660 1646 4672 1680
rect 4706 1646 4744 1680
rect 4778 1646 4926 1680
rect 4660 1640 4926 1646
rect 4927 1641 4965 1691
rect 4966 1680 6185 1692
rect 6187 1691 6223 1692
rect 4966 1646 5117 1680
rect 5151 1646 5189 1680
rect 5223 1646 6185 1680
rect 4928 1640 4964 1641
rect 4966 1640 6185 1646
rect 6186 1641 6224 1691
rect 6225 1680 7474 1692
rect 7476 1691 7512 1692
rect 6225 1646 6376 1680
rect 6410 1646 6448 1680
rect 6482 1646 7474 1680
rect 6187 1640 6223 1641
rect 6225 1640 7474 1646
rect 7475 1641 7513 1691
rect 7514 1680 8419 1692
rect 8421 1691 8457 1692
rect 7514 1646 7635 1680
rect 7669 1646 7707 1680
rect 7741 1646 8419 1680
rect 7476 1640 7512 1641
rect 7514 1640 8419 1646
rect 8420 1641 8458 1691
rect 8459 1684 9012 1692
rect 8459 1650 8894 1684
rect 8928 1650 8966 1684
rect 9000 1650 9012 1684
rect 8421 1640 8457 1641
rect 8459 1640 9012 1650
rect 3530 1547 3576 1559
rect 3530 1513 3536 1547
rect 3570 1513 3576 1547
rect 4660 1557 4926 1567
rect 4928 1566 4964 1567
rect 4660 1523 4672 1557
rect 4706 1523 4744 1557
rect 4778 1523 4926 1557
rect 4660 1515 4926 1523
rect 4927 1516 4965 1566
rect 4966 1556 6185 1567
rect 6187 1566 6223 1567
rect 4966 1522 5117 1556
rect 5151 1522 5189 1556
rect 5223 1522 6185 1556
rect 4928 1515 4964 1516
rect 4966 1515 6185 1522
rect 6186 1516 6224 1566
rect 6225 1557 7474 1567
rect 6225 1523 6376 1557
rect 6410 1523 6448 1557
rect 6482 1523 7474 1557
rect 6187 1515 6223 1516
rect 6225 1515 7474 1523
rect 7475 1516 7476 1566
rect 7512 1516 7513 1566
rect 7514 1555 8419 1567
rect 7514 1521 7635 1555
rect 7669 1521 7707 1555
rect 7741 1521 8419 1555
rect 7514 1515 8419 1521
rect 8420 1516 8421 1566
rect 8457 1516 8458 1566
rect 8459 1556 9012 1567
rect 8459 1522 8894 1556
rect 8928 1522 8966 1556
rect 9000 1522 9012 1556
rect 8459 1515 9012 1522
rect 9175 1552 9221 1892
rect 10118 1552 10124 1558
rect 3530 1428 3576 1513
rect 9175 1506 10124 1552
rect 10176 1506 10196 1558
rect 10248 1506 10268 1558
rect 10320 1506 10340 1558
rect 10392 1506 10412 1558
rect 10464 1506 10470 1558
tri 3356 1422 3362 1428 se
rect 3362 1422 3576 1428
tri 3322 1388 3356 1422 se
rect 3356 1388 3422 1422
rect 3456 1388 3498 1422
rect 3532 1388 3576 1422
tri 3321 1387 3322 1388 se
rect 3322 1387 3576 1388
tri 3292 1358 3321 1387 se
rect 3321 1382 3576 1387
rect 5472 1421 6023 1432
rect 5472 1387 5485 1421
rect 5519 1387 5557 1421
rect 5591 1387 6023 1421
rect 3321 1358 3388 1382
rect 3292 129 3388 1358
tri 3388 1338 3432 1382 nw
rect 5472 1380 6023 1387
rect 6024 1381 6025 1431
rect 6061 1381 6062 1431
rect 6063 1421 10768 1432
rect 6063 1387 10650 1421
rect 10684 1387 10722 1421
rect 10756 1387 10768 1421
rect 6063 1380 10768 1387
rect 3516 1303 5438 1309
rect 3516 1269 3528 1303
rect 3562 1269 3600 1303
rect 3634 1269 4235 1303
rect 4269 1269 4307 1303
rect 4341 1269 5221 1303
rect 5255 1269 5293 1303
rect 5327 1269 5438 1303
rect 3516 1263 5438 1269
tri 4227 1262 4228 1263 ne
rect 4228 1262 4346 1263
tri 4346 1262 4347 1263 nw
tri 5358 1262 5359 1263 ne
rect 5359 1262 5438 1263
tri 4228 1229 4261 1262 ne
rect 4261 169 4313 1262
tri 4313 1229 4346 1262 nw
tri 5359 1229 5392 1262 ne
rect 4364 1172 4759 1182
rect 4364 1138 4376 1172
rect 4410 1138 4448 1172
rect 4482 1138 4759 1172
rect 4364 1130 4759 1138
rect 4760 1131 4761 1181
rect 4797 1131 4798 1181
rect 4799 1172 5356 1182
rect 4799 1138 5238 1172
rect 5272 1138 5310 1172
rect 5344 1138 5356 1172
rect 4799 1130 5356 1138
rect 4364 1046 4759 1054
rect 4364 1012 4376 1046
rect 4410 1012 4448 1046
rect 4482 1012 4759 1046
rect 4364 1002 4759 1012
rect 4760 1003 4761 1053
rect 4797 1003 4798 1053
rect 4799 1046 5356 1054
rect 4799 1012 5238 1046
rect 5272 1012 5310 1046
rect 5344 1012 5356 1046
rect 4799 1002 5356 1012
rect 4364 920 4763 928
rect 4364 886 4376 920
rect 4410 886 4448 920
rect 4482 886 4763 920
rect 4364 876 4763 886
rect 4764 877 4765 927
rect 4801 877 4802 927
rect 4803 920 5356 928
rect 4803 886 5238 920
rect 5272 886 5310 920
rect 5344 886 5356 920
rect 4803 876 5356 886
rect 4364 794 4763 802
rect 4364 760 4376 794
rect 4410 760 4448 794
rect 4482 760 4763 794
rect 4364 750 4763 760
rect 4764 751 4765 801
rect 4801 751 4802 801
rect 4803 794 5356 802
rect 4803 760 5238 794
rect 5272 760 5310 794
rect 5344 760 5356 794
rect 4803 750 5356 760
rect 5392 797 5438 1262
rect 5473 1296 6024 1308
rect 5473 1262 5485 1296
rect 5519 1262 5557 1296
rect 5591 1262 6024 1296
rect 5473 1256 6024 1262
rect 6025 1257 6026 1307
rect 6062 1257 6063 1307
rect 6064 1299 10768 1308
rect 6064 1265 10650 1299
rect 10684 1265 10722 1299
rect 10756 1265 10768 1299
rect 6064 1256 10768 1265
rect 5472 1169 6024 1178
rect 5472 1135 5485 1169
rect 5519 1135 5557 1169
rect 5591 1135 6024 1169
rect 5472 1126 6024 1135
rect 6025 1127 6026 1177
rect 6062 1127 6063 1177
rect 6064 1169 10768 1178
rect 6064 1135 10650 1169
rect 10684 1135 10722 1169
rect 10756 1135 10768 1169
rect 6064 1126 10768 1135
rect 5472 1043 6024 1055
rect 5472 1009 5485 1043
rect 5519 1009 5557 1043
rect 5591 1009 6024 1043
rect 5472 1003 6024 1009
rect 6025 1004 6026 1054
rect 6062 1004 6063 1054
rect 6064 1043 10768 1055
rect 6064 1009 10650 1043
rect 10684 1009 10722 1043
rect 10756 1009 10768 1043
rect 6064 1003 10768 1009
rect 5472 917 6024 929
rect 5472 883 5485 917
rect 5519 883 5557 917
rect 5591 883 6024 917
rect 5472 877 6024 883
rect 6025 878 6026 928
rect 6062 878 6063 928
rect 6064 917 10768 929
rect 6064 883 10650 917
rect 10684 883 10722 917
rect 10756 883 10768 917
rect 6064 877 10768 883
tri 5438 797 5472 831 sw
rect 5392 791 10768 797
rect 5392 757 5485 791
rect 5519 757 5557 791
rect 5591 757 10650 791
rect 10684 757 10722 791
rect 10756 757 10768 791
rect 5392 751 10768 757
rect 4364 668 4764 678
rect 4364 634 4376 668
rect 4410 634 4448 668
rect 4482 634 4764 668
rect 4364 626 4764 634
rect 4765 627 4766 677
rect 4802 627 4803 677
rect 4804 668 5356 678
rect 4804 634 5238 668
rect 5272 634 5310 668
rect 5344 634 5356 668
rect 4804 626 5356 634
rect 5471 667 10862 673
rect 5471 633 5483 667
rect 5517 633 5556 667
rect 5590 633 5629 667
rect 5663 633 5702 667
rect 5736 633 5775 667
rect 5809 633 5848 667
rect 5882 633 5920 667
rect 5954 633 5992 667
rect 6026 633 6064 667
rect 6098 633 6136 667
rect 6170 633 6208 667
rect 6242 633 6280 667
rect 6314 633 6352 667
rect 6386 633 6424 667
rect 6458 633 6496 667
rect 6530 633 6568 667
rect 6602 633 6640 667
rect 6674 633 6712 667
rect 6746 633 6784 667
rect 6818 633 6856 667
rect 6890 633 6928 667
rect 6962 633 7000 667
rect 7034 633 7072 667
rect 7106 633 7144 667
rect 7178 633 7216 667
rect 7250 633 7288 667
rect 7322 633 7360 667
rect 7394 633 7432 667
rect 7466 633 7504 667
rect 7538 633 7576 667
rect 7610 633 7648 667
rect 7682 633 7720 667
rect 7754 633 7792 667
rect 7826 633 7864 667
rect 7898 633 7936 667
rect 7970 633 8008 667
rect 8042 633 8080 667
rect 8114 633 8152 667
rect 8186 633 8224 667
rect 8258 633 8296 667
rect 8330 633 8368 667
rect 8402 633 8440 667
rect 8474 633 8512 667
rect 8546 633 8584 667
rect 8618 633 8656 667
rect 8690 633 8728 667
rect 8762 633 8800 667
rect 8834 633 8872 667
rect 8906 633 8944 667
rect 8978 633 9016 667
rect 9050 633 9088 667
rect 9122 633 9160 667
rect 9194 633 9232 667
rect 9266 633 9304 667
rect 9338 633 9376 667
rect 9410 633 9448 667
rect 9482 633 9520 667
rect 9554 633 9592 667
rect 9626 633 9664 667
rect 9698 633 9736 667
rect 9770 633 9808 667
rect 9842 633 9880 667
rect 9914 633 9952 667
rect 9986 633 10024 667
rect 10058 633 10096 667
rect 10130 633 10168 667
rect 10202 633 10240 667
rect 10274 633 10312 667
rect 10346 633 10384 667
rect 10418 633 10456 667
rect 10490 633 10528 667
rect 10562 633 10600 667
rect 10634 633 10672 667
rect 10706 633 10744 667
rect 10778 633 10816 667
rect 10850 633 10862 667
rect 5471 627 10862 633
rect 4364 542 4764 548
rect 4364 508 4376 542
rect 4410 508 4448 542
rect 4482 508 4764 542
rect 4364 496 4764 508
rect 4765 497 4766 547
rect 4802 497 4803 547
rect 4804 542 5358 548
rect 4804 508 5238 542
rect 5272 508 5310 542
rect 5344 508 5358 542
rect 4804 496 5358 508
rect 4364 416 4763 425
rect 4364 382 4376 416
rect 4410 382 4448 416
rect 4482 382 4763 416
rect 4364 373 4763 382
rect 4764 374 4765 424
rect 4801 374 4802 424
rect 4803 416 5356 425
rect 4803 382 5238 416
rect 5272 382 5310 416
rect 5344 382 5356 416
rect 4803 373 5356 382
rect 4364 290 4763 299
rect 4765 298 4801 299
rect 4364 256 4376 290
rect 4410 256 4448 290
rect 4482 256 4763 290
rect 4364 247 4763 256
rect 4764 248 4802 298
rect 4803 290 5356 299
rect 4803 256 5238 290
rect 5272 256 5310 290
rect 5344 256 5356 290
rect 4765 247 4801 248
rect 4803 247 5356 256
rect 3516 163 5344 169
tri 3388 129 3402 143 sw
rect 3516 129 3528 163
rect 3562 129 3600 163
rect 3634 129 4235 163
rect 4269 129 4307 163
rect 4341 129 5226 163
rect 5260 129 5298 163
rect 5332 129 5344 163
rect 3292 46 3402 129
tri 3402 46 3485 129 sw
rect 3516 123 5344 129
rect 3292 40 5468 46
rect 3292 6 3422 40
rect 3456 6 3496 40
rect 3530 6 3570 40
rect 3604 6 3644 40
rect 3678 6 3718 40
rect 3752 6 3792 40
rect 3826 6 3866 40
rect 3900 6 3940 40
rect 3974 6 4014 40
rect 4048 6 4088 40
rect 4122 6 4162 40
rect 4196 6 4236 40
rect 4270 6 4310 40
rect 4344 6 4384 40
rect 4418 6 4458 40
rect 4492 6 4532 40
rect 4566 6 4606 40
rect 4640 6 4680 40
rect 4714 6 4754 40
rect 4788 6 4828 40
rect 4862 6 4902 40
rect 4936 6 4976 40
rect 5010 6 5050 40
rect 5084 6 5124 40
rect 5158 6 5198 40
rect 5232 6 5272 40
rect 5306 6 5347 40
rect 5381 6 5422 40
rect 5456 6 5468 40
rect 3292 0 5468 6
<< rmetal1 >>
rect 4294 1817 4296 1818
rect 4294 1767 4295 1817
rect 4294 1766 4296 1767
rect 4332 1817 4334 1818
rect 4333 1767 4334 1817
rect 5302 1817 5304 1818
rect 5340 1817 5342 1818
rect 4332 1766 4334 1767
rect 5302 1767 5303 1817
rect 5341 1767 5342 1817
rect 6204 1817 6206 1818
rect 6242 1817 6244 1818
rect 5302 1766 5304 1767
rect 5340 1766 5342 1767
rect 6204 1767 6205 1817
rect 6243 1767 6244 1817
rect 7463 1817 7465 1818
rect 7501 1817 7503 1818
rect 6204 1766 6206 1767
rect 6242 1766 6244 1767
rect 7463 1767 7464 1817
rect 7502 1767 7503 1817
rect 8422 1817 8424 1818
rect 8460 1817 8462 1818
rect 7463 1766 7465 1767
rect 7501 1766 7503 1767
rect 8422 1767 8423 1817
rect 8461 1767 8462 1817
rect 8422 1766 8424 1767
rect 8460 1766 8462 1767
rect 4926 1691 4928 1692
rect 4964 1691 4966 1692
rect 4926 1641 4927 1691
rect 4965 1641 4966 1691
rect 6185 1691 6187 1692
rect 6223 1691 6225 1692
rect 4926 1640 4928 1641
rect 4964 1640 4966 1641
rect 6185 1641 6186 1691
rect 6224 1641 6225 1691
rect 7474 1691 7476 1692
rect 7512 1691 7514 1692
rect 6185 1640 6187 1641
rect 6223 1640 6225 1641
rect 7474 1641 7475 1691
rect 7513 1641 7514 1691
rect 8419 1691 8421 1692
rect 8457 1691 8459 1692
rect 7474 1640 7476 1641
rect 7512 1640 7514 1641
rect 8419 1641 8420 1691
rect 8458 1641 8459 1691
rect 8419 1640 8421 1641
rect 8457 1640 8459 1641
rect 4926 1566 4928 1567
rect 4964 1566 4966 1567
rect 4926 1516 4927 1566
rect 4965 1516 4966 1566
rect 6185 1566 6187 1567
rect 6223 1566 6225 1567
rect 4926 1515 4928 1516
rect 4964 1515 4966 1516
rect 6185 1516 6186 1566
rect 6224 1516 6225 1566
rect 7474 1566 7476 1567
rect 6185 1515 6187 1516
rect 6223 1515 6225 1516
rect 7474 1516 7475 1566
rect 7474 1515 7476 1516
rect 7512 1566 7514 1567
rect 7513 1516 7514 1566
rect 8419 1566 8421 1567
rect 7512 1515 7514 1516
rect 8419 1516 8420 1566
rect 8419 1515 8421 1516
rect 8457 1566 8459 1567
rect 8458 1516 8459 1566
rect 8457 1515 8459 1516
rect 6023 1431 6025 1432
rect 6023 1381 6024 1431
rect 6023 1380 6025 1381
rect 6061 1431 6063 1432
rect 6062 1381 6063 1431
rect 6061 1380 6063 1381
rect 4759 1181 4761 1182
rect 4759 1131 4760 1181
rect 4759 1130 4761 1131
rect 4797 1181 4799 1182
rect 4798 1131 4799 1181
rect 4797 1130 4799 1131
rect 4759 1053 4761 1054
rect 4759 1003 4760 1053
rect 4759 1002 4761 1003
rect 4797 1053 4799 1054
rect 4798 1003 4799 1053
rect 4797 1002 4799 1003
rect 4763 927 4765 928
rect 4763 877 4764 927
rect 4763 876 4765 877
rect 4801 927 4803 928
rect 4802 877 4803 927
rect 4801 876 4803 877
rect 4763 801 4765 802
rect 4763 751 4764 801
rect 4763 750 4765 751
rect 4801 801 4803 802
rect 4802 751 4803 801
rect 4801 750 4803 751
rect 6024 1307 6026 1308
rect 6024 1257 6025 1307
rect 6024 1256 6026 1257
rect 6062 1307 6064 1308
rect 6063 1257 6064 1307
rect 6062 1256 6064 1257
rect 6024 1177 6026 1178
rect 6024 1127 6025 1177
rect 6024 1126 6026 1127
rect 6062 1177 6064 1178
rect 6063 1127 6064 1177
rect 6062 1126 6064 1127
rect 6024 1054 6026 1055
rect 6024 1004 6025 1054
rect 6024 1003 6026 1004
rect 6062 1054 6064 1055
rect 6063 1004 6064 1054
rect 6062 1003 6064 1004
rect 6024 928 6026 929
rect 6024 878 6025 928
rect 6024 877 6026 878
rect 6062 928 6064 929
rect 6063 878 6064 928
rect 6062 877 6064 878
rect 4764 677 4766 678
rect 4764 627 4765 677
rect 4764 626 4766 627
rect 4802 677 4804 678
rect 4803 627 4804 677
rect 4802 626 4804 627
rect 4764 547 4766 548
rect 4764 497 4765 547
rect 4764 496 4766 497
rect 4802 547 4804 548
rect 4803 497 4804 547
rect 4802 496 4804 497
rect 4763 424 4765 425
rect 4763 374 4764 424
rect 4763 373 4765 374
rect 4801 424 4803 425
rect 4802 374 4803 424
rect 4801 373 4803 374
rect 4763 298 4765 299
rect 4801 298 4803 299
rect 4763 248 4764 298
rect 4802 248 4803 298
rect 4763 247 4765 248
rect 4801 247 4803 248
<< via1 >>
rect 3551 2055 3603 2105
rect 3551 2053 3570 2055
rect 3570 2053 3603 2055
rect 3615 2093 3667 2105
rect 3679 2093 3731 2105
rect 4191 2093 4243 2105
rect 4256 2093 4308 2105
rect 4321 2093 4373 2105
rect 4386 2093 4438 2105
rect 3615 2059 3648 2093
rect 3648 2059 3667 2093
rect 3679 2059 3682 2093
rect 3682 2059 3721 2093
rect 3721 2059 3731 2093
rect 4191 2059 4193 2093
rect 4193 2059 4232 2093
rect 4232 2059 4243 2093
rect 4256 2059 4266 2093
rect 4266 2059 4305 2093
rect 4305 2059 4308 2093
rect 4321 2059 4339 2093
rect 4339 2059 4373 2093
rect 4386 2059 4412 2093
rect 4412 2059 4438 2093
rect 3615 2053 3667 2059
rect 3679 2053 3731 2059
rect 4191 2053 4243 2059
rect 4256 2053 4308 2059
rect 4321 2053 4373 2059
rect 4386 2053 4438 2059
rect 4450 2093 4502 2105
rect 4450 2059 4451 2093
rect 4451 2059 4485 2093
rect 4485 2059 4502 2093
rect 4450 2053 4502 2059
rect 4514 2093 4566 2105
rect 4514 2059 4524 2093
rect 4524 2059 4558 2093
rect 4558 2059 4566 2093
rect 4514 2053 4566 2059
rect 4578 2093 4630 2105
rect 4578 2059 4597 2093
rect 4597 2059 4630 2093
rect 4578 2053 4630 2059
rect 10124 1506 10176 1558
rect 10196 1506 10248 1558
rect 10268 1506 10320 1558
rect 10340 1506 10392 1558
rect 10412 1506 10464 1558
<< metal2 >>
rect 3545 2053 3551 2105
rect 3603 2053 3615 2105
rect 3667 2053 3679 2105
rect 3731 2053 3737 2105
rect 4185 2053 4191 2105
rect 4243 2053 4256 2105
rect 4308 2053 4321 2105
rect 4373 2053 4386 2105
rect 4438 2053 4450 2105
rect 4502 2053 4514 2105
rect 4566 2053 4578 2105
rect 4630 2053 4636 2105
rect 10118 1506 10124 1558
rect 10176 1506 10196 1558
rect 10248 1506 10268 1558
rect 10320 1506 10340 1558
rect 10392 1506 10412 1558
rect 10464 1506 10470 1558
use nDFres_CDNS_524688791851256  nDFres_CDNS_524688791851256_0
timestamp 1704896540
transform -1 0 8896 0 -1 1573
box -68 -26 1225 92
use nDFres_CDNS_524688791851256  nDFres_CDNS_524688791851256_1
timestamp 1704896540
transform -1 0 7637 0 -1 1573
box -68 -26 1225 92
use nDFres_CDNS_524688791851256  nDFres_CDNS_524688791851256_2
timestamp 1704896540
transform -1 0 6378 0 -1 1573
box -68 -26 1225 92
use nDFres_CDNS_524688791851256  nDFres_CDNS_524688791851256_3
timestamp 1704896540
transform -1 0 8896 0 -1 1825
box -68 -26 1225 92
use nDFres_CDNS_524688791851256  nDFres_CDNS_524688791851256_4
timestamp 1704896540
transform -1 0 7637 0 -1 1825
box -68 -26 1225 92
use nDFres_CDNS_524688791851256  nDFres_CDNS_524688791851256_5
timestamp 1704896540
transform 1 0 5221 0 -1 1699
box -68 -26 1225 92
use nDFres_CDNS_524688791851256  nDFres_CDNS_524688791851256_6
timestamp 1704896540
transform 1 0 6480 0 -1 1699
box -68 -26 1225 92
use nDFres_CDNS_524688791851256  nDFres_CDNS_524688791851256_7
timestamp 1704896540
transform 1 0 7739 0 -1 1699
box -68 -26 1225 92
use nDFres_CDNS_524688791851257  nDFres_CDNS_524688791851257_0
timestamp 1704896540
transform -1 0 8896 0 1 1885
box -68 -26 5131 92
use nDFres_CDNS_524688791851257  nDFres_CDNS_524688791851257_1
timestamp 1704896540
transform -1 0 10652 0 1 744
box -68 -26 5131 92
use nDFres_CDNS_524688791851257  nDFres_CDNS_524688791851257_2
timestamp 1704896540
transform -1 0 10652 0 1 870
box -68 -26 5131 92
use nDFres_CDNS_524688791851257  nDFres_CDNS_524688791851257_3
timestamp 1704896540
transform -1 0 5240 0 -1 180
box -68 -26 5131 92
use nDFres_CDNS_524688791851257  nDFres_CDNS_524688791851257_4
timestamp 1704896540
transform -1 0 5240 0 -1 1188
box -68 -26 5131 92
use nDFres_CDNS_524688791851257  nDFres_CDNS_524688791851257_5
timestamp 1704896540
transform -1 0 10652 0 -1 1188
box -68 -26 5131 92
use nDFres_CDNS_524688791851257  nDFres_CDNS_524688791851257_6
timestamp 1704896540
transform -1 0 5240 0 -1 936
box -68 -26 5131 92
use nDFres_CDNS_524688791851257  nDFres_CDNS_524688791851257_7
timestamp 1704896540
transform -1 0 5240 0 -1 558
box -68 -26 5131 92
use nDFres_CDNS_524688791851257  nDFres_CDNS_524688791851257_8
timestamp 1704896540
transform -1 0 5240 0 -1 1314
box -68 -26 5131 92
use nDFres_CDNS_524688791851257  nDFres_CDNS_524688791851257_9
timestamp 1704896540
transform -1 0 5240 0 -1 306
box -68 -26 5131 92
use nDFres_CDNS_524688791851257  nDFres_CDNS_524688791851257_10
timestamp 1704896540
transform 1 0 5589 0 -1 1062
box -68 -26 5131 92
use nDFres_CDNS_524688791851257  nDFres_CDNS_524688791851257_11
timestamp 1704896540
transform 1 0 177 0 -1 1062
box -68 -26 5131 92
use nDFres_CDNS_524688791851257  nDFres_CDNS_524688791851257_12
timestamp 1704896540
transform 1 0 177 0 -1 810
box -68 -26 5131 92
use nDFres_CDNS_524688791851257  nDFres_CDNS_524688791851257_13
timestamp 1704896540
transform 1 0 177 0 -1 684
box -68 -26 5131 92
use nDFres_CDNS_524688791851257  nDFres_CDNS_524688791851257_14
timestamp 1704896540
transform 1 0 5589 0 -1 1440
box -68 -26 5131 92
use nDFres_CDNS_524688791851257  nDFres_CDNS_524688791851257_15
timestamp 1704896540
transform 1 0 5589 0 -1 1314
box -68 -26 5131 92
use nDFres_CDNS_524688791851257  nDFres_CDNS_524688791851257_16
timestamp 1704896540
transform 1 0 177 0 -1 432
box -68 -26 5131 92
use nDFres_CDNS_524688791851258  nDFres_CDNS_524688791851258_0
timestamp 1704896540
transform -1 0 5119 0 -1 1573
box -68 -26 1354 92
use nDFres_CDNS_524688791851258  nDFres_CDNS_524688791851258_1
timestamp 1704896540
transform 1 0 3833 0 -1 1699
box -68 -26 1354 92
use nDFres_CDNS_524688791851259  nDFres_CDNS_524688791851259_0
timestamp 1704896540
transform -1 0 6378 0 -1 1825
box -68 -26 868 92
use nDFres_CDNS_524688791851259  nDFres_CDNS_524688791851259_1
timestamp 1704896540
transform -1 0 5476 0 -1 1825
box -68 -26 868 92
use nDFres_CDNS_524688791851260  nDFres_CDNS_524688791851260_0
timestamp 1704896540
transform -1 0 4574 0 -1 1825
box -68 -26 809 92
use pfet_CDNS_524688791851261  pfet_CDNS_524688791851261_0
timestamp 1704896540
transform 0 -1 8800 -1 0 2602
box -89 -36 245 1036
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851254  sky130_fd_io__sio_tk_em1o_CDNS_524688791851254_0
timestamp 1704896540
transform -1 0 6116 0 1 877
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851254  sky130_fd_io__sio_tk_em1o_CDNS_524688791851254_1
timestamp 1704896540
transform -1 0 8511 0 -1 1567
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851254  sky130_fd_io__sio_tk_em1o_CDNS_524688791851254_2
timestamp 1704896540
transform -1 0 4851 0 -1 1054
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851254  sky130_fd_io__sio_tk_em1o_CDNS_524688791851254_3
timestamp 1704896540
transform -1 0 6116 0 -1 1178
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851254  sky130_fd_io__sio_tk_em1o_CDNS_524688791851254_4
timestamp 1704896540
transform -1 0 7566 0 -1 1567
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851254  sky130_fd_io__sio_tk_em1o_CDNS_524688791851254_5
timestamp 1704896540
transform -1 0 4855 0 -1 928
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851254  sky130_fd_io__sio_tk_em1o_CDNS_524688791851254_6
timestamp 1704896540
transform -1 0 4856 0 -1 548
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851254  sky130_fd_io__sio_tk_em1o_CDNS_524688791851254_7
timestamp 1704896540
transform -1 0 4386 0 -1 1818
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851254  sky130_fd_io__sio_tk_em1o_CDNS_524688791851254_8
timestamp 1704896540
transform 1 0 5972 0 -1 1055
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851254  sky130_fd_io__sio_tk_em1o_CDNS_524688791851254_9
timestamp 1704896540
transform 1 0 4707 0 -1 1182
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851254  sky130_fd_io__sio_tk_em1o_CDNS_524688791851254_10
timestamp 1704896540
transform 1 0 4712 0 -1 678
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851254  sky130_fd_io__sio_tk_em1o_CDNS_524688791851254_11
timestamp 1704896540
transform 1 0 4711 0 -1 802
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851254  sky130_fd_io__sio_tk_em1o_CDNS_524688791851254_12
timestamp 1704896540
transform 1 0 5971 0 -1 1432
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851254  sky130_fd_io__sio_tk_em1o_CDNS_524688791851254_13
timestamp 1704896540
transform 1 0 5972 0 -1 1308
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851254  sky130_fd_io__sio_tk_em1o_CDNS_524688791851254_14
timestamp 1704896540
transform 1 0 4711 0 -1 425
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851255  sky130_fd_io__sio_tk_em1s_CDNS_524688791851255_0
timestamp 1704896540
transform -1 0 6277 0 -1 1567
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851255  sky130_fd_io__sio_tk_em1s_CDNS_524688791851255_1
timestamp 1704896540
transform -1 0 8514 0 -1 1818
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851255  sky130_fd_io__sio_tk_em1s_CDNS_524688791851255_2
timestamp 1704896540
transform -1 0 5018 0 -1 1567
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851255  sky130_fd_io__sio_tk_em1s_CDNS_524688791851255_3
timestamp 1704896540
transform -1 0 7555 0 -1 1818
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851255  sky130_fd_io__sio_tk_em1s_CDNS_524688791851255_4
timestamp 1704896540
transform -1 0 5394 0 -1 1818
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851255  sky130_fd_io__sio_tk_em1s_CDNS_524688791851255_5
timestamp 1704896540
transform -1 0 6296 0 -1 1818
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851255  sky130_fd_io__sio_tk_em1s_CDNS_524688791851255_6
timestamp 1704896540
transform -1 0 4855 0 -1 299
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851255  sky130_fd_io__sio_tk_em1s_CDNS_524688791851255_7
timestamp 1704896540
transform 1 0 6133 0 -1 1692
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851255  sky130_fd_io__sio_tk_em1s_CDNS_524688791851255_8
timestamp 1704896540
transform 1 0 7422 0 -1 1692
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851255  sky130_fd_io__sio_tk_em1s_CDNS_524688791851255_9
timestamp 1704896540
transform 1 0 8367 0 -1 1692
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851255  sky130_fd_io__sio_tk_em1s_CDNS_524688791851255_10
timestamp 1704896540
transform 1 0 4874 0 -1 1692
box 0 0 1 1
<< labels >>
flabel comment s 9129 2090 9129 2090 3 FreeSans 400 270 0 0 vcc_io
flabel comment s 4782 397 4782 397 0 FreeSans 400 90 0 0 o21
flabel metal1 s 6713 2053 6784 2099 3 FreeSans 520 0 0 0 vgnd
port 1 nsew
flabel metal1 s 7842 2293 8046 2386 3 FreeSans 520 0 0 0 vpwr
port 2 nsew
flabel metal1 s 5190 248 5356 298 3 FreeSans 520 0 0 0 ngate
port 3 nsew
<< properties >>
string GDS_END 86588158
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86503836
string path 104.625 51.975 115.900 51.975 
<< end >>
