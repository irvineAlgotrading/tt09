magic
tech sky130A
timestamp 1704896540
<< metal1 >>
rect 0 0 3 218
rect 285 0 288 218
<< via1 >>
rect 3 0 285 218
<< metal2 >>
rect 0 0 3 218
rect 285 0 288 218
<< properties >>
string GDS_END 93931994
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 93927830
<< end >>
