magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect 0 1165 2135 1333
<< pwell >>
rect 60 14 2069 100
<< mvpsubdiff >>
rect 86 40 110 74
rect 144 40 180 74
rect 214 40 250 74
rect 284 40 320 74
rect 354 40 390 74
rect 424 40 460 74
rect 494 40 530 74
rect 564 40 600 74
rect 634 40 670 74
rect 704 40 740 74
rect 774 40 810 74
rect 844 40 880 74
rect 914 40 950 74
rect 984 40 1019 74
rect 1053 40 1088 74
rect 1122 40 1157 74
rect 1191 40 1226 74
rect 1260 40 1295 74
rect 1329 40 1364 74
rect 1398 40 1433 74
rect 1467 40 1502 74
rect 1536 40 1571 74
rect 1605 40 1640 74
rect 1674 40 1709 74
rect 1743 40 1778 74
rect 1812 40 1847 74
rect 1881 40 1916 74
rect 1950 40 1985 74
rect 2019 40 2043 74
<< mvnsubdiff >>
rect 67 1232 101 1266
rect 135 1232 169 1266
rect 203 1232 237 1266
rect 271 1232 305 1266
rect 339 1232 373 1266
rect 407 1232 441 1266
rect 475 1232 509 1266
rect 543 1232 577 1266
rect 611 1232 645 1266
rect 679 1232 713 1266
rect 747 1232 781 1266
rect 815 1232 849 1266
rect 883 1232 917 1266
rect 951 1232 985 1266
rect 1019 1232 1053 1266
rect 1087 1232 1121 1266
rect 1155 1232 1189 1266
rect 1223 1232 1257 1266
rect 1291 1232 1325 1266
rect 1359 1232 1393 1266
rect 1427 1232 1461 1266
rect 1495 1232 1529 1266
rect 1563 1232 1597 1266
rect 1631 1232 1665 1266
rect 1699 1232 1733 1266
rect 1767 1232 1801 1266
rect 1835 1232 1869 1266
rect 1903 1232 1937 1266
rect 1971 1232 2068 1266
<< mvpsubdiffcont >>
rect 110 40 144 74
rect 180 40 214 74
rect 250 40 284 74
rect 320 40 354 74
rect 390 40 424 74
rect 460 40 494 74
rect 530 40 564 74
rect 600 40 634 74
rect 670 40 704 74
rect 740 40 774 74
rect 810 40 844 74
rect 880 40 914 74
rect 950 40 984 74
rect 1019 40 1053 74
rect 1088 40 1122 74
rect 1157 40 1191 74
rect 1226 40 1260 74
rect 1295 40 1329 74
rect 1364 40 1398 74
rect 1433 40 1467 74
rect 1502 40 1536 74
rect 1571 40 1605 74
rect 1640 40 1674 74
rect 1709 40 1743 74
rect 1778 40 1812 74
rect 1847 40 1881 74
rect 1916 40 1950 74
rect 1985 40 2019 74
<< mvnsubdiffcont >>
rect 101 1232 135 1266
rect 169 1232 203 1266
rect 237 1232 271 1266
rect 305 1232 339 1266
rect 373 1232 407 1266
rect 441 1232 475 1266
rect 509 1232 543 1266
rect 577 1232 611 1266
rect 645 1232 679 1266
rect 713 1232 747 1266
rect 781 1232 815 1266
rect 849 1232 883 1266
rect 917 1232 951 1266
rect 985 1232 1019 1266
rect 1053 1232 1087 1266
rect 1121 1232 1155 1266
rect 1189 1232 1223 1266
rect 1257 1232 1291 1266
rect 1325 1232 1359 1266
rect 1393 1232 1427 1266
rect 1461 1232 1495 1266
rect 1529 1232 1563 1266
rect 1597 1232 1631 1266
rect 1665 1232 1699 1266
rect 1733 1232 1767 1266
rect 1801 1232 1835 1266
rect 1869 1232 1903 1266
rect 1937 1232 1971 1266
<< poly >>
rect 119 504 239 521
rect 119 470 158 504
rect 192 470 239 504
rect 119 436 239 470
rect 119 402 158 436
rect 192 402 239 436
rect 119 385 239 402
rect 295 504 415 521
rect 295 470 334 504
rect 368 470 415 504
rect 295 436 415 470
rect 295 402 334 436
rect 368 402 415 436
rect 295 385 415 402
rect 471 504 591 521
rect 471 470 510 504
rect 544 470 591 504
rect 471 436 591 470
rect 471 402 510 436
rect 544 402 591 436
rect 471 385 591 402
rect 647 504 767 521
rect 647 470 686 504
rect 720 470 767 504
rect 647 436 767 470
rect 647 402 686 436
rect 720 402 767 436
rect 647 385 767 402
rect 823 504 943 521
rect 823 470 862 504
rect 896 470 943 504
rect 823 436 943 470
rect 823 402 862 436
rect 896 402 943 436
rect 823 385 943 402
rect 999 504 1119 521
rect 999 470 1038 504
rect 1072 470 1119 504
rect 999 436 1119 470
rect 999 402 1038 436
rect 1072 402 1119 436
rect 999 385 1119 402
rect 1285 504 1405 521
rect 1285 470 1324 504
rect 1358 470 1405 504
rect 1285 436 1405 470
rect 1285 402 1324 436
rect 1358 402 1405 436
rect 1285 385 1405 402
<< polycont >>
rect 158 470 192 504
rect 158 402 192 436
rect 334 470 368 504
rect 334 402 368 436
rect 510 470 544 504
rect 510 402 544 436
rect 686 470 720 504
rect 686 402 720 436
rect 862 470 896 504
rect 862 402 896 436
rect 1038 470 1072 504
rect 1038 402 1072 436
rect 1324 470 1358 504
rect 1324 402 1358 436
<< locali >>
rect 67 1232 79 1266
rect 135 1232 154 1266
rect 203 1232 229 1266
rect 271 1232 304 1266
rect 339 1232 373 1266
rect 413 1232 441 1266
rect 488 1232 509 1266
rect 563 1232 577 1266
rect 638 1232 645 1266
rect 747 1232 754 1266
rect 815 1232 829 1266
rect 883 1232 904 1266
rect 951 1232 979 1266
rect 1019 1232 1053 1266
rect 1088 1232 1121 1266
rect 1163 1232 1189 1266
rect 1238 1232 1257 1266
rect 1313 1232 1325 1266
rect 1388 1232 1393 1266
rect 1427 1232 1429 1266
rect 1495 1232 1504 1266
rect 1563 1232 1578 1266
rect 1631 1232 1652 1266
rect 1699 1232 1726 1266
rect 1767 1232 1800 1266
rect 1835 1232 1869 1266
rect 1908 1232 1937 1266
rect 1982 1232 2022 1266
rect 2056 1232 2068 1266
rect 250 1072 284 1123
rect 250 987 284 1038
rect 74 896 108 944
rect 74 814 108 862
rect 74 732 108 780
rect 602 1072 636 1123
rect 602 987 636 1038
rect 250 902 284 953
rect 250 817 284 868
rect 250 732 284 783
rect 426 896 460 944
rect 426 814 460 862
rect 426 732 460 780
rect 954 1072 988 1123
rect 954 987 988 1038
rect 602 902 636 953
rect 602 817 636 868
rect 602 732 636 783
rect 778 896 812 944
rect 778 814 812 862
rect 778 732 812 780
rect 1416 1072 1450 1123
rect 1416 987 1450 1038
rect 954 902 988 953
rect 954 817 988 868
rect 954 732 988 783
rect 1130 896 1164 944
rect 1130 814 1164 862
rect 1130 732 1164 780
rect 74 649 108 698
rect 426 649 460 698
rect 778 649 812 698
rect 1130 649 1164 698
rect 1240 896 1274 944
rect 1240 814 1274 862
rect 1240 732 1274 780
rect 1416 902 1450 953
rect 1416 817 1450 868
rect 1416 732 1450 783
rect 1240 649 1274 698
rect 158 507 192 520
rect 158 436 192 470
rect 158 386 192 401
rect 334 507 368 520
rect 334 436 368 470
rect 334 386 368 401
rect 510 507 544 520
rect 510 436 544 470
rect 510 386 544 401
rect 686 507 720 520
rect 686 436 720 470
rect 686 386 720 401
rect 862 507 896 520
rect 862 436 896 470
rect 862 386 896 401
rect 1038 507 1072 520
rect 1038 436 1072 470
rect 1038 386 1072 401
rect 1324 507 1358 520
rect 1324 436 1358 470
rect 1707 437 1741 475
rect 1910 449 1944 487
rect 1324 386 1358 401
rect 74 274 108 312
rect 426 274 460 312
rect 778 274 812 312
rect 250 188 284 226
rect 1130 274 1164 312
rect 602 188 636 226
rect 1240 274 1274 312
rect 954 188 988 226
rect 1416 188 1450 226
rect 144 40 160 74
rect 214 40 234 74
rect 284 40 308 74
rect 354 40 382 74
rect 424 40 456 74
rect 494 40 530 74
rect 564 40 600 74
rect 638 40 670 74
rect 712 40 740 74
rect 786 40 810 74
rect 860 40 880 74
rect 934 40 950 74
rect 1008 40 1019 74
rect 1082 40 1088 74
rect 1155 40 1157 74
rect 1191 40 1194 74
rect 1260 40 1267 74
rect 1329 40 1340 74
rect 1398 40 1413 74
rect 1467 40 1486 74
rect 1536 40 1559 74
rect 1605 40 1632 74
rect 1674 40 1705 74
rect 1743 40 1778 74
rect 1812 40 1847 74
rect 1885 40 1916 74
rect 1958 40 1985 74
rect 2031 40 2043 74
<< viali >>
rect 79 1232 101 1266
rect 101 1232 113 1266
rect 154 1232 169 1266
rect 169 1232 188 1266
rect 229 1232 237 1266
rect 237 1232 263 1266
rect 304 1232 305 1266
rect 305 1232 338 1266
rect 379 1232 407 1266
rect 407 1232 413 1266
rect 454 1232 475 1266
rect 475 1232 488 1266
rect 529 1232 543 1266
rect 543 1232 563 1266
rect 604 1232 611 1266
rect 611 1232 638 1266
rect 679 1232 713 1266
rect 754 1232 781 1266
rect 781 1232 788 1266
rect 829 1232 849 1266
rect 849 1232 863 1266
rect 904 1232 917 1266
rect 917 1232 938 1266
rect 979 1232 985 1266
rect 985 1232 1013 1266
rect 1054 1232 1087 1266
rect 1087 1232 1088 1266
rect 1129 1232 1155 1266
rect 1155 1232 1163 1266
rect 1204 1232 1223 1266
rect 1223 1232 1238 1266
rect 1279 1232 1291 1266
rect 1291 1232 1313 1266
rect 1354 1232 1359 1266
rect 1359 1232 1388 1266
rect 1429 1232 1461 1266
rect 1461 1232 1463 1266
rect 1504 1232 1529 1266
rect 1529 1232 1538 1266
rect 1578 1232 1597 1266
rect 1597 1232 1612 1266
rect 1652 1232 1665 1266
rect 1665 1232 1686 1266
rect 1726 1232 1733 1266
rect 1733 1232 1760 1266
rect 1800 1232 1801 1266
rect 1801 1232 1834 1266
rect 1874 1232 1903 1266
rect 1903 1232 1908 1266
rect 1948 1232 1971 1266
rect 1971 1232 1982 1266
rect 2022 1232 2056 1266
rect 250 1123 284 1157
rect 250 1038 284 1072
rect 74 944 108 978
rect 74 862 108 896
rect 74 780 108 814
rect 74 698 108 732
rect 250 953 284 987
rect 602 1123 636 1157
rect 602 1038 636 1072
rect 250 868 284 902
rect 250 783 284 817
rect 250 698 284 732
rect 426 944 460 978
rect 426 862 460 896
rect 426 780 460 814
rect 426 698 460 732
rect 602 953 636 987
rect 954 1123 988 1157
rect 954 1038 988 1072
rect 602 868 636 902
rect 602 783 636 817
rect 602 698 636 732
rect 778 944 812 978
rect 778 862 812 896
rect 778 780 812 814
rect 778 698 812 732
rect 954 953 988 987
rect 1416 1123 1450 1157
rect 1416 1038 1450 1072
rect 954 868 988 902
rect 954 783 988 817
rect 954 698 988 732
rect 1130 944 1164 978
rect 1130 862 1164 896
rect 1130 780 1164 814
rect 1130 698 1164 732
rect 74 615 108 649
rect 426 615 460 649
rect 778 615 812 649
rect 1130 615 1164 649
rect 1240 944 1274 978
rect 1240 862 1274 896
rect 1240 780 1274 814
rect 1240 698 1274 732
rect 1416 953 1450 987
rect 1416 868 1450 902
rect 1416 783 1450 817
rect 1416 698 1450 732
rect 1240 615 1274 649
rect 158 504 192 507
rect 158 473 192 504
rect 158 402 192 435
rect 158 401 192 402
rect 334 504 368 507
rect 334 473 368 504
rect 334 402 368 435
rect 334 401 368 402
rect 510 504 544 507
rect 510 473 544 504
rect 510 402 544 435
rect 510 401 544 402
rect 686 504 720 507
rect 686 473 720 504
rect 686 402 720 435
rect 686 401 720 402
rect 862 504 896 507
rect 862 473 896 504
rect 862 402 896 435
rect 862 401 896 402
rect 1038 504 1072 507
rect 1038 473 1072 504
rect 1038 402 1072 435
rect 1038 401 1072 402
rect 1324 504 1358 507
rect 1324 473 1358 504
rect 1324 402 1358 435
rect 1707 475 1741 509
rect 1707 403 1741 437
rect 1910 487 1944 521
rect 1910 415 1944 449
rect 1324 401 1358 402
rect 74 312 108 346
rect 74 240 108 274
rect 426 312 460 346
rect 250 226 284 260
rect 426 240 460 274
rect 778 312 812 346
rect 250 154 284 188
rect 602 226 636 260
rect 778 240 812 274
rect 1130 312 1164 346
rect 602 154 636 188
rect 954 226 988 260
rect 1130 240 1164 274
rect 1240 312 1274 346
rect 1240 240 1274 274
rect 954 154 988 188
rect 1416 226 1450 260
rect 1416 154 1450 188
rect 86 40 110 74
rect 110 40 120 74
rect 160 40 180 74
rect 180 40 194 74
rect 234 40 250 74
rect 250 40 268 74
rect 308 40 320 74
rect 320 40 342 74
rect 382 40 390 74
rect 390 40 416 74
rect 456 40 460 74
rect 460 40 490 74
rect 530 40 564 74
rect 604 40 634 74
rect 634 40 638 74
rect 678 40 704 74
rect 704 40 712 74
rect 752 40 774 74
rect 774 40 786 74
rect 826 40 844 74
rect 844 40 860 74
rect 900 40 914 74
rect 914 40 934 74
rect 974 40 984 74
rect 984 40 1008 74
rect 1048 40 1053 74
rect 1053 40 1082 74
rect 1121 40 1122 74
rect 1122 40 1155 74
rect 1194 40 1226 74
rect 1226 40 1228 74
rect 1267 40 1295 74
rect 1295 40 1301 74
rect 1340 40 1364 74
rect 1364 40 1374 74
rect 1413 40 1433 74
rect 1433 40 1447 74
rect 1486 40 1502 74
rect 1502 40 1520 74
rect 1559 40 1571 74
rect 1571 40 1593 74
rect 1632 40 1640 74
rect 1640 40 1666 74
rect 1705 40 1709 74
rect 1709 40 1739 74
rect 1778 40 1812 74
rect 1851 40 1881 74
rect 1881 40 1885 74
rect 1924 40 1950 74
rect 1950 40 1958 74
rect 1997 40 2019 74
rect 2019 40 2031 74
<< metal1 >>
rect 67 1266 2069 1333
rect 67 1232 79 1266
rect 113 1232 154 1266
rect 188 1232 229 1266
rect 263 1232 304 1266
rect 338 1232 379 1266
rect 413 1232 454 1266
rect 488 1232 529 1266
rect 563 1232 604 1266
rect 638 1232 679 1266
rect 713 1232 754 1266
rect 788 1232 829 1266
rect 863 1232 904 1266
rect 938 1232 979 1266
rect 1013 1232 1054 1266
rect 1088 1232 1129 1266
rect 1163 1232 1204 1266
rect 1238 1232 1279 1266
rect 1313 1232 1354 1266
rect 1388 1232 1429 1266
rect 1463 1232 1504 1266
rect 1538 1232 1578 1266
rect 1612 1232 1652 1266
rect 1686 1232 1726 1266
rect 1760 1232 1800 1266
rect 1834 1232 1874 1266
rect 1908 1232 1948 1266
rect 1982 1232 2022 1266
rect 2056 1232 2069 1266
rect 67 1157 2069 1232
rect 67 1123 250 1157
rect 284 1123 602 1157
rect 636 1123 954 1157
rect 988 1123 1416 1157
rect 1450 1123 2069 1157
rect 67 1072 2069 1123
rect 67 1038 250 1072
rect 284 1038 602 1072
rect 636 1038 954 1072
rect 988 1038 1416 1072
rect 1450 1038 2069 1072
rect 67 1033 2069 1038
tri 210 999 244 1033 ne
rect 68 978 114 990
rect 68 944 74 978
rect 108 944 114 978
rect 68 896 114 944
rect 68 862 74 896
rect 108 862 114 896
rect 68 814 114 862
rect 68 780 74 814
rect 108 780 114 814
rect 68 732 114 780
rect 68 698 74 732
rect 108 698 114 732
rect 68 649 114 698
rect 244 987 290 1033
tri 290 999 324 1033 nw
tri 562 999 596 1033 ne
rect 244 953 250 987
rect 284 953 290 987
rect 244 902 290 953
rect 244 868 250 902
rect 284 868 290 902
rect 244 817 290 868
rect 244 783 250 817
rect 284 783 290 817
rect 244 732 290 783
rect 244 698 250 732
rect 284 698 290 732
rect 244 686 290 698
rect 417 978 469 990
rect 417 944 426 978
rect 460 944 469 978
rect 417 896 469 944
rect 417 862 426 896
rect 460 862 469 896
rect 417 819 469 862
rect 417 740 469 767
tri 114 649 148 683 sw
rect 417 661 469 688
rect 596 987 642 1033
tri 642 999 676 1033 nw
tri 914 999 948 1033 ne
rect 596 953 602 987
rect 636 953 642 987
rect 596 902 642 953
rect 596 868 602 902
rect 636 868 642 902
rect 596 817 642 868
rect 596 783 602 817
rect 636 783 642 817
rect 596 732 642 783
rect 596 698 602 732
rect 636 698 642 732
rect 596 686 642 698
rect 769 978 821 990
rect 769 944 778 978
rect 812 944 821 978
rect 769 896 821 944
rect 769 862 778 896
rect 812 862 821 896
rect 769 814 821 862
rect 769 780 778 814
rect 812 780 821 814
rect 769 732 821 780
rect 769 725 778 732
rect 812 725 821 732
rect 68 615 74 649
rect 108 615 374 649
rect 68 603 374 615
rect 417 603 469 609
rect 948 987 994 1033
tri 994 999 1028 1033 nw
tri 1376 999 1410 1033 ne
rect 948 953 954 987
rect 988 953 994 987
rect 948 902 994 953
rect 948 868 954 902
rect 988 868 994 902
rect 948 817 994 868
rect 948 783 954 817
rect 988 783 994 817
rect 948 732 994 783
rect 948 698 954 732
rect 988 698 994 732
rect 948 686 994 698
rect 1124 978 1170 990
rect 1124 944 1130 978
rect 1164 944 1170 978
rect 1124 896 1170 944
rect 1124 862 1130 896
rect 1164 862 1170 896
rect 1124 814 1170 862
rect 1124 780 1130 814
rect 1164 780 1170 814
rect 1124 732 1170 780
rect 1124 698 1130 732
rect 1164 698 1170 732
rect 769 661 821 673
rect 769 603 821 609
rect 1124 649 1170 698
rect 1124 615 1130 649
rect 1164 615 1170 649
rect 68 346 114 603
tri 114 569 148 603 nw
tri 294 569 328 603 ne
rect 328 521 374 603
tri 374 521 406 553 sw
rect 328 519 406 521
tri 406 519 408 521 sw
rect 152 507 198 519
rect 152 473 158 507
rect 192 473 198 507
rect 152 435 198 473
rect 152 401 158 435
rect 192 401 198 435
rect 152 389 198 401
rect 328 507 550 519
rect 328 473 334 507
rect 368 473 510 507
rect 544 473 550 507
rect 328 435 550 473
rect 328 401 334 435
rect 368 401 510 435
rect 544 401 550 435
rect 328 389 550 401
rect 680 507 902 519
rect 680 473 686 507
rect 720 473 862 507
rect 896 473 902 507
rect 680 435 902 473
rect 680 401 686 435
rect 720 401 862 435
rect 896 401 902 435
rect 680 397 902 401
rect 680 389 726 397
tri 726 389 734 397 nw
tri 822 389 830 397 ne
rect 830 389 902 397
rect 1032 507 1078 519
rect 1032 473 1038 507
rect 1072 473 1078 507
rect 1032 435 1078 473
rect 1032 401 1038 435
rect 1072 401 1078 435
rect 1032 389 1078 401
tri 830 363 856 389 ne
rect 68 312 74 346
rect 108 312 114 346
rect 68 274 114 312
rect 68 240 74 274
rect 108 240 114 274
rect 417 352 469 358
rect 417 288 469 300
rect 68 228 114 240
rect 244 260 290 272
tri 238 228 244 234 se
rect 244 228 250 260
tri 236 226 238 228 se
rect 238 226 250 228
rect 284 226 290 260
rect 769 350 821 358
rect 856 350 902 389
tri 902 350 936 384 sw
tri 1090 350 1124 384 se
rect 1124 350 1170 615
rect 856 346 1170 350
rect 856 312 1130 346
rect 1164 312 1170 346
rect 856 304 1170 312
rect 769 286 821 298
tri 1090 274 1120 304 ne
rect 1120 274 1170 304
tri 290 226 298 234 sw
rect 417 228 469 236
rect 596 260 642 272
tri 590 228 596 234 se
rect 596 228 602 260
tri 588 226 590 228 se
rect 590 226 602 228
rect 636 226 642 260
tri 1120 272 1122 274 ne
rect 1122 272 1130 274
rect 948 260 994 272
tri 1122 270 1124 272 ne
tri 642 226 650 234 sw
rect 769 228 821 234
tri 942 228 948 234 se
rect 948 228 954 260
tri 940 226 942 228 se
rect 942 226 954 228
rect 988 226 994 260
rect 1124 240 1130 272
rect 1164 240 1170 274
tri 994 226 1002 234 sw
rect 1124 228 1170 240
rect 1231 984 1283 990
rect 1231 920 1283 932
rect 1231 862 1240 868
rect 1274 862 1283 868
rect 1231 814 1283 862
rect 1231 780 1240 814
rect 1274 780 1283 814
rect 1231 732 1283 780
rect 1231 698 1240 732
rect 1274 698 1283 732
rect 1231 649 1283 698
rect 1410 987 1456 1033
tri 1456 999 1490 1033 nw
tri 1557 999 1591 1033 ne
rect 1410 953 1416 987
rect 1450 953 1456 987
tri 1600 961 1634 995 ne
tri 1680 961 1714 995 nw
tri 1952 961 1986 995 ne
tri 2032 961 2066 995 nw
rect 1410 902 1456 953
rect 1410 868 1416 902
rect 1450 868 1456 902
rect 1410 817 1456 868
tri 1776 865 1810 899 ne
tri 1856 865 1890 899 nw
rect 1410 783 1416 817
rect 1450 783 1456 817
rect 1410 732 1456 783
rect 1410 698 1416 732
rect 1450 698 1456 732
rect 1410 686 1456 698
rect 1231 615 1240 649
rect 1274 615 1283 649
tri 1769 625 1810 666 se
rect 1231 346 1283 615
rect 1318 579 1849 625
rect 1318 507 1370 579
tri 1370 551 1398 579 nw
tri 1776 551 1804 579 ne
rect 1804 551 1810 579
tri 1804 545 1810 551 ne
rect 1901 525 1953 533
rect 1318 473 1324 507
rect 1358 473 1370 507
rect 1318 435 1370 473
rect 1318 401 1324 435
rect 1358 401 1370 435
rect 1318 389 1370 401
rect 1698 513 1750 521
rect 1698 449 1750 461
rect 1901 461 1953 473
rect 1901 403 1953 409
rect 1698 391 1750 397
tri 1856 391 1864 399 sw
rect 1856 389 1864 391
tri 1864 389 1866 391 sw
rect 1856 365 1866 389
tri 1866 365 1890 389 sw
rect 1231 312 1240 346
rect 1274 312 1283 346
rect 1231 274 1283 312
rect 1231 240 1240 274
rect 1274 240 1283 274
rect 1231 228 1283 240
rect 1410 260 1456 272
tri 1404 228 1410 234 se
rect 1410 228 1416 260
tri 1402 226 1404 228 se
rect 1404 226 1416 228
rect 1450 226 1456 260
tri 210 200 236 226 se
rect 236 200 298 226
tri 298 200 324 226 sw
tri 562 200 588 226 se
rect 588 200 650 226
tri 650 200 676 226 sw
tri 914 200 940 226 se
rect 940 200 1002 226
tri 1002 200 1028 226 sw
tri 1376 200 1402 226 se
rect 1402 200 1456 226
tri 1456 200 1490 234 sw
tri 1556 200 1590 234 se
rect 74 188 2069 200
rect 74 154 250 188
rect 284 154 602 188
rect 636 154 954 188
rect 988 154 1416 188
rect 1450 154 2069 188
rect 74 74 2069 154
rect 74 40 86 74
rect 120 40 160 74
rect 194 40 234 74
rect 268 40 308 74
rect 342 40 382 74
rect 416 40 456 74
rect 490 40 530 74
rect 564 40 604 74
rect 638 40 678 74
rect 712 40 752 74
rect 786 40 826 74
rect 860 40 900 74
rect 934 40 974 74
rect 1008 40 1048 74
rect 1082 40 1121 74
rect 1155 40 1194 74
rect 1228 40 1267 74
rect 1301 40 1340 74
rect 1374 40 1413 74
rect 1447 40 1486 74
rect 1520 40 1559 74
rect 1593 40 1632 74
rect 1666 40 1705 74
rect 1739 40 1778 74
rect 1812 40 1851 74
rect 1885 40 1924 74
rect 1958 40 1997 74
rect 2031 40 2069 74
rect 74 0 2069 40
<< via1 >>
rect 417 814 469 819
rect 417 780 426 814
rect 426 780 460 814
rect 460 780 469 814
rect 417 767 469 780
rect 417 732 469 740
rect 417 698 426 732
rect 426 698 460 732
rect 460 698 469 732
rect 417 688 469 698
rect 769 698 778 725
rect 778 698 812 725
rect 812 698 821 725
rect 417 649 469 661
rect 417 615 426 649
rect 426 615 460 649
rect 460 615 469 649
rect 417 609 469 615
rect 769 673 821 698
rect 769 649 821 661
rect 769 615 778 649
rect 778 615 812 649
rect 812 615 821 649
rect 769 609 821 615
rect 417 346 469 352
rect 417 312 426 346
rect 426 312 460 346
rect 460 312 469 346
rect 417 300 469 312
rect 417 274 469 288
rect 417 240 426 274
rect 426 240 460 274
rect 460 240 469 274
rect 769 346 821 350
rect 769 312 778 346
rect 778 312 812 346
rect 812 312 821 346
rect 769 298 821 312
rect 769 274 821 286
rect 417 236 469 240
rect 769 240 778 274
rect 778 240 812 274
rect 812 240 821 274
rect 769 234 821 240
rect 1231 978 1283 984
rect 1231 944 1240 978
rect 1240 944 1274 978
rect 1274 944 1283 978
rect 1231 932 1283 944
rect 1231 896 1283 920
rect 1231 868 1240 896
rect 1240 868 1274 896
rect 1274 868 1283 896
rect 1901 521 1953 525
rect 1698 509 1750 513
rect 1698 475 1707 509
rect 1707 475 1741 509
rect 1741 475 1750 509
rect 1698 461 1750 475
rect 1698 437 1750 449
rect 1698 403 1707 437
rect 1707 403 1741 437
rect 1741 403 1750 437
rect 1901 487 1910 521
rect 1910 487 1944 521
rect 1944 487 1953 521
rect 1901 473 1953 487
rect 1901 449 1953 461
rect 1901 415 1910 449
rect 1910 415 1944 449
rect 1944 415 1953 449
rect 1901 409 1953 415
rect 1698 397 1750 403
<< metal2 >>
rect 1231 984 1283 990
rect 1231 920 1283 932
rect 1231 862 1283 868
rect 417 824 1878 825
tri 1878 824 1879 825 sw
rect 417 819 1879 824
rect 469 773 1879 819
rect 417 740 469 767
tri 469 739 503 773 nw
tri 1856 750 1879 773 ne
tri 1879 750 1953 824 sw
tri 1879 739 1890 750 ne
rect 1890 739 1953 750
tri 1890 731 1898 739 ne
rect 1898 731 1953 739
rect 417 661 469 688
rect 417 352 469 609
rect 417 288 469 300
rect 417 230 469 236
rect 769 730 1675 731
tri 1675 730 1676 731 sw
tri 1898 730 1899 731 ne
rect 1899 730 1953 731
rect 769 725 1676 730
rect 821 679 1676 725
rect 769 661 821 673
tri 821 645 855 679 nw
tri 1653 656 1676 679 ne
tri 1676 656 1750 730 sw
tri 1899 728 1901 730 ne
tri 1676 645 1687 656 ne
rect 1687 645 1750 656
tri 1687 634 1698 645 ne
rect 769 350 821 609
rect 1698 513 1750 645
rect 1698 449 1750 461
rect 1901 525 1953 730
rect 1901 461 1953 473
rect 1901 403 1953 409
rect 1698 391 1750 397
rect 769 286 821 298
rect 769 228 821 234
use nfet_CDNS_5595914180814  nfet_CDNS_5595914180814_0
timestamp 1704896540
transform 1 0 295 0 1 154
box -79 -32 375 232
use nfet_CDNS_5595914180814  nfet_CDNS_5595914180814_1
timestamp 1704896540
transform -1 0 943 0 1 154
box -79 -32 375 232
use nfet_CDNS_5595914180817  nfet_CDNS_5595914180817_0
timestamp 1704896540
transform 1 0 119 0 1 154
box -79 -32 199 232
use nfet_CDNS_5595914180817  nfet_CDNS_5595914180817_1
timestamp 1704896540
transform -1 0 1119 0 1 154
box -79 -32 199 232
use nfet_CDNS_5595914180817  nfet_CDNS_5595914180817_2
timestamp 1704896540
transform 1 0 1285 0 1 154
box -79 -32 199 232
use pfet_CDNS_5595914180810  pfet_CDNS_5595914180810_0
timestamp 1704896540
transform 1 0 295 0 -1 1153
box -119 -66 415 666
use pfet_CDNS_5595914180810  pfet_CDNS_5595914180810_1
timestamp 1704896540
transform -1 0 943 0 -1 1153
box -119 -66 415 666
use pfet_CDNS_5595914180813  pfet_CDNS_5595914180813_0
timestamp 1704896540
transform 1 0 119 0 -1 1153
box -119 -66 239 666
use pfet_CDNS_5595914180813  pfet_CDNS_5595914180813_1
timestamp 1704896540
transform -1 0 1119 0 -1 1153
box -119 -66 239 666
use pfet_CDNS_5595914180813  pfet_CDNS_5595914180813_2
timestamp 1704896540
transform 1 0 1285 0 -1 1153
box -119 -66 239 666
use sky130_fd_io__amuxsplitv2_hvsbt_nand2  sky130_fd_io__amuxsplitv2_hvsbt_nand2_0
timestamp 1704896540
transform 1 0 1566 0 1 71
box -42 24 569 1127
<< labels >>
flabel metal1 s 1039 411 1068 498 3 FreeSans 200 0 0 0 enable_vdda_h
port 2 nsew
flabel metal1 s 1242 533 1270 640 3 FreeSans 200 0 0 0 hold
port 3 nsew
flabel metal1 s 1326 418 1352 500 3 FreeSans 200 0 0 0 reset
port 4 nsew
flabel metal1 s 134 1156 381 1297 3 FreeSans 200 0 0 0 vcc_io
port 5 nsew
flabel metal1 s 123 19 366 137 3 FreeSans 200 0 0 0 vgnd
port 6 nsew
flabel metal1 s 159 403 192 504 3 FreeSans 100 0 0 0 hld_vdda_h_n
port 7 nsew
<< properties >>
string GDS_END 829548
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 804242
<< end >>
