/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */

`ifndef SKY130_FD_IO__TOP_GPIO_OVTV2_PP_BLACKBOX_V
`define SKY130_FD_IO__TOP_GPIO_OVTV2_PP_BLACKBOX_V

/**
 * top_gpio_ovtv2: General Purpose I/0.
 *
 * Verilog stub definition (black box with power pins).
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none

(* blackbox *)
module sky130_fd_io__top_gpio_ovtv2 (
           OUT             ,
           OE_N            ,
           HLD_H_N         ,
           ENABLE_H        ,
           ENABLE_INP_H    ,
           ENABLE_VDDA_H   ,
           ENABLE_VDDIO    ,
           ENABLE_VSWITCH_H,
           INP_DIS         ,
           VTRIP_SEL       ,
           HYS_TRIM        ,
           SLOW            ,
           SLEW_CTL        ,
           HLD_OVR         ,
           ANALOG_EN       ,
           ANALOG_SEL      ,
           ANALOG_POL      ,
           DM              ,
           IB_MODE_SEL     ,
           VINREF          ,
           PAD             ,
           PAD_A_NOESD_H   ,
           PAD_A_ESD_0_H   ,
           PAD_A_ESD_1_H   ,
           AMUXBUS_A       ,
           AMUXBUS_B       ,
           IN              ,
           IN_H            ,
           TIE_HI_ESD      ,
           TIE_LO_ESD      ,
           VDDIO           ,
           VDDIO_Q         ,
           VDDA            ,
           VCCD            ,
           VSWITCH         ,
           VCCHIB          ,
           VSSA            ,
           VSSD            ,
           VSSIO_Q         ,
           VSSIO
       );

input        OUT             ;
input        OE_N            ;
input        HLD_H_N         ;
input        ENABLE_H        ;
input        ENABLE_INP_H    ;
input        ENABLE_VDDA_H   ;
input        ENABLE_VDDIO    ;
input        ENABLE_VSWITCH_H;
input        INP_DIS         ;
input        VTRIP_SEL       ;
input        HYS_TRIM        ;
input        SLOW            ;
input  [1:0] SLEW_CTL        ;
input        HLD_OVR         ;
input        ANALOG_EN       ;
input        ANALOG_SEL      ;
input        ANALOG_POL      ;
input  [2:0] DM              ;
input  [1:0] IB_MODE_SEL     ;
input        VINREF          ;
inout        PAD             ;
inout        PAD_A_NOESD_H   ;
inout        PAD_A_ESD_0_H   ;
inout        PAD_A_ESD_1_H   ;
inout        AMUXBUS_A       ;
inout        AMUXBUS_B       ;
output       IN              ;
output       IN_H            ;
output       TIE_HI_ESD      ;
output       TIE_LO_ESD      ;
inout        VDDIO           ;
inout        VDDIO_Q         ;
inout        VDDA            ;
inout        VCCD            ;
inout        VSWITCH         ;
inout        VCCHIB          ;
inout        VSSA            ;
inout        VSSD            ;
inout        VSSIO_Q         ;
inout        VSSIO           ;
endmodule

`default_nettype wire
`endif  // SKY130_FD_IO__TOP_GPIO_OVTV2_PP_BLACKBOX_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */

`ifndef SKY130_FD_IO__TOP_GPIOV2_PP_BLACKBOX_V
`define SKY130_FD_IO__TOP_GPIOV2_PP_BLACKBOX_V

/**
 * top_gpiov2: General Purpose I/0.
 *
 * Verilog stub definition (black box with power pins).
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none

(* blackbox *)
module sky130_fd_io__top_gpiov2 (
           OUT             ,
           OE_N            ,
           HLD_H_N         ,
           ENABLE_H        ,
           ENABLE_INP_H    ,
           ENABLE_VDDA_H   ,
           ENABLE_VSWITCH_H,
           ENABLE_VDDIO    ,
           INP_DIS         ,
           IB_MODE_SEL     ,
           VTRIP_SEL       ,
           SLOW            ,
           HLD_OVR         ,
           ANALOG_EN       ,
           ANALOG_SEL      ,
           ANALOG_POL      ,
           DM              ,
           PAD             ,
           PAD_A_NOESD_H   ,
           PAD_A_ESD_0_H   ,
           PAD_A_ESD_1_H   ,
           AMUXBUS_A       ,
           AMUXBUS_B       ,
           IN              ,
           IN_H            ,
           TIE_HI_ESD      ,
           TIE_LO_ESD      ,
           VDDIO           ,
           VDDIO_Q         ,
           VDDA            ,
           VCCD            ,
           VSWITCH         ,
           VCCHIB          ,
           VSSA            ,
           VSSD            ,
           VSSIO_Q         ,
           VSSIO
       );

input        OUT             ;
input        OE_N            ;
input        HLD_H_N         ;
input        ENABLE_H        ;
input        ENABLE_INP_H    ;
input        ENABLE_VDDA_H   ;
input        ENABLE_VSWITCH_H;
input        ENABLE_VDDIO    ;
input        INP_DIS         ;
input        IB_MODE_SEL     ;
input        VTRIP_SEL       ;
input        SLOW            ;
input        HLD_OVR         ;
input        ANALOG_EN       ;
input        ANALOG_SEL      ;
input        ANALOG_POL      ;
input  [2:0] DM              ;
inout        PAD             ;
inout        PAD_A_NOESD_H   ;
inout        PAD_A_ESD_0_H   ;
inout        PAD_A_ESD_1_H   ;
inout        AMUXBUS_A       ;
inout        AMUXBUS_B       ;
output       IN              ;
output       IN_H            ;
output       TIE_HI_ESD      ;
output       TIE_LO_ESD      ;
inout        VDDIO           ;
inout        VDDIO_Q         ;
inout        VDDA            ;
inout        VCCD            ;
inout        VSWITCH         ;
inout        VCCHIB          ;
inout        VSSA            ;
inout        VSSD            ;
inout        VSSIO_Q         ;
inout        VSSIO           ;
endmodule

`default_nettype wire
`endif  // SKY130_FD_IO__TOP_GPIOV2_PP_BLACKBOX_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */

`ifndef SKY130_FD_IO__TOP_GROUND_HVC_WPAD_PP_BLACKBOX_V
`define SKY130_FD_IO__TOP_GROUND_HVC_WPAD_PP_BLACKBOX_V

/**
 * top_ground_hvc_wpad: Ground pad.
 *
 * Verilog stub definition (black box with power pins).
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none

(* blackbox *)
module sky130_fd_io__top_ground_hvc_wpad (
           G_PAD      ,
           AMUXBUS_A  ,
           AMUXBUS_B  ,
           OGC_HVC    ,
           DRN_HVC    ,
           SRC_BDY_HVC,
           G_CORE     ,
           VDDIO      ,
           VDDIO_Q    ,
           VDDA       ,
           VCCD       ,
           VSWITCH    ,
           VCCHIB     ,
           VSSA       ,
           VSSD       ,
           VSSIO_Q    ,
           VSSIO
       );

inout G_PAD      ;
inout AMUXBUS_A  ;
inout AMUXBUS_B  ;
inout OGC_HVC    ;
inout DRN_HVC    ;
inout SRC_BDY_HVC;
inout G_CORE     ;
inout VDDIO      ;
inout VDDIO_Q    ;
inout VDDA       ;
inout VCCD       ;
inout VSWITCH    ;
inout VCCHIB     ;
inout VSSA       ;
inout VSSD       ;
inout VSSIO_Q    ;
inout VSSIO      ;
endmodule

`default_nettype wire
`endif  // SKY130_FD_IO__TOP_GROUND_HVC_WPAD_PP_BLACKBOX_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */

`ifndef SKY130_FD_IO__TOP_GROUND_LVC_WPAD_PP_BLACKBOX_V
`define SKY130_FD_IO__TOP_GROUND_LVC_WPAD_PP_BLACKBOX_V

/**
 * top_ground_lvc_wpad: Base ground I/O pad with low voltage clamp.
 *
 * Verilog stub definition (black box with power pins).
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none

(* blackbox *)
module sky130_fd_io__top_ground_lvc_wpad (
           G_PAD       ,
           AMUXBUS_A   ,
           AMUXBUS_B   ,
           SRC_BDY_LVC1,
           SRC_BDY_LVC2,
           OGC_LVC     ,
           DRN_LVC1    ,
           BDY2_B2B    ,
           DRN_LVC2    ,
           G_CORE      ,
           VDDIO       ,
           VDDIO_Q     ,
           VDDA        ,
           VCCD        ,
           VSWITCH     ,
           VCCHIB      ,
           VSSA        ,
           VSSD        ,
           VSSIO_Q     ,
           VSSIO
       );

inout G_PAD       ;
inout AMUXBUS_A   ;
inout AMUXBUS_B   ;
inout SRC_BDY_LVC1;
inout SRC_BDY_LVC2;
inout OGC_LVC     ;
inout DRN_LVC1    ;
inout BDY2_B2B    ;
inout DRN_LVC2    ;
inout G_CORE      ;
inout VDDIO       ;
inout VDDIO_Q     ;
inout VDDA        ;
inout VCCD        ;
inout VSWITCH     ;
inout VCCHIB      ;
inout VSSA        ;
inout VSSD        ;
inout VSSIO_Q     ;
inout VSSIO       ;
endmodule

`default_nettype wire
`endif  // SKY130_FD_IO__TOP_GROUND_LVC_WPAD_PP_BLACKBOX_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */

`ifndef SKY130_FD_IO__TOP_POWER_HVC_WPAD_PP_BLACKBOX_V
`define SKY130_FD_IO__TOP_POWER_HVC_WPAD_PP_BLACKBOX_V

/**
 * top_power_hvc_wpad: A power pad with an ESD high-voltage clamp.
 *
 * Verilog stub definition (black box with power pins).
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none

(* blackbox *)
module sky130_fd_io__top_power_hvc_wpad (
           P_PAD      ,
           AMUXBUS_A  ,
           AMUXBUS_B  ,
           OGC_HVC    ,
           DRN_HVC    ,
           SRC_BDY_HVC,
           P_CORE     ,
           VDDIO      ,
           VDDIO_Q    ,
           VDDA       ,
           VCCD       ,
           VSWITCH    ,
           VCCHIB     ,
           VSSA       ,
           VSSD       ,
           VSSIO_Q    ,
           VSSIO
       );

inout P_PAD      ;
inout AMUXBUS_A  ;
inout AMUXBUS_B  ;
inout OGC_HVC    ;
inout DRN_HVC    ;
inout SRC_BDY_HVC;
inout P_CORE     ;
inout VDDIO      ;
inout VDDIO_Q    ;
inout VDDA       ;
inout VCCD       ;
inout VSWITCH    ;
inout VCCHIB     ;
inout VSSA       ;
inout VSSD       ;
inout VSSIO_Q    ;
inout VSSIO      ;
endmodule

`default_nettype wire
`endif  // SKY130_FD_IO__TOP_POWER_HVC_WPAD_PP_BLACKBOX_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */

`ifndef SKY130_FD_IO__TOP_POWER_HVC_WPADV2_PP_BLACKBOX_V
`define SKY130_FD_IO__TOP_POWER_HVC_WPADV2_PP_BLACKBOX_V

/**
 * top_power_hvc_wpadv2: A power pad with an ESD high-voltage clamp.
 *
 * Verilog stub definition (black box with power pins).
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none

(* blackbox *)
module sky130_fd_io__top_power_hvc_wpadv2 (
           P_PAD      ,
           AMUXBUS_A  ,
           AMUXBUS_B  ,
           OGC_HVC    ,
           DRN_HVC    ,
           SRC_BDY_HVC,
           P_CORE     ,
           VDDIO      ,
           VDDIO_Q    ,
           VDDA       ,
           VCCD       ,
           VSWITCH    ,
           VCCHIB     ,
           VSSA       ,
           VSSD       ,
           VSSIO_Q    ,
           VSSIO
       );

inout P_PAD      ;
inout AMUXBUS_A  ;
inout AMUXBUS_B  ;
inout OGC_HVC    ;
inout DRN_HVC    ;
inout SRC_BDY_HVC;
inout P_CORE     ;
inout VDDIO      ;
inout VDDIO_Q    ;
inout VDDA       ;
inout VCCD       ;
inout VSWITCH    ;
inout VCCHIB     ;
inout VSSA       ;
inout VSSD       ;
inout VSSIO_Q    ;
inout VSSIO      ;
endmodule

`default_nettype wire
`endif  // SKY130_FD_IO__TOP_POWER_HVC_WPADV2_PP_BLACKBOX_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */

`ifndef SKY130_FD_IO__TOP_POWER_LVC_WPAD_PP_BLACKBOX_V
`define SKY130_FD_IO__TOP_POWER_LVC_WPAD_PP_BLACKBOX_V

/**
 * top_power_lvc_wpad: A power pad with an ESD low-voltage clamp.
 *
 * Verilog stub definition (black box with power pins).
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none

(* blackbox *)
module sky130_fd_io__top_power_lvc_wpad (
           P_PAD       ,
           AMUXBUS_A   ,
           AMUXBUS_B   ,
           SRC_BDY_LVC1,
           SRC_BDY_LVC2,
           OGC_LVC     ,
           DRN_LVC1    ,
           BDY2_B2B    ,
           DRN_LVC2    ,
           P_CORE      ,
           VDDIO       ,
           VDDIO_Q     ,
           VDDA        ,
           VCCD        ,
           VSWITCH     ,
           VCCHIB      ,
           VSSA        ,
           VSSD        ,
           VSSIO_Q     ,
           VSSIO
       );

inout P_PAD       ;
inout AMUXBUS_A   ;
inout AMUXBUS_B   ;
inout SRC_BDY_LVC1;
inout SRC_BDY_LVC2;
inout OGC_LVC     ;
inout DRN_LVC1    ;
inout BDY2_B2B    ;
inout DRN_LVC2    ;
inout P_CORE      ;
inout VDDIO       ;
inout VDDIO_Q     ;
inout VDDA        ;
inout VCCD        ;
inout VSWITCH     ;
inout VCCHIB      ;
inout VSSA        ;
inout VSSD        ;
inout VSSIO_Q     ;
inout VSSIO       ;
endmodule

`default_nettype wire
`endif  // SKY130_FD_IO__TOP_POWER_LVC_WPAD_PP_BLACKBOX_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */

`ifndef SKY130_FD_IO__TOP_REFGEN_PP_BLACKBOX_V
`define SKY130_FD_IO__TOP_REFGEN_PP_BLACKBOX_V

/**
 * top_refgen: The REFGEN block (sky130_fd_io__top_refgen) is used to
 *             provide the input trip point (VINREF) for the
 *             differential input buffer in SIO and also
 *             the output buffer regulated output level (VOUTREF).
 *             Verilog HDL for "sky130_fd_io",
 *             "sky130_fd_io_top_refgen" "timing_tmp".
 *
 * Verilog stub definition (black box with power pins).
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none

(* blackbox *)
module sky130_fd_io__top_refgen (
           VINREF      ,
           VOUTREF     ,
           REFLEAK_BIAS,
           HLD_H_N     ,
           IBUF_SEL    ,
           OD_H        ,
           VOHREF      ,
           VREF_SEL    ,
           VREG_EN     ,
           VTRIP_SEL   ,
           VCCD        ,
           VCCHIB      ,
           VDDA        ,
           VDDIO       ,
           VDDIO_Q     ,
           VSSD        ,
           VSSIO       ,
           VSSIO_Q
       );

output VINREF      ;
output VOUTREF     ;
inout  REFLEAK_BIAS;
input  HLD_H_N     ;
input  IBUF_SEL    ;
input  OD_H        ;
input  VOHREF      ;
input  VREF_SEL    ;
input  VREG_EN     ;
input  VTRIP_SEL   ;
inout  VCCD        ;
inout  VCCHIB      ;
inout  VDDA        ;
inout  VDDIO       ;
inout  VDDIO_Q     ;
inout  VSSD        ;
inout  VSSIO       ;
inout  VSSIO_Q     ;
endmodule

`default_nettype wire
`endif  // SKY130_FD_IO__TOP_REFGEN_PP_BLACKBOX_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */

`ifndef SKY130_FD_IO__TOP_REFGEN_NEW_PP_BLACKBOX_V
`define SKY130_FD_IO__TOP_REFGEN_NEW_PP_BLACKBOX_V

/**
 * top_refgen_new: The REFGEN block (sky130_fd_io__top_refgen) is used
 *                 to provide the input trip point (VINREF) for the
 *                 differential input buffer in SIO and also
 *                 the output buffer regulated output level (VOUTREF).
 *
 * Verilog stub definition (black box with power pins).
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none

(* blackbox *)
module sky130_fd_io__top_refgen_new (
           VINREF       ,
           VOUTREF      ,
           REFLEAK_BIAS ,
           AMUXBUS_A    ,
           AMUXBUS_B    ,
           DFT_REFGEN   ,
           HLD_H_N      ,
           IBUF_SEL     ,
           ENABLE_H     ,
           ENABLE_VDDA_H,
           VOH_SEL      ,
           VOHREF       ,
           VREF_SEL     ,
           VREG_EN      ,
           VTRIP_SEL    ,
           VOUTREF_DFT  ,
           VINREF_DFT   ,
           VCCD         ,
           VCCHIB       ,
           VDDA         ,
           VDDIO        ,
           VDDIO_Q      ,
           VSSD         ,
           VSSIO        ,
           VSSIO_Q      ,
           VSWITCH      ,
           VSSA
       );

output       VINREF       ;
output       VOUTREF      ;
inout        REFLEAK_BIAS ;
inout        AMUXBUS_A    ;
inout        AMUXBUS_B    ;
input        DFT_REFGEN   ;
input        HLD_H_N      ;
input        IBUF_SEL     ;
input        ENABLE_H     ;
input        ENABLE_VDDA_H;
input  [2:0] VOH_SEL      ;
input        VOHREF       ;
input  [1:0] VREF_SEL     ;
input        VREG_EN      ;
input        VTRIP_SEL    ;
inout        VOUTREF_DFT  ;
inout        VINREF_DFT   ;
inout        VCCD         ;
inout        VCCHIB       ;
inout        VDDA         ;
inout        VDDIO        ;
inout        VDDIO_Q      ;
inout        VSSD         ;
inout        VSSIO        ;
inout        VSSIO_Q      ;
inout        VSWITCH      ;
inout        VSSA         ;
endmodule

`default_nettype wire
`endif  // SKY130_FD_IO__TOP_REFGEN_NEW_PP_BLACKBOX_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */

`ifndef SKY130_FD_IO__TOP_SIO_PP_BLACKBOX_V
`define SKY130_FD_IO__TOP_SIO_PP_BLACKBOX_V

/**
 * top_sio: Special I/O PAD that provides additionally a
 *          regulated output buffer and a differential input buffer.
 *          SIO cells are ONLY available IN pairs (see top_sio_macro).
 *
 * Verilog stub definition (black box with power pins).
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none

(* blackbox *)
module sky130_fd_io__top_sio (
           IN_H         ,
           PAD_A_NOESD_H,
           PAD          ,
           DM           ,
           HLD_H_N      ,
           INP_DIS      ,
           IN           ,
           ENABLE_H     ,
           OE_N         ,
           SLOW         ,
           VTRIP_SEL    ,
           VINREF       ,
           VOUTREF      ,
           VREG_EN      ,
           IBUF_SEL     ,
           REFLEAK_BIAS ,
           PAD_A_ESD_0_H,
           TIE_LO_ESD   ,
           HLD_OVR      ,
           OUT          ,
           PAD_A_ESD_1_H,
           VSSIO        ,
           VSSIO_Q      ,
           VSSD         ,
           VCCD         ,
           VDDIO        ,
           VCCHIB       ,
           VDDIO_Q
       );

output       IN_H         ;
inout        PAD_A_NOESD_H;
inout        PAD          ;
input  [2:0] DM           ;
input        HLD_H_N      ;
input        INP_DIS      ;
output       IN           ;
input        ENABLE_H     ;
input        OE_N         ;
input        SLOW         ;
input        VTRIP_SEL    ;
input        VINREF       ;
input        VOUTREF      ;
input        VREG_EN      ;
input        IBUF_SEL     ;
input        REFLEAK_BIAS ;
inout        PAD_A_ESD_0_H;
output       TIE_LO_ESD   ;
input        HLD_OVR      ;
input        OUT          ;
inout        PAD_A_ESD_1_H;
inout        VSSIO        ;
inout        VSSIO_Q      ;
inout        VSSD         ;
inout        VCCD         ;
inout        VDDIO        ;
inout        VCCHIB       ;
inout        VDDIO_Q      ;
endmodule

`default_nettype wire
`endif  // SKY130_FD_IO__TOP_SIO_PP_BLACKBOX_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */

`ifndef SKY130_FD_IO__TOP_SIO_MACRO_PP_BLACKBOX_V
`define SKY130_FD_IO__TOP_SIO_MACRO_PP_BLACKBOX_V

/**
 * top_sio_macro: sky130_fd_io__sio_macro consists of two SIO cells
 *                and a reference generator cell.
 *
 * Verilog stub definition (black box with power pins).
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none

(* blackbox *)
module sky130_fd_io__top_sio_macro (
           AMUXBUS_A       ,
           AMUXBUS_B       ,
           VINREF_DFT      ,
           VOUTREF_DFT     ,
           DFT_REFGEN      ,
           HLD_H_N_REFGEN  ,
           IBUF_SEL_REFGEN ,
           ENABLE_VDDA_H   ,
           ENABLE_H        ,
           VOHREF          ,
           VREG_EN_REFGEN  ,
           VTRIP_SEL_REFGEN,
           TIE_LO_ESD      ,
           IN_H            ,
           IN              ,
           PAD_A_NOESD_H   ,
           PAD             ,
           PAD_A_ESD_1_H   ,
           PAD_A_ESD_0_H   ,
           SLOW            ,
           VTRIP_SEL       ,
           HLD_H_N         ,
           VREG_EN         ,
           VOH_SEL         ,
           INP_DIS         ,
           HLD_OVR         ,
           OE_N            ,
           VREF_SEL        ,
           IBUF_SEL        ,
           DM0             ,
           DM1             ,
           OUT             ,
           VCCD            ,
           VCCHIB          ,
           VDDA            ,
           VDDIO           ,
           VDDIO_Q         ,
           VSSD            ,
           VSSIO           ,
           VSSIO_Q         ,
           VSWITCH         ,
           VSSA
       );

inout        AMUXBUS_A       ;
inout        AMUXBUS_B       ;
inout        VINREF_DFT      ;
inout        VOUTREF_DFT     ;
input        DFT_REFGEN      ;
input        HLD_H_N_REFGEN  ;
input        IBUF_SEL_REFGEN ;
input        ENABLE_VDDA_H   ;
input        ENABLE_H        ;
input        VOHREF          ;
input        VREG_EN_REFGEN  ;
input        VTRIP_SEL_REFGEN;
output [1:0] TIE_LO_ESD      ;
output [1:0] IN_H            ;
output [1:0] IN              ;
inout  [1:0] PAD_A_NOESD_H   ;
inout  [1:0] PAD             ;
inout  [1:0] PAD_A_ESD_1_H   ;
inout  [1:0] PAD_A_ESD_0_H   ;
input  [1:0] SLOW            ;
input  [1:0] VTRIP_SEL       ;
input  [1:0] HLD_H_N         ;
input  [1:0] VREG_EN         ;
input  [2:0] VOH_SEL         ;
input  [1:0] INP_DIS         ;
input  [1:0] HLD_OVR         ;
input  [1:0] OE_N            ;
input  [1:0] VREF_SEL        ;
input  [1:0] IBUF_SEL        ;
input  [2:0] DM0             ;
input  [2:0] DM1             ;
input  [1:0] OUT             ;
inout        VCCD            ;
inout        VCCHIB          ;
inout        VDDA            ;
inout        VDDIO           ;
inout        VDDIO_Q         ;
inout        VSSD            ;
inout        VSSIO           ;
inout        VSSIO_Q         ;
inout        VSWITCH         ;
inout        VSSA            ;
endmodule

`default_nettype wire
`endif  // SKY130_FD_IO__TOP_SIO_MACRO_PP_BLACKBOX_V


//--------EOF---------

/**
 * Copyright 2020 The SkyWater PDK Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     https://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */

`ifndef SKY130_FD_IO__TOP_XRES4V2_PP_BLACKBOX_V
`define SKY130_FD_IO__TOP_XRES4V2_PP_BLACKBOX_V

/**
 * top_xres4v2: XRES (Input buffer with Glitch filter).
 *
 * Verilog stub definition (black box with power pins).
 *
 * WARNING: This file is autogenerated, do not modify directly!
 */

`timescale 1ns / 1ps
`default_nettype none

(* blackbox *)
module sky130_fd_io__top_xres4v2 (
           XRES_H_N        ,
           AMUXBUS_A       ,
           AMUXBUS_B       ,
           PAD             ,
           DISABLE_PULLUP_H,
           ENABLE_H        ,
           EN_VDDIO_SIG_H  ,
           INP_SEL_H       ,
           FILT_IN_H       ,
           PULLUP_H        ,
           ENABLE_VDDIO    ,
           PAD_A_ESD_H     ,
           TIE_HI_ESD      ,
           TIE_LO_ESD      ,
           TIE_WEAK_HI_H   ,
           VCCD            ,
           VCCHIB          ,
           VDDA            ,
           VDDIO           ,
           VDDIO_Q         ,
           VSSA            ,
           VSSD            ,
           VSSIO           ,
           VSSIO_Q         ,
           VSWITCH
       );

output XRES_H_N        ;
inout  AMUXBUS_A       ;
inout  AMUXBUS_B       ;
inout  PAD             ;
input  DISABLE_PULLUP_H;
input  ENABLE_H        ;
input  EN_VDDIO_SIG_H  ;
input  INP_SEL_H       ;
input  FILT_IN_H       ;
inout  PULLUP_H        ;
input  ENABLE_VDDIO    ;
inout  PAD_A_ESD_H     ;
output TIE_HI_ESD      ;
output TIE_LO_ESD      ;
inout  TIE_WEAK_HI_H   ;
input  VCCD            ;
input  VCCHIB          ;
input  VDDA            ;
input  VDDIO           ;
input  VDDIO_Q         ;
input  VSSA            ;
input  VSSD            ;
input  VSSIO           ;
input  VSSIO_Q         ;
input  VSWITCH         ;
endmodule

`default_nettype wire
`endif  // SKY130_FD_IO__TOP_XRES4V2_PP_BLACKBOX_V


//--------EOF---------

