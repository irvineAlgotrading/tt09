magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< dnwell >>
rect 1746 1768 89244 87496
<< nwell >>
rect 1662 87412 89328 87580
rect 1662 1852 1830 87412
rect 89160 1852 89328 87412
rect 1662 1684 89328 1852
<< nsubdiff >>
rect 2057 87513 2107 87537
rect 2057 87479 2065 87513
rect 2099 87479 2107 87513
rect 2057 87455 2107 87479
rect 2393 87513 2443 87537
rect 2393 87479 2401 87513
rect 2435 87479 2443 87513
rect 2393 87455 2443 87479
rect 2729 87513 2779 87537
rect 2729 87479 2737 87513
rect 2771 87479 2779 87513
rect 2729 87455 2779 87479
rect 3065 87513 3115 87537
rect 3065 87479 3073 87513
rect 3107 87479 3115 87513
rect 3065 87455 3115 87479
rect 3401 87513 3451 87537
rect 3401 87479 3409 87513
rect 3443 87479 3451 87513
rect 3401 87455 3451 87479
rect 3737 87513 3787 87537
rect 3737 87479 3745 87513
rect 3779 87479 3787 87513
rect 3737 87455 3787 87479
rect 4073 87513 4123 87537
rect 4073 87479 4081 87513
rect 4115 87479 4123 87513
rect 4073 87455 4123 87479
rect 4409 87513 4459 87537
rect 4409 87479 4417 87513
rect 4451 87479 4459 87513
rect 4409 87455 4459 87479
rect 4745 87513 4795 87537
rect 4745 87479 4753 87513
rect 4787 87479 4795 87513
rect 4745 87455 4795 87479
rect 5081 87513 5131 87537
rect 5081 87479 5089 87513
rect 5123 87479 5131 87513
rect 5081 87455 5131 87479
rect 5417 87513 5467 87537
rect 5417 87479 5425 87513
rect 5459 87479 5467 87513
rect 5417 87455 5467 87479
rect 5753 87513 5803 87537
rect 5753 87479 5761 87513
rect 5795 87479 5803 87513
rect 5753 87455 5803 87479
rect 6089 87513 6139 87537
rect 6089 87479 6097 87513
rect 6131 87479 6139 87513
rect 6089 87455 6139 87479
rect 6425 87513 6475 87537
rect 6425 87479 6433 87513
rect 6467 87479 6475 87513
rect 6425 87455 6475 87479
rect 6761 87513 6811 87537
rect 6761 87479 6769 87513
rect 6803 87479 6811 87513
rect 6761 87455 6811 87479
rect 7097 87513 7147 87537
rect 7097 87479 7105 87513
rect 7139 87479 7147 87513
rect 7097 87455 7147 87479
rect 7433 87513 7483 87537
rect 7433 87479 7441 87513
rect 7475 87479 7483 87513
rect 7433 87455 7483 87479
rect 7769 87513 7819 87537
rect 7769 87479 7777 87513
rect 7811 87479 7819 87513
rect 7769 87455 7819 87479
rect 8105 87513 8155 87537
rect 8105 87479 8113 87513
rect 8147 87479 8155 87513
rect 8105 87455 8155 87479
rect 8441 87513 8491 87537
rect 8441 87479 8449 87513
rect 8483 87479 8491 87513
rect 8441 87455 8491 87479
rect 8777 87513 8827 87537
rect 8777 87479 8785 87513
rect 8819 87479 8827 87513
rect 8777 87455 8827 87479
rect 9113 87513 9163 87537
rect 9113 87479 9121 87513
rect 9155 87479 9163 87513
rect 9113 87455 9163 87479
rect 9449 87513 9499 87537
rect 9449 87479 9457 87513
rect 9491 87479 9499 87513
rect 9449 87455 9499 87479
rect 9785 87513 9835 87537
rect 9785 87479 9793 87513
rect 9827 87479 9835 87513
rect 9785 87455 9835 87479
rect 10121 87513 10171 87537
rect 10121 87479 10129 87513
rect 10163 87479 10171 87513
rect 10121 87455 10171 87479
rect 10457 87513 10507 87537
rect 10457 87479 10465 87513
rect 10499 87479 10507 87513
rect 10457 87455 10507 87479
rect 10793 87513 10843 87537
rect 10793 87479 10801 87513
rect 10835 87479 10843 87513
rect 10793 87455 10843 87479
rect 11129 87513 11179 87537
rect 11129 87479 11137 87513
rect 11171 87479 11179 87513
rect 11129 87455 11179 87479
rect 11465 87513 11515 87537
rect 11465 87479 11473 87513
rect 11507 87479 11515 87513
rect 11465 87455 11515 87479
rect 11801 87513 11851 87537
rect 11801 87479 11809 87513
rect 11843 87479 11851 87513
rect 11801 87455 11851 87479
rect 12137 87513 12187 87537
rect 12137 87479 12145 87513
rect 12179 87479 12187 87513
rect 12137 87455 12187 87479
rect 12473 87513 12523 87537
rect 12473 87479 12481 87513
rect 12515 87479 12523 87513
rect 12473 87455 12523 87479
rect 12809 87513 12859 87537
rect 12809 87479 12817 87513
rect 12851 87479 12859 87513
rect 12809 87455 12859 87479
rect 13145 87513 13195 87537
rect 13145 87479 13153 87513
rect 13187 87479 13195 87513
rect 13145 87455 13195 87479
rect 13481 87513 13531 87537
rect 13481 87479 13489 87513
rect 13523 87479 13531 87513
rect 13481 87455 13531 87479
rect 13817 87513 13867 87537
rect 13817 87479 13825 87513
rect 13859 87479 13867 87513
rect 13817 87455 13867 87479
rect 14153 87513 14203 87537
rect 14153 87479 14161 87513
rect 14195 87479 14203 87513
rect 14153 87455 14203 87479
rect 14489 87513 14539 87537
rect 14489 87479 14497 87513
rect 14531 87479 14539 87513
rect 14489 87455 14539 87479
rect 14825 87513 14875 87537
rect 14825 87479 14833 87513
rect 14867 87479 14875 87513
rect 14825 87455 14875 87479
rect 15161 87513 15211 87537
rect 15161 87479 15169 87513
rect 15203 87479 15211 87513
rect 15161 87455 15211 87479
rect 15497 87513 15547 87537
rect 15497 87479 15505 87513
rect 15539 87479 15547 87513
rect 15497 87455 15547 87479
rect 15833 87513 15883 87537
rect 15833 87479 15841 87513
rect 15875 87479 15883 87513
rect 15833 87455 15883 87479
rect 16169 87513 16219 87537
rect 16169 87479 16177 87513
rect 16211 87479 16219 87513
rect 16169 87455 16219 87479
rect 16505 87513 16555 87537
rect 16505 87479 16513 87513
rect 16547 87479 16555 87513
rect 16505 87455 16555 87479
rect 16841 87513 16891 87537
rect 16841 87479 16849 87513
rect 16883 87479 16891 87513
rect 16841 87455 16891 87479
rect 17177 87513 17227 87537
rect 17177 87479 17185 87513
rect 17219 87479 17227 87513
rect 17177 87455 17227 87479
rect 17513 87513 17563 87537
rect 17513 87479 17521 87513
rect 17555 87479 17563 87513
rect 17513 87455 17563 87479
rect 17849 87513 17899 87537
rect 17849 87479 17857 87513
rect 17891 87479 17899 87513
rect 17849 87455 17899 87479
rect 18185 87513 18235 87537
rect 18185 87479 18193 87513
rect 18227 87479 18235 87513
rect 18185 87455 18235 87479
rect 18521 87513 18571 87537
rect 18521 87479 18529 87513
rect 18563 87479 18571 87513
rect 18521 87455 18571 87479
rect 18857 87513 18907 87537
rect 18857 87479 18865 87513
rect 18899 87479 18907 87513
rect 18857 87455 18907 87479
rect 19193 87513 19243 87537
rect 19193 87479 19201 87513
rect 19235 87479 19243 87513
rect 19193 87455 19243 87479
rect 19529 87513 19579 87537
rect 19529 87479 19537 87513
rect 19571 87479 19579 87513
rect 19529 87455 19579 87479
rect 19865 87513 19915 87537
rect 19865 87479 19873 87513
rect 19907 87479 19915 87513
rect 19865 87455 19915 87479
rect 20201 87513 20251 87537
rect 20201 87479 20209 87513
rect 20243 87479 20251 87513
rect 20201 87455 20251 87479
rect 20537 87513 20587 87537
rect 20537 87479 20545 87513
rect 20579 87479 20587 87513
rect 20537 87455 20587 87479
rect 20873 87513 20923 87537
rect 20873 87479 20881 87513
rect 20915 87479 20923 87513
rect 20873 87455 20923 87479
rect 21209 87513 21259 87537
rect 21209 87479 21217 87513
rect 21251 87479 21259 87513
rect 21209 87455 21259 87479
rect 21545 87513 21595 87537
rect 21545 87479 21553 87513
rect 21587 87479 21595 87513
rect 21545 87455 21595 87479
rect 21881 87513 21931 87537
rect 21881 87479 21889 87513
rect 21923 87479 21931 87513
rect 21881 87455 21931 87479
rect 22217 87513 22267 87537
rect 22217 87479 22225 87513
rect 22259 87479 22267 87513
rect 22217 87455 22267 87479
rect 22553 87513 22603 87537
rect 22553 87479 22561 87513
rect 22595 87479 22603 87513
rect 22553 87455 22603 87479
rect 22889 87513 22939 87537
rect 22889 87479 22897 87513
rect 22931 87479 22939 87513
rect 22889 87455 22939 87479
rect 23225 87513 23275 87537
rect 23225 87479 23233 87513
rect 23267 87479 23275 87513
rect 23225 87455 23275 87479
rect 23561 87513 23611 87537
rect 23561 87479 23569 87513
rect 23603 87479 23611 87513
rect 23561 87455 23611 87479
rect 23897 87513 23947 87537
rect 23897 87479 23905 87513
rect 23939 87479 23947 87513
rect 23897 87455 23947 87479
rect 24233 87513 24283 87537
rect 24233 87479 24241 87513
rect 24275 87479 24283 87513
rect 24233 87455 24283 87479
rect 24569 87513 24619 87537
rect 24569 87479 24577 87513
rect 24611 87479 24619 87513
rect 24569 87455 24619 87479
rect 24905 87513 24955 87537
rect 24905 87479 24913 87513
rect 24947 87479 24955 87513
rect 24905 87455 24955 87479
rect 25241 87513 25291 87537
rect 25241 87479 25249 87513
rect 25283 87479 25291 87513
rect 25241 87455 25291 87479
rect 25577 87513 25627 87537
rect 25577 87479 25585 87513
rect 25619 87479 25627 87513
rect 25577 87455 25627 87479
rect 25913 87513 25963 87537
rect 25913 87479 25921 87513
rect 25955 87479 25963 87513
rect 25913 87455 25963 87479
rect 26249 87513 26299 87537
rect 26249 87479 26257 87513
rect 26291 87479 26299 87513
rect 26249 87455 26299 87479
rect 26585 87513 26635 87537
rect 26585 87479 26593 87513
rect 26627 87479 26635 87513
rect 26585 87455 26635 87479
rect 26921 87513 26971 87537
rect 26921 87479 26929 87513
rect 26963 87479 26971 87513
rect 26921 87455 26971 87479
rect 27257 87513 27307 87537
rect 27257 87479 27265 87513
rect 27299 87479 27307 87513
rect 27257 87455 27307 87479
rect 27593 87513 27643 87537
rect 27593 87479 27601 87513
rect 27635 87479 27643 87513
rect 27593 87455 27643 87479
rect 27929 87513 27979 87537
rect 27929 87479 27937 87513
rect 27971 87479 27979 87513
rect 27929 87455 27979 87479
rect 28265 87513 28315 87537
rect 28265 87479 28273 87513
rect 28307 87479 28315 87513
rect 28265 87455 28315 87479
rect 28601 87513 28651 87537
rect 28601 87479 28609 87513
rect 28643 87479 28651 87513
rect 28601 87455 28651 87479
rect 28937 87513 28987 87537
rect 28937 87479 28945 87513
rect 28979 87479 28987 87513
rect 28937 87455 28987 87479
rect 29273 87513 29323 87537
rect 29273 87479 29281 87513
rect 29315 87479 29323 87513
rect 29273 87455 29323 87479
rect 29609 87513 29659 87537
rect 29609 87479 29617 87513
rect 29651 87479 29659 87513
rect 29609 87455 29659 87479
rect 29945 87513 29995 87537
rect 29945 87479 29953 87513
rect 29987 87479 29995 87513
rect 29945 87455 29995 87479
rect 30281 87513 30331 87537
rect 30281 87479 30289 87513
rect 30323 87479 30331 87513
rect 30281 87455 30331 87479
rect 30617 87513 30667 87537
rect 30617 87479 30625 87513
rect 30659 87479 30667 87513
rect 30617 87455 30667 87479
rect 30953 87513 31003 87537
rect 30953 87479 30961 87513
rect 30995 87479 31003 87513
rect 30953 87455 31003 87479
rect 31289 87513 31339 87537
rect 31289 87479 31297 87513
rect 31331 87479 31339 87513
rect 31289 87455 31339 87479
rect 31625 87513 31675 87537
rect 31625 87479 31633 87513
rect 31667 87479 31675 87513
rect 31625 87455 31675 87479
rect 31961 87513 32011 87537
rect 31961 87479 31969 87513
rect 32003 87479 32011 87513
rect 31961 87455 32011 87479
rect 32297 87513 32347 87537
rect 32297 87479 32305 87513
rect 32339 87479 32347 87513
rect 32297 87455 32347 87479
rect 32633 87513 32683 87537
rect 32633 87479 32641 87513
rect 32675 87479 32683 87513
rect 32633 87455 32683 87479
rect 32969 87513 33019 87537
rect 32969 87479 32977 87513
rect 33011 87479 33019 87513
rect 32969 87455 33019 87479
rect 33305 87513 33355 87537
rect 33305 87479 33313 87513
rect 33347 87479 33355 87513
rect 33305 87455 33355 87479
rect 33641 87513 33691 87537
rect 33641 87479 33649 87513
rect 33683 87479 33691 87513
rect 33641 87455 33691 87479
rect 33977 87513 34027 87537
rect 33977 87479 33985 87513
rect 34019 87479 34027 87513
rect 33977 87455 34027 87479
rect 34313 87513 34363 87537
rect 34313 87479 34321 87513
rect 34355 87479 34363 87513
rect 34313 87455 34363 87479
rect 34649 87513 34699 87537
rect 34649 87479 34657 87513
rect 34691 87479 34699 87513
rect 34649 87455 34699 87479
rect 34985 87513 35035 87537
rect 34985 87479 34993 87513
rect 35027 87479 35035 87513
rect 34985 87455 35035 87479
rect 35321 87513 35371 87537
rect 35321 87479 35329 87513
rect 35363 87479 35371 87513
rect 35321 87455 35371 87479
rect 35657 87513 35707 87537
rect 35657 87479 35665 87513
rect 35699 87479 35707 87513
rect 35657 87455 35707 87479
rect 35993 87513 36043 87537
rect 35993 87479 36001 87513
rect 36035 87479 36043 87513
rect 35993 87455 36043 87479
rect 36329 87513 36379 87537
rect 36329 87479 36337 87513
rect 36371 87479 36379 87513
rect 36329 87455 36379 87479
rect 36665 87513 36715 87537
rect 36665 87479 36673 87513
rect 36707 87479 36715 87513
rect 36665 87455 36715 87479
rect 37001 87513 37051 87537
rect 37001 87479 37009 87513
rect 37043 87479 37051 87513
rect 37001 87455 37051 87479
rect 37337 87513 37387 87537
rect 37337 87479 37345 87513
rect 37379 87479 37387 87513
rect 37337 87455 37387 87479
rect 37673 87513 37723 87537
rect 37673 87479 37681 87513
rect 37715 87479 37723 87513
rect 37673 87455 37723 87479
rect 38009 87513 38059 87537
rect 38009 87479 38017 87513
rect 38051 87479 38059 87513
rect 38009 87455 38059 87479
rect 38345 87513 38395 87537
rect 38345 87479 38353 87513
rect 38387 87479 38395 87513
rect 38345 87455 38395 87479
rect 38681 87513 38731 87537
rect 38681 87479 38689 87513
rect 38723 87479 38731 87513
rect 38681 87455 38731 87479
rect 39017 87513 39067 87537
rect 39017 87479 39025 87513
rect 39059 87479 39067 87513
rect 39017 87455 39067 87479
rect 39353 87513 39403 87537
rect 39353 87479 39361 87513
rect 39395 87479 39403 87513
rect 39353 87455 39403 87479
rect 39689 87513 39739 87537
rect 39689 87479 39697 87513
rect 39731 87479 39739 87513
rect 39689 87455 39739 87479
rect 40025 87513 40075 87537
rect 40025 87479 40033 87513
rect 40067 87479 40075 87513
rect 40025 87455 40075 87479
rect 40361 87513 40411 87537
rect 40361 87479 40369 87513
rect 40403 87479 40411 87513
rect 40361 87455 40411 87479
rect 40697 87513 40747 87537
rect 40697 87479 40705 87513
rect 40739 87479 40747 87513
rect 40697 87455 40747 87479
rect 41033 87513 41083 87537
rect 41033 87479 41041 87513
rect 41075 87479 41083 87513
rect 41033 87455 41083 87479
rect 41369 87513 41419 87537
rect 41369 87479 41377 87513
rect 41411 87479 41419 87513
rect 41369 87455 41419 87479
rect 41705 87513 41755 87537
rect 41705 87479 41713 87513
rect 41747 87479 41755 87513
rect 41705 87455 41755 87479
rect 42041 87513 42091 87537
rect 42041 87479 42049 87513
rect 42083 87479 42091 87513
rect 42041 87455 42091 87479
rect 42377 87513 42427 87537
rect 42377 87479 42385 87513
rect 42419 87479 42427 87513
rect 42377 87455 42427 87479
rect 42713 87513 42763 87537
rect 42713 87479 42721 87513
rect 42755 87479 42763 87513
rect 42713 87455 42763 87479
rect 43049 87513 43099 87537
rect 43049 87479 43057 87513
rect 43091 87479 43099 87513
rect 43049 87455 43099 87479
rect 43385 87513 43435 87537
rect 43385 87479 43393 87513
rect 43427 87479 43435 87513
rect 43385 87455 43435 87479
rect 43721 87513 43771 87537
rect 43721 87479 43729 87513
rect 43763 87479 43771 87513
rect 43721 87455 43771 87479
rect 44057 87513 44107 87537
rect 44057 87479 44065 87513
rect 44099 87479 44107 87513
rect 44057 87455 44107 87479
rect 44393 87513 44443 87537
rect 44393 87479 44401 87513
rect 44435 87479 44443 87513
rect 44393 87455 44443 87479
rect 44729 87513 44779 87537
rect 44729 87479 44737 87513
rect 44771 87479 44779 87513
rect 44729 87455 44779 87479
rect 45065 87513 45115 87537
rect 45065 87479 45073 87513
rect 45107 87479 45115 87513
rect 45065 87455 45115 87479
rect 45401 87513 45451 87537
rect 45401 87479 45409 87513
rect 45443 87479 45451 87513
rect 45401 87455 45451 87479
rect 45737 87513 45787 87537
rect 45737 87479 45745 87513
rect 45779 87479 45787 87513
rect 45737 87455 45787 87479
rect 46073 87513 46123 87537
rect 46073 87479 46081 87513
rect 46115 87479 46123 87513
rect 46073 87455 46123 87479
rect 46409 87513 46459 87537
rect 46409 87479 46417 87513
rect 46451 87479 46459 87513
rect 46409 87455 46459 87479
rect 46745 87513 46795 87537
rect 46745 87479 46753 87513
rect 46787 87479 46795 87513
rect 46745 87455 46795 87479
rect 47081 87513 47131 87537
rect 47081 87479 47089 87513
rect 47123 87479 47131 87513
rect 47081 87455 47131 87479
rect 47417 87513 47467 87537
rect 47417 87479 47425 87513
rect 47459 87479 47467 87513
rect 47417 87455 47467 87479
rect 47753 87513 47803 87537
rect 47753 87479 47761 87513
rect 47795 87479 47803 87513
rect 47753 87455 47803 87479
rect 48089 87513 48139 87537
rect 48089 87479 48097 87513
rect 48131 87479 48139 87513
rect 48089 87455 48139 87479
rect 48425 87513 48475 87537
rect 48425 87479 48433 87513
rect 48467 87479 48475 87513
rect 48425 87455 48475 87479
rect 48761 87513 48811 87537
rect 48761 87479 48769 87513
rect 48803 87479 48811 87513
rect 48761 87455 48811 87479
rect 49097 87513 49147 87537
rect 49097 87479 49105 87513
rect 49139 87479 49147 87513
rect 49097 87455 49147 87479
rect 49433 87513 49483 87537
rect 49433 87479 49441 87513
rect 49475 87479 49483 87513
rect 49433 87455 49483 87479
rect 49769 87513 49819 87537
rect 49769 87479 49777 87513
rect 49811 87479 49819 87513
rect 49769 87455 49819 87479
rect 50105 87513 50155 87537
rect 50105 87479 50113 87513
rect 50147 87479 50155 87513
rect 50105 87455 50155 87479
rect 50441 87513 50491 87537
rect 50441 87479 50449 87513
rect 50483 87479 50491 87513
rect 50441 87455 50491 87479
rect 50777 87513 50827 87537
rect 50777 87479 50785 87513
rect 50819 87479 50827 87513
rect 50777 87455 50827 87479
rect 51113 87513 51163 87537
rect 51113 87479 51121 87513
rect 51155 87479 51163 87513
rect 51113 87455 51163 87479
rect 51449 87513 51499 87537
rect 51449 87479 51457 87513
rect 51491 87479 51499 87513
rect 51449 87455 51499 87479
rect 51785 87513 51835 87537
rect 51785 87479 51793 87513
rect 51827 87479 51835 87513
rect 51785 87455 51835 87479
rect 52121 87513 52171 87537
rect 52121 87479 52129 87513
rect 52163 87479 52171 87513
rect 52121 87455 52171 87479
rect 52457 87513 52507 87537
rect 52457 87479 52465 87513
rect 52499 87479 52507 87513
rect 52457 87455 52507 87479
rect 52793 87513 52843 87537
rect 52793 87479 52801 87513
rect 52835 87479 52843 87513
rect 52793 87455 52843 87479
rect 53129 87513 53179 87537
rect 53129 87479 53137 87513
rect 53171 87479 53179 87513
rect 53129 87455 53179 87479
rect 53465 87513 53515 87537
rect 53465 87479 53473 87513
rect 53507 87479 53515 87513
rect 53465 87455 53515 87479
rect 53801 87513 53851 87537
rect 53801 87479 53809 87513
rect 53843 87479 53851 87513
rect 53801 87455 53851 87479
rect 54137 87513 54187 87537
rect 54137 87479 54145 87513
rect 54179 87479 54187 87513
rect 54137 87455 54187 87479
rect 54473 87513 54523 87537
rect 54473 87479 54481 87513
rect 54515 87479 54523 87513
rect 54473 87455 54523 87479
rect 54809 87513 54859 87537
rect 54809 87479 54817 87513
rect 54851 87479 54859 87513
rect 54809 87455 54859 87479
rect 55145 87513 55195 87537
rect 55145 87479 55153 87513
rect 55187 87479 55195 87513
rect 55145 87455 55195 87479
rect 55481 87513 55531 87537
rect 55481 87479 55489 87513
rect 55523 87479 55531 87513
rect 55481 87455 55531 87479
rect 55817 87513 55867 87537
rect 55817 87479 55825 87513
rect 55859 87479 55867 87513
rect 55817 87455 55867 87479
rect 56153 87513 56203 87537
rect 56153 87479 56161 87513
rect 56195 87479 56203 87513
rect 56153 87455 56203 87479
rect 56489 87513 56539 87537
rect 56489 87479 56497 87513
rect 56531 87479 56539 87513
rect 56489 87455 56539 87479
rect 56825 87513 56875 87537
rect 56825 87479 56833 87513
rect 56867 87479 56875 87513
rect 56825 87455 56875 87479
rect 57161 87513 57211 87537
rect 57161 87479 57169 87513
rect 57203 87479 57211 87513
rect 57161 87455 57211 87479
rect 57497 87513 57547 87537
rect 57497 87479 57505 87513
rect 57539 87479 57547 87513
rect 57497 87455 57547 87479
rect 57833 87513 57883 87537
rect 57833 87479 57841 87513
rect 57875 87479 57883 87513
rect 57833 87455 57883 87479
rect 58169 87513 58219 87537
rect 58169 87479 58177 87513
rect 58211 87479 58219 87513
rect 58169 87455 58219 87479
rect 58505 87513 58555 87537
rect 58505 87479 58513 87513
rect 58547 87479 58555 87513
rect 58505 87455 58555 87479
rect 58841 87513 58891 87537
rect 58841 87479 58849 87513
rect 58883 87479 58891 87513
rect 58841 87455 58891 87479
rect 59177 87513 59227 87537
rect 59177 87479 59185 87513
rect 59219 87479 59227 87513
rect 59177 87455 59227 87479
rect 59513 87513 59563 87537
rect 59513 87479 59521 87513
rect 59555 87479 59563 87513
rect 59513 87455 59563 87479
rect 59849 87513 59899 87537
rect 59849 87479 59857 87513
rect 59891 87479 59899 87513
rect 59849 87455 59899 87479
rect 60185 87513 60235 87537
rect 60185 87479 60193 87513
rect 60227 87479 60235 87513
rect 60185 87455 60235 87479
rect 60521 87513 60571 87537
rect 60521 87479 60529 87513
rect 60563 87479 60571 87513
rect 60521 87455 60571 87479
rect 60857 87513 60907 87537
rect 60857 87479 60865 87513
rect 60899 87479 60907 87513
rect 60857 87455 60907 87479
rect 61193 87513 61243 87537
rect 61193 87479 61201 87513
rect 61235 87479 61243 87513
rect 61193 87455 61243 87479
rect 61529 87513 61579 87537
rect 61529 87479 61537 87513
rect 61571 87479 61579 87513
rect 61529 87455 61579 87479
rect 61865 87513 61915 87537
rect 61865 87479 61873 87513
rect 61907 87479 61915 87513
rect 61865 87455 61915 87479
rect 62201 87513 62251 87537
rect 62201 87479 62209 87513
rect 62243 87479 62251 87513
rect 62201 87455 62251 87479
rect 62537 87513 62587 87537
rect 62537 87479 62545 87513
rect 62579 87479 62587 87513
rect 62537 87455 62587 87479
rect 62873 87513 62923 87537
rect 62873 87479 62881 87513
rect 62915 87479 62923 87513
rect 62873 87455 62923 87479
rect 63209 87513 63259 87537
rect 63209 87479 63217 87513
rect 63251 87479 63259 87513
rect 63209 87455 63259 87479
rect 63545 87513 63595 87537
rect 63545 87479 63553 87513
rect 63587 87479 63595 87513
rect 63545 87455 63595 87479
rect 63881 87513 63931 87537
rect 63881 87479 63889 87513
rect 63923 87479 63931 87513
rect 63881 87455 63931 87479
rect 64217 87513 64267 87537
rect 64217 87479 64225 87513
rect 64259 87479 64267 87513
rect 64217 87455 64267 87479
rect 64553 87513 64603 87537
rect 64553 87479 64561 87513
rect 64595 87479 64603 87513
rect 64553 87455 64603 87479
rect 64889 87513 64939 87537
rect 64889 87479 64897 87513
rect 64931 87479 64939 87513
rect 64889 87455 64939 87479
rect 65225 87513 65275 87537
rect 65225 87479 65233 87513
rect 65267 87479 65275 87513
rect 65225 87455 65275 87479
rect 65561 87513 65611 87537
rect 65561 87479 65569 87513
rect 65603 87479 65611 87513
rect 65561 87455 65611 87479
rect 65897 87513 65947 87537
rect 65897 87479 65905 87513
rect 65939 87479 65947 87513
rect 65897 87455 65947 87479
rect 66233 87513 66283 87537
rect 66233 87479 66241 87513
rect 66275 87479 66283 87513
rect 66233 87455 66283 87479
rect 66569 87513 66619 87537
rect 66569 87479 66577 87513
rect 66611 87479 66619 87513
rect 66569 87455 66619 87479
rect 66905 87513 66955 87537
rect 66905 87479 66913 87513
rect 66947 87479 66955 87513
rect 66905 87455 66955 87479
rect 67241 87513 67291 87537
rect 67241 87479 67249 87513
rect 67283 87479 67291 87513
rect 67241 87455 67291 87479
rect 67577 87513 67627 87537
rect 67577 87479 67585 87513
rect 67619 87479 67627 87513
rect 67577 87455 67627 87479
rect 67913 87513 67963 87537
rect 67913 87479 67921 87513
rect 67955 87479 67963 87513
rect 67913 87455 67963 87479
rect 68249 87513 68299 87537
rect 68249 87479 68257 87513
rect 68291 87479 68299 87513
rect 68249 87455 68299 87479
rect 68585 87513 68635 87537
rect 68585 87479 68593 87513
rect 68627 87479 68635 87513
rect 68585 87455 68635 87479
rect 68921 87513 68971 87537
rect 68921 87479 68929 87513
rect 68963 87479 68971 87513
rect 68921 87455 68971 87479
rect 69257 87513 69307 87537
rect 69257 87479 69265 87513
rect 69299 87479 69307 87513
rect 69257 87455 69307 87479
rect 69593 87513 69643 87537
rect 69593 87479 69601 87513
rect 69635 87479 69643 87513
rect 69593 87455 69643 87479
rect 69929 87513 69979 87537
rect 69929 87479 69937 87513
rect 69971 87479 69979 87513
rect 69929 87455 69979 87479
rect 70265 87513 70315 87537
rect 70265 87479 70273 87513
rect 70307 87479 70315 87513
rect 70265 87455 70315 87479
rect 70601 87513 70651 87537
rect 70601 87479 70609 87513
rect 70643 87479 70651 87513
rect 70601 87455 70651 87479
rect 70937 87513 70987 87537
rect 70937 87479 70945 87513
rect 70979 87479 70987 87513
rect 70937 87455 70987 87479
rect 71273 87513 71323 87537
rect 71273 87479 71281 87513
rect 71315 87479 71323 87513
rect 71273 87455 71323 87479
rect 71609 87513 71659 87537
rect 71609 87479 71617 87513
rect 71651 87479 71659 87513
rect 71609 87455 71659 87479
rect 71945 87513 71995 87537
rect 71945 87479 71953 87513
rect 71987 87479 71995 87513
rect 71945 87455 71995 87479
rect 72281 87513 72331 87537
rect 72281 87479 72289 87513
rect 72323 87479 72331 87513
rect 72281 87455 72331 87479
rect 72617 87513 72667 87537
rect 72617 87479 72625 87513
rect 72659 87479 72667 87513
rect 72617 87455 72667 87479
rect 72953 87513 73003 87537
rect 72953 87479 72961 87513
rect 72995 87479 73003 87513
rect 72953 87455 73003 87479
rect 73289 87513 73339 87537
rect 73289 87479 73297 87513
rect 73331 87479 73339 87513
rect 73289 87455 73339 87479
rect 73625 87513 73675 87537
rect 73625 87479 73633 87513
rect 73667 87479 73675 87513
rect 73625 87455 73675 87479
rect 73961 87513 74011 87537
rect 73961 87479 73969 87513
rect 74003 87479 74011 87513
rect 73961 87455 74011 87479
rect 74297 87513 74347 87537
rect 74297 87479 74305 87513
rect 74339 87479 74347 87513
rect 74297 87455 74347 87479
rect 74633 87513 74683 87537
rect 74633 87479 74641 87513
rect 74675 87479 74683 87513
rect 74633 87455 74683 87479
rect 74969 87513 75019 87537
rect 74969 87479 74977 87513
rect 75011 87479 75019 87513
rect 74969 87455 75019 87479
rect 75305 87513 75355 87537
rect 75305 87479 75313 87513
rect 75347 87479 75355 87513
rect 75305 87455 75355 87479
rect 75641 87513 75691 87537
rect 75641 87479 75649 87513
rect 75683 87479 75691 87513
rect 75641 87455 75691 87479
rect 75977 87513 76027 87537
rect 75977 87479 75985 87513
rect 76019 87479 76027 87513
rect 75977 87455 76027 87479
rect 76313 87513 76363 87537
rect 76313 87479 76321 87513
rect 76355 87479 76363 87513
rect 76313 87455 76363 87479
rect 76649 87513 76699 87537
rect 76649 87479 76657 87513
rect 76691 87479 76699 87513
rect 76649 87455 76699 87479
rect 76985 87513 77035 87537
rect 76985 87479 76993 87513
rect 77027 87479 77035 87513
rect 76985 87455 77035 87479
rect 77321 87513 77371 87537
rect 77321 87479 77329 87513
rect 77363 87479 77371 87513
rect 77321 87455 77371 87479
rect 77657 87513 77707 87537
rect 77657 87479 77665 87513
rect 77699 87479 77707 87513
rect 77657 87455 77707 87479
rect 77993 87513 78043 87537
rect 77993 87479 78001 87513
rect 78035 87479 78043 87513
rect 77993 87455 78043 87479
rect 78329 87513 78379 87537
rect 78329 87479 78337 87513
rect 78371 87479 78379 87513
rect 78329 87455 78379 87479
rect 78665 87513 78715 87537
rect 78665 87479 78673 87513
rect 78707 87479 78715 87513
rect 78665 87455 78715 87479
rect 79001 87513 79051 87537
rect 79001 87479 79009 87513
rect 79043 87479 79051 87513
rect 79001 87455 79051 87479
rect 79337 87513 79387 87537
rect 79337 87479 79345 87513
rect 79379 87479 79387 87513
rect 79337 87455 79387 87479
rect 79673 87513 79723 87537
rect 79673 87479 79681 87513
rect 79715 87479 79723 87513
rect 79673 87455 79723 87479
rect 80009 87513 80059 87537
rect 80009 87479 80017 87513
rect 80051 87479 80059 87513
rect 80009 87455 80059 87479
rect 80345 87513 80395 87537
rect 80345 87479 80353 87513
rect 80387 87479 80395 87513
rect 80345 87455 80395 87479
rect 80681 87513 80731 87537
rect 80681 87479 80689 87513
rect 80723 87479 80731 87513
rect 80681 87455 80731 87479
rect 81017 87513 81067 87537
rect 81017 87479 81025 87513
rect 81059 87479 81067 87513
rect 81017 87455 81067 87479
rect 81353 87513 81403 87537
rect 81353 87479 81361 87513
rect 81395 87479 81403 87513
rect 81353 87455 81403 87479
rect 81689 87513 81739 87537
rect 81689 87479 81697 87513
rect 81731 87479 81739 87513
rect 81689 87455 81739 87479
rect 82025 87513 82075 87537
rect 82025 87479 82033 87513
rect 82067 87479 82075 87513
rect 82025 87455 82075 87479
rect 82361 87513 82411 87537
rect 82361 87479 82369 87513
rect 82403 87479 82411 87513
rect 82361 87455 82411 87479
rect 82697 87513 82747 87537
rect 82697 87479 82705 87513
rect 82739 87479 82747 87513
rect 82697 87455 82747 87479
rect 83033 87513 83083 87537
rect 83033 87479 83041 87513
rect 83075 87479 83083 87513
rect 83033 87455 83083 87479
rect 83369 87513 83419 87537
rect 83369 87479 83377 87513
rect 83411 87479 83419 87513
rect 83369 87455 83419 87479
rect 83705 87513 83755 87537
rect 83705 87479 83713 87513
rect 83747 87479 83755 87513
rect 83705 87455 83755 87479
rect 84041 87513 84091 87537
rect 84041 87479 84049 87513
rect 84083 87479 84091 87513
rect 84041 87455 84091 87479
rect 84377 87513 84427 87537
rect 84377 87479 84385 87513
rect 84419 87479 84427 87513
rect 84377 87455 84427 87479
rect 84713 87513 84763 87537
rect 84713 87479 84721 87513
rect 84755 87479 84763 87513
rect 84713 87455 84763 87479
rect 85049 87513 85099 87537
rect 85049 87479 85057 87513
rect 85091 87479 85099 87513
rect 85049 87455 85099 87479
rect 85385 87513 85435 87537
rect 85385 87479 85393 87513
rect 85427 87479 85435 87513
rect 85385 87455 85435 87479
rect 85721 87513 85771 87537
rect 85721 87479 85729 87513
rect 85763 87479 85771 87513
rect 85721 87455 85771 87479
rect 86057 87513 86107 87537
rect 86057 87479 86065 87513
rect 86099 87479 86107 87513
rect 86057 87455 86107 87479
rect 86393 87513 86443 87537
rect 86393 87479 86401 87513
rect 86435 87479 86443 87513
rect 86393 87455 86443 87479
rect 86729 87513 86779 87537
rect 86729 87479 86737 87513
rect 86771 87479 86779 87513
rect 86729 87455 86779 87479
rect 87065 87513 87115 87537
rect 87065 87479 87073 87513
rect 87107 87479 87115 87513
rect 87065 87455 87115 87479
rect 87401 87513 87451 87537
rect 87401 87479 87409 87513
rect 87443 87479 87451 87513
rect 87401 87455 87451 87479
rect 87737 87513 87787 87537
rect 87737 87479 87745 87513
rect 87779 87479 87787 87513
rect 87737 87455 87787 87479
rect 88073 87513 88123 87537
rect 88073 87479 88081 87513
rect 88115 87479 88123 87513
rect 88073 87455 88123 87479
rect 88409 87513 88459 87537
rect 88409 87479 88417 87513
rect 88451 87479 88459 87513
rect 88409 87455 88459 87479
rect 88745 87513 88795 87537
rect 88745 87479 88753 87513
rect 88787 87479 88795 87513
rect 88745 87455 88795 87479
rect 1721 87129 1771 87153
rect 1721 87095 1729 87129
rect 1763 87095 1771 87129
rect 1721 87071 1771 87095
rect 89219 87129 89269 87153
rect 89219 87095 89227 87129
rect 89261 87095 89269 87129
rect 89219 87071 89269 87095
rect 1721 86793 1771 86817
rect 1721 86759 1729 86793
rect 1763 86759 1771 86793
rect 1721 86735 1771 86759
rect 89219 86793 89269 86817
rect 89219 86759 89227 86793
rect 89261 86759 89269 86793
rect 89219 86735 89269 86759
rect 1721 86457 1771 86481
rect 1721 86423 1729 86457
rect 1763 86423 1771 86457
rect 1721 86399 1771 86423
rect 89219 86457 89269 86481
rect 89219 86423 89227 86457
rect 89261 86423 89269 86457
rect 89219 86399 89269 86423
rect 1721 86121 1771 86145
rect 1721 86087 1729 86121
rect 1763 86087 1771 86121
rect 1721 86063 1771 86087
rect 89219 86121 89269 86145
rect 89219 86087 89227 86121
rect 89261 86087 89269 86121
rect 89219 86063 89269 86087
rect 1721 85785 1771 85809
rect 1721 85751 1729 85785
rect 1763 85751 1771 85785
rect 1721 85727 1771 85751
rect 89219 85785 89269 85809
rect 89219 85751 89227 85785
rect 89261 85751 89269 85785
rect 89219 85727 89269 85751
rect 1721 85449 1771 85473
rect 1721 85415 1729 85449
rect 1763 85415 1771 85449
rect 1721 85391 1771 85415
rect 89219 85449 89269 85473
rect 89219 85415 89227 85449
rect 89261 85415 89269 85449
rect 89219 85391 89269 85415
rect 1721 85113 1771 85137
rect 1721 85079 1729 85113
rect 1763 85079 1771 85113
rect 1721 85055 1771 85079
rect 89219 85113 89269 85137
rect 89219 85079 89227 85113
rect 89261 85079 89269 85113
rect 89219 85055 89269 85079
rect 1721 84777 1771 84801
rect 1721 84743 1729 84777
rect 1763 84743 1771 84777
rect 1721 84719 1771 84743
rect 89219 84777 89269 84801
rect 89219 84743 89227 84777
rect 89261 84743 89269 84777
rect 89219 84719 89269 84743
rect 1721 84441 1771 84465
rect 1721 84407 1729 84441
rect 1763 84407 1771 84441
rect 1721 84383 1771 84407
rect 89219 84441 89269 84465
rect 89219 84407 89227 84441
rect 89261 84407 89269 84441
rect 89219 84383 89269 84407
rect 1721 84105 1771 84129
rect 1721 84071 1729 84105
rect 1763 84071 1771 84105
rect 1721 84047 1771 84071
rect 89219 84105 89269 84129
rect 89219 84071 89227 84105
rect 89261 84071 89269 84105
rect 89219 84047 89269 84071
rect 1721 83769 1771 83793
rect 1721 83735 1729 83769
rect 1763 83735 1771 83769
rect 1721 83711 1771 83735
rect 89219 83769 89269 83793
rect 89219 83735 89227 83769
rect 89261 83735 89269 83769
rect 89219 83711 89269 83735
rect 1721 83433 1771 83457
rect 1721 83399 1729 83433
rect 1763 83399 1771 83433
rect 1721 83375 1771 83399
rect 89219 83433 89269 83457
rect 89219 83399 89227 83433
rect 89261 83399 89269 83433
rect 89219 83375 89269 83399
rect 1721 83097 1771 83121
rect 1721 83063 1729 83097
rect 1763 83063 1771 83097
rect 1721 83039 1771 83063
rect 89219 83097 89269 83121
rect 89219 83063 89227 83097
rect 89261 83063 89269 83097
rect 89219 83039 89269 83063
rect 1721 82761 1771 82785
rect 1721 82727 1729 82761
rect 1763 82727 1771 82761
rect 1721 82703 1771 82727
rect 89219 82761 89269 82785
rect 89219 82727 89227 82761
rect 89261 82727 89269 82761
rect 89219 82703 89269 82727
rect 1721 82425 1771 82449
rect 1721 82391 1729 82425
rect 1763 82391 1771 82425
rect 1721 82367 1771 82391
rect 89219 82425 89269 82449
rect 89219 82391 89227 82425
rect 89261 82391 89269 82425
rect 89219 82367 89269 82391
rect 1721 82089 1771 82113
rect 1721 82055 1729 82089
rect 1763 82055 1771 82089
rect 1721 82031 1771 82055
rect 89219 82089 89269 82113
rect 89219 82055 89227 82089
rect 89261 82055 89269 82089
rect 89219 82031 89269 82055
rect 1721 81753 1771 81777
rect 1721 81719 1729 81753
rect 1763 81719 1771 81753
rect 1721 81695 1771 81719
rect 89219 81753 89269 81777
rect 89219 81719 89227 81753
rect 89261 81719 89269 81753
rect 89219 81695 89269 81719
rect 1721 81417 1771 81441
rect 1721 81383 1729 81417
rect 1763 81383 1771 81417
rect 1721 81359 1771 81383
rect 89219 81417 89269 81441
rect 89219 81383 89227 81417
rect 89261 81383 89269 81417
rect 89219 81359 89269 81383
rect 1721 81081 1771 81105
rect 1721 81047 1729 81081
rect 1763 81047 1771 81081
rect 1721 81023 1771 81047
rect 89219 81081 89269 81105
rect 89219 81047 89227 81081
rect 89261 81047 89269 81081
rect 89219 81023 89269 81047
rect 1721 80745 1771 80769
rect 1721 80711 1729 80745
rect 1763 80711 1771 80745
rect 1721 80687 1771 80711
rect 89219 80745 89269 80769
rect 89219 80711 89227 80745
rect 89261 80711 89269 80745
rect 89219 80687 89269 80711
rect 1721 80409 1771 80433
rect 1721 80375 1729 80409
rect 1763 80375 1771 80409
rect 1721 80351 1771 80375
rect 89219 80409 89269 80433
rect 89219 80375 89227 80409
rect 89261 80375 89269 80409
rect 89219 80351 89269 80375
rect 1721 80073 1771 80097
rect 1721 80039 1729 80073
rect 1763 80039 1771 80073
rect 1721 80015 1771 80039
rect 89219 80073 89269 80097
rect 89219 80039 89227 80073
rect 89261 80039 89269 80073
rect 89219 80015 89269 80039
rect 1721 79737 1771 79761
rect 1721 79703 1729 79737
rect 1763 79703 1771 79737
rect 1721 79679 1771 79703
rect 89219 79737 89269 79761
rect 89219 79703 89227 79737
rect 89261 79703 89269 79737
rect 89219 79679 89269 79703
rect 1721 79401 1771 79425
rect 1721 79367 1729 79401
rect 1763 79367 1771 79401
rect 1721 79343 1771 79367
rect 89219 79401 89269 79425
rect 89219 79367 89227 79401
rect 89261 79367 89269 79401
rect 89219 79343 89269 79367
rect 1721 79065 1771 79089
rect 1721 79031 1729 79065
rect 1763 79031 1771 79065
rect 1721 79007 1771 79031
rect 89219 79065 89269 79089
rect 89219 79031 89227 79065
rect 89261 79031 89269 79065
rect 89219 79007 89269 79031
rect 1721 78729 1771 78753
rect 1721 78695 1729 78729
rect 1763 78695 1771 78729
rect 1721 78671 1771 78695
rect 89219 78729 89269 78753
rect 89219 78695 89227 78729
rect 89261 78695 89269 78729
rect 89219 78671 89269 78695
rect 1721 78393 1771 78417
rect 1721 78359 1729 78393
rect 1763 78359 1771 78393
rect 1721 78335 1771 78359
rect 89219 78393 89269 78417
rect 89219 78359 89227 78393
rect 89261 78359 89269 78393
rect 89219 78335 89269 78359
rect 1721 78057 1771 78081
rect 1721 78023 1729 78057
rect 1763 78023 1771 78057
rect 1721 77999 1771 78023
rect 89219 78057 89269 78081
rect 89219 78023 89227 78057
rect 89261 78023 89269 78057
rect 89219 77999 89269 78023
rect 1721 77721 1771 77745
rect 1721 77687 1729 77721
rect 1763 77687 1771 77721
rect 1721 77663 1771 77687
rect 89219 77721 89269 77745
rect 89219 77687 89227 77721
rect 89261 77687 89269 77721
rect 89219 77663 89269 77687
rect 1721 77385 1771 77409
rect 1721 77351 1729 77385
rect 1763 77351 1771 77385
rect 1721 77327 1771 77351
rect 89219 77385 89269 77409
rect 89219 77351 89227 77385
rect 89261 77351 89269 77385
rect 89219 77327 89269 77351
rect 1721 77049 1771 77073
rect 1721 77015 1729 77049
rect 1763 77015 1771 77049
rect 1721 76991 1771 77015
rect 89219 77049 89269 77073
rect 89219 77015 89227 77049
rect 89261 77015 89269 77049
rect 89219 76991 89269 77015
rect 1721 76713 1771 76737
rect 1721 76679 1729 76713
rect 1763 76679 1771 76713
rect 1721 76655 1771 76679
rect 89219 76713 89269 76737
rect 89219 76679 89227 76713
rect 89261 76679 89269 76713
rect 89219 76655 89269 76679
rect 1721 76377 1771 76401
rect 1721 76343 1729 76377
rect 1763 76343 1771 76377
rect 1721 76319 1771 76343
rect 89219 76377 89269 76401
rect 89219 76343 89227 76377
rect 89261 76343 89269 76377
rect 89219 76319 89269 76343
rect 1721 76041 1771 76065
rect 1721 76007 1729 76041
rect 1763 76007 1771 76041
rect 1721 75983 1771 76007
rect 89219 76041 89269 76065
rect 89219 76007 89227 76041
rect 89261 76007 89269 76041
rect 89219 75983 89269 76007
rect 1721 75705 1771 75729
rect 1721 75671 1729 75705
rect 1763 75671 1771 75705
rect 1721 75647 1771 75671
rect 89219 75705 89269 75729
rect 89219 75671 89227 75705
rect 89261 75671 89269 75705
rect 89219 75647 89269 75671
rect 1721 75369 1771 75393
rect 1721 75335 1729 75369
rect 1763 75335 1771 75369
rect 1721 75311 1771 75335
rect 89219 75369 89269 75393
rect 89219 75335 89227 75369
rect 89261 75335 89269 75369
rect 89219 75311 89269 75335
rect 1721 75033 1771 75057
rect 1721 74999 1729 75033
rect 1763 74999 1771 75033
rect 1721 74975 1771 74999
rect 89219 75033 89269 75057
rect 89219 74999 89227 75033
rect 89261 74999 89269 75033
rect 89219 74975 89269 74999
rect 1721 74697 1771 74721
rect 1721 74663 1729 74697
rect 1763 74663 1771 74697
rect 1721 74639 1771 74663
rect 89219 74697 89269 74721
rect 89219 74663 89227 74697
rect 89261 74663 89269 74697
rect 89219 74639 89269 74663
rect 1721 74361 1771 74385
rect 1721 74327 1729 74361
rect 1763 74327 1771 74361
rect 1721 74303 1771 74327
rect 89219 74361 89269 74385
rect 89219 74327 89227 74361
rect 89261 74327 89269 74361
rect 89219 74303 89269 74327
rect 1721 74025 1771 74049
rect 1721 73991 1729 74025
rect 1763 73991 1771 74025
rect 1721 73967 1771 73991
rect 89219 74025 89269 74049
rect 89219 73991 89227 74025
rect 89261 73991 89269 74025
rect 89219 73967 89269 73991
rect 1721 73689 1771 73713
rect 1721 73655 1729 73689
rect 1763 73655 1771 73689
rect 1721 73631 1771 73655
rect 89219 73689 89269 73713
rect 89219 73655 89227 73689
rect 89261 73655 89269 73689
rect 89219 73631 89269 73655
rect 1721 73353 1771 73377
rect 1721 73319 1729 73353
rect 1763 73319 1771 73353
rect 1721 73295 1771 73319
rect 89219 73353 89269 73377
rect 89219 73319 89227 73353
rect 89261 73319 89269 73353
rect 89219 73295 89269 73319
rect 1721 73017 1771 73041
rect 1721 72983 1729 73017
rect 1763 72983 1771 73017
rect 1721 72959 1771 72983
rect 89219 73017 89269 73041
rect 89219 72983 89227 73017
rect 89261 72983 89269 73017
rect 89219 72959 89269 72983
rect 1721 72681 1771 72705
rect 1721 72647 1729 72681
rect 1763 72647 1771 72681
rect 1721 72623 1771 72647
rect 89219 72681 89269 72705
rect 89219 72647 89227 72681
rect 89261 72647 89269 72681
rect 89219 72623 89269 72647
rect 1721 72345 1771 72369
rect 1721 72311 1729 72345
rect 1763 72311 1771 72345
rect 1721 72287 1771 72311
rect 89219 72345 89269 72369
rect 89219 72311 89227 72345
rect 89261 72311 89269 72345
rect 89219 72287 89269 72311
rect 1721 72009 1771 72033
rect 1721 71975 1729 72009
rect 1763 71975 1771 72009
rect 1721 71951 1771 71975
rect 89219 72009 89269 72033
rect 89219 71975 89227 72009
rect 89261 71975 89269 72009
rect 89219 71951 89269 71975
rect 1721 71673 1771 71697
rect 1721 71639 1729 71673
rect 1763 71639 1771 71673
rect 1721 71615 1771 71639
rect 89219 71673 89269 71697
rect 89219 71639 89227 71673
rect 89261 71639 89269 71673
rect 89219 71615 89269 71639
rect 1721 71337 1771 71361
rect 1721 71303 1729 71337
rect 1763 71303 1771 71337
rect 1721 71279 1771 71303
rect 89219 71337 89269 71361
rect 89219 71303 89227 71337
rect 89261 71303 89269 71337
rect 89219 71279 89269 71303
rect 1721 71001 1771 71025
rect 1721 70967 1729 71001
rect 1763 70967 1771 71001
rect 1721 70943 1771 70967
rect 89219 71001 89269 71025
rect 89219 70967 89227 71001
rect 89261 70967 89269 71001
rect 89219 70943 89269 70967
rect 1721 70665 1771 70689
rect 1721 70631 1729 70665
rect 1763 70631 1771 70665
rect 1721 70607 1771 70631
rect 89219 70665 89269 70689
rect 89219 70631 89227 70665
rect 89261 70631 89269 70665
rect 89219 70607 89269 70631
rect 1721 70329 1771 70353
rect 1721 70295 1729 70329
rect 1763 70295 1771 70329
rect 1721 70271 1771 70295
rect 89219 70329 89269 70353
rect 89219 70295 89227 70329
rect 89261 70295 89269 70329
rect 89219 70271 89269 70295
rect 1721 69993 1771 70017
rect 1721 69959 1729 69993
rect 1763 69959 1771 69993
rect 1721 69935 1771 69959
rect 89219 69993 89269 70017
rect 89219 69959 89227 69993
rect 89261 69959 89269 69993
rect 89219 69935 89269 69959
rect 1721 69657 1771 69681
rect 1721 69623 1729 69657
rect 1763 69623 1771 69657
rect 1721 69599 1771 69623
rect 89219 69657 89269 69681
rect 89219 69623 89227 69657
rect 89261 69623 89269 69657
rect 89219 69599 89269 69623
rect 1721 69321 1771 69345
rect 1721 69287 1729 69321
rect 1763 69287 1771 69321
rect 1721 69263 1771 69287
rect 89219 69321 89269 69345
rect 89219 69287 89227 69321
rect 89261 69287 89269 69321
rect 89219 69263 89269 69287
rect 1721 68985 1771 69009
rect 1721 68951 1729 68985
rect 1763 68951 1771 68985
rect 1721 68927 1771 68951
rect 89219 68985 89269 69009
rect 89219 68951 89227 68985
rect 89261 68951 89269 68985
rect 89219 68927 89269 68951
rect 1721 68649 1771 68673
rect 1721 68615 1729 68649
rect 1763 68615 1771 68649
rect 1721 68591 1771 68615
rect 89219 68649 89269 68673
rect 89219 68615 89227 68649
rect 89261 68615 89269 68649
rect 89219 68591 89269 68615
rect 1721 68313 1771 68337
rect 1721 68279 1729 68313
rect 1763 68279 1771 68313
rect 1721 68255 1771 68279
rect 89219 68313 89269 68337
rect 89219 68279 89227 68313
rect 89261 68279 89269 68313
rect 89219 68255 89269 68279
rect 1721 67977 1771 68001
rect 1721 67943 1729 67977
rect 1763 67943 1771 67977
rect 1721 67919 1771 67943
rect 89219 67977 89269 68001
rect 89219 67943 89227 67977
rect 89261 67943 89269 67977
rect 89219 67919 89269 67943
rect 1721 67641 1771 67665
rect 1721 67607 1729 67641
rect 1763 67607 1771 67641
rect 1721 67583 1771 67607
rect 89219 67641 89269 67665
rect 89219 67607 89227 67641
rect 89261 67607 89269 67641
rect 89219 67583 89269 67607
rect 1721 67305 1771 67329
rect 1721 67271 1729 67305
rect 1763 67271 1771 67305
rect 1721 67247 1771 67271
rect 89219 67305 89269 67329
rect 89219 67271 89227 67305
rect 89261 67271 89269 67305
rect 89219 67247 89269 67271
rect 1721 66969 1771 66993
rect 1721 66935 1729 66969
rect 1763 66935 1771 66969
rect 1721 66911 1771 66935
rect 89219 66969 89269 66993
rect 89219 66935 89227 66969
rect 89261 66935 89269 66969
rect 89219 66911 89269 66935
rect 1721 66633 1771 66657
rect 1721 66599 1729 66633
rect 1763 66599 1771 66633
rect 1721 66575 1771 66599
rect 89219 66633 89269 66657
rect 89219 66599 89227 66633
rect 89261 66599 89269 66633
rect 89219 66575 89269 66599
rect 1721 66297 1771 66321
rect 1721 66263 1729 66297
rect 1763 66263 1771 66297
rect 1721 66239 1771 66263
rect 89219 66297 89269 66321
rect 89219 66263 89227 66297
rect 89261 66263 89269 66297
rect 89219 66239 89269 66263
rect 1721 65961 1771 65985
rect 1721 65927 1729 65961
rect 1763 65927 1771 65961
rect 1721 65903 1771 65927
rect 89219 65961 89269 65985
rect 89219 65927 89227 65961
rect 89261 65927 89269 65961
rect 89219 65903 89269 65927
rect 1721 65625 1771 65649
rect 1721 65591 1729 65625
rect 1763 65591 1771 65625
rect 1721 65567 1771 65591
rect 89219 65625 89269 65649
rect 89219 65591 89227 65625
rect 89261 65591 89269 65625
rect 89219 65567 89269 65591
rect 1721 65289 1771 65313
rect 1721 65255 1729 65289
rect 1763 65255 1771 65289
rect 1721 65231 1771 65255
rect 89219 65289 89269 65313
rect 89219 65255 89227 65289
rect 89261 65255 89269 65289
rect 89219 65231 89269 65255
rect 1721 64953 1771 64977
rect 1721 64919 1729 64953
rect 1763 64919 1771 64953
rect 1721 64895 1771 64919
rect 89219 64953 89269 64977
rect 89219 64919 89227 64953
rect 89261 64919 89269 64953
rect 89219 64895 89269 64919
rect 1721 64617 1771 64641
rect 1721 64583 1729 64617
rect 1763 64583 1771 64617
rect 1721 64559 1771 64583
rect 89219 64617 89269 64641
rect 89219 64583 89227 64617
rect 89261 64583 89269 64617
rect 89219 64559 89269 64583
rect 1721 64281 1771 64305
rect 1721 64247 1729 64281
rect 1763 64247 1771 64281
rect 1721 64223 1771 64247
rect 89219 64281 89269 64305
rect 89219 64247 89227 64281
rect 89261 64247 89269 64281
rect 89219 64223 89269 64247
rect 1721 63945 1771 63969
rect 1721 63911 1729 63945
rect 1763 63911 1771 63945
rect 1721 63887 1771 63911
rect 89219 63945 89269 63969
rect 89219 63911 89227 63945
rect 89261 63911 89269 63945
rect 89219 63887 89269 63911
rect 1721 63609 1771 63633
rect 1721 63575 1729 63609
rect 1763 63575 1771 63609
rect 1721 63551 1771 63575
rect 89219 63609 89269 63633
rect 89219 63575 89227 63609
rect 89261 63575 89269 63609
rect 89219 63551 89269 63575
rect 1721 63273 1771 63297
rect 1721 63239 1729 63273
rect 1763 63239 1771 63273
rect 1721 63215 1771 63239
rect 89219 63273 89269 63297
rect 89219 63239 89227 63273
rect 89261 63239 89269 63273
rect 89219 63215 89269 63239
rect 1721 62937 1771 62961
rect 1721 62903 1729 62937
rect 1763 62903 1771 62937
rect 1721 62879 1771 62903
rect 89219 62937 89269 62961
rect 89219 62903 89227 62937
rect 89261 62903 89269 62937
rect 89219 62879 89269 62903
rect 1721 62601 1771 62625
rect 1721 62567 1729 62601
rect 1763 62567 1771 62601
rect 1721 62543 1771 62567
rect 89219 62601 89269 62625
rect 89219 62567 89227 62601
rect 89261 62567 89269 62601
rect 89219 62543 89269 62567
rect 1721 62265 1771 62289
rect 1721 62231 1729 62265
rect 1763 62231 1771 62265
rect 1721 62207 1771 62231
rect 89219 62265 89269 62289
rect 89219 62231 89227 62265
rect 89261 62231 89269 62265
rect 89219 62207 89269 62231
rect 1721 61929 1771 61953
rect 1721 61895 1729 61929
rect 1763 61895 1771 61929
rect 1721 61871 1771 61895
rect 89219 61929 89269 61953
rect 89219 61895 89227 61929
rect 89261 61895 89269 61929
rect 89219 61871 89269 61895
rect 1721 61593 1771 61617
rect 1721 61559 1729 61593
rect 1763 61559 1771 61593
rect 1721 61535 1771 61559
rect 89219 61593 89269 61617
rect 89219 61559 89227 61593
rect 89261 61559 89269 61593
rect 89219 61535 89269 61559
rect 1721 61257 1771 61281
rect 1721 61223 1729 61257
rect 1763 61223 1771 61257
rect 1721 61199 1771 61223
rect 89219 61257 89269 61281
rect 89219 61223 89227 61257
rect 89261 61223 89269 61257
rect 89219 61199 89269 61223
rect 1721 60921 1771 60945
rect 1721 60887 1729 60921
rect 1763 60887 1771 60921
rect 1721 60863 1771 60887
rect 89219 60921 89269 60945
rect 89219 60887 89227 60921
rect 89261 60887 89269 60921
rect 89219 60863 89269 60887
rect 1721 60585 1771 60609
rect 1721 60551 1729 60585
rect 1763 60551 1771 60585
rect 1721 60527 1771 60551
rect 89219 60585 89269 60609
rect 89219 60551 89227 60585
rect 89261 60551 89269 60585
rect 89219 60527 89269 60551
rect 1721 60249 1771 60273
rect 1721 60215 1729 60249
rect 1763 60215 1771 60249
rect 1721 60191 1771 60215
rect 89219 60249 89269 60273
rect 89219 60215 89227 60249
rect 89261 60215 89269 60249
rect 89219 60191 89269 60215
rect 1721 59913 1771 59937
rect 1721 59879 1729 59913
rect 1763 59879 1771 59913
rect 1721 59855 1771 59879
rect 89219 59913 89269 59937
rect 89219 59879 89227 59913
rect 89261 59879 89269 59913
rect 89219 59855 89269 59879
rect 1721 59577 1771 59601
rect 1721 59543 1729 59577
rect 1763 59543 1771 59577
rect 1721 59519 1771 59543
rect 89219 59577 89269 59601
rect 89219 59543 89227 59577
rect 89261 59543 89269 59577
rect 89219 59519 89269 59543
rect 1721 59241 1771 59265
rect 1721 59207 1729 59241
rect 1763 59207 1771 59241
rect 1721 59183 1771 59207
rect 89219 59241 89269 59265
rect 89219 59207 89227 59241
rect 89261 59207 89269 59241
rect 89219 59183 89269 59207
rect 1721 58905 1771 58929
rect 1721 58871 1729 58905
rect 1763 58871 1771 58905
rect 1721 58847 1771 58871
rect 89219 58905 89269 58929
rect 89219 58871 89227 58905
rect 89261 58871 89269 58905
rect 89219 58847 89269 58871
rect 1721 58569 1771 58593
rect 1721 58535 1729 58569
rect 1763 58535 1771 58569
rect 1721 58511 1771 58535
rect 89219 58569 89269 58593
rect 89219 58535 89227 58569
rect 89261 58535 89269 58569
rect 89219 58511 89269 58535
rect 1721 58233 1771 58257
rect 1721 58199 1729 58233
rect 1763 58199 1771 58233
rect 1721 58175 1771 58199
rect 89219 58233 89269 58257
rect 89219 58199 89227 58233
rect 89261 58199 89269 58233
rect 89219 58175 89269 58199
rect 1721 57897 1771 57921
rect 1721 57863 1729 57897
rect 1763 57863 1771 57897
rect 1721 57839 1771 57863
rect 89219 57897 89269 57921
rect 89219 57863 89227 57897
rect 89261 57863 89269 57897
rect 89219 57839 89269 57863
rect 1721 57561 1771 57585
rect 1721 57527 1729 57561
rect 1763 57527 1771 57561
rect 1721 57503 1771 57527
rect 89219 57561 89269 57585
rect 89219 57527 89227 57561
rect 89261 57527 89269 57561
rect 89219 57503 89269 57527
rect 1721 57225 1771 57249
rect 1721 57191 1729 57225
rect 1763 57191 1771 57225
rect 1721 57167 1771 57191
rect 89219 57225 89269 57249
rect 89219 57191 89227 57225
rect 89261 57191 89269 57225
rect 89219 57167 89269 57191
rect 1721 56889 1771 56913
rect 1721 56855 1729 56889
rect 1763 56855 1771 56889
rect 1721 56831 1771 56855
rect 89219 56889 89269 56913
rect 89219 56855 89227 56889
rect 89261 56855 89269 56889
rect 89219 56831 89269 56855
rect 1721 56553 1771 56577
rect 1721 56519 1729 56553
rect 1763 56519 1771 56553
rect 1721 56495 1771 56519
rect 89219 56553 89269 56577
rect 89219 56519 89227 56553
rect 89261 56519 89269 56553
rect 89219 56495 89269 56519
rect 1721 56217 1771 56241
rect 1721 56183 1729 56217
rect 1763 56183 1771 56217
rect 1721 56159 1771 56183
rect 89219 56217 89269 56241
rect 89219 56183 89227 56217
rect 89261 56183 89269 56217
rect 89219 56159 89269 56183
rect 1721 55881 1771 55905
rect 1721 55847 1729 55881
rect 1763 55847 1771 55881
rect 1721 55823 1771 55847
rect 89219 55881 89269 55905
rect 89219 55847 89227 55881
rect 89261 55847 89269 55881
rect 89219 55823 89269 55847
rect 1721 55545 1771 55569
rect 1721 55511 1729 55545
rect 1763 55511 1771 55545
rect 1721 55487 1771 55511
rect 89219 55545 89269 55569
rect 89219 55511 89227 55545
rect 89261 55511 89269 55545
rect 89219 55487 89269 55511
rect 1721 55209 1771 55233
rect 1721 55175 1729 55209
rect 1763 55175 1771 55209
rect 1721 55151 1771 55175
rect 89219 55209 89269 55233
rect 89219 55175 89227 55209
rect 89261 55175 89269 55209
rect 89219 55151 89269 55175
rect 1721 54873 1771 54897
rect 1721 54839 1729 54873
rect 1763 54839 1771 54873
rect 1721 54815 1771 54839
rect 89219 54873 89269 54897
rect 89219 54839 89227 54873
rect 89261 54839 89269 54873
rect 89219 54815 89269 54839
rect 1721 54537 1771 54561
rect 1721 54503 1729 54537
rect 1763 54503 1771 54537
rect 1721 54479 1771 54503
rect 89219 54537 89269 54561
rect 89219 54503 89227 54537
rect 89261 54503 89269 54537
rect 89219 54479 89269 54503
rect 1721 54201 1771 54225
rect 1721 54167 1729 54201
rect 1763 54167 1771 54201
rect 1721 54143 1771 54167
rect 89219 54201 89269 54225
rect 89219 54167 89227 54201
rect 89261 54167 89269 54201
rect 89219 54143 89269 54167
rect 1721 53865 1771 53889
rect 1721 53831 1729 53865
rect 1763 53831 1771 53865
rect 1721 53807 1771 53831
rect 89219 53865 89269 53889
rect 89219 53831 89227 53865
rect 89261 53831 89269 53865
rect 89219 53807 89269 53831
rect 1721 53529 1771 53553
rect 1721 53495 1729 53529
rect 1763 53495 1771 53529
rect 1721 53471 1771 53495
rect 89219 53529 89269 53553
rect 89219 53495 89227 53529
rect 89261 53495 89269 53529
rect 89219 53471 89269 53495
rect 1721 53193 1771 53217
rect 1721 53159 1729 53193
rect 1763 53159 1771 53193
rect 1721 53135 1771 53159
rect 89219 53193 89269 53217
rect 89219 53159 89227 53193
rect 89261 53159 89269 53193
rect 89219 53135 89269 53159
rect 1721 52857 1771 52881
rect 1721 52823 1729 52857
rect 1763 52823 1771 52857
rect 1721 52799 1771 52823
rect 89219 52857 89269 52881
rect 89219 52823 89227 52857
rect 89261 52823 89269 52857
rect 89219 52799 89269 52823
rect 1721 52521 1771 52545
rect 1721 52487 1729 52521
rect 1763 52487 1771 52521
rect 1721 52463 1771 52487
rect 89219 52521 89269 52545
rect 89219 52487 89227 52521
rect 89261 52487 89269 52521
rect 89219 52463 89269 52487
rect 1721 52185 1771 52209
rect 1721 52151 1729 52185
rect 1763 52151 1771 52185
rect 1721 52127 1771 52151
rect 89219 52185 89269 52209
rect 89219 52151 89227 52185
rect 89261 52151 89269 52185
rect 89219 52127 89269 52151
rect 1721 51849 1771 51873
rect 1721 51815 1729 51849
rect 1763 51815 1771 51849
rect 1721 51791 1771 51815
rect 89219 51849 89269 51873
rect 89219 51815 89227 51849
rect 89261 51815 89269 51849
rect 89219 51791 89269 51815
rect 1721 51513 1771 51537
rect 1721 51479 1729 51513
rect 1763 51479 1771 51513
rect 1721 51455 1771 51479
rect 89219 51513 89269 51537
rect 89219 51479 89227 51513
rect 89261 51479 89269 51513
rect 89219 51455 89269 51479
rect 1721 51177 1771 51201
rect 1721 51143 1729 51177
rect 1763 51143 1771 51177
rect 1721 51119 1771 51143
rect 89219 51177 89269 51201
rect 89219 51143 89227 51177
rect 89261 51143 89269 51177
rect 89219 51119 89269 51143
rect 1721 50841 1771 50865
rect 1721 50807 1729 50841
rect 1763 50807 1771 50841
rect 1721 50783 1771 50807
rect 89219 50841 89269 50865
rect 89219 50807 89227 50841
rect 89261 50807 89269 50841
rect 89219 50783 89269 50807
rect 1721 50505 1771 50529
rect 1721 50471 1729 50505
rect 1763 50471 1771 50505
rect 1721 50447 1771 50471
rect 89219 50505 89269 50529
rect 89219 50471 89227 50505
rect 89261 50471 89269 50505
rect 89219 50447 89269 50471
rect 1721 50169 1771 50193
rect 1721 50135 1729 50169
rect 1763 50135 1771 50169
rect 1721 50111 1771 50135
rect 89219 50169 89269 50193
rect 89219 50135 89227 50169
rect 89261 50135 89269 50169
rect 89219 50111 89269 50135
rect 1721 49833 1771 49857
rect 1721 49799 1729 49833
rect 1763 49799 1771 49833
rect 1721 49775 1771 49799
rect 89219 49833 89269 49857
rect 89219 49799 89227 49833
rect 89261 49799 89269 49833
rect 89219 49775 89269 49799
rect 1721 49497 1771 49521
rect 1721 49463 1729 49497
rect 1763 49463 1771 49497
rect 1721 49439 1771 49463
rect 89219 49497 89269 49521
rect 89219 49463 89227 49497
rect 89261 49463 89269 49497
rect 89219 49439 89269 49463
rect 1721 49161 1771 49185
rect 1721 49127 1729 49161
rect 1763 49127 1771 49161
rect 1721 49103 1771 49127
rect 89219 49161 89269 49185
rect 89219 49127 89227 49161
rect 89261 49127 89269 49161
rect 89219 49103 89269 49127
rect 1721 48825 1771 48849
rect 1721 48791 1729 48825
rect 1763 48791 1771 48825
rect 1721 48767 1771 48791
rect 89219 48825 89269 48849
rect 89219 48791 89227 48825
rect 89261 48791 89269 48825
rect 89219 48767 89269 48791
rect 1721 48489 1771 48513
rect 1721 48455 1729 48489
rect 1763 48455 1771 48489
rect 1721 48431 1771 48455
rect 89219 48489 89269 48513
rect 89219 48455 89227 48489
rect 89261 48455 89269 48489
rect 89219 48431 89269 48455
rect 1721 48153 1771 48177
rect 1721 48119 1729 48153
rect 1763 48119 1771 48153
rect 1721 48095 1771 48119
rect 89219 48153 89269 48177
rect 89219 48119 89227 48153
rect 89261 48119 89269 48153
rect 89219 48095 89269 48119
rect 1721 47817 1771 47841
rect 1721 47783 1729 47817
rect 1763 47783 1771 47817
rect 1721 47759 1771 47783
rect 89219 47817 89269 47841
rect 89219 47783 89227 47817
rect 89261 47783 89269 47817
rect 89219 47759 89269 47783
rect 1721 47481 1771 47505
rect 1721 47447 1729 47481
rect 1763 47447 1771 47481
rect 1721 47423 1771 47447
rect 89219 47481 89269 47505
rect 89219 47447 89227 47481
rect 89261 47447 89269 47481
rect 89219 47423 89269 47447
rect 1721 47145 1771 47169
rect 1721 47111 1729 47145
rect 1763 47111 1771 47145
rect 1721 47087 1771 47111
rect 89219 47145 89269 47169
rect 89219 47111 89227 47145
rect 89261 47111 89269 47145
rect 89219 47087 89269 47111
rect 1721 46809 1771 46833
rect 1721 46775 1729 46809
rect 1763 46775 1771 46809
rect 1721 46751 1771 46775
rect 89219 46809 89269 46833
rect 89219 46775 89227 46809
rect 89261 46775 89269 46809
rect 89219 46751 89269 46775
rect 1721 46473 1771 46497
rect 1721 46439 1729 46473
rect 1763 46439 1771 46473
rect 1721 46415 1771 46439
rect 89219 46473 89269 46497
rect 89219 46439 89227 46473
rect 89261 46439 89269 46473
rect 89219 46415 89269 46439
rect 1721 46137 1771 46161
rect 1721 46103 1729 46137
rect 1763 46103 1771 46137
rect 1721 46079 1771 46103
rect 89219 46137 89269 46161
rect 89219 46103 89227 46137
rect 89261 46103 89269 46137
rect 89219 46079 89269 46103
rect 1721 45801 1771 45825
rect 1721 45767 1729 45801
rect 1763 45767 1771 45801
rect 1721 45743 1771 45767
rect 89219 45801 89269 45825
rect 89219 45767 89227 45801
rect 89261 45767 89269 45801
rect 89219 45743 89269 45767
rect 1721 45465 1771 45489
rect 1721 45431 1729 45465
rect 1763 45431 1771 45465
rect 1721 45407 1771 45431
rect 89219 45465 89269 45489
rect 89219 45431 89227 45465
rect 89261 45431 89269 45465
rect 89219 45407 89269 45431
rect 1721 45129 1771 45153
rect 1721 45095 1729 45129
rect 1763 45095 1771 45129
rect 1721 45071 1771 45095
rect 89219 45129 89269 45153
rect 89219 45095 89227 45129
rect 89261 45095 89269 45129
rect 89219 45071 89269 45095
rect 1721 44793 1771 44817
rect 1721 44759 1729 44793
rect 1763 44759 1771 44793
rect 1721 44735 1771 44759
rect 89219 44793 89269 44817
rect 89219 44759 89227 44793
rect 89261 44759 89269 44793
rect 89219 44735 89269 44759
rect 1721 44457 1771 44481
rect 1721 44423 1729 44457
rect 1763 44423 1771 44457
rect 1721 44399 1771 44423
rect 89219 44457 89269 44481
rect 89219 44423 89227 44457
rect 89261 44423 89269 44457
rect 89219 44399 89269 44423
rect 1721 44121 1771 44145
rect 1721 44087 1729 44121
rect 1763 44087 1771 44121
rect 1721 44063 1771 44087
rect 89219 44121 89269 44145
rect 89219 44087 89227 44121
rect 89261 44087 89269 44121
rect 89219 44063 89269 44087
rect 1721 43785 1771 43809
rect 1721 43751 1729 43785
rect 1763 43751 1771 43785
rect 1721 43727 1771 43751
rect 89219 43785 89269 43809
rect 89219 43751 89227 43785
rect 89261 43751 89269 43785
rect 89219 43727 89269 43751
rect 1721 43449 1771 43473
rect 1721 43415 1729 43449
rect 1763 43415 1771 43449
rect 1721 43391 1771 43415
rect 89219 43449 89269 43473
rect 89219 43415 89227 43449
rect 89261 43415 89269 43449
rect 89219 43391 89269 43415
rect 1721 43113 1771 43137
rect 1721 43079 1729 43113
rect 1763 43079 1771 43113
rect 1721 43055 1771 43079
rect 89219 43113 89269 43137
rect 89219 43079 89227 43113
rect 89261 43079 89269 43113
rect 89219 43055 89269 43079
rect 1721 42777 1771 42801
rect 1721 42743 1729 42777
rect 1763 42743 1771 42777
rect 1721 42719 1771 42743
rect 89219 42777 89269 42801
rect 89219 42743 89227 42777
rect 89261 42743 89269 42777
rect 89219 42719 89269 42743
rect 1721 42441 1771 42465
rect 1721 42407 1729 42441
rect 1763 42407 1771 42441
rect 1721 42383 1771 42407
rect 89219 42441 89269 42465
rect 89219 42407 89227 42441
rect 89261 42407 89269 42441
rect 89219 42383 89269 42407
rect 1721 42105 1771 42129
rect 1721 42071 1729 42105
rect 1763 42071 1771 42105
rect 1721 42047 1771 42071
rect 89219 42105 89269 42129
rect 89219 42071 89227 42105
rect 89261 42071 89269 42105
rect 89219 42047 89269 42071
rect 1721 41769 1771 41793
rect 1721 41735 1729 41769
rect 1763 41735 1771 41769
rect 1721 41711 1771 41735
rect 89219 41769 89269 41793
rect 89219 41735 89227 41769
rect 89261 41735 89269 41769
rect 89219 41711 89269 41735
rect 1721 41433 1771 41457
rect 1721 41399 1729 41433
rect 1763 41399 1771 41433
rect 1721 41375 1771 41399
rect 89219 41433 89269 41457
rect 89219 41399 89227 41433
rect 89261 41399 89269 41433
rect 89219 41375 89269 41399
rect 1721 41097 1771 41121
rect 1721 41063 1729 41097
rect 1763 41063 1771 41097
rect 1721 41039 1771 41063
rect 89219 41097 89269 41121
rect 89219 41063 89227 41097
rect 89261 41063 89269 41097
rect 89219 41039 89269 41063
rect 1721 40761 1771 40785
rect 1721 40727 1729 40761
rect 1763 40727 1771 40761
rect 1721 40703 1771 40727
rect 89219 40761 89269 40785
rect 89219 40727 89227 40761
rect 89261 40727 89269 40761
rect 89219 40703 89269 40727
rect 1721 40425 1771 40449
rect 1721 40391 1729 40425
rect 1763 40391 1771 40425
rect 1721 40367 1771 40391
rect 89219 40425 89269 40449
rect 89219 40391 89227 40425
rect 89261 40391 89269 40425
rect 89219 40367 89269 40391
rect 1721 40089 1771 40113
rect 1721 40055 1729 40089
rect 1763 40055 1771 40089
rect 1721 40031 1771 40055
rect 89219 40089 89269 40113
rect 89219 40055 89227 40089
rect 89261 40055 89269 40089
rect 89219 40031 89269 40055
rect 1721 39753 1771 39777
rect 1721 39719 1729 39753
rect 1763 39719 1771 39753
rect 1721 39695 1771 39719
rect 89219 39753 89269 39777
rect 89219 39719 89227 39753
rect 89261 39719 89269 39753
rect 89219 39695 89269 39719
rect 1721 39417 1771 39441
rect 1721 39383 1729 39417
rect 1763 39383 1771 39417
rect 1721 39359 1771 39383
rect 89219 39417 89269 39441
rect 89219 39383 89227 39417
rect 89261 39383 89269 39417
rect 89219 39359 89269 39383
rect 1721 39081 1771 39105
rect 1721 39047 1729 39081
rect 1763 39047 1771 39081
rect 1721 39023 1771 39047
rect 89219 39081 89269 39105
rect 89219 39047 89227 39081
rect 89261 39047 89269 39081
rect 89219 39023 89269 39047
rect 1721 38745 1771 38769
rect 1721 38711 1729 38745
rect 1763 38711 1771 38745
rect 1721 38687 1771 38711
rect 89219 38745 89269 38769
rect 89219 38711 89227 38745
rect 89261 38711 89269 38745
rect 89219 38687 89269 38711
rect 1721 38409 1771 38433
rect 1721 38375 1729 38409
rect 1763 38375 1771 38409
rect 1721 38351 1771 38375
rect 89219 38409 89269 38433
rect 89219 38375 89227 38409
rect 89261 38375 89269 38409
rect 89219 38351 89269 38375
rect 1721 38073 1771 38097
rect 1721 38039 1729 38073
rect 1763 38039 1771 38073
rect 1721 38015 1771 38039
rect 89219 38073 89269 38097
rect 89219 38039 89227 38073
rect 89261 38039 89269 38073
rect 89219 38015 89269 38039
rect 1721 37737 1771 37761
rect 1721 37703 1729 37737
rect 1763 37703 1771 37737
rect 1721 37679 1771 37703
rect 89219 37737 89269 37761
rect 89219 37703 89227 37737
rect 89261 37703 89269 37737
rect 89219 37679 89269 37703
rect 1721 37401 1771 37425
rect 1721 37367 1729 37401
rect 1763 37367 1771 37401
rect 1721 37343 1771 37367
rect 89219 37401 89269 37425
rect 89219 37367 89227 37401
rect 89261 37367 89269 37401
rect 89219 37343 89269 37367
rect 1721 37065 1771 37089
rect 1721 37031 1729 37065
rect 1763 37031 1771 37065
rect 1721 37007 1771 37031
rect 89219 37065 89269 37089
rect 89219 37031 89227 37065
rect 89261 37031 89269 37065
rect 89219 37007 89269 37031
rect 1721 36729 1771 36753
rect 1721 36695 1729 36729
rect 1763 36695 1771 36729
rect 1721 36671 1771 36695
rect 89219 36729 89269 36753
rect 89219 36695 89227 36729
rect 89261 36695 89269 36729
rect 89219 36671 89269 36695
rect 1721 36393 1771 36417
rect 1721 36359 1729 36393
rect 1763 36359 1771 36393
rect 1721 36335 1771 36359
rect 89219 36393 89269 36417
rect 89219 36359 89227 36393
rect 89261 36359 89269 36393
rect 89219 36335 89269 36359
rect 1721 36057 1771 36081
rect 1721 36023 1729 36057
rect 1763 36023 1771 36057
rect 1721 35999 1771 36023
rect 89219 36057 89269 36081
rect 89219 36023 89227 36057
rect 89261 36023 89269 36057
rect 89219 35999 89269 36023
rect 1721 35721 1771 35745
rect 1721 35687 1729 35721
rect 1763 35687 1771 35721
rect 1721 35663 1771 35687
rect 89219 35721 89269 35745
rect 89219 35687 89227 35721
rect 89261 35687 89269 35721
rect 89219 35663 89269 35687
rect 1721 35385 1771 35409
rect 1721 35351 1729 35385
rect 1763 35351 1771 35385
rect 1721 35327 1771 35351
rect 89219 35385 89269 35409
rect 89219 35351 89227 35385
rect 89261 35351 89269 35385
rect 89219 35327 89269 35351
rect 1721 35049 1771 35073
rect 1721 35015 1729 35049
rect 1763 35015 1771 35049
rect 1721 34991 1771 35015
rect 89219 35049 89269 35073
rect 89219 35015 89227 35049
rect 89261 35015 89269 35049
rect 89219 34991 89269 35015
rect 1721 34713 1771 34737
rect 1721 34679 1729 34713
rect 1763 34679 1771 34713
rect 1721 34655 1771 34679
rect 89219 34713 89269 34737
rect 89219 34679 89227 34713
rect 89261 34679 89269 34713
rect 89219 34655 89269 34679
rect 1721 34377 1771 34401
rect 1721 34343 1729 34377
rect 1763 34343 1771 34377
rect 1721 34319 1771 34343
rect 89219 34377 89269 34401
rect 89219 34343 89227 34377
rect 89261 34343 89269 34377
rect 89219 34319 89269 34343
rect 1721 34041 1771 34065
rect 1721 34007 1729 34041
rect 1763 34007 1771 34041
rect 1721 33983 1771 34007
rect 89219 34041 89269 34065
rect 89219 34007 89227 34041
rect 89261 34007 89269 34041
rect 89219 33983 89269 34007
rect 1721 33705 1771 33729
rect 1721 33671 1729 33705
rect 1763 33671 1771 33705
rect 1721 33647 1771 33671
rect 89219 33705 89269 33729
rect 89219 33671 89227 33705
rect 89261 33671 89269 33705
rect 89219 33647 89269 33671
rect 1721 33369 1771 33393
rect 1721 33335 1729 33369
rect 1763 33335 1771 33369
rect 1721 33311 1771 33335
rect 89219 33369 89269 33393
rect 89219 33335 89227 33369
rect 89261 33335 89269 33369
rect 89219 33311 89269 33335
rect 1721 33033 1771 33057
rect 1721 32999 1729 33033
rect 1763 32999 1771 33033
rect 1721 32975 1771 32999
rect 89219 33033 89269 33057
rect 89219 32999 89227 33033
rect 89261 32999 89269 33033
rect 89219 32975 89269 32999
rect 1721 32697 1771 32721
rect 1721 32663 1729 32697
rect 1763 32663 1771 32697
rect 1721 32639 1771 32663
rect 89219 32697 89269 32721
rect 89219 32663 89227 32697
rect 89261 32663 89269 32697
rect 89219 32639 89269 32663
rect 1721 32361 1771 32385
rect 1721 32327 1729 32361
rect 1763 32327 1771 32361
rect 1721 32303 1771 32327
rect 89219 32361 89269 32385
rect 89219 32327 89227 32361
rect 89261 32327 89269 32361
rect 89219 32303 89269 32327
rect 1721 32025 1771 32049
rect 1721 31991 1729 32025
rect 1763 31991 1771 32025
rect 1721 31967 1771 31991
rect 89219 32025 89269 32049
rect 89219 31991 89227 32025
rect 89261 31991 89269 32025
rect 89219 31967 89269 31991
rect 1721 31689 1771 31713
rect 1721 31655 1729 31689
rect 1763 31655 1771 31689
rect 1721 31631 1771 31655
rect 89219 31689 89269 31713
rect 89219 31655 89227 31689
rect 89261 31655 89269 31689
rect 89219 31631 89269 31655
rect 1721 31353 1771 31377
rect 1721 31319 1729 31353
rect 1763 31319 1771 31353
rect 1721 31295 1771 31319
rect 89219 31353 89269 31377
rect 89219 31319 89227 31353
rect 89261 31319 89269 31353
rect 89219 31295 89269 31319
rect 1721 31017 1771 31041
rect 1721 30983 1729 31017
rect 1763 30983 1771 31017
rect 1721 30959 1771 30983
rect 89219 31017 89269 31041
rect 89219 30983 89227 31017
rect 89261 30983 89269 31017
rect 89219 30959 89269 30983
rect 1721 30681 1771 30705
rect 1721 30647 1729 30681
rect 1763 30647 1771 30681
rect 1721 30623 1771 30647
rect 89219 30681 89269 30705
rect 89219 30647 89227 30681
rect 89261 30647 89269 30681
rect 89219 30623 89269 30647
rect 1721 30345 1771 30369
rect 1721 30311 1729 30345
rect 1763 30311 1771 30345
rect 1721 30287 1771 30311
rect 89219 30345 89269 30369
rect 89219 30311 89227 30345
rect 89261 30311 89269 30345
rect 89219 30287 89269 30311
rect 1721 30009 1771 30033
rect 1721 29975 1729 30009
rect 1763 29975 1771 30009
rect 1721 29951 1771 29975
rect 89219 30009 89269 30033
rect 89219 29975 89227 30009
rect 89261 29975 89269 30009
rect 89219 29951 89269 29975
rect 1721 29673 1771 29697
rect 1721 29639 1729 29673
rect 1763 29639 1771 29673
rect 1721 29615 1771 29639
rect 89219 29673 89269 29697
rect 89219 29639 89227 29673
rect 89261 29639 89269 29673
rect 89219 29615 89269 29639
rect 1721 29337 1771 29361
rect 1721 29303 1729 29337
rect 1763 29303 1771 29337
rect 1721 29279 1771 29303
rect 89219 29337 89269 29361
rect 89219 29303 89227 29337
rect 89261 29303 89269 29337
rect 89219 29279 89269 29303
rect 1721 29001 1771 29025
rect 1721 28967 1729 29001
rect 1763 28967 1771 29001
rect 1721 28943 1771 28967
rect 89219 29001 89269 29025
rect 89219 28967 89227 29001
rect 89261 28967 89269 29001
rect 89219 28943 89269 28967
rect 1721 28665 1771 28689
rect 1721 28631 1729 28665
rect 1763 28631 1771 28665
rect 1721 28607 1771 28631
rect 89219 28665 89269 28689
rect 89219 28631 89227 28665
rect 89261 28631 89269 28665
rect 89219 28607 89269 28631
rect 1721 28329 1771 28353
rect 1721 28295 1729 28329
rect 1763 28295 1771 28329
rect 1721 28271 1771 28295
rect 89219 28329 89269 28353
rect 89219 28295 89227 28329
rect 89261 28295 89269 28329
rect 89219 28271 89269 28295
rect 1721 27993 1771 28017
rect 1721 27959 1729 27993
rect 1763 27959 1771 27993
rect 1721 27935 1771 27959
rect 89219 27993 89269 28017
rect 89219 27959 89227 27993
rect 89261 27959 89269 27993
rect 89219 27935 89269 27959
rect 1721 27657 1771 27681
rect 1721 27623 1729 27657
rect 1763 27623 1771 27657
rect 1721 27599 1771 27623
rect 89219 27657 89269 27681
rect 89219 27623 89227 27657
rect 89261 27623 89269 27657
rect 89219 27599 89269 27623
rect 1721 27321 1771 27345
rect 1721 27287 1729 27321
rect 1763 27287 1771 27321
rect 1721 27263 1771 27287
rect 89219 27321 89269 27345
rect 89219 27287 89227 27321
rect 89261 27287 89269 27321
rect 89219 27263 89269 27287
rect 1721 26985 1771 27009
rect 1721 26951 1729 26985
rect 1763 26951 1771 26985
rect 1721 26927 1771 26951
rect 89219 26985 89269 27009
rect 89219 26951 89227 26985
rect 89261 26951 89269 26985
rect 89219 26927 89269 26951
rect 1721 26649 1771 26673
rect 1721 26615 1729 26649
rect 1763 26615 1771 26649
rect 1721 26591 1771 26615
rect 89219 26649 89269 26673
rect 89219 26615 89227 26649
rect 89261 26615 89269 26649
rect 89219 26591 89269 26615
rect 1721 26313 1771 26337
rect 1721 26279 1729 26313
rect 1763 26279 1771 26313
rect 1721 26255 1771 26279
rect 89219 26313 89269 26337
rect 89219 26279 89227 26313
rect 89261 26279 89269 26313
rect 89219 26255 89269 26279
rect 1721 25977 1771 26001
rect 1721 25943 1729 25977
rect 1763 25943 1771 25977
rect 1721 25919 1771 25943
rect 89219 25977 89269 26001
rect 89219 25943 89227 25977
rect 89261 25943 89269 25977
rect 89219 25919 89269 25943
rect 1721 25641 1771 25665
rect 1721 25607 1729 25641
rect 1763 25607 1771 25641
rect 1721 25583 1771 25607
rect 89219 25641 89269 25665
rect 89219 25607 89227 25641
rect 89261 25607 89269 25641
rect 89219 25583 89269 25607
rect 1721 25305 1771 25329
rect 1721 25271 1729 25305
rect 1763 25271 1771 25305
rect 1721 25247 1771 25271
rect 89219 25305 89269 25329
rect 89219 25271 89227 25305
rect 89261 25271 89269 25305
rect 89219 25247 89269 25271
rect 1721 24969 1771 24993
rect 1721 24935 1729 24969
rect 1763 24935 1771 24969
rect 1721 24911 1771 24935
rect 89219 24969 89269 24993
rect 89219 24935 89227 24969
rect 89261 24935 89269 24969
rect 89219 24911 89269 24935
rect 1721 24633 1771 24657
rect 1721 24599 1729 24633
rect 1763 24599 1771 24633
rect 1721 24575 1771 24599
rect 89219 24633 89269 24657
rect 89219 24599 89227 24633
rect 89261 24599 89269 24633
rect 89219 24575 89269 24599
rect 1721 24297 1771 24321
rect 1721 24263 1729 24297
rect 1763 24263 1771 24297
rect 1721 24239 1771 24263
rect 89219 24297 89269 24321
rect 89219 24263 89227 24297
rect 89261 24263 89269 24297
rect 89219 24239 89269 24263
rect 1721 23961 1771 23985
rect 1721 23927 1729 23961
rect 1763 23927 1771 23961
rect 1721 23903 1771 23927
rect 89219 23961 89269 23985
rect 89219 23927 89227 23961
rect 89261 23927 89269 23961
rect 89219 23903 89269 23927
rect 1721 23625 1771 23649
rect 1721 23591 1729 23625
rect 1763 23591 1771 23625
rect 1721 23567 1771 23591
rect 89219 23625 89269 23649
rect 89219 23591 89227 23625
rect 89261 23591 89269 23625
rect 89219 23567 89269 23591
rect 1721 23289 1771 23313
rect 1721 23255 1729 23289
rect 1763 23255 1771 23289
rect 1721 23231 1771 23255
rect 89219 23289 89269 23313
rect 89219 23255 89227 23289
rect 89261 23255 89269 23289
rect 89219 23231 89269 23255
rect 1721 22953 1771 22977
rect 1721 22919 1729 22953
rect 1763 22919 1771 22953
rect 1721 22895 1771 22919
rect 89219 22953 89269 22977
rect 89219 22919 89227 22953
rect 89261 22919 89269 22953
rect 89219 22895 89269 22919
rect 1721 22617 1771 22641
rect 1721 22583 1729 22617
rect 1763 22583 1771 22617
rect 1721 22559 1771 22583
rect 89219 22617 89269 22641
rect 89219 22583 89227 22617
rect 89261 22583 89269 22617
rect 89219 22559 89269 22583
rect 1721 22281 1771 22305
rect 1721 22247 1729 22281
rect 1763 22247 1771 22281
rect 1721 22223 1771 22247
rect 89219 22281 89269 22305
rect 89219 22247 89227 22281
rect 89261 22247 89269 22281
rect 89219 22223 89269 22247
rect 1721 21945 1771 21969
rect 1721 21911 1729 21945
rect 1763 21911 1771 21945
rect 1721 21887 1771 21911
rect 89219 21945 89269 21969
rect 89219 21911 89227 21945
rect 89261 21911 89269 21945
rect 89219 21887 89269 21911
rect 1721 21609 1771 21633
rect 1721 21575 1729 21609
rect 1763 21575 1771 21609
rect 1721 21551 1771 21575
rect 89219 21609 89269 21633
rect 89219 21575 89227 21609
rect 89261 21575 89269 21609
rect 89219 21551 89269 21575
rect 1721 21273 1771 21297
rect 1721 21239 1729 21273
rect 1763 21239 1771 21273
rect 1721 21215 1771 21239
rect 89219 21273 89269 21297
rect 89219 21239 89227 21273
rect 89261 21239 89269 21273
rect 89219 21215 89269 21239
rect 1721 20937 1771 20961
rect 1721 20903 1729 20937
rect 1763 20903 1771 20937
rect 1721 20879 1771 20903
rect 89219 20937 89269 20961
rect 89219 20903 89227 20937
rect 89261 20903 89269 20937
rect 89219 20879 89269 20903
rect 1721 20601 1771 20625
rect 1721 20567 1729 20601
rect 1763 20567 1771 20601
rect 1721 20543 1771 20567
rect 89219 20601 89269 20625
rect 89219 20567 89227 20601
rect 89261 20567 89269 20601
rect 89219 20543 89269 20567
rect 1721 20265 1771 20289
rect 1721 20231 1729 20265
rect 1763 20231 1771 20265
rect 1721 20207 1771 20231
rect 89219 20265 89269 20289
rect 89219 20231 89227 20265
rect 89261 20231 89269 20265
rect 89219 20207 89269 20231
rect 1721 19929 1771 19953
rect 1721 19895 1729 19929
rect 1763 19895 1771 19929
rect 1721 19871 1771 19895
rect 89219 19929 89269 19953
rect 89219 19895 89227 19929
rect 89261 19895 89269 19929
rect 89219 19871 89269 19895
rect 1721 19593 1771 19617
rect 1721 19559 1729 19593
rect 1763 19559 1771 19593
rect 1721 19535 1771 19559
rect 89219 19593 89269 19617
rect 89219 19559 89227 19593
rect 89261 19559 89269 19593
rect 89219 19535 89269 19559
rect 1721 19257 1771 19281
rect 1721 19223 1729 19257
rect 1763 19223 1771 19257
rect 1721 19199 1771 19223
rect 89219 19257 89269 19281
rect 89219 19223 89227 19257
rect 89261 19223 89269 19257
rect 89219 19199 89269 19223
rect 1721 18921 1771 18945
rect 1721 18887 1729 18921
rect 1763 18887 1771 18921
rect 1721 18863 1771 18887
rect 89219 18921 89269 18945
rect 89219 18887 89227 18921
rect 89261 18887 89269 18921
rect 89219 18863 89269 18887
rect 1721 18585 1771 18609
rect 1721 18551 1729 18585
rect 1763 18551 1771 18585
rect 1721 18527 1771 18551
rect 89219 18585 89269 18609
rect 89219 18551 89227 18585
rect 89261 18551 89269 18585
rect 89219 18527 89269 18551
rect 1721 18249 1771 18273
rect 1721 18215 1729 18249
rect 1763 18215 1771 18249
rect 1721 18191 1771 18215
rect 89219 18249 89269 18273
rect 89219 18215 89227 18249
rect 89261 18215 89269 18249
rect 89219 18191 89269 18215
rect 1721 17913 1771 17937
rect 1721 17879 1729 17913
rect 1763 17879 1771 17913
rect 1721 17855 1771 17879
rect 89219 17913 89269 17937
rect 89219 17879 89227 17913
rect 89261 17879 89269 17913
rect 89219 17855 89269 17879
rect 1721 17577 1771 17601
rect 1721 17543 1729 17577
rect 1763 17543 1771 17577
rect 1721 17519 1771 17543
rect 89219 17577 89269 17601
rect 89219 17543 89227 17577
rect 89261 17543 89269 17577
rect 89219 17519 89269 17543
rect 1721 17241 1771 17265
rect 1721 17207 1729 17241
rect 1763 17207 1771 17241
rect 1721 17183 1771 17207
rect 89219 17241 89269 17265
rect 89219 17207 89227 17241
rect 89261 17207 89269 17241
rect 89219 17183 89269 17207
rect 1721 16905 1771 16929
rect 1721 16871 1729 16905
rect 1763 16871 1771 16905
rect 1721 16847 1771 16871
rect 89219 16905 89269 16929
rect 89219 16871 89227 16905
rect 89261 16871 89269 16905
rect 89219 16847 89269 16871
rect 1721 16569 1771 16593
rect 1721 16535 1729 16569
rect 1763 16535 1771 16569
rect 1721 16511 1771 16535
rect 89219 16569 89269 16593
rect 89219 16535 89227 16569
rect 89261 16535 89269 16569
rect 89219 16511 89269 16535
rect 1721 16233 1771 16257
rect 1721 16199 1729 16233
rect 1763 16199 1771 16233
rect 1721 16175 1771 16199
rect 89219 16233 89269 16257
rect 89219 16199 89227 16233
rect 89261 16199 89269 16233
rect 89219 16175 89269 16199
rect 1721 15897 1771 15921
rect 1721 15863 1729 15897
rect 1763 15863 1771 15897
rect 1721 15839 1771 15863
rect 89219 15897 89269 15921
rect 89219 15863 89227 15897
rect 89261 15863 89269 15897
rect 89219 15839 89269 15863
rect 1721 15561 1771 15585
rect 1721 15527 1729 15561
rect 1763 15527 1771 15561
rect 1721 15503 1771 15527
rect 89219 15561 89269 15585
rect 89219 15527 89227 15561
rect 89261 15527 89269 15561
rect 89219 15503 89269 15527
rect 1721 15225 1771 15249
rect 1721 15191 1729 15225
rect 1763 15191 1771 15225
rect 1721 15167 1771 15191
rect 89219 15225 89269 15249
rect 89219 15191 89227 15225
rect 89261 15191 89269 15225
rect 89219 15167 89269 15191
rect 1721 14889 1771 14913
rect 1721 14855 1729 14889
rect 1763 14855 1771 14889
rect 1721 14831 1771 14855
rect 89219 14889 89269 14913
rect 89219 14855 89227 14889
rect 89261 14855 89269 14889
rect 89219 14831 89269 14855
rect 1721 14553 1771 14577
rect 1721 14519 1729 14553
rect 1763 14519 1771 14553
rect 1721 14495 1771 14519
rect 89219 14553 89269 14577
rect 89219 14519 89227 14553
rect 89261 14519 89269 14553
rect 89219 14495 89269 14519
rect 1721 14217 1771 14241
rect 1721 14183 1729 14217
rect 1763 14183 1771 14217
rect 1721 14159 1771 14183
rect 89219 14217 89269 14241
rect 89219 14183 89227 14217
rect 89261 14183 89269 14217
rect 89219 14159 89269 14183
rect 1721 13881 1771 13905
rect 1721 13847 1729 13881
rect 1763 13847 1771 13881
rect 1721 13823 1771 13847
rect 89219 13881 89269 13905
rect 89219 13847 89227 13881
rect 89261 13847 89269 13881
rect 89219 13823 89269 13847
rect 1721 13545 1771 13569
rect 1721 13511 1729 13545
rect 1763 13511 1771 13545
rect 1721 13487 1771 13511
rect 89219 13545 89269 13569
rect 89219 13511 89227 13545
rect 89261 13511 89269 13545
rect 89219 13487 89269 13511
rect 1721 13209 1771 13233
rect 1721 13175 1729 13209
rect 1763 13175 1771 13209
rect 1721 13151 1771 13175
rect 89219 13209 89269 13233
rect 89219 13175 89227 13209
rect 89261 13175 89269 13209
rect 89219 13151 89269 13175
rect 1721 12873 1771 12897
rect 1721 12839 1729 12873
rect 1763 12839 1771 12873
rect 1721 12815 1771 12839
rect 89219 12873 89269 12897
rect 89219 12839 89227 12873
rect 89261 12839 89269 12873
rect 89219 12815 89269 12839
rect 1721 12537 1771 12561
rect 1721 12503 1729 12537
rect 1763 12503 1771 12537
rect 1721 12479 1771 12503
rect 89219 12537 89269 12561
rect 89219 12503 89227 12537
rect 89261 12503 89269 12537
rect 89219 12479 89269 12503
rect 1721 12201 1771 12225
rect 1721 12167 1729 12201
rect 1763 12167 1771 12201
rect 1721 12143 1771 12167
rect 89219 12201 89269 12225
rect 89219 12167 89227 12201
rect 89261 12167 89269 12201
rect 89219 12143 89269 12167
rect 1721 11865 1771 11889
rect 1721 11831 1729 11865
rect 1763 11831 1771 11865
rect 1721 11807 1771 11831
rect 89219 11865 89269 11889
rect 89219 11831 89227 11865
rect 89261 11831 89269 11865
rect 89219 11807 89269 11831
rect 1721 11529 1771 11553
rect 1721 11495 1729 11529
rect 1763 11495 1771 11529
rect 1721 11471 1771 11495
rect 89219 11529 89269 11553
rect 89219 11495 89227 11529
rect 89261 11495 89269 11529
rect 89219 11471 89269 11495
rect 1721 11193 1771 11217
rect 1721 11159 1729 11193
rect 1763 11159 1771 11193
rect 1721 11135 1771 11159
rect 89219 11193 89269 11217
rect 89219 11159 89227 11193
rect 89261 11159 89269 11193
rect 89219 11135 89269 11159
rect 1721 10857 1771 10881
rect 1721 10823 1729 10857
rect 1763 10823 1771 10857
rect 1721 10799 1771 10823
rect 89219 10857 89269 10881
rect 89219 10823 89227 10857
rect 89261 10823 89269 10857
rect 89219 10799 89269 10823
rect 1721 10521 1771 10545
rect 1721 10487 1729 10521
rect 1763 10487 1771 10521
rect 1721 10463 1771 10487
rect 89219 10521 89269 10545
rect 89219 10487 89227 10521
rect 89261 10487 89269 10521
rect 89219 10463 89269 10487
rect 1721 10185 1771 10209
rect 1721 10151 1729 10185
rect 1763 10151 1771 10185
rect 1721 10127 1771 10151
rect 89219 10185 89269 10209
rect 89219 10151 89227 10185
rect 89261 10151 89269 10185
rect 89219 10127 89269 10151
rect 1721 9849 1771 9873
rect 1721 9815 1729 9849
rect 1763 9815 1771 9849
rect 1721 9791 1771 9815
rect 89219 9849 89269 9873
rect 89219 9815 89227 9849
rect 89261 9815 89269 9849
rect 89219 9791 89269 9815
rect 1721 9513 1771 9537
rect 1721 9479 1729 9513
rect 1763 9479 1771 9513
rect 1721 9455 1771 9479
rect 89219 9513 89269 9537
rect 89219 9479 89227 9513
rect 89261 9479 89269 9513
rect 89219 9455 89269 9479
rect 1721 9177 1771 9201
rect 1721 9143 1729 9177
rect 1763 9143 1771 9177
rect 1721 9119 1771 9143
rect 89219 9177 89269 9201
rect 89219 9143 89227 9177
rect 89261 9143 89269 9177
rect 89219 9119 89269 9143
rect 1721 8841 1771 8865
rect 1721 8807 1729 8841
rect 1763 8807 1771 8841
rect 1721 8783 1771 8807
rect 89219 8841 89269 8865
rect 89219 8807 89227 8841
rect 89261 8807 89269 8841
rect 89219 8783 89269 8807
rect 1721 8505 1771 8529
rect 1721 8471 1729 8505
rect 1763 8471 1771 8505
rect 1721 8447 1771 8471
rect 89219 8505 89269 8529
rect 89219 8471 89227 8505
rect 89261 8471 89269 8505
rect 89219 8447 89269 8471
rect 1721 8169 1771 8193
rect 1721 8135 1729 8169
rect 1763 8135 1771 8169
rect 1721 8111 1771 8135
rect 89219 8169 89269 8193
rect 89219 8135 89227 8169
rect 89261 8135 89269 8169
rect 89219 8111 89269 8135
rect 1721 7833 1771 7857
rect 1721 7799 1729 7833
rect 1763 7799 1771 7833
rect 1721 7775 1771 7799
rect 89219 7833 89269 7857
rect 89219 7799 89227 7833
rect 89261 7799 89269 7833
rect 89219 7775 89269 7799
rect 1721 7497 1771 7521
rect 1721 7463 1729 7497
rect 1763 7463 1771 7497
rect 1721 7439 1771 7463
rect 89219 7497 89269 7521
rect 89219 7463 89227 7497
rect 89261 7463 89269 7497
rect 89219 7439 89269 7463
rect 1721 7161 1771 7185
rect 1721 7127 1729 7161
rect 1763 7127 1771 7161
rect 1721 7103 1771 7127
rect 89219 7161 89269 7185
rect 89219 7127 89227 7161
rect 89261 7127 89269 7161
rect 89219 7103 89269 7127
rect 1721 6825 1771 6849
rect 1721 6791 1729 6825
rect 1763 6791 1771 6825
rect 1721 6767 1771 6791
rect 89219 6825 89269 6849
rect 89219 6791 89227 6825
rect 89261 6791 89269 6825
rect 89219 6767 89269 6791
rect 1721 6489 1771 6513
rect 1721 6455 1729 6489
rect 1763 6455 1771 6489
rect 1721 6431 1771 6455
rect 89219 6489 89269 6513
rect 89219 6455 89227 6489
rect 89261 6455 89269 6489
rect 89219 6431 89269 6455
rect 1721 6153 1771 6177
rect 1721 6119 1729 6153
rect 1763 6119 1771 6153
rect 1721 6095 1771 6119
rect 89219 6153 89269 6177
rect 89219 6119 89227 6153
rect 89261 6119 89269 6153
rect 89219 6095 89269 6119
rect 1721 5817 1771 5841
rect 1721 5783 1729 5817
rect 1763 5783 1771 5817
rect 1721 5759 1771 5783
rect 89219 5817 89269 5841
rect 89219 5783 89227 5817
rect 89261 5783 89269 5817
rect 89219 5759 89269 5783
rect 1721 5481 1771 5505
rect 1721 5447 1729 5481
rect 1763 5447 1771 5481
rect 1721 5423 1771 5447
rect 89219 5481 89269 5505
rect 89219 5447 89227 5481
rect 89261 5447 89269 5481
rect 89219 5423 89269 5447
rect 1721 5145 1771 5169
rect 1721 5111 1729 5145
rect 1763 5111 1771 5145
rect 1721 5087 1771 5111
rect 89219 5145 89269 5169
rect 89219 5111 89227 5145
rect 89261 5111 89269 5145
rect 89219 5087 89269 5111
rect 1721 4809 1771 4833
rect 1721 4775 1729 4809
rect 1763 4775 1771 4809
rect 1721 4751 1771 4775
rect 89219 4809 89269 4833
rect 89219 4775 89227 4809
rect 89261 4775 89269 4809
rect 89219 4751 89269 4775
rect 1721 4473 1771 4497
rect 1721 4439 1729 4473
rect 1763 4439 1771 4473
rect 1721 4415 1771 4439
rect 89219 4473 89269 4497
rect 89219 4439 89227 4473
rect 89261 4439 89269 4473
rect 89219 4415 89269 4439
rect 1721 4137 1771 4161
rect 1721 4103 1729 4137
rect 1763 4103 1771 4137
rect 1721 4079 1771 4103
rect 89219 4137 89269 4161
rect 89219 4103 89227 4137
rect 89261 4103 89269 4137
rect 89219 4079 89269 4103
rect 1721 3801 1771 3825
rect 1721 3767 1729 3801
rect 1763 3767 1771 3801
rect 1721 3743 1771 3767
rect 89219 3801 89269 3825
rect 89219 3767 89227 3801
rect 89261 3767 89269 3801
rect 89219 3743 89269 3767
rect 1721 3465 1771 3489
rect 1721 3431 1729 3465
rect 1763 3431 1771 3465
rect 1721 3407 1771 3431
rect 89219 3465 89269 3489
rect 89219 3431 89227 3465
rect 89261 3431 89269 3465
rect 89219 3407 89269 3431
rect 1721 3129 1771 3153
rect 1721 3095 1729 3129
rect 1763 3095 1771 3129
rect 1721 3071 1771 3095
rect 89219 3129 89269 3153
rect 89219 3095 89227 3129
rect 89261 3095 89269 3129
rect 89219 3071 89269 3095
rect 1721 2793 1771 2817
rect 1721 2759 1729 2793
rect 1763 2759 1771 2793
rect 1721 2735 1771 2759
rect 89219 2793 89269 2817
rect 89219 2759 89227 2793
rect 89261 2759 89269 2793
rect 89219 2735 89269 2759
rect 1721 2457 1771 2481
rect 1721 2423 1729 2457
rect 1763 2423 1771 2457
rect 1721 2399 1771 2423
rect 89219 2457 89269 2481
rect 89219 2423 89227 2457
rect 89261 2423 89269 2457
rect 89219 2399 89269 2423
rect 1721 2121 1771 2145
rect 1721 2087 1729 2121
rect 1763 2087 1771 2121
rect 1721 2063 1771 2087
rect 89219 2121 89269 2145
rect 89219 2087 89227 2121
rect 89261 2087 89269 2121
rect 89219 2063 89269 2087
rect 2057 1785 2107 1809
rect 2057 1751 2065 1785
rect 2099 1751 2107 1785
rect 2057 1727 2107 1751
rect 2393 1785 2443 1809
rect 2393 1751 2401 1785
rect 2435 1751 2443 1785
rect 2393 1727 2443 1751
rect 2729 1785 2779 1809
rect 2729 1751 2737 1785
rect 2771 1751 2779 1785
rect 2729 1727 2779 1751
rect 3065 1785 3115 1809
rect 3065 1751 3073 1785
rect 3107 1751 3115 1785
rect 3065 1727 3115 1751
rect 3401 1785 3451 1809
rect 3401 1751 3409 1785
rect 3443 1751 3451 1785
rect 3401 1727 3451 1751
rect 3737 1785 3787 1809
rect 3737 1751 3745 1785
rect 3779 1751 3787 1785
rect 3737 1727 3787 1751
rect 4073 1785 4123 1809
rect 4073 1751 4081 1785
rect 4115 1751 4123 1785
rect 4073 1727 4123 1751
rect 4409 1785 4459 1809
rect 4409 1751 4417 1785
rect 4451 1751 4459 1785
rect 4409 1727 4459 1751
rect 4745 1785 4795 1809
rect 4745 1751 4753 1785
rect 4787 1751 4795 1785
rect 4745 1727 4795 1751
rect 5081 1785 5131 1809
rect 5081 1751 5089 1785
rect 5123 1751 5131 1785
rect 5081 1727 5131 1751
rect 5417 1785 5467 1809
rect 5417 1751 5425 1785
rect 5459 1751 5467 1785
rect 5417 1727 5467 1751
rect 5753 1785 5803 1809
rect 5753 1751 5761 1785
rect 5795 1751 5803 1785
rect 5753 1727 5803 1751
rect 6089 1785 6139 1809
rect 6089 1751 6097 1785
rect 6131 1751 6139 1785
rect 6089 1727 6139 1751
rect 6425 1785 6475 1809
rect 6425 1751 6433 1785
rect 6467 1751 6475 1785
rect 6425 1727 6475 1751
rect 6761 1785 6811 1809
rect 6761 1751 6769 1785
rect 6803 1751 6811 1785
rect 6761 1727 6811 1751
rect 7097 1785 7147 1809
rect 7097 1751 7105 1785
rect 7139 1751 7147 1785
rect 7097 1727 7147 1751
rect 7433 1785 7483 1809
rect 7433 1751 7441 1785
rect 7475 1751 7483 1785
rect 7433 1727 7483 1751
rect 7769 1785 7819 1809
rect 7769 1751 7777 1785
rect 7811 1751 7819 1785
rect 7769 1727 7819 1751
rect 8105 1785 8155 1809
rect 8105 1751 8113 1785
rect 8147 1751 8155 1785
rect 8105 1727 8155 1751
rect 8441 1785 8491 1809
rect 8441 1751 8449 1785
rect 8483 1751 8491 1785
rect 8441 1727 8491 1751
rect 8777 1785 8827 1809
rect 8777 1751 8785 1785
rect 8819 1751 8827 1785
rect 8777 1727 8827 1751
rect 9113 1785 9163 1809
rect 9113 1751 9121 1785
rect 9155 1751 9163 1785
rect 9113 1727 9163 1751
rect 9449 1785 9499 1809
rect 9449 1751 9457 1785
rect 9491 1751 9499 1785
rect 9449 1727 9499 1751
rect 9785 1785 9835 1809
rect 9785 1751 9793 1785
rect 9827 1751 9835 1785
rect 9785 1727 9835 1751
rect 10121 1785 10171 1809
rect 10121 1751 10129 1785
rect 10163 1751 10171 1785
rect 10121 1727 10171 1751
rect 10457 1785 10507 1809
rect 10457 1751 10465 1785
rect 10499 1751 10507 1785
rect 10457 1727 10507 1751
rect 10793 1785 10843 1809
rect 10793 1751 10801 1785
rect 10835 1751 10843 1785
rect 10793 1727 10843 1751
rect 11129 1785 11179 1809
rect 11129 1751 11137 1785
rect 11171 1751 11179 1785
rect 11129 1727 11179 1751
rect 11465 1785 11515 1809
rect 11465 1751 11473 1785
rect 11507 1751 11515 1785
rect 11465 1727 11515 1751
rect 11801 1785 11851 1809
rect 11801 1751 11809 1785
rect 11843 1751 11851 1785
rect 11801 1727 11851 1751
rect 12137 1785 12187 1809
rect 12137 1751 12145 1785
rect 12179 1751 12187 1785
rect 12137 1727 12187 1751
rect 12473 1785 12523 1809
rect 12473 1751 12481 1785
rect 12515 1751 12523 1785
rect 12473 1727 12523 1751
rect 12809 1785 12859 1809
rect 12809 1751 12817 1785
rect 12851 1751 12859 1785
rect 12809 1727 12859 1751
rect 13145 1785 13195 1809
rect 13145 1751 13153 1785
rect 13187 1751 13195 1785
rect 13145 1727 13195 1751
rect 13481 1785 13531 1809
rect 13481 1751 13489 1785
rect 13523 1751 13531 1785
rect 13481 1727 13531 1751
rect 13817 1785 13867 1809
rect 13817 1751 13825 1785
rect 13859 1751 13867 1785
rect 13817 1727 13867 1751
rect 14153 1785 14203 1809
rect 14153 1751 14161 1785
rect 14195 1751 14203 1785
rect 14153 1727 14203 1751
rect 14489 1785 14539 1809
rect 14489 1751 14497 1785
rect 14531 1751 14539 1785
rect 14489 1727 14539 1751
rect 14825 1785 14875 1809
rect 14825 1751 14833 1785
rect 14867 1751 14875 1785
rect 14825 1727 14875 1751
rect 15161 1785 15211 1809
rect 15161 1751 15169 1785
rect 15203 1751 15211 1785
rect 15161 1727 15211 1751
rect 15497 1785 15547 1809
rect 15497 1751 15505 1785
rect 15539 1751 15547 1785
rect 15497 1727 15547 1751
rect 15833 1785 15883 1809
rect 15833 1751 15841 1785
rect 15875 1751 15883 1785
rect 15833 1727 15883 1751
rect 16169 1785 16219 1809
rect 16169 1751 16177 1785
rect 16211 1751 16219 1785
rect 16169 1727 16219 1751
rect 16505 1785 16555 1809
rect 16505 1751 16513 1785
rect 16547 1751 16555 1785
rect 16505 1727 16555 1751
rect 16841 1785 16891 1809
rect 16841 1751 16849 1785
rect 16883 1751 16891 1785
rect 16841 1727 16891 1751
rect 17177 1785 17227 1809
rect 17177 1751 17185 1785
rect 17219 1751 17227 1785
rect 17177 1727 17227 1751
rect 17513 1785 17563 1809
rect 17513 1751 17521 1785
rect 17555 1751 17563 1785
rect 17513 1727 17563 1751
rect 17849 1785 17899 1809
rect 17849 1751 17857 1785
rect 17891 1751 17899 1785
rect 17849 1727 17899 1751
rect 18185 1785 18235 1809
rect 18185 1751 18193 1785
rect 18227 1751 18235 1785
rect 18185 1727 18235 1751
rect 18521 1785 18571 1809
rect 18521 1751 18529 1785
rect 18563 1751 18571 1785
rect 18521 1727 18571 1751
rect 18857 1785 18907 1809
rect 18857 1751 18865 1785
rect 18899 1751 18907 1785
rect 18857 1727 18907 1751
rect 19193 1785 19243 1809
rect 19193 1751 19201 1785
rect 19235 1751 19243 1785
rect 19193 1727 19243 1751
rect 19529 1785 19579 1809
rect 19529 1751 19537 1785
rect 19571 1751 19579 1785
rect 19529 1727 19579 1751
rect 19865 1785 19915 1809
rect 19865 1751 19873 1785
rect 19907 1751 19915 1785
rect 19865 1727 19915 1751
rect 20201 1785 20251 1809
rect 20201 1751 20209 1785
rect 20243 1751 20251 1785
rect 20201 1727 20251 1751
rect 20537 1785 20587 1809
rect 20537 1751 20545 1785
rect 20579 1751 20587 1785
rect 20537 1727 20587 1751
rect 20873 1785 20923 1809
rect 20873 1751 20881 1785
rect 20915 1751 20923 1785
rect 20873 1727 20923 1751
rect 21209 1785 21259 1809
rect 21209 1751 21217 1785
rect 21251 1751 21259 1785
rect 21209 1727 21259 1751
rect 21545 1785 21595 1809
rect 21545 1751 21553 1785
rect 21587 1751 21595 1785
rect 21545 1727 21595 1751
rect 21881 1785 21931 1809
rect 21881 1751 21889 1785
rect 21923 1751 21931 1785
rect 21881 1727 21931 1751
rect 22217 1785 22267 1809
rect 22217 1751 22225 1785
rect 22259 1751 22267 1785
rect 22217 1727 22267 1751
rect 22553 1785 22603 1809
rect 22553 1751 22561 1785
rect 22595 1751 22603 1785
rect 22553 1727 22603 1751
rect 22889 1785 22939 1809
rect 22889 1751 22897 1785
rect 22931 1751 22939 1785
rect 22889 1727 22939 1751
rect 23225 1785 23275 1809
rect 23225 1751 23233 1785
rect 23267 1751 23275 1785
rect 23225 1727 23275 1751
rect 23561 1785 23611 1809
rect 23561 1751 23569 1785
rect 23603 1751 23611 1785
rect 23561 1727 23611 1751
rect 23897 1785 23947 1809
rect 23897 1751 23905 1785
rect 23939 1751 23947 1785
rect 23897 1727 23947 1751
rect 24233 1785 24283 1809
rect 24233 1751 24241 1785
rect 24275 1751 24283 1785
rect 24233 1727 24283 1751
rect 24569 1785 24619 1809
rect 24569 1751 24577 1785
rect 24611 1751 24619 1785
rect 24569 1727 24619 1751
rect 24905 1785 24955 1809
rect 24905 1751 24913 1785
rect 24947 1751 24955 1785
rect 24905 1727 24955 1751
rect 25241 1785 25291 1809
rect 25241 1751 25249 1785
rect 25283 1751 25291 1785
rect 25241 1727 25291 1751
rect 25577 1785 25627 1809
rect 25577 1751 25585 1785
rect 25619 1751 25627 1785
rect 25577 1727 25627 1751
rect 25913 1785 25963 1809
rect 25913 1751 25921 1785
rect 25955 1751 25963 1785
rect 25913 1727 25963 1751
rect 26249 1785 26299 1809
rect 26249 1751 26257 1785
rect 26291 1751 26299 1785
rect 26249 1727 26299 1751
rect 26585 1785 26635 1809
rect 26585 1751 26593 1785
rect 26627 1751 26635 1785
rect 26585 1727 26635 1751
rect 26921 1785 26971 1809
rect 26921 1751 26929 1785
rect 26963 1751 26971 1785
rect 26921 1727 26971 1751
rect 27257 1785 27307 1809
rect 27257 1751 27265 1785
rect 27299 1751 27307 1785
rect 27257 1727 27307 1751
rect 27593 1785 27643 1809
rect 27593 1751 27601 1785
rect 27635 1751 27643 1785
rect 27593 1727 27643 1751
rect 27929 1785 27979 1809
rect 27929 1751 27937 1785
rect 27971 1751 27979 1785
rect 27929 1727 27979 1751
rect 28265 1785 28315 1809
rect 28265 1751 28273 1785
rect 28307 1751 28315 1785
rect 28265 1727 28315 1751
rect 28601 1785 28651 1809
rect 28601 1751 28609 1785
rect 28643 1751 28651 1785
rect 28601 1727 28651 1751
rect 28937 1785 28987 1809
rect 28937 1751 28945 1785
rect 28979 1751 28987 1785
rect 28937 1727 28987 1751
rect 29273 1785 29323 1809
rect 29273 1751 29281 1785
rect 29315 1751 29323 1785
rect 29273 1727 29323 1751
rect 29609 1785 29659 1809
rect 29609 1751 29617 1785
rect 29651 1751 29659 1785
rect 29609 1727 29659 1751
rect 29945 1785 29995 1809
rect 29945 1751 29953 1785
rect 29987 1751 29995 1785
rect 29945 1727 29995 1751
rect 30281 1785 30331 1809
rect 30281 1751 30289 1785
rect 30323 1751 30331 1785
rect 30281 1727 30331 1751
rect 30617 1785 30667 1809
rect 30617 1751 30625 1785
rect 30659 1751 30667 1785
rect 30617 1727 30667 1751
rect 30953 1785 31003 1809
rect 30953 1751 30961 1785
rect 30995 1751 31003 1785
rect 30953 1727 31003 1751
rect 31289 1785 31339 1809
rect 31289 1751 31297 1785
rect 31331 1751 31339 1785
rect 31289 1727 31339 1751
rect 31625 1785 31675 1809
rect 31625 1751 31633 1785
rect 31667 1751 31675 1785
rect 31625 1727 31675 1751
rect 31961 1785 32011 1809
rect 31961 1751 31969 1785
rect 32003 1751 32011 1785
rect 31961 1727 32011 1751
rect 32297 1785 32347 1809
rect 32297 1751 32305 1785
rect 32339 1751 32347 1785
rect 32297 1727 32347 1751
rect 32633 1785 32683 1809
rect 32633 1751 32641 1785
rect 32675 1751 32683 1785
rect 32633 1727 32683 1751
rect 32969 1785 33019 1809
rect 32969 1751 32977 1785
rect 33011 1751 33019 1785
rect 32969 1727 33019 1751
rect 33305 1785 33355 1809
rect 33305 1751 33313 1785
rect 33347 1751 33355 1785
rect 33305 1727 33355 1751
rect 33641 1785 33691 1809
rect 33641 1751 33649 1785
rect 33683 1751 33691 1785
rect 33641 1727 33691 1751
rect 33977 1785 34027 1809
rect 33977 1751 33985 1785
rect 34019 1751 34027 1785
rect 33977 1727 34027 1751
rect 34313 1785 34363 1809
rect 34313 1751 34321 1785
rect 34355 1751 34363 1785
rect 34313 1727 34363 1751
rect 34649 1785 34699 1809
rect 34649 1751 34657 1785
rect 34691 1751 34699 1785
rect 34649 1727 34699 1751
rect 34985 1785 35035 1809
rect 34985 1751 34993 1785
rect 35027 1751 35035 1785
rect 34985 1727 35035 1751
rect 35321 1785 35371 1809
rect 35321 1751 35329 1785
rect 35363 1751 35371 1785
rect 35321 1727 35371 1751
rect 35657 1785 35707 1809
rect 35657 1751 35665 1785
rect 35699 1751 35707 1785
rect 35657 1727 35707 1751
rect 35993 1785 36043 1809
rect 35993 1751 36001 1785
rect 36035 1751 36043 1785
rect 35993 1727 36043 1751
rect 36329 1785 36379 1809
rect 36329 1751 36337 1785
rect 36371 1751 36379 1785
rect 36329 1727 36379 1751
rect 36665 1785 36715 1809
rect 36665 1751 36673 1785
rect 36707 1751 36715 1785
rect 36665 1727 36715 1751
rect 37001 1785 37051 1809
rect 37001 1751 37009 1785
rect 37043 1751 37051 1785
rect 37001 1727 37051 1751
rect 37337 1785 37387 1809
rect 37337 1751 37345 1785
rect 37379 1751 37387 1785
rect 37337 1727 37387 1751
rect 37673 1785 37723 1809
rect 37673 1751 37681 1785
rect 37715 1751 37723 1785
rect 37673 1727 37723 1751
rect 38009 1785 38059 1809
rect 38009 1751 38017 1785
rect 38051 1751 38059 1785
rect 38009 1727 38059 1751
rect 38345 1785 38395 1809
rect 38345 1751 38353 1785
rect 38387 1751 38395 1785
rect 38345 1727 38395 1751
rect 38681 1785 38731 1809
rect 38681 1751 38689 1785
rect 38723 1751 38731 1785
rect 38681 1727 38731 1751
rect 39017 1785 39067 1809
rect 39017 1751 39025 1785
rect 39059 1751 39067 1785
rect 39017 1727 39067 1751
rect 39353 1785 39403 1809
rect 39353 1751 39361 1785
rect 39395 1751 39403 1785
rect 39353 1727 39403 1751
rect 39689 1785 39739 1809
rect 39689 1751 39697 1785
rect 39731 1751 39739 1785
rect 39689 1727 39739 1751
rect 40025 1785 40075 1809
rect 40025 1751 40033 1785
rect 40067 1751 40075 1785
rect 40025 1727 40075 1751
rect 40361 1785 40411 1809
rect 40361 1751 40369 1785
rect 40403 1751 40411 1785
rect 40361 1727 40411 1751
rect 40697 1785 40747 1809
rect 40697 1751 40705 1785
rect 40739 1751 40747 1785
rect 40697 1727 40747 1751
rect 41033 1785 41083 1809
rect 41033 1751 41041 1785
rect 41075 1751 41083 1785
rect 41033 1727 41083 1751
rect 41369 1785 41419 1809
rect 41369 1751 41377 1785
rect 41411 1751 41419 1785
rect 41369 1727 41419 1751
rect 41705 1785 41755 1809
rect 41705 1751 41713 1785
rect 41747 1751 41755 1785
rect 41705 1727 41755 1751
rect 42041 1785 42091 1809
rect 42041 1751 42049 1785
rect 42083 1751 42091 1785
rect 42041 1727 42091 1751
rect 42377 1785 42427 1809
rect 42377 1751 42385 1785
rect 42419 1751 42427 1785
rect 42377 1727 42427 1751
rect 42713 1785 42763 1809
rect 42713 1751 42721 1785
rect 42755 1751 42763 1785
rect 42713 1727 42763 1751
rect 43049 1785 43099 1809
rect 43049 1751 43057 1785
rect 43091 1751 43099 1785
rect 43049 1727 43099 1751
rect 43385 1785 43435 1809
rect 43385 1751 43393 1785
rect 43427 1751 43435 1785
rect 43385 1727 43435 1751
rect 43721 1785 43771 1809
rect 43721 1751 43729 1785
rect 43763 1751 43771 1785
rect 43721 1727 43771 1751
rect 44057 1785 44107 1809
rect 44057 1751 44065 1785
rect 44099 1751 44107 1785
rect 44057 1727 44107 1751
rect 44393 1785 44443 1809
rect 44393 1751 44401 1785
rect 44435 1751 44443 1785
rect 44393 1727 44443 1751
rect 44729 1785 44779 1809
rect 44729 1751 44737 1785
rect 44771 1751 44779 1785
rect 44729 1727 44779 1751
rect 45065 1785 45115 1809
rect 45065 1751 45073 1785
rect 45107 1751 45115 1785
rect 45065 1727 45115 1751
rect 45401 1785 45451 1809
rect 45401 1751 45409 1785
rect 45443 1751 45451 1785
rect 45401 1727 45451 1751
rect 45737 1785 45787 1809
rect 45737 1751 45745 1785
rect 45779 1751 45787 1785
rect 45737 1727 45787 1751
rect 46073 1785 46123 1809
rect 46073 1751 46081 1785
rect 46115 1751 46123 1785
rect 46073 1727 46123 1751
rect 46409 1785 46459 1809
rect 46409 1751 46417 1785
rect 46451 1751 46459 1785
rect 46409 1727 46459 1751
rect 46745 1785 46795 1809
rect 46745 1751 46753 1785
rect 46787 1751 46795 1785
rect 46745 1727 46795 1751
rect 47081 1785 47131 1809
rect 47081 1751 47089 1785
rect 47123 1751 47131 1785
rect 47081 1727 47131 1751
rect 47417 1785 47467 1809
rect 47417 1751 47425 1785
rect 47459 1751 47467 1785
rect 47417 1727 47467 1751
rect 47753 1785 47803 1809
rect 47753 1751 47761 1785
rect 47795 1751 47803 1785
rect 47753 1727 47803 1751
rect 48089 1785 48139 1809
rect 48089 1751 48097 1785
rect 48131 1751 48139 1785
rect 48089 1727 48139 1751
rect 48425 1785 48475 1809
rect 48425 1751 48433 1785
rect 48467 1751 48475 1785
rect 48425 1727 48475 1751
rect 48761 1785 48811 1809
rect 48761 1751 48769 1785
rect 48803 1751 48811 1785
rect 48761 1727 48811 1751
rect 49097 1785 49147 1809
rect 49097 1751 49105 1785
rect 49139 1751 49147 1785
rect 49097 1727 49147 1751
rect 49433 1785 49483 1809
rect 49433 1751 49441 1785
rect 49475 1751 49483 1785
rect 49433 1727 49483 1751
rect 49769 1785 49819 1809
rect 49769 1751 49777 1785
rect 49811 1751 49819 1785
rect 49769 1727 49819 1751
rect 50105 1785 50155 1809
rect 50105 1751 50113 1785
rect 50147 1751 50155 1785
rect 50105 1727 50155 1751
rect 50441 1785 50491 1809
rect 50441 1751 50449 1785
rect 50483 1751 50491 1785
rect 50441 1727 50491 1751
rect 50777 1785 50827 1809
rect 50777 1751 50785 1785
rect 50819 1751 50827 1785
rect 50777 1727 50827 1751
rect 51113 1785 51163 1809
rect 51113 1751 51121 1785
rect 51155 1751 51163 1785
rect 51113 1727 51163 1751
rect 51449 1785 51499 1809
rect 51449 1751 51457 1785
rect 51491 1751 51499 1785
rect 51449 1727 51499 1751
rect 51785 1785 51835 1809
rect 51785 1751 51793 1785
rect 51827 1751 51835 1785
rect 51785 1727 51835 1751
rect 52121 1785 52171 1809
rect 52121 1751 52129 1785
rect 52163 1751 52171 1785
rect 52121 1727 52171 1751
rect 52457 1785 52507 1809
rect 52457 1751 52465 1785
rect 52499 1751 52507 1785
rect 52457 1727 52507 1751
rect 52793 1785 52843 1809
rect 52793 1751 52801 1785
rect 52835 1751 52843 1785
rect 52793 1727 52843 1751
rect 53129 1785 53179 1809
rect 53129 1751 53137 1785
rect 53171 1751 53179 1785
rect 53129 1727 53179 1751
rect 53465 1785 53515 1809
rect 53465 1751 53473 1785
rect 53507 1751 53515 1785
rect 53465 1727 53515 1751
rect 53801 1785 53851 1809
rect 53801 1751 53809 1785
rect 53843 1751 53851 1785
rect 53801 1727 53851 1751
rect 54137 1785 54187 1809
rect 54137 1751 54145 1785
rect 54179 1751 54187 1785
rect 54137 1727 54187 1751
rect 54473 1785 54523 1809
rect 54473 1751 54481 1785
rect 54515 1751 54523 1785
rect 54473 1727 54523 1751
rect 54809 1785 54859 1809
rect 54809 1751 54817 1785
rect 54851 1751 54859 1785
rect 54809 1727 54859 1751
rect 55145 1785 55195 1809
rect 55145 1751 55153 1785
rect 55187 1751 55195 1785
rect 55145 1727 55195 1751
rect 55481 1785 55531 1809
rect 55481 1751 55489 1785
rect 55523 1751 55531 1785
rect 55481 1727 55531 1751
rect 55817 1785 55867 1809
rect 55817 1751 55825 1785
rect 55859 1751 55867 1785
rect 55817 1727 55867 1751
rect 56153 1785 56203 1809
rect 56153 1751 56161 1785
rect 56195 1751 56203 1785
rect 56153 1727 56203 1751
rect 56489 1785 56539 1809
rect 56489 1751 56497 1785
rect 56531 1751 56539 1785
rect 56489 1727 56539 1751
rect 56825 1785 56875 1809
rect 56825 1751 56833 1785
rect 56867 1751 56875 1785
rect 56825 1727 56875 1751
rect 57161 1785 57211 1809
rect 57161 1751 57169 1785
rect 57203 1751 57211 1785
rect 57161 1727 57211 1751
rect 57497 1785 57547 1809
rect 57497 1751 57505 1785
rect 57539 1751 57547 1785
rect 57497 1727 57547 1751
rect 57833 1785 57883 1809
rect 57833 1751 57841 1785
rect 57875 1751 57883 1785
rect 57833 1727 57883 1751
rect 58169 1785 58219 1809
rect 58169 1751 58177 1785
rect 58211 1751 58219 1785
rect 58169 1727 58219 1751
rect 58505 1785 58555 1809
rect 58505 1751 58513 1785
rect 58547 1751 58555 1785
rect 58505 1727 58555 1751
rect 58841 1785 58891 1809
rect 58841 1751 58849 1785
rect 58883 1751 58891 1785
rect 58841 1727 58891 1751
rect 59177 1785 59227 1809
rect 59177 1751 59185 1785
rect 59219 1751 59227 1785
rect 59177 1727 59227 1751
rect 59513 1785 59563 1809
rect 59513 1751 59521 1785
rect 59555 1751 59563 1785
rect 59513 1727 59563 1751
rect 59849 1785 59899 1809
rect 59849 1751 59857 1785
rect 59891 1751 59899 1785
rect 59849 1727 59899 1751
rect 60185 1785 60235 1809
rect 60185 1751 60193 1785
rect 60227 1751 60235 1785
rect 60185 1727 60235 1751
rect 60521 1785 60571 1809
rect 60521 1751 60529 1785
rect 60563 1751 60571 1785
rect 60521 1727 60571 1751
rect 60857 1785 60907 1809
rect 60857 1751 60865 1785
rect 60899 1751 60907 1785
rect 60857 1727 60907 1751
rect 61193 1785 61243 1809
rect 61193 1751 61201 1785
rect 61235 1751 61243 1785
rect 61193 1727 61243 1751
rect 61529 1785 61579 1809
rect 61529 1751 61537 1785
rect 61571 1751 61579 1785
rect 61529 1727 61579 1751
rect 61865 1785 61915 1809
rect 61865 1751 61873 1785
rect 61907 1751 61915 1785
rect 61865 1727 61915 1751
rect 62201 1785 62251 1809
rect 62201 1751 62209 1785
rect 62243 1751 62251 1785
rect 62201 1727 62251 1751
rect 62537 1785 62587 1809
rect 62537 1751 62545 1785
rect 62579 1751 62587 1785
rect 62537 1727 62587 1751
rect 62873 1785 62923 1809
rect 62873 1751 62881 1785
rect 62915 1751 62923 1785
rect 62873 1727 62923 1751
rect 63209 1785 63259 1809
rect 63209 1751 63217 1785
rect 63251 1751 63259 1785
rect 63209 1727 63259 1751
rect 63545 1785 63595 1809
rect 63545 1751 63553 1785
rect 63587 1751 63595 1785
rect 63545 1727 63595 1751
rect 63881 1785 63931 1809
rect 63881 1751 63889 1785
rect 63923 1751 63931 1785
rect 63881 1727 63931 1751
rect 64217 1785 64267 1809
rect 64217 1751 64225 1785
rect 64259 1751 64267 1785
rect 64217 1727 64267 1751
rect 64553 1785 64603 1809
rect 64553 1751 64561 1785
rect 64595 1751 64603 1785
rect 64553 1727 64603 1751
rect 64889 1785 64939 1809
rect 64889 1751 64897 1785
rect 64931 1751 64939 1785
rect 64889 1727 64939 1751
rect 65225 1785 65275 1809
rect 65225 1751 65233 1785
rect 65267 1751 65275 1785
rect 65225 1727 65275 1751
rect 65561 1785 65611 1809
rect 65561 1751 65569 1785
rect 65603 1751 65611 1785
rect 65561 1727 65611 1751
rect 65897 1785 65947 1809
rect 65897 1751 65905 1785
rect 65939 1751 65947 1785
rect 65897 1727 65947 1751
rect 66233 1785 66283 1809
rect 66233 1751 66241 1785
rect 66275 1751 66283 1785
rect 66233 1727 66283 1751
rect 66569 1785 66619 1809
rect 66569 1751 66577 1785
rect 66611 1751 66619 1785
rect 66569 1727 66619 1751
rect 66905 1785 66955 1809
rect 66905 1751 66913 1785
rect 66947 1751 66955 1785
rect 66905 1727 66955 1751
rect 67241 1785 67291 1809
rect 67241 1751 67249 1785
rect 67283 1751 67291 1785
rect 67241 1727 67291 1751
rect 67577 1785 67627 1809
rect 67577 1751 67585 1785
rect 67619 1751 67627 1785
rect 67577 1727 67627 1751
rect 67913 1785 67963 1809
rect 67913 1751 67921 1785
rect 67955 1751 67963 1785
rect 67913 1727 67963 1751
rect 68249 1785 68299 1809
rect 68249 1751 68257 1785
rect 68291 1751 68299 1785
rect 68249 1727 68299 1751
rect 68585 1785 68635 1809
rect 68585 1751 68593 1785
rect 68627 1751 68635 1785
rect 68585 1727 68635 1751
rect 68921 1785 68971 1809
rect 68921 1751 68929 1785
rect 68963 1751 68971 1785
rect 68921 1727 68971 1751
rect 69257 1785 69307 1809
rect 69257 1751 69265 1785
rect 69299 1751 69307 1785
rect 69257 1727 69307 1751
rect 69593 1785 69643 1809
rect 69593 1751 69601 1785
rect 69635 1751 69643 1785
rect 69593 1727 69643 1751
rect 69929 1785 69979 1809
rect 69929 1751 69937 1785
rect 69971 1751 69979 1785
rect 69929 1727 69979 1751
rect 70265 1785 70315 1809
rect 70265 1751 70273 1785
rect 70307 1751 70315 1785
rect 70265 1727 70315 1751
rect 70601 1785 70651 1809
rect 70601 1751 70609 1785
rect 70643 1751 70651 1785
rect 70601 1727 70651 1751
rect 70937 1785 70987 1809
rect 70937 1751 70945 1785
rect 70979 1751 70987 1785
rect 70937 1727 70987 1751
rect 71273 1785 71323 1809
rect 71273 1751 71281 1785
rect 71315 1751 71323 1785
rect 71273 1727 71323 1751
rect 71609 1785 71659 1809
rect 71609 1751 71617 1785
rect 71651 1751 71659 1785
rect 71609 1727 71659 1751
rect 71945 1785 71995 1809
rect 71945 1751 71953 1785
rect 71987 1751 71995 1785
rect 71945 1727 71995 1751
rect 72281 1785 72331 1809
rect 72281 1751 72289 1785
rect 72323 1751 72331 1785
rect 72281 1727 72331 1751
rect 72617 1785 72667 1809
rect 72617 1751 72625 1785
rect 72659 1751 72667 1785
rect 72617 1727 72667 1751
rect 72953 1785 73003 1809
rect 72953 1751 72961 1785
rect 72995 1751 73003 1785
rect 72953 1727 73003 1751
rect 73289 1785 73339 1809
rect 73289 1751 73297 1785
rect 73331 1751 73339 1785
rect 73289 1727 73339 1751
rect 73625 1785 73675 1809
rect 73625 1751 73633 1785
rect 73667 1751 73675 1785
rect 73625 1727 73675 1751
rect 73961 1785 74011 1809
rect 73961 1751 73969 1785
rect 74003 1751 74011 1785
rect 73961 1727 74011 1751
rect 74297 1785 74347 1809
rect 74297 1751 74305 1785
rect 74339 1751 74347 1785
rect 74297 1727 74347 1751
rect 74633 1785 74683 1809
rect 74633 1751 74641 1785
rect 74675 1751 74683 1785
rect 74633 1727 74683 1751
rect 74969 1785 75019 1809
rect 74969 1751 74977 1785
rect 75011 1751 75019 1785
rect 74969 1727 75019 1751
rect 75305 1785 75355 1809
rect 75305 1751 75313 1785
rect 75347 1751 75355 1785
rect 75305 1727 75355 1751
rect 75641 1785 75691 1809
rect 75641 1751 75649 1785
rect 75683 1751 75691 1785
rect 75641 1727 75691 1751
rect 75977 1785 76027 1809
rect 75977 1751 75985 1785
rect 76019 1751 76027 1785
rect 75977 1727 76027 1751
rect 76313 1785 76363 1809
rect 76313 1751 76321 1785
rect 76355 1751 76363 1785
rect 76313 1727 76363 1751
rect 76649 1785 76699 1809
rect 76649 1751 76657 1785
rect 76691 1751 76699 1785
rect 76649 1727 76699 1751
rect 76985 1785 77035 1809
rect 76985 1751 76993 1785
rect 77027 1751 77035 1785
rect 76985 1727 77035 1751
rect 77321 1785 77371 1809
rect 77321 1751 77329 1785
rect 77363 1751 77371 1785
rect 77321 1727 77371 1751
rect 77657 1785 77707 1809
rect 77657 1751 77665 1785
rect 77699 1751 77707 1785
rect 77657 1727 77707 1751
rect 77993 1785 78043 1809
rect 77993 1751 78001 1785
rect 78035 1751 78043 1785
rect 77993 1727 78043 1751
rect 78329 1785 78379 1809
rect 78329 1751 78337 1785
rect 78371 1751 78379 1785
rect 78329 1727 78379 1751
rect 78665 1785 78715 1809
rect 78665 1751 78673 1785
rect 78707 1751 78715 1785
rect 78665 1727 78715 1751
rect 79001 1785 79051 1809
rect 79001 1751 79009 1785
rect 79043 1751 79051 1785
rect 79001 1727 79051 1751
rect 79337 1785 79387 1809
rect 79337 1751 79345 1785
rect 79379 1751 79387 1785
rect 79337 1727 79387 1751
rect 79673 1785 79723 1809
rect 79673 1751 79681 1785
rect 79715 1751 79723 1785
rect 79673 1727 79723 1751
rect 80009 1785 80059 1809
rect 80009 1751 80017 1785
rect 80051 1751 80059 1785
rect 80009 1727 80059 1751
rect 80345 1785 80395 1809
rect 80345 1751 80353 1785
rect 80387 1751 80395 1785
rect 80345 1727 80395 1751
rect 80681 1785 80731 1809
rect 80681 1751 80689 1785
rect 80723 1751 80731 1785
rect 80681 1727 80731 1751
rect 81017 1785 81067 1809
rect 81017 1751 81025 1785
rect 81059 1751 81067 1785
rect 81017 1727 81067 1751
rect 81353 1785 81403 1809
rect 81353 1751 81361 1785
rect 81395 1751 81403 1785
rect 81353 1727 81403 1751
rect 81689 1785 81739 1809
rect 81689 1751 81697 1785
rect 81731 1751 81739 1785
rect 81689 1727 81739 1751
rect 82025 1785 82075 1809
rect 82025 1751 82033 1785
rect 82067 1751 82075 1785
rect 82025 1727 82075 1751
rect 82361 1785 82411 1809
rect 82361 1751 82369 1785
rect 82403 1751 82411 1785
rect 82361 1727 82411 1751
rect 82697 1785 82747 1809
rect 82697 1751 82705 1785
rect 82739 1751 82747 1785
rect 82697 1727 82747 1751
rect 83033 1785 83083 1809
rect 83033 1751 83041 1785
rect 83075 1751 83083 1785
rect 83033 1727 83083 1751
rect 83369 1785 83419 1809
rect 83369 1751 83377 1785
rect 83411 1751 83419 1785
rect 83369 1727 83419 1751
rect 83705 1785 83755 1809
rect 83705 1751 83713 1785
rect 83747 1751 83755 1785
rect 83705 1727 83755 1751
rect 84041 1785 84091 1809
rect 84041 1751 84049 1785
rect 84083 1751 84091 1785
rect 84041 1727 84091 1751
rect 84377 1785 84427 1809
rect 84377 1751 84385 1785
rect 84419 1751 84427 1785
rect 84377 1727 84427 1751
rect 84713 1785 84763 1809
rect 84713 1751 84721 1785
rect 84755 1751 84763 1785
rect 84713 1727 84763 1751
rect 85049 1785 85099 1809
rect 85049 1751 85057 1785
rect 85091 1751 85099 1785
rect 85049 1727 85099 1751
rect 85385 1785 85435 1809
rect 85385 1751 85393 1785
rect 85427 1751 85435 1785
rect 85385 1727 85435 1751
rect 85721 1785 85771 1809
rect 85721 1751 85729 1785
rect 85763 1751 85771 1785
rect 85721 1727 85771 1751
rect 86057 1785 86107 1809
rect 86057 1751 86065 1785
rect 86099 1751 86107 1785
rect 86057 1727 86107 1751
rect 86393 1785 86443 1809
rect 86393 1751 86401 1785
rect 86435 1751 86443 1785
rect 86393 1727 86443 1751
rect 86729 1785 86779 1809
rect 86729 1751 86737 1785
rect 86771 1751 86779 1785
rect 86729 1727 86779 1751
rect 87065 1785 87115 1809
rect 87065 1751 87073 1785
rect 87107 1751 87115 1785
rect 87065 1727 87115 1751
rect 87401 1785 87451 1809
rect 87401 1751 87409 1785
rect 87443 1751 87451 1785
rect 87401 1727 87451 1751
rect 87737 1785 87787 1809
rect 87737 1751 87745 1785
rect 87779 1751 87787 1785
rect 87737 1727 87787 1751
rect 88073 1785 88123 1809
rect 88073 1751 88081 1785
rect 88115 1751 88123 1785
rect 88073 1727 88123 1751
rect 88409 1785 88459 1809
rect 88409 1751 88417 1785
rect 88451 1751 88459 1785
rect 88409 1727 88459 1751
rect 88745 1785 88795 1809
rect 88745 1751 88753 1785
rect 88787 1751 88795 1785
rect 88745 1727 88795 1751
<< nsubdiffcont >>
rect 2065 87479 2099 87513
rect 2401 87479 2435 87513
rect 2737 87479 2771 87513
rect 3073 87479 3107 87513
rect 3409 87479 3443 87513
rect 3745 87479 3779 87513
rect 4081 87479 4115 87513
rect 4417 87479 4451 87513
rect 4753 87479 4787 87513
rect 5089 87479 5123 87513
rect 5425 87479 5459 87513
rect 5761 87479 5795 87513
rect 6097 87479 6131 87513
rect 6433 87479 6467 87513
rect 6769 87479 6803 87513
rect 7105 87479 7139 87513
rect 7441 87479 7475 87513
rect 7777 87479 7811 87513
rect 8113 87479 8147 87513
rect 8449 87479 8483 87513
rect 8785 87479 8819 87513
rect 9121 87479 9155 87513
rect 9457 87479 9491 87513
rect 9793 87479 9827 87513
rect 10129 87479 10163 87513
rect 10465 87479 10499 87513
rect 10801 87479 10835 87513
rect 11137 87479 11171 87513
rect 11473 87479 11507 87513
rect 11809 87479 11843 87513
rect 12145 87479 12179 87513
rect 12481 87479 12515 87513
rect 12817 87479 12851 87513
rect 13153 87479 13187 87513
rect 13489 87479 13523 87513
rect 13825 87479 13859 87513
rect 14161 87479 14195 87513
rect 14497 87479 14531 87513
rect 14833 87479 14867 87513
rect 15169 87479 15203 87513
rect 15505 87479 15539 87513
rect 15841 87479 15875 87513
rect 16177 87479 16211 87513
rect 16513 87479 16547 87513
rect 16849 87479 16883 87513
rect 17185 87479 17219 87513
rect 17521 87479 17555 87513
rect 17857 87479 17891 87513
rect 18193 87479 18227 87513
rect 18529 87479 18563 87513
rect 18865 87479 18899 87513
rect 19201 87479 19235 87513
rect 19537 87479 19571 87513
rect 19873 87479 19907 87513
rect 20209 87479 20243 87513
rect 20545 87479 20579 87513
rect 20881 87479 20915 87513
rect 21217 87479 21251 87513
rect 21553 87479 21587 87513
rect 21889 87479 21923 87513
rect 22225 87479 22259 87513
rect 22561 87479 22595 87513
rect 22897 87479 22931 87513
rect 23233 87479 23267 87513
rect 23569 87479 23603 87513
rect 23905 87479 23939 87513
rect 24241 87479 24275 87513
rect 24577 87479 24611 87513
rect 24913 87479 24947 87513
rect 25249 87479 25283 87513
rect 25585 87479 25619 87513
rect 25921 87479 25955 87513
rect 26257 87479 26291 87513
rect 26593 87479 26627 87513
rect 26929 87479 26963 87513
rect 27265 87479 27299 87513
rect 27601 87479 27635 87513
rect 27937 87479 27971 87513
rect 28273 87479 28307 87513
rect 28609 87479 28643 87513
rect 28945 87479 28979 87513
rect 29281 87479 29315 87513
rect 29617 87479 29651 87513
rect 29953 87479 29987 87513
rect 30289 87479 30323 87513
rect 30625 87479 30659 87513
rect 30961 87479 30995 87513
rect 31297 87479 31331 87513
rect 31633 87479 31667 87513
rect 31969 87479 32003 87513
rect 32305 87479 32339 87513
rect 32641 87479 32675 87513
rect 32977 87479 33011 87513
rect 33313 87479 33347 87513
rect 33649 87479 33683 87513
rect 33985 87479 34019 87513
rect 34321 87479 34355 87513
rect 34657 87479 34691 87513
rect 34993 87479 35027 87513
rect 35329 87479 35363 87513
rect 35665 87479 35699 87513
rect 36001 87479 36035 87513
rect 36337 87479 36371 87513
rect 36673 87479 36707 87513
rect 37009 87479 37043 87513
rect 37345 87479 37379 87513
rect 37681 87479 37715 87513
rect 38017 87479 38051 87513
rect 38353 87479 38387 87513
rect 38689 87479 38723 87513
rect 39025 87479 39059 87513
rect 39361 87479 39395 87513
rect 39697 87479 39731 87513
rect 40033 87479 40067 87513
rect 40369 87479 40403 87513
rect 40705 87479 40739 87513
rect 41041 87479 41075 87513
rect 41377 87479 41411 87513
rect 41713 87479 41747 87513
rect 42049 87479 42083 87513
rect 42385 87479 42419 87513
rect 42721 87479 42755 87513
rect 43057 87479 43091 87513
rect 43393 87479 43427 87513
rect 43729 87479 43763 87513
rect 44065 87479 44099 87513
rect 44401 87479 44435 87513
rect 44737 87479 44771 87513
rect 45073 87479 45107 87513
rect 45409 87479 45443 87513
rect 45745 87479 45779 87513
rect 46081 87479 46115 87513
rect 46417 87479 46451 87513
rect 46753 87479 46787 87513
rect 47089 87479 47123 87513
rect 47425 87479 47459 87513
rect 47761 87479 47795 87513
rect 48097 87479 48131 87513
rect 48433 87479 48467 87513
rect 48769 87479 48803 87513
rect 49105 87479 49139 87513
rect 49441 87479 49475 87513
rect 49777 87479 49811 87513
rect 50113 87479 50147 87513
rect 50449 87479 50483 87513
rect 50785 87479 50819 87513
rect 51121 87479 51155 87513
rect 51457 87479 51491 87513
rect 51793 87479 51827 87513
rect 52129 87479 52163 87513
rect 52465 87479 52499 87513
rect 52801 87479 52835 87513
rect 53137 87479 53171 87513
rect 53473 87479 53507 87513
rect 53809 87479 53843 87513
rect 54145 87479 54179 87513
rect 54481 87479 54515 87513
rect 54817 87479 54851 87513
rect 55153 87479 55187 87513
rect 55489 87479 55523 87513
rect 55825 87479 55859 87513
rect 56161 87479 56195 87513
rect 56497 87479 56531 87513
rect 56833 87479 56867 87513
rect 57169 87479 57203 87513
rect 57505 87479 57539 87513
rect 57841 87479 57875 87513
rect 58177 87479 58211 87513
rect 58513 87479 58547 87513
rect 58849 87479 58883 87513
rect 59185 87479 59219 87513
rect 59521 87479 59555 87513
rect 59857 87479 59891 87513
rect 60193 87479 60227 87513
rect 60529 87479 60563 87513
rect 60865 87479 60899 87513
rect 61201 87479 61235 87513
rect 61537 87479 61571 87513
rect 61873 87479 61907 87513
rect 62209 87479 62243 87513
rect 62545 87479 62579 87513
rect 62881 87479 62915 87513
rect 63217 87479 63251 87513
rect 63553 87479 63587 87513
rect 63889 87479 63923 87513
rect 64225 87479 64259 87513
rect 64561 87479 64595 87513
rect 64897 87479 64931 87513
rect 65233 87479 65267 87513
rect 65569 87479 65603 87513
rect 65905 87479 65939 87513
rect 66241 87479 66275 87513
rect 66577 87479 66611 87513
rect 66913 87479 66947 87513
rect 67249 87479 67283 87513
rect 67585 87479 67619 87513
rect 67921 87479 67955 87513
rect 68257 87479 68291 87513
rect 68593 87479 68627 87513
rect 68929 87479 68963 87513
rect 69265 87479 69299 87513
rect 69601 87479 69635 87513
rect 69937 87479 69971 87513
rect 70273 87479 70307 87513
rect 70609 87479 70643 87513
rect 70945 87479 70979 87513
rect 71281 87479 71315 87513
rect 71617 87479 71651 87513
rect 71953 87479 71987 87513
rect 72289 87479 72323 87513
rect 72625 87479 72659 87513
rect 72961 87479 72995 87513
rect 73297 87479 73331 87513
rect 73633 87479 73667 87513
rect 73969 87479 74003 87513
rect 74305 87479 74339 87513
rect 74641 87479 74675 87513
rect 74977 87479 75011 87513
rect 75313 87479 75347 87513
rect 75649 87479 75683 87513
rect 75985 87479 76019 87513
rect 76321 87479 76355 87513
rect 76657 87479 76691 87513
rect 76993 87479 77027 87513
rect 77329 87479 77363 87513
rect 77665 87479 77699 87513
rect 78001 87479 78035 87513
rect 78337 87479 78371 87513
rect 78673 87479 78707 87513
rect 79009 87479 79043 87513
rect 79345 87479 79379 87513
rect 79681 87479 79715 87513
rect 80017 87479 80051 87513
rect 80353 87479 80387 87513
rect 80689 87479 80723 87513
rect 81025 87479 81059 87513
rect 81361 87479 81395 87513
rect 81697 87479 81731 87513
rect 82033 87479 82067 87513
rect 82369 87479 82403 87513
rect 82705 87479 82739 87513
rect 83041 87479 83075 87513
rect 83377 87479 83411 87513
rect 83713 87479 83747 87513
rect 84049 87479 84083 87513
rect 84385 87479 84419 87513
rect 84721 87479 84755 87513
rect 85057 87479 85091 87513
rect 85393 87479 85427 87513
rect 85729 87479 85763 87513
rect 86065 87479 86099 87513
rect 86401 87479 86435 87513
rect 86737 87479 86771 87513
rect 87073 87479 87107 87513
rect 87409 87479 87443 87513
rect 87745 87479 87779 87513
rect 88081 87479 88115 87513
rect 88417 87479 88451 87513
rect 88753 87479 88787 87513
rect 1729 87095 1763 87129
rect 89227 87095 89261 87129
rect 1729 86759 1763 86793
rect 89227 86759 89261 86793
rect 1729 86423 1763 86457
rect 89227 86423 89261 86457
rect 1729 86087 1763 86121
rect 89227 86087 89261 86121
rect 1729 85751 1763 85785
rect 89227 85751 89261 85785
rect 1729 85415 1763 85449
rect 89227 85415 89261 85449
rect 1729 85079 1763 85113
rect 89227 85079 89261 85113
rect 1729 84743 1763 84777
rect 89227 84743 89261 84777
rect 1729 84407 1763 84441
rect 89227 84407 89261 84441
rect 1729 84071 1763 84105
rect 89227 84071 89261 84105
rect 1729 83735 1763 83769
rect 89227 83735 89261 83769
rect 1729 83399 1763 83433
rect 89227 83399 89261 83433
rect 1729 83063 1763 83097
rect 89227 83063 89261 83097
rect 1729 82727 1763 82761
rect 89227 82727 89261 82761
rect 1729 82391 1763 82425
rect 89227 82391 89261 82425
rect 1729 82055 1763 82089
rect 89227 82055 89261 82089
rect 1729 81719 1763 81753
rect 89227 81719 89261 81753
rect 1729 81383 1763 81417
rect 89227 81383 89261 81417
rect 1729 81047 1763 81081
rect 89227 81047 89261 81081
rect 1729 80711 1763 80745
rect 89227 80711 89261 80745
rect 1729 80375 1763 80409
rect 89227 80375 89261 80409
rect 1729 80039 1763 80073
rect 89227 80039 89261 80073
rect 1729 79703 1763 79737
rect 89227 79703 89261 79737
rect 1729 79367 1763 79401
rect 89227 79367 89261 79401
rect 1729 79031 1763 79065
rect 89227 79031 89261 79065
rect 1729 78695 1763 78729
rect 89227 78695 89261 78729
rect 1729 78359 1763 78393
rect 89227 78359 89261 78393
rect 1729 78023 1763 78057
rect 89227 78023 89261 78057
rect 1729 77687 1763 77721
rect 89227 77687 89261 77721
rect 1729 77351 1763 77385
rect 89227 77351 89261 77385
rect 1729 77015 1763 77049
rect 89227 77015 89261 77049
rect 1729 76679 1763 76713
rect 89227 76679 89261 76713
rect 1729 76343 1763 76377
rect 89227 76343 89261 76377
rect 1729 76007 1763 76041
rect 89227 76007 89261 76041
rect 1729 75671 1763 75705
rect 89227 75671 89261 75705
rect 1729 75335 1763 75369
rect 89227 75335 89261 75369
rect 1729 74999 1763 75033
rect 89227 74999 89261 75033
rect 1729 74663 1763 74697
rect 89227 74663 89261 74697
rect 1729 74327 1763 74361
rect 89227 74327 89261 74361
rect 1729 73991 1763 74025
rect 89227 73991 89261 74025
rect 1729 73655 1763 73689
rect 89227 73655 89261 73689
rect 1729 73319 1763 73353
rect 89227 73319 89261 73353
rect 1729 72983 1763 73017
rect 89227 72983 89261 73017
rect 1729 72647 1763 72681
rect 89227 72647 89261 72681
rect 1729 72311 1763 72345
rect 89227 72311 89261 72345
rect 1729 71975 1763 72009
rect 89227 71975 89261 72009
rect 1729 71639 1763 71673
rect 89227 71639 89261 71673
rect 1729 71303 1763 71337
rect 89227 71303 89261 71337
rect 1729 70967 1763 71001
rect 89227 70967 89261 71001
rect 1729 70631 1763 70665
rect 89227 70631 89261 70665
rect 1729 70295 1763 70329
rect 89227 70295 89261 70329
rect 1729 69959 1763 69993
rect 89227 69959 89261 69993
rect 1729 69623 1763 69657
rect 89227 69623 89261 69657
rect 1729 69287 1763 69321
rect 89227 69287 89261 69321
rect 1729 68951 1763 68985
rect 89227 68951 89261 68985
rect 1729 68615 1763 68649
rect 89227 68615 89261 68649
rect 1729 68279 1763 68313
rect 89227 68279 89261 68313
rect 1729 67943 1763 67977
rect 89227 67943 89261 67977
rect 1729 67607 1763 67641
rect 89227 67607 89261 67641
rect 1729 67271 1763 67305
rect 89227 67271 89261 67305
rect 1729 66935 1763 66969
rect 89227 66935 89261 66969
rect 1729 66599 1763 66633
rect 89227 66599 89261 66633
rect 1729 66263 1763 66297
rect 89227 66263 89261 66297
rect 1729 65927 1763 65961
rect 89227 65927 89261 65961
rect 1729 65591 1763 65625
rect 89227 65591 89261 65625
rect 1729 65255 1763 65289
rect 89227 65255 89261 65289
rect 1729 64919 1763 64953
rect 89227 64919 89261 64953
rect 1729 64583 1763 64617
rect 89227 64583 89261 64617
rect 1729 64247 1763 64281
rect 89227 64247 89261 64281
rect 1729 63911 1763 63945
rect 89227 63911 89261 63945
rect 1729 63575 1763 63609
rect 89227 63575 89261 63609
rect 1729 63239 1763 63273
rect 89227 63239 89261 63273
rect 1729 62903 1763 62937
rect 89227 62903 89261 62937
rect 1729 62567 1763 62601
rect 89227 62567 89261 62601
rect 1729 62231 1763 62265
rect 89227 62231 89261 62265
rect 1729 61895 1763 61929
rect 89227 61895 89261 61929
rect 1729 61559 1763 61593
rect 89227 61559 89261 61593
rect 1729 61223 1763 61257
rect 89227 61223 89261 61257
rect 1729 60887 1763 60921
rect 89227 60887 89261 60921
rect 1729 60551 1763 60585
rect 89227 60551 89261 60585
rect 1729 60215 1763 60249
rect 89227 60215 89261 60249
rect 1729 59879 1763 59913
rect 89227 59879 89261 59913
rect 1729 59543 1763 59577
rect 89227 59543 89261 59577
rect 1729 59207 1763 59241
rect 89227 59207 89261 59241
rect 1729 58871 1763 58905
rect 89227 58871 89261 58905
rect 1729 58535 1763 58569
rect 89227 58535 89261 58569
rect 1729 58199 1763 58233
rect 89227 58199 89261 58233
rect 1729 57863 1763 57897
rect 89227 57863 89261 57897
rect 1729 57527 1763 57561
rect 89227 57527 89261 57561
rect 1729 57191 1763 57225
rect 89227 57191 89261 57225
rect 1729 56855 1763 56889
rect 89227 56855 89261 56889
rect 1729 56519 1763 56553
rect 89227 56519 89261 56553
rect 1729 56183 1763 56217
rect 89227 56183 89261 56217
rect 1729 55847 1763 55881
rect 89227 55847 89261 55881
rect 1729 55511 1763 55545
rect 89227 55511 89261 55545
rect 1729 55175 1763 55209
rect 89227 55175 89261 55209
rect 1729 54839 1763 54873
rect 89227 54839 89261 54873
rect 1729 54503 1763 54537
rect 89227 54503 89261 54537
rect 1729 54167 1763 54201
rect 89227 54167 89261 54201
rect 1729 53831 1763 53865
rect 89227 53831 89261 53865
rect 1729 53495 1763 53529
rect 89227 53495 89261 53529
rect 1729 53159 1763 53193
rect 89227 53159 89261 53193
rect 1729 52823 1763 52857
rect 89227 52823 89261 52857
rect 1729 52487 1763 52521
rect 89227 52487 89261 52521
rect 1729 52151 1763 52185
rect 89227 52151 89261 52185
rect 1729 51815 1763 51849
rect 89227 51815 89261 51849
rect 1729 51479 1763 51513
rect 89227 51479 89261 51513
rect 1729 51143 1763 51177
rect 89227 51143 89261 51177
rect 1729 50807 1763 50841
rect 89227 50807 89261 50841
rect 1729 50471 1763 50505
rect 89227 50471 89261 50505
rect 1729 50135 1763 50169
rect 89227 50135 89261 50169
rect 1729 49799 1763 49833
rect 89227 49799 89261 49833
rect 1729 49463 1763 49497
rect 89227 49463 89261 49497
rect 1729 49127 1763 49161
rect 89227 49127 89261 49161
rect 1729 48791 1763 48825
rect 89227 48791 89261 48825
rect 1729 48455 1763 48489
rect 89227 48455 89261 48489
rect 1729 48119 1763 48153
rect 89227 48119 89261 48153
rect 1729 47783 1763 47817
rect 89227 47783 89261 47817
rect 1729 47447 1763 47481
rect 89227 47447 89261 47481
rect 1729 47111 1763 47145
rect 89227 47111 89261 47145
rect 1729 46775 1763 46809
rect 89227 46775 89261 46809
rect 1729 46439 1763 46473
rect 89227 46439 89261 46473
rect 1729 46103 1763 46137
rect 89227 46103 89261 46137
rect 1729 45767 1763 45801
rect 89227 45767 89261 45801
rect 1729 45431 1763 45465
rect 89227 45431 89261 45465
rect 1729 45095 1763 45129
rect 89227 45095 89261 45129
rect 1729 44759 1763 44793
rect 89227 44759 89261 44793
rect 1729 44423 1763 44457
rect 89227 44423 89261 44457
rect 1729 44087 1763 44121
rect 89227 44087 89261 44121
rect 1729 43751 1763 43785
rect 89227 43751 89261 43785
rect 1729 43415 1763 43449
rect 89227 43415 89261 43449
rect 1729 43079 1763 43113
rect 89227 43079 89261 43113
rect 1729 42743 1763 42777
rect 89227 42743 89261 42777
rect 1729 42407 1763 42441
rect 89227 42407 89261 42441
rect 1729 42071 1763 42105
rect 89227 42071 89261 42105
rect 1729 41735 1763 41769
rect 89227 41735 89261 41769
rect 1729 41399 1763 41433
rect 89227 41399 89261 41433
rect 1729 41063 1763 41097
rect 89227 41063 89261 41097
rect 1729 40727 1763 40761
rect 89227 40727 89261 40761
rect 1729 40391 1763 40425
rect 89227 40391 89261 40425
rect 1729 40055 1763 40089
rect 89227 40055 89261 40089
rect 1729 39719 1763 39753
rect 89227 39719 89261 39753
rect 1729 39383 1763 39417
rect 89227 39383 89261 39417
rect 1729 39047 1763 39081
rect 89227 39047 89261 39081
rect 1729 38711 1763 38745
rect 89227 38711 89261 38745
rect 1729 38375 1763 38409
rect 89227 38375 89261 38409
rect 1729 38039 1763 38073
rect 89227 38039 89261 38073
rect 1729 37703 1763 37737
rect 89227 37703 89261 37737
rect 1729 37367 1763 37401
rect 89227 37367 89261 37401
rect 1729 37031 1763 37065
rect 89227 37031 89261 37065
rect 1729 36695 1763 36729
rect 89227 36695 89261 36729
rect 1729 36359 1763 36393
rect 89227 36359 89261 36393
rect 1729 36023 1763 36057
rect 89227 36023 89261 36057
rect 1729 35687 1763 35721
rect 89227 35687 89261 35721
rect 1729 35351 1763 35385
rect 89227 35351 89261 35385
rect 1729 35015 1763 35049
rect 89227 35015 89261 35049
rect 1729 34679 1763 34713
rect 89227 34679 89261 34713
rect 1729 34343 1763 34377
rect 89227 34343 89261 34377
rect 1729 34007 1763 34041
rect 89227 34007 89261 34041
rect 1729 33671 1763 33705
rect 89227 33671 89261 33705
rect 1729 33335 1763 33369
rect 89227 33335 89261 33369
rect 1729 32999 1763 33033
rect 89227 32999 89261 33033
rect 1729 32663 1763 32697
rect 89227 32663 89261 32697
rect 1729 32327 1763 32361
rect 89227 32327 89261 32361
rect 1729 31991 1763 32025
rect 89227 31991 89261 32025
rect 1729 31655 1763 31689
rect 89227 31655 89261 31689
rect 1729 31319 1763 31353
rect 89227 31319 89261 31353
rect 1729 30983 1763 31017
rect 89227 30983 89261 31017
rect 1729 30647 1763 30681
rect 89227 30647 89261 30681
rect 1729 30311 1763 30345
rect 89227 30311 89261 30345
rect 1729 29975 1763 30009
rect 89227 29975 89261 30009
rect 1729 29639 1763 29673
rect 89227 29639 89261 29673
rect 1729 29303 1763 29337
rect 89227 29303 89261 29337
rect 1729 28967 1763 29001
rect 89227 28967 89261 29001
rect 1729 28631 1763 28665
rect 89227 28631 89261 28665
rect 1729 28295 1763 28329
rect 89227 28295 89261 28329
rect 1729 27959 1763 27993
rect 89227 27959 89261 27993
rect 1729 27623 1763 27657
rect 89227 27623 89261 27657
rect 1729 27287 1763 27321
rect 89227 27287 89261 27321
rect 1729 26951 1763 26985
rect 89227 26951 89261 26985
rect 1729 26615 1763 26649
rect 89227 26615 89261 26649
rect 1729 26279 1763 26313
rect 89227 26279 89261 26313
rect 1729 25943 1763 25977
rect 89227 25943 89261 25977
rect 1729 25607 1763 25641
rect 89227 25607 89261 25641
rect 1729 25271 1763 25305
rect 89227 25271 89261 25305
rect 1729 24935 1763 24969
rect 89227 24935 89261 24969
rect 1729 24599 1763 24633
rect 89227 24599 89261 24633
rect 1729 24263 1763 24297
rect 89227 24263 89261 24297
rect 1729 23927 1763 23961
rect 89227 23927 89261 23961
rect 1729 23591 1763 23625
rect 89227 23591 89261 23625
rect 1729 23255 1763 23289
rect 89227 23255 89261 23289
rect 1729 22919 1763 22953
rect 89227 22919 89261 22953
rect 1729 22583 1763 22617
rect 89227 22583 89261 22617
rect 1729 22247 1763 22281
rect 89227 22247 89261 22281
rect 1729 21911 1763 21945
rect 89227 21911 89261 21945
rect 1729 21575 1763 21609
rect 89227 21575 89261 21609
rect 1729 21239 1763 21273
rect 89227 21239 89261 21273
rect 1729 20903 1763 20937
rect 89227 20903 89261 20937
rect 1729 20567 1763 20601
rect 89227 20567 89261 20601
rect 1729 20231 1763 20265
rect 89227 20231 89261 20265
rect 1729 19895 1763 19929
rect 89227 19895 89261 19929
rect 1729 19559 1763 19593
rect 89227 19559 89261 19593
rect 1729 19223 1763 19257
rect 89227 19223 89261 19257
rect 1729 18887 1763 18921
rect 89227 18887 89261 18921
rect 1729 18551 1763 18585
rect 89227 18551 89261 18585
rect 1729 18215 1763 18249
rect 89227 18215 89261 18249
rect 1729 17879 1763 17913
rect 89227 17879 89261 17913
rect 1729 17543 1763 17577
rect 89227 17543 89261 17577
rect 1729 17207 1763 17241
rect 89227 17207 89261 17241
rect 1729 16871 1763 16905
rect 89227 16871 89261 16905
rect 1729 16535 1763 16569
rect 89227 16535 89261 16569
rect 1729 16199 1763 16233
rect 89227 16199 89261 16233
rect 1729 15863 1763 15897
rect 89227 15863 89261 15897
rect 1729 15527 1763 15561
rect 89227 15527 89261 15561
rect 1729 15191 1763 15225
rect 89227 15191 89261 15225
rect 1729 14855 1763 14889
rect 89227 14855 89261 14889
rect 1729 14519 1763 14553
rect 89227 14519 89261 14553
rect 1729 14183 1763 14217
rect 89227 14183 89261 14217
rect 1729 13847 1763 13881
rect 89227 13847 89261 13881
rect 1729 13511 1763 13545
rect 89227 13511 89261 13545
rect 1729 13175 1763 13209
rect 89227 13175 89261 13209
rect 1729 12839 1763 12873
rect 89227 12839 89261 12873
rect 1729 12503 1763 12537
rect 89227 12503 89261 12537
rect 1729 12167 1763 12201
rect 89227 12167 89261 12201
rect 1729 11831 1763 11865
rect 89227 11831 89261 11865
rect 1729 11495 1763 11529
rect 89227 11495 89261 11529
rect 1729 11159 1763 11193
rect 89227 11159 89261 11193
rect 1729 10823 1763 10857
rect 89227 10823 89261 10857
rect 1729 10487 1763 10521
rect 89227 10487 89261 10521
rect 1729 10151 1763 10185
rect 89227 10151 89261 10185
rect 1729 9815 1763 9849
rect 89227 9815 89261 9849
rect 1729 9479 1763 9513
rect 89227 9479 89261 9513
rect 1729 9143 1763 9177
rect 89227 9143 89261 9177
rect 1729 8807 1763 8841
rect 89227 8807 89261 8841
rect 1729 8471 1763 8505
rect 89227 8471 89261 8505
rect 1729 8135 1763 8169
rect 89227 8135 89261 8169
rect 1729 7799 1763 7833
rect 89227 7799 89261 7833
rect 1729 7463 1763 7497
rect 89227 7463 89261 7497
rect 1729 7127 1763 7161
rect 89227 7127 89261 7161
rect 1729 6791 1763 6825
rect 89227 6791 89261 6825
rect 1729 6455 1763 6489
rect 89227 6455 89261 6489
rect 1729 6119 1763 6153
rect 89227 6119 89261 6153
rect 1729 5783 1763 5817
rect 89227 5783 89261 5817
rect 1729 5447 1763 5481
rect 89227 5447 89261 5481
rect 1729 5111 1763 5145
rect 89227 5111 89261 5145
rect 1729 4775 1763 4809
rect 89227 4775 89261 4809
rect 1729 4439 1763 4473
rect 89227 4439 89261 4473
rect 1729 4103 1763 4137
rect 89227 4103 89261 4137
rect 1729 3767 1763 3801
rect 89227 3767 89261 3801
rect 1729 3431 1763 3465
rect 89227 3431 89261 3465
rect 1729 3095 1763 3129
rect 89227 3095 89261 3129
rect 1729 2759 1763 2793
rect 89227 2759 89261 2793
rect 1729 2423 1763 2457
rect 89227 2423 89261 2457
rect 1729 2087 1763 2121
rect 89227 2087 89261 2121
rect 2065 1751 2099 1785
rect 2401 1751 2435 1785
rect 2737 1751 2771 1785
rect 3073 1751 3107 1785
rect 3409 1751 3443 1785
rect 3745 1751 3779 1785
rect 4081 1751 4115 1785
rect 4417 1751 4451 1785
rect 4753 1751 4787 1785
rect 5089 1751 5123 1785
rect 5425 1751 5459 1785
rect 5761 1751 5795 1785
rect 6097 1751 6131 1785
rect 6433 1751 6467 1785
rect 6769 1751 6803 1785
rect 7105 1751 7139 1785
rect 7441 1751 7475 1785
rect 7777 1751 7811 1785
rect 8113 1751 8147 1785
rect 8449 1751 8483 1785
rect 8785 1751 8819 1785
rect 9121 1751 9155 1785
rect 9457 1751 9491 1785
rect 9793 1751 9827 1785
rect 10129 1751 10163 1785
rect 10465 1751 10499 1785
rect 10801 1751 10835 1785
rect 11137 1751 11171 1785
rect 11473 1751 11507 1785
rect 11809 1751 11843 1785
rect 12145 1751 12179 1785
rect 12481 1751 12515 1785
rect 12817 1751 12851 1785
rect 13153 1751 13187 1785
rect 13489 1751 13523 1785
rect 13825 1751 13859 1785
rect 14161 1751 14195 1785
rect 14497 1751 14531 1785
rect 14833 1751 14867 1785
rect 15169 1751 15203 1785
rect 15505 1751 15539 1785
rect 15841 1751 15875 1785
rect 16177 1751 16211 1785
rect 16513 1751 16547 1785
rect 16849 1751 16883 1785
rect 17185 1751 17219 1785
rect 17521 1751 17555 1785
rect 17857 1751 17891 1785
rect 18193 1751 18227 1785
rect 18529 1751 18563 1785
rect 18865 1751 18899 1785
rect 19201 1751 19235 1785
rect 19537 1751 19571 1785
rect 19873 1751 19907 1785
rect 20209 1751 20243 1785
rect 20545 1751 20579 1785
rect 20881 1751 20915 1785
rect 21217 1751 21251 1785
rect 21553 1751 21587 1785
rect 21889 1751 21923 1785
rect 22225 1751 22259 1785
rect 22561 1751 22595 1785
rect 22897 1751 22931 1785
rect 23233 1751 23267 1785
rect 23569 1751 23603 1785
rect 23905 1751 23939 1785
rect 24241 1751 24275 1785
rect 24577 1751 24611 1785
rect 24913 1751 24947 1785
rect 25249 1751 25283 1785
rect 25585 1751 25619 1785
rect 25921 1751 25955 1785
rect 26257 1751 26291 1785
rect 26593 1751 26627 1785
rect 26929 1751 26963 1785
rect 27265 1751 27299 1785
rect 27601 1751 27635 1785
rect 27937 1751 27971 1785
rect 28273 1751 28307 1785
rect 28609 1751 28643 1785
rect 28945 1751 28979 1785
rect 29281 1751 29315 1785
rect 29617 1751 29651 1785
rect 29953 1751 29987 1785
rect 30289 1751 30323 1785
rect 30625 1751 30659 1785
rect 30961 1751 30995 1785
rect 31297 1751 31331 1785
rect 31633 1751 31667 1785
rect 31969 1751 32003 1785
rect 32305 1751 32339 1785
rect 32641 1751 32675 1785
rect 32977 1751 33011 1785
rect 33313 1751 33347 1785
rect 33649 1751 33683 1785
rect 33985 1751 34019 1785
rect 34321 1751 34355 1785
rect 34657 1751 34691 1785
rect 34993 1751 35027 1785
rect 35329 1751 35363 1785
rect 35665 1751 35699 1785
rect 36001 1751 36035 1785
rect 36337 1751 36371 1785
rect 36673 1751 36707 1785
rect 37009 1751 37043 1785
rect 37345 1751 37379 1785
rect 37681 1751 37715 1785
rect 38017 1751 38051 1785
rect 38353 1751 38387 1785
rect 38689 1751 38723 1785
rect 39025 1751 39059 1785
rect 39361 1751 39395 1785
rect 39697 1751 39731 1785
rect 40033 1751 40067 1785
rect 40369 1751 40403 1785
rect 40705 1751 40739 1785
rect 41041 1751 41075 1785
rect 41377 1751 41411 1785
rect 41713 1751 41747 1785
rect 42049 1751 42083 1785
rect 42385 1751 42419 1785
rect 42721 1751 42755 1785
rect 43057 1751 43091 1785
rect 43393 1751 43427 1785
rect 43729 1751 43763 1785
rect 44065 1751 44099 1785
rect 44401 1751 44435 1785
rect 44737 1751 44771 1785
rect 45073 1751 45107 1785
rect 45409 1751 45443 1785
rect 45745 1751 45779 1785
rect 46081 1751 46115 1785
rect 46417 1751 46451 1785
rect 46753 1751 46787 1785
rect 47089 1751 47123 1785
rect 47425 1751 47459 1785
rect 47761 1751 47795 1785
rect 48097 1751 48131 1785
rect 48433 1751 48467 1785
rect 48769 1751 48803 1785
rect 49105 1751 49139 1785
rect 49441 1751 49475 1785
rect 49777 1751 49811 1785
rect 50113 1751 50147 1785
rect 50449 1751 50483 1785
rect 50785 1751 50819 1785
rect 51121 1751 51155 1785
rect 51457 1751 51491 1785
rect 51793 1751 51827 1785
rect 52129 1751 52163 1785
rect 52465 1751 52499 1785
rect 52801 1751 52835 1785
rect 53137 1751 53171 1785
rect 53473 1751 53507 1785
rect 53809 1751 53843 1785
rect 54145 1751 54179 1785
rect 54481 1751 54515 1785
rect 54817 1751 54851 1785
rect 55153 1751 55187 1785
rect 55489 1751 55523 1785
rect 55825 1751 55859 1785
rect 56161 1751 56195 1785
rect 56497 1751 56531 1785
rect 56833 1751 56867 1785
rect 57169 1751 57203 1785
rect 57505 1751 57539 1785
rect 57841 1751 57875 1785
rect 58177 1751 58211 1785
rect 58513 1751 58547 1785
rect 58849 1751 58883 1785
rect 59185 1751 59219 1785
rect 59521 1751 59555 1785
rect 59857 1751 59891 1785
rect 60193 1751 60227 1785
rect 60529 1751 60563 1785
rect 60865 1751 60899 1785
rect 61201 1751 61235 1785
rect 61537 1751 61571 1785
rect 61873 1751 61907 1785
rect 62209 1751 62243 1785
rect 62545 1751 62579 1785
rect 62881 1751 62915 1785
rect 63217 1751 63251 1785
rect 63553 1751 63587 1785
rect 63889 1751 63923 1785
rect 64225 1751 64259 1785
rect 64561 1751 64595 1785
rect 64897 1751 64931 1785
rect 65233 1751 65267 1785
rect 65569 1751 65603 1785
rect 65905 1751 65939 1785
rect 66241 1751 66275 1785
rect 66577 1751 66611 1785
rect 66913 1751 66947 1785
rect 67249 1751 67283 1785
rect 67585 1751 67619 1785
rect 67921 1751 67955 1785
rect 68257 1751 68291 1785
rect 68593 1751 68627 1785
rect 68929 1751 68963 1785
rect 69265 1751 69299 1785
rect 69601 1751 69635 1785
rect 69937 1751 69971 1785
rect 70273 1751 70307 1785
rect 70609 1751 70643 1785
rect 70945 1751 70979 1785
rect 71281 1751 71315 1785
rect 71617 1751 71651 1785
rect 71953 1751 71987 1785
rect 72289 1751 72323 1785
rect 72625 1751 72659 1785
rect 72961 1751 72995 1785
rect 73297 1751 73331 1785
rect 73633 1751 73667 1785
rect 73969 1751 74003 1785
rect 74305 1751 74339 1785
rect 74641 1751 74675 1785
rect 74977 1751 75011 1785
rect 75313 1751 75347 1785
rect 75649 1751 75683 1785
rect 75985 1751 76019 1785
rect 76321 1751 76355 1785
rect 76657 1751 76691 1785
rect 76993 1751 77027 1785
rect 77329 1751 77363 1785
rect 77665 1751 77699 1785
rect 78001 1751 78035 1785
rect 78337 1751 78371 1785
rect 78673 1751 78707 1785
rect 79009 1751 79043 1785
rect 79345 1751 79379 1785
rect 79681 1751 79715 1785
rect 80017 1751 80051 1785
rect 80353 1751 80387 1785
rect 80689 1751 80723 1785
rect 81025 1751 81059 1785
rect 81361 1751 81395 1785
rect 81697 1751 81731 1785
rect 82033 1751 82067 1785
rect 82369 1751 82403 1785
rect 82705 1751 82739 1785
rect 83041 1751 83075 1785
rect 83377 1751 83411 1785
rect 83713 1751 83747 1785
rect 84049 1751 84083 1785
rect 84385 1751 84419 1785
rect 84721 1751 84755 1785
rect 85057 1751 85091 1785
rect 85393 1751 85427 1785
rect 85729 1751 85763 1785
rect 86065 1751 86099 1785
rect 86401 1751 86435 1785
rect 86737 1751 86771 1785
rect 87073 1751 87107 1785
rect 87409 1751 87443 1785
rect 87745 1751 87779 1785
rect 88081 1751 88115 1785
rect 88417 1751 88451 1785
rect 88753 1751 88787 1785
<< locali >>
rect 2065 87513 2099 87529
rect 2065 87463 2099 87479
rect 2401 87513 2435 87529
rect 2401 87463 2435 87479
rect 2737 87513 2771 87529
rect 2737 87463 2771 87479
rect 3073 87513 3107 87529
rect 3073 87463 3107 87479
rect 3409 87513 3443 87529
rect 3409 87463 3443 87479
rect 3745 87513 3779 87529
rect 3745 87463 3779 87479
rect 4081 87513 4115 87529
rect 4081 87463 4115 87479
rect 4417 87513 4451 87529
rect 4417 87463 4451 87479
rect 4753 87513 4787 87529
rect 4753 87463 4787 87479
rect 5089 87513 5123 87529
rect 5089 87463 5123 87479
rect 5425 87513 5459 87529
rect 5425 87463 5459 87479
rect 5761 87513 5795 87529
rect 5761 87463 5795 87479
rect 6097 87513 6131 87529
rect 6097 87463 6131 87479
rect 6433 87513 6467 87529
rect 6433 87463 6467 87479
rect 6769 87513 6803 87529
rect 6769 87463 6803 87479
rect 7105 87513 7139 87529
rect 7105 87463 7139 87479
rect 7441 87513 7475 87529
rect 7441 87463 7475 87479
rect 7777 87513 7811 87529
rect 7777 87463 7811 87479
rect 8113 87513 8147 87529
rect 8113 87463 8147 87479
rect 8449 87513 8483 87529
rect 8449 87463 8483 87479
rect 8785 87513 8819 87529
rect 8785 87463 8819 87479
rect 9121 87513 9155 87529
rect 9121 87463 9155 87479
rect 9457 87513 9491 87529
rect 9457 87463 9491 87479
rect 9793 87513 9827 87529
rect 9793 87463 9827 87479
rect 10129 87513 10163 87529
rect 10129 87463 10163 87479
rect 10465 87513 10499 87529
rect 10465 87463 10499 87479
rect 10801 87513 10835 87529
rect 10801 87463 10835 87479
rect 11137 87513 11171 87529
rect 11137 87463 11171 87479
rect 11473 87513 11507 87529
rect 11473 87463 11507 87479
rect 11809 87513 11843 87529
rect 11809 87463 11843 87479
rect 12145 87513 12179 87529
rect 12145 87463 12179 87479
rect 12481 87513 12515 87529
rect 12481 87463 12515 87479
rect 12817 87513 12851 87529
rect 12817 87463 12851 87479
rect 13153 87513 13187 87529
rect 13153 87463 13187 87479
rect 13489 87513 13523 87529
rect 13489 87463 13523 87479
rect 13825 87513 13859 87529
rect 13825 87463 13859 87479
rect 14161 87513 14195 87529
rect 14161 87463 14195 87479
rect 14497 87513 14531 87529
rect 14497 87463 14531 87479
rect 14833 87513 14867 87529
rect 14833 87463 14867 87479
rect 15169 87513 15203 87529
rect 15169 87463 15203 87479
rect 15505 87513 15539 87529
rect 15505 87463 15539 87479
rect 15841 87513 15875 87529
rect 15841 87463 15875 87479
rect 16177 87513 16211 87529
rect 16177 87463 16211 87479
rect 16513 87513 16547 87529
rect 16513 87463 16547 87479
rect 16849 87513 16883 87529
rect 16849 87463 16883 87479
rect 17185 87513 17219 87529
rect 17185 87463 17219 87479
rect 17521 87513 17555 87529
rect 17521 87463 17555 87479
rect 17857 87513 17891 87529
rect 17857 87463 17891 87479
rect 18193 87513 18227 87529
rect 18193 87463 18227 87479
rect 18529 87513 18563 87529
rect 18529 87463 18563 87479
rect 18865 87513 18899 87529
rect 18865 87463 18899 87479
rect 19201 87513 19235 87529
rect 19201 87463 19235 87479
rect 19537 87513 19571 87529
rect 19537 87463 19571 87479
rect 19873 87513 19907 87529
rect 19873 87463 19907 87479
rect 20209 87513 20243 87529
rect 20209 87463 20243 87479
rect 20545 87513 20579 87529
rect 20545 87463 20579 87479
rect 20881 87513 20915 87529
rect 20881 87463 20915 87479
rect 21217 87513 21251 87529
rect 21217 87463 21251 87479
rect 21553 87513 21587 87529
rect 21553 87463 21587 87479
rect 21889 87513 21923 87529
rect 21889 87463 21923 87479
rect 22225 87513 22259 87529
rect 22225 87463 22259 87479
rect 22561 87513 22595 87529
rect 22561 87463 22595 87479
rect 22897 87513 22931 87529
rect 22897 87463 22931 87479
rect 23233 87513 23267 87529
rect 23233 87463 23267 87479
rect 23569 87513 23603 87529
rect 23569 87463 23603 87479
rect 23905 87513 23939 87529
rect 23905 87463 23939 87479
rect 24241 87513 24275 87529
rect 24241 87463 24275 87479
rect 24577 87513 24611 87529
rect 24577 87463 24611 87479
rect 24913 87513 24947 87529
rect 24913 87463 24947 87479
rect 25249 87513 25283 87529
rect 25249 87463 25283 87479
rect 25585 87513 25619 87529
rect 25585 87463 25619 87479
rect 25921 87513 25955 87529
rect 25921 87463 25955 87479
rect 26257 87513 26291 87529
rect 26257 87463 26291 87479
rect 26593 87513 26627 87529
rect 26593 87463 26627 87479
rect 26929 87513 26963 87529
rect 26929 87463 26963 87479
rect 27265 87513 27299 87529
rect 27265 87463 27299 87479
rect 27601 87513 27635 87529
rect 27601 87463 27635 87479
rect 27937 87513 27971 87529
rect 27937 87463 27971 87479
rect 28273 87513 28307 87529
rect 28273 87463 28307 87479
rect 28609 87513 28643 87529
rect 28609 87463 28643 87479
rect 28945 87513 28979 87529
rect 28945 87463 28979 87479
rect 29281 87513 29315 87529
rect 29281 87463 29315 87479
rect 29617 87513 29651 87529
rect 29617 87463 29651 87479
rect 29953 87513 29987 87529
rect 29953 87463 29987 87479
rect 30289 87513 30323 87529
rect 30289 87463 30323 87479
rect 30625 87513 30659 87529
rect 30625 87463 30659 87479
rect 30961 87513 30995 87529
rect 30961 87463 30995 87479
rect 31297 87513 31331 87529
rect 31297 87463 31331 87479
rect 31633 87513 31667 87529
rect 31633 87463 31667 87479
rect 31969 87513 32003 87529
rect 31969 87463 32003 87479
rect 32305 87513 32339 87529
rect 32305 87463 32339 87479
rect 32641 87513 32675 87529
rect 32641 87463 32675 87479
rect 32977 87513 33011 87529
rect 32977 87463 33011 87479
rect 33313 87513 33347 87529
rect 33313 87463 33347 87479
rect 33649 87513 33683 87529
rect 33649 87463 33683 87479
rect 33985 87513 34019 87529
rect 33985 87463 34019 87479
rect 34321 87513 34355 87529
rect 34321 87463 34355 87479
rect 34657 87513 34691 87529
rect 34657 87463 34691 87479
rect 34993 87513 35027 87529
rect 34993 87463 35027 87479
rect 35329 87513 35363 87529
rect 35329 87463 35363 87479
rect 35665 87513 35699 87529
rect 35665 87463 35699 87479
rect 36001 87513 36035 87529
rect 36001 87463 36035 87479
rect 36337 87513 36371 87529
rect 36337 87463 36371 87479
rect 36673 87513 36707 87529
rect 36673 87463 36707 87479
rect 37009 87513 37043 87529
rect 37009 87463 37043 87479
rect 37345 87513 37379 87529
rect 37345 87463 37379 87479
rect 37681 87513 37715 87529
rect 37681 87463 37715 87479
rect 38017 87513 38051 87529
rect 38017 87463 38051 87479
rect 38353 87513 38387 87529
rect 38353 87463 38387 87479
rect 38689 87513 38723 87529
rect 38689 87463 38723 87479
rect 39025 87513 39059 87529
rect 39025 87463 39059 87479
rect 39361 87513 39395 87529
rect 39361 87463 39395 87479
rect 39697 87513 39731 87529
rect 39697 87463 39731 87479
rect 40033 87513 40067 87529
rect 40033 87463 40067 87479
rect 40369 87513 40403 87529
rect 40369 87463 40403 87479
rect 40705 87513 40739 87529
rect 40705 87463 40739 87479
rect 41041 87513 41075 87529
rect 41041 87463 41075 87479
rect 41377 87513 41411 87529
rect 41377 87463 41411 87479
rect 41713 87513 41747 87529
rect 41713 87463 41747 87479
rect 42049 87513 42083 87529
rect 42049 87463 42083 87479
rect 42385 87513 42419 87529
rect 42385 87463 42419 87479
rect 42721 87513 42755 87529
rect 42721 87463 42755 87479
rect 43057 87513 43091 87529
rect 43057 87463 43091 87479
rect 43393 87513 43427 87529
rect 43393 87463 43427 87479
rect 43729 87513 43763 87529
rect 43729 87463 43763 87479
rect 44065 87513 44099 87529
rect 44065 87463 44099 87479
rect 44401 87513 44435 87529
rect 44401 87463 44435 87479
rect 44737 87513 44771 87529
rect 44737 87463 44771 87479
rect 45073 87513 45107 87529
rect 45073 87463 45107 87479
rect 45409 87513 45443 87529
rect 45409 87463 45443 87479
rect 45745 87513 45779 87529
rect 45745 87463 45779 87479
rect 46081 87513 46115 87529
rect 46081 87463 46115 87479
rect 46417 87513 46451 87529
rect 46417 87463 46451 87479
rect 46753 87513 46787 87529
rect 46753 87463 46787 87479
rect 47089 87513 47123 87529
rect 47089 87463 47123 87479
rect 47425 87513 47459 87529
rect 47425 87463 47459 87479
rect 47761 87513 47795 87529
rect 47761 87463 47795 87479
rect 48097 87513 48131 87529
rect 48097 87463 48131 87479
rect 48433 87513 48467 87529
rect 48433 87463 48467 87479
rect 48769 87513 48803 87529
rect 48769 87463 48803 87479
rect 49105 87513 49139 87529
rect 49105 87463 49139 87479
rect 49441 87513 49475 87529
rect 49441 87463 49475 87479
rect 49777 87513 49811 87529
rect 49777 87463 49811 87479
rect 50113 87513 50147 87529
rect 50113 87463 50147 87479
rect 50449 87513 50483 87529
rect 50449 87463 50483 87479
rect 50785 87513 50819 87529
rect 50785 87463 50819 87479
rect 51121 87513 51155 87529
rect 51121 87463 51155 87479
rect 51457 87513 51491 87529
rect 51457 87463 51491 87479
rect 51793 87513 51827 87529
rect 51793 87463 51827 87479
rect 52129 87513 52163 87529
rect 52129 87463 52163 87479
rect 52465 87513 52499 87529
rect 52465 87463 52499 87479
rect 52801 87513 52835 87529
rect 52801 87463 52835 87479
rect 53137 87513 53171 87529
rect 53137 87463 53171 87479
rect 53473 87513 53507 87529
rect 53473 87463 53507 87479
rect 53809 87513 53843 87529
rect 53809 87463 53843 87479
rect 54145 87513 54179 87529
rect 54145 87463 54179 87479
rect 54481 87513 54515 87529
rect 54481 87463 54515 87479
rect 54817 87513 54851 87529
rect 54817 87463 54851 87479
rect 55153 87513 55187 87529
rect 55153 87463 55187 87479
rect 55489 87513 55523 87529
rect 55489 87463 55523 87479
rect 55825 87513 55859 87529
rect 55825 87463 55859 87479
rect 56161 87513 56195 87529
rect 56161 87463 56195 87479
rect 56497 87513 56531 87529
rect 56497 87463 56531 87479
rect 56833 87513 56867 87529
rect 56833 87463 56867 87479
rect 57169 87513 57203 87529
rect 57169 87463 57203 87479
rect 57505 87513 57539 87529
rect 57505 87463 57539 87479
rect 57841 87513 57875 87529
rect 57841 87463 57875 87479
rect 58177 87513 58211 87529
rect 58177 87463 58211 87479
rect 58513 87513 58547 87529
rect 58513 87463 58547 87479
rect 58849 87513 58883 87529
rect 58849 87463 58883 87479
rect 59185 87513 59219 87529
rect 59185 87463 59219 87479
rect 59521 87513 59555 87529
rect 59521 87463 59555 87479
rect 59857 87513 59891 87529
rect 59857 87463 59891 87479
rect 60193 87513 60227 87529
rect 60193 87463 60227 87479
rect 60529 87513 60563 87529
rect 60529 87463 60563 87479
rect 60865 87513 60899 87529
rect 60865 87463 60899 87479
rect 61201 87513 61235 87529
rect 61201 87463 61235 87479
rect 61537 87513 61571 87529
rect 61537 87463 61571 87479
rect 61873 87513 61907 87529
rect 61873 87463 61907 87479
rect 62209 87513 62243 87529
rect 62209 87463 62243 87479
rect 62545 87513 62579 87529
rect 62545 87463 62579 87479
rect 62881 87513 62915 87529
rect 62881 87463 62915 87479
rect 63217 87513 63251 87529
rect 63217 87463 63251 87479
rect 63553 87513 63587 87529
rect 63553 87463 63587 87479
rect 63889 87513 63923 87529
rect 63889 87463 63923 87479
rect 64225 87513 64259 87529
rect 64225 87463 64259 87479
rect 64561 87513 64595 87529
rect 64561 87463 64595 87479
rect 64897 87513 64931 87529
rect 64897 87463 64931 87479
rect 65233 87513 65267 87529
rect 65233 87463 65267 87479
rect 65569 87513 65603 87529
rect 65569 87463 65603 87479
rect 65905 87513 65939 87529
rect 65905 87463 65939 87479
rect 66241 87513 66275 87529
rect 66241 87463 66275 87479
rect 66577 87513 66611 87529
rect 66577 87463 66611 87479
rect 66913 87513 66947 87529
rect 66913 87463 66947 87479
rect 67249 87513 67283 87529
rect 67249 87463 67283 87479
rect 67585 87513 67619 87529
rect 67585 87463 67619 87479
rect 67921 87513 67955 87529
rect 67921 87463 67955 87479
rect 68257 87513 68291 87529
rect 68257 87463 68291 87479
rect 68593 87513 68627 87529
rect 68593 87463 68627 87479
rect 68929 87513 68963 87529
rect 68929 87463 68963 87479
rect 69265 87513 69299 87529
rect 69265 87463 69299 87479
rect 69601 87513 69635 87529
rect 69601 87463 69635 87479
rect 69937 87513 69971 87529
rect 69937 87463 69971 87479
rect 70273 87513 70307 87529
rect 70273 87463 70307 87479
rect 70609 87513 70643 87529
rect 70609 87463 70643 87479
rect 70945 87513 70979 87529
rect 70945 87463 70979 87479
rect 71281 87513 71315 87529
rect 71281 87463 71315 87479
rect 71617 87513 71651 87529
rect 71617 87463 71651 87479
rect 71953 87513 71987 87529
rect 71953 87463 71987 87479
rect 72289 87513 72323 87529
rect 72289 87463 72323 87479
rect 72625 87513 72659 87529
rect 72625 87463 72659 87479
rect 72961 87513 72995 87529
rect 72961 87463 72995 87479
rect 73297 87513 73331 87529
rect 73297 87463 73331 87479
rect 73633 87513 73667 87529
rect 73633 87463 73667 87479
rect 73969 87513 74003 87529
rect 73969 87463 74003 87479
rect 74305 87513 74339 87529
rect 74305 87463 74339 87479
rect 74641 87513 74675 87529
rect 74641 87463 74675 87479
rect 74977 87513 75011 87529
rect 74977 87463 75011 87479
rect 75313 87513 75347 87529
rect 75313 87463 75347 87479
rect 75649 87513 75683 87529
rect 75649 87463 75683 87479
rect 75985 87513 76019 87529
rect 75985 87463 76019 87479
rect 76321 87513 76355 87529
rect 76321 87463 76355 87479
rect 76657 87513 76691 87529
rect 76657 87463 76691 87479
rect 76993 87513 77027 87529
rect 76993 87463 77027 87479
rect 77329 87513 77363 87529
rect 77329 87463 77363 87479
rect 77665 87513 77699 87529
rect 77665 87463 77699 87479
rect 78001 87513 78035 87529
rect 78001 87463 78035 87479
rect 78337 87513 78371 87529
rect 78337 87463 78371 87479
rect 78673 87513 78707 87529
rect 78673 87463 78707 87479
rect 79009 87513 79043 87529
rect 79009 87463 79043 87479
rect 79345 87513 79379 87529
rect 79345 87463 79379 87479
rect 79681 87513 79715 87529
rect 79681 87463 79715 87479
rect 80017 87513 80051 87529
rect 80017 87463 80051 87479
rect 80353 87513 80387 87529
rect 80353 87463 80387 87479
rect 80689 87513 80723 87529
rect 80689 87463 80723 87479
rect 81025 87513 81059 87529
rect 81025 87463 81059 87479
rect 81361 87513 81395 87529
rect 81361 87463 81395 87479
rect 81697 87513 81731 87529
rect 81697 87463 81731 87479
rect 82033 87513 82067 87529
rect 82033 87463 82067 87479
rect 82369 87513 82403 87529
rect 82369 87463 82403 87479
rect 82705 87513 82739 87529
rect 82705 87463 82739 87479
rect 83041 87513 83075 87529
rect 83041 87463 83075 87479
rect 83377 87513 83411 87529
rect 83377 87463 83411 87479
rect 83713 87513 83747 87529
rect 83713 87463 83747 87479
rect 84049 87513 84083 87529
rect 84049 87463 84083 87479
rect 84385 87513 84419 87529
rect 84385 87463 84419 87479
rect 84721 87513 84755 87529
rect 84721 87463 84755 87479
rect 85057 87513 85091 87529
rect 85057 87463 85091 87479
rect 85393 87513 85427 87529
rect 85393 87463 85427 87479
rect 85729 87513 85763 87529
rect 85729 87463 85763 87479
rect 86065 87513 86099 87529
rect 86065 87463 86099 87479
rect 86401 87513 86435 87529
rect 86401 87463 86435 87479
rect 86737 87513 86771 87529
rect 86737 87463 86771 87479
rect 87073 87513 87107 87529
rect 87073 87463 87107 87479
rect 87409 87513 87443 87529
rect 87409 87463 87443 87479
rect 87745 87513 87779 87529
rect 87745 87463 87779 87479
rect 88081 87513 88115 87529
rect 88081 87463 88115 87479
rect 88417 87513 88451 87529
rect 88417 87463 88451 87479
rect 88753 87513 88787 87529
rect 88753 87463 88787 87479
rect 1729 87129 1763 87145
rect 1729 87079 1763 87095
rect 89227 87129 89261 87145
rect 89227 87079 89261 87095
rect 1729 86793 1763 86809
rect 1729 86743 1763 86759
rect 89227 86793 89261 86809
rect 89227 86743 89261 86759
rect 1729 86457 1763 86473
rect 1729 86407 1763 86423
rect 89227 86457 89261 86473
rect 89227 86407 89261 86423
rect 1729 86121 1763 86137
rect 1729 86071 1763 86087
rect 89227 86121 89261 86137
rect 89227 86071 89261 86087
rect 1729 85785 1763 85801
rect 1729 85735 1763 85751
rect 89227 85785 89261 85801
rect 89227 85735 89261 85751
rect 1729 85449 1763 85465
rect 1729 85399 1763 85415
rect 89227 85449 89261 85465
rect 89227 85399 89261 85415
rect 1729 85113 1763 85129
rect 1729 85063 1763 85079
rect 89227 85113 89261 85129
rect 89227 85063 89261 85079
rect 1729 84777 1763 84793
rect 1729 84727 1763 84743
rect 89227 84777 89261 84793
rect 89227 84727 89261 84743
rect 1729 84441 1763 84457
rect 1729 84391 1763 84407
rect 89227 84441 89261 84457
rect 89227 84391 89261 84407
rect 1729 84105 1763 84121
rect 1729 84055 1763 84071
rect 89227 84105 89261 84121
rect 89227 84055 89261 84071
rect 1729 83769 1763 83785
rect 1729 83719 1763 83735
rect 89227 83769 89261 83785
rect 89227 83719 89261 83735
rect 1729 83433 1763 83449
rect 1729 83383 1763 83399
rect 89227 83433 89261 83449
rect 89227 83383 89261 83399
rect 1729 83097 1763 83113
rect 1729 83047 1763 83063
rect 89227 83097 89261 83113
rect 89227 83047 89261 83063
rect 1729 82761 1763 82777
rect 1729 82711 1763 82727
rect 89227 82761 89261 82777
rect 89227 82711 89261 82727
rect 1729 82425 1763 82441
rect 1729 82375 1763 82391
rect 89227 82425 89261 82441
rect 89227 82375 89261 82391
rect 1729 82089 1763 82105
rect 1729 82039 1763 82055
rect 89227 82089 89261 82105
rect 89227 82039 89261 82055
rect 1729 81753 1763 81769
rect 1729 81703 1763 81719
rect 89227 81753 89261 81769
rect 89227 81703 89261 81719
rect 1729 81417 1763 81433
rect 1729 81367 1763 81383
rect 89227 81417 89261 81433
rect 89227 81367 89261 81383
rect 1729 81081 1763 81097
rect 1729 81031 1763 81047
rect 89227 81081 89261 81097
rect 89227 81031 89261 81047
rect 1729 80745 1763 80761
rect 1729 80695 1763 80711
rect 89227 80745 89261 80761
rect 89227 80695 89261 80711
rect 1729 80409 1763 80425
rect 1729 80359 1763 80375
rect 89227 80409 89261 80425
rect 89227 80359 89261 80375
rect 1729 80073 1763 80089
rect 1729 80023 1763 80039
rect 89227 80073 89261 80089
rect 89227 80023 89261 80039
rect 1729 79737 1763 79753
rect 1729 79687 1763 79703
rect 89227 79737 89261 79753
rect 89227 79687 89261 79703
rect 1729 79401 1763 79417
rect 1729 79351 1763 79367
rect 89227 79401 89261 79417
rect 89227 79351 89261 79367
rect 1729 79065 1763 79081
rect 1729 79015 1763 79031
rect 89227 79065 89261 79081
rect 89227 79015 89261 79031
rect 1729 78729 1763 78745
rect 1729 78679 1763 78695
rect 89227 78729 89261 78745
rect 89227 78679 89261 78695
rect 1729 78393 1763 78409
rect 1729 78343 1763 78359
rect 89227 78393 89261 78409
rect 89227 78343 89261 78359
rect 1729 78057 1763 78073
rect 1729 78007 1763 78023
rect 89227 78057 89261 78073
rect 89227 78007 89261 78023
rect 1729 77721 1763 77737
rect 1729 77671 1763 77687
rect 89227 77721 89261 77737
rect 89227 77671 89261 77687
rect 1729 77385 1763 77401
rect 1729 77335 1763 77351
rect 89227 77385 89261 77401
rect 89227 77335 89261 77351
rect 1729 77049 1763 77065
rect 1729 76999 1763 77015
rect 89227 77049 89261 77065
rect 89227 76999 89261 77015
rect 1729 76713 1763 76729
rect 1729 76663 1763 76679
rect 89227 76713 89261 76729
rect 89227 76663 89261 76679
rect 1729 76377 1763 76393
rect 1729 76327 1763 76343
rect 89227 76377 89261 76393
rect 89227 76327 89261 76343
rect 1729 76041 1763 76057
rect 1729 75991 1763 76007
rect 89227 76041 89261 76057
rect 89227 75991 89261 76007
rect 1729 75705 1763 75721
rect 1729 75655 1763 75671
rect 89227 75705 89261 75721
rect 89227 75655 89261 75671
rect 1729 75369 1763 75385
rect 1729 75319 1763 75335
rect 89227 75369 89261 75385
rect 89227 75319 89261 75335
rect 1729 75033 1763 75049
rect 1729 74983 1763 74999
rect 89227 75033 89261 75049
rect 89227 74983 89261 74999
rect 1729 74697 1763 74713
rect 1729 74647 1763 74663
rect 89227 74697 89261 74713
rect 89227 74647 89261 74663
rect 1729 74361 1763 74377
rect 1729 74311 1763 74327
rect 89227 74361 89261 74377
rect 89227 74311 89261 74327
rect 1729 74025 1763 74041
rect 1729 73975 1763 73991
rect 89227 74025 89261 74041
rect 89227 73975 89261 73991
rect 1729 73689 1763 73705
rect 1729 73639 1763 73655
rect 89227 73689 89261 73705
rect 89227 73639 89261 73655
rect 1729 73353 1763 73369
rect 1729 73303 1763 73319
rect 89227 73353 89261 73369
rect 89227 73303 89261 73319
rect 1729 73017 1763 73033
rect 1729 72967 1763 72983
rect 89227 73017 89261 73033
rect 89227 72967 89261 72983
rect 1729 72681 1763 72697
rect 1729 72631 1763 72647
rect 89227 72681 89261 72697
rect 89227 72631 89261 72647
rect 1729 72345 1763 72361
rect 1729 72295 1763 72311
rect 89227 72345 89261 72361
rect 89227 72295 89261 72311
rect 1729 72009 1763 72025
rect 1729 71959 1763 71975
rect 89227 72009 89261 72025
rect 89227 71959 89261 71975
rect 1729 71673 1763 71689
rect 1729 71623 1763 71639
rect 89227 71673 89261 71689
rect 89227 71623 89261 71639
rect 1729 71337 1763 71353
rect 1729 71287 1763 71303
rect 89227 71337 89261 71353
rect 89227 71287 89261 71303
rect 1729 71001 1763 71017
rect 1729 70951 1763 70967
rect 89227 71001 89261 71017
rect 89227 70951 89261 70967
rect 1729 70665 1763 70681
rect 1729 70615 1763 70631
rect 89227 70665 89261 70681
rect 89227 70615 89261 70631
rect 1729 70329 1763 70345
rect 1729 70279 1763 70295
rect 89227 70329 89261 70345
rect 89227 70279 89261 70295
rect 1729 69993 1763 70009
rect 1729 69943 1763 69959
rect 89227 69993 89261 70009
rect 89227 69943 89261 69959
rect 1729 69657 1763 69673
rect 1729 69607 1763 69623
rect 89227 69657 89261 69673
rect 89227 69607 89261 69623
rect 1729 69321 1763 69337
rect 1729 69271 1763 69287
rect 89227 69321 89261 69337
rect 89227 69271 89261 69287
rect 1729 68985 1763 69001
rect 1729 68935 1763 68951
rect 89227 68985 89261 69001
rect 89227 68935 89261 68951
rect 1729 68649 1763 68665
rect 1729 68599 1763 68615
rect 89227 68649 89261 68665
rect 89227 68599 89261 68615
rect 1729 68313 1763 68329
rect 1729 68263 1763 68279
rect 89227 68313 89261 68329
rect 89227 68263 89261 68279
rect 1729 67977 1763 67993
rect 1729 67927 1763 67943
rect 89227 67977 89261 67993
rect 89227 67927 89261 67943
rect 1729 67641 1763 67657
rect 1729 67591 1763 67607
rect 89227 67641 89261 67657
rect 89227 67591 89261 67607
rect 1729 67305 1763 67321
rect 1729 67255 1763 67271
rect 89227 67305 89261 67321
rect 89227 67255 89261 67271
rect 1729 66969 1763 66985
rect 1729 66919 1763 66935
rect 89227 66969 89261 66985
rect 89227 66919 89261 66935
rect 1729 66633 1763 66649
rect 1729 66583 1763 66599
rect 89227 66633 89261 66649
rect 89227 66583 89261 66599
rect 1729 66297 1763 66313
rect 1729 66247 1763 66263
rect 89227 66297 89261 66313
rect 89227 66247 89261 66263
rect 1729 65961 1763 65977
rect 1729 65911 1763 65927
rect 89227 65961 89261 65977
rect 89227 65911 89261 65927
rect 1729 65625 1763 65641
rect 1729 65575 1763 65591
rect 89227 65625 89261 65641
rect 89227 65575 89261 65591
rect 1729 65289 1763 65305
rect 1729 65239 1763 65255
rect 89227 65289 89261 65305
rect 89227 65239 89261 65255
rect 1729 64953 1763 64969
rect 1729 64903 1763 64919
rect 89227 64953 89261 64969
rect 89227 64903 89261 64919
rect 1729 64617 1763 64633
rect 1729 64567 1763 64583
rect 89227 64617 89261 64633
rect 89227 64567 89261 64583
rect 1729 64281 1763 64297
rect 1729 64231 1763 64247
rect 89227 64281 89261 64297
rect 89227 64231 89261 64247
rect 1729 63945 1763 63961
rect 1729 63895 1763 63911
rect 89227 63945 89261 63961
rect 89227 63895 89261 63911
rect 1729 63609 1763 63625
rect 1729 63559 1763 63575
rect 89227 63609 89261 63625
rect 89227 63559 89261 63575
rect 1729 63273 1763 63289
rect 1729 63223 1763 63239
rect 89227 63273 89261 63289
rect 89227 63223 89261 63239
rect 1729 62937 1763 62953
rect 1729 62887 1763 62903
rect 89227 62937 89261 62953
rect 89227 62887 89261 62903
rect 1729 62601 1763 62617
rect 1729 62551 1763 62567
rect 89227 62601 89261 62617
rect 89227 62551 89261 62567
rect 1729 62265 1763 62281
rect 1729 62215 1763 62231
rect 89227 62265 89261 62281
rect 89227 62215 89261 62231
rect 1729 61929 1763 61945
rect 1729 61879 1763 61895
rect 89227 61929 89261 61945
rect 89227 61879 89261 61895
rect 1729 61593 1763 61609
rect 1729 61543 1763 61559
rect 89227 61593 89261 61609
rect 89227 61543 89261 61559
rect 1729 61257 1763 61273
rect 1729 61207 1763 61223
rect 89227 61257 89261 61273
rect 89227 61207 89261 61223
rect 1729 60921 1763 60937
rect 1729 60871 1763 60887
rect 89227 60921 89261 60937
rect 89227 60871 89261 60887
rect 1729 60585 1763 60601
rect 1729 60535 1763 60551
rect 89227 60585 89261 60601
rect 89227 60535 89261 60551
rect 1729 60249 1763 60265
rect 1729 60199 1763 60215
rect 89227 60249 89261 60265
rect 89227 60199 89261 60215
rect 1729 59913 1763 59929
rect 1729 59863 1763 59879
rect 89227 59913 89261 59929
rect 89227 59863 89261 59879
rect 1729 59577 1763 59593
rect 1729 59527 1763 59543
rect 89227 59577 89261 59593
rect 89227 59527 89261 59543
rect 1729 59241 1763 59257
rect 1729 59191 1763 59207
rect 89227 59241 89261 59257
rect 89227 59191 89261 59207
rect 1729 58905 1763 58921
rect 1729 58855 1763 58871
rect 89227 58905 89261 58921
rect 89227 58855 89261 58871
rect 1729 58569 1763 58585
rect 1729 58519 1763 58535
rect 89227 58569 89261 58585
rect 89227 58519 89261 58535
rect 1729 58233 1763 58249
rect 1729 58183 1763 58199
rect 89227 58233 89261 58249
rect 89227 58183 89261 58199
rect 1729 57897 1763 57913
rect 1729 57847 1763 57863
rect 89227 57897 89261 57913
rect 89227 57847 89261 57863
rect 1729 57561 1763 57577
rect 1729 57511 1763 57527
rect 89227 57561 89261 57577
rect 89227 57511 89261 57527
rect 1729 57225 1763 57241
rect 1729 57175 1763 57191
rect 89227 57225 89261 57241
rect 89227 57175 89261 57191
rect 1729 56889 1763 56905
rect 1729 56839 1763 56855
rect 89227 56889 89261 56905
rect 89227 56839 89261 56855
rect 1729 56553 1763 56569
rect 1729 56503 1763 56519
rect 89227 56553 89261 56569
rect 89227 56503 89261 56519
rect 1729 56217 1763 56233
rect 1729 56167 1763 56183
rect 89227 56217 89261 56233
rect 89227 56167 89261 56183
rect 1729 55881 1763 55897
rect 1729 55831 1763 55847
rect 89227 55881 89261 55897
rect 89227 55831 89261 55847
rect 1729 55545 1763 55561
rect 1729 55495 1763 55511
rect 89227 55545 89261 55561
rect 89227 55495 89261 55511
rect 1729 55209 1763 55225
rect 1729 55159 1763 55175
rect 89227 55209 89261 55225
rect 89227 55159 89261 55175
rect 1729 54873 1763 54889
rect 1729 54823 1763 54839
rect 89227 54873 89261 54889
rect 89227 54823 89261 54839
rect 1729 54537 1763 54553
rect 1729 54487 1763 54503
rect 89227 54537 89261 54553
rect 89227 54487 89261 54503
rect 1729 54201 1763 54217
rect 1729 54151 1763 54167
rect 89227 54201 89261 54217
rect 89227 54151 89261 54167
rect 1729 53865 1763 53881
rect 1729 53815 1763 53831
rect 89227 53865 89261 53881
rect 89227 53815 89261 53831
rect 1729 53529 1763 53545
rect 1729 53479 1763 53495
rect 89227 53529 89261 53545
rect 89227 53479 89261 53495
rect 1729 53193 1763 53209
rect 1729 53143 1763 53159
rect 89227 53193 89261 53209
rect 89227 53143 89261 53159
rect 1729 52857 1763 52873
rect 1729 52807 1763 52823
rect 89227 52857 89261 52873
rect 89227 52807 89261 52823
rect 1729 52521 1763 52537
rect 1729 52471 1763 52487
rect 89227 52521 89261 52537
rect 89227 52471 89261 52487
rect 1729 52185 1763 52201
rect 1729 52135 1763 52151
rect 89227 52185 89261 52201
rect 89227 52135 89261 52151
rect 1729 51849 1763 51865
rect 1729 51799 1763 51815
rect 89227 51849 89261 51865
rect 89227 51799 89261 51815
rect 1729 51513 1763 51529
rect 1729 51463 1763 51479
rect 89227 51513 89261 51529
rect 89227 51463 89261 51479
rect 1729 51177 1763 51193
rect 1729 51127 1763 51143
rect 89227 51177 89261 51193
rect 89227 51127 89261 51143
rect 1729 50841 1763 50857
rect 1729 50791 1763 50807
rect 89227 50841 89261 50857
rect 89227 50791 89261 50807
rect 1729 50505 1763 50521
rect 1729 50455 1763 50471
rect 89227 50505 89261 50521
rect 89227 50455 89261 50471
rect 1729 50169 1763 50185
rect 1729 50119 1763 50135
rect 89227 50169 89261 50185
rect 89227 50119 89261 50135
rect 1729 49833 1763 49849
rect 1729 49783 1763 49799
rect 89227 49833 89261 49849
rect 89227 49783 89261 49799
rect 1729 49497 1763 49513
rect 1729 49447 1763 49463
rect 89227 49497 89261 49513
rect 89227 49447 89261 49463
rect 1729 49161 1763 49177
rect 1729 49111 1763 49127
rect 89227 49161 89261 49177
rect 89227 49111 89261 49127
rect 1729 48825 1763 48841
rect 1729 48775 1763 48791
rect 89227 48825 89261 48841
rect 89227 48775 89261 48791
rect 1729 48489 1763 48505
rect 1729 48439 1763 48455
rect 89227 48489 89261 48505
rect 89227 48439 89261 48455
rect 1729 48153 1763 48169
rect 1729 48103 1763 48119
rect 89227 48153 89261 48169
rect 89227 48103 89261 48119
rect 1729 47817 1763 47833
rect 1729 47767 1763 47783
rect 89227 47817 89261 47833
rect 89227 47767 89261 47783
rect 1729 47481 1763 47497
rect 1729 47431 1763 47447
rect 89227 47481 89261 47497
rect 89227 47431 89261 47447
rect 1729 47145 1763 47161
rect 1729 47095 1763 47111
rect 89227 47145 89261 47161
rect 89227 47095 89261 47111
rect 1729 46809 1763 46825
rect 1729 46759 1763 46775
rect 89227 46809 89261 46825
rect 89227 46759 89261 46775
rect 1729 46473 1763 46489
rect 1729 46423 1763 46439
rect 89227 46473 89261 46489
rect 89227 46423 89261 46439
rect 1729 46137 1763 46153
rect 1729 46087 1763 46103
rect 89227 46137 89261 46153
rect 89227 46087 89261 46103
rect 1729 45801 1763 45817
rect 1729 45751 1763 45767
rect 89227 45801 89261 45817
rect 89227 45751 89261 45767
rect 1729 45465 1763 45481
rect 1729 45415 1763 45431
rect 89227 45465 89261 45481
rect 89227 45415 89261 45431
rect 1729 45129 1763 45145
rect 1729 45079 1763 45095
rect 89227 45129 89261 45145
rect 89227 45079 89261 45095
rect 1729 44793 1763 44809
rect 1729 44743 1763 44759
rect 89227 44793 89261 44809
rect 89227 44743 89261 44759
rect 1729 44457 1763 44473
rect 1729 44407 1763 44423
rect 89227 44457 89261 44473
rect 89227 44407 89261 44423
rect 1729 44121 1763 44137
rect 1729 44071 1763 44087
rect 89227 44121 89261 44137
rect 89227 44071 89261 44087
rect 1729 43785 1763 43801
rect 1729 43735 1763 43751
rect 89227 43785 89261 43801
rect 89227 43735 89261 43751
rect 1729 43449 1763 43465
rect 1729 43399 1763 43415
rect 89227 43449 89261 43465
rect 89227 43399 89261 43415
rect 1729 43113 1763 43129
rect 1729 43063 1763 43079
rect 89227 43113 89261 43129
rect 89227 43063 89261 43079
rect 1729 42777 1763 42793
rect 1729 42727 1763 42743
rect 89227 42777 89261 42793
rect 89227 42727 89261 42743
rect 1729 42441 1763 42457
rect 1729 42391 1763 42407
rect 89227 42441 89261 42457
rect 89227 42391 89261 42407
rect 1729 42105 1763 42121
rect 1729 42055 1763 42071
rect 89227 42105 89261 42121
rect 89227 42055 89261 42071
rect 1729 41769 1763 41785
rect 1729 41719 1763 41735
rect 89227 41769 89261 41785
rect 89227 41719 89261 41735
rect 1729 41433 1763 41449
rect 1729 41383 1763 41399
rect 89227 41433 89261 41449
rect 89227 41383 89261 41399
rect 1729 41097 1763 41113
rect 1729 41047 1763 41063
rect 89227 41097 89261 41113
rect 89227 41047 89261 41063
rect 1729 40761 1763 40777
rect 1729 40711 1763 40727
rect 89227 40761 89261 40777
rect 89227 40711 89261 40727
rect 1729 40425 1763 40441
rect 1729 40375 1763 40391
rect 89227 40425 89261 40441
rect 89227 40375 89261 40391
rect 1729 40089 1763 40105
rect 1729 40039 1763 40055
rect 89227 40089 89261 40105
rect 89227 40039 89261 40055
rect 1729 39753 1763 39769
rect 1729 39703 1763 39719
rect 89227 39753 89261 39769
rect 89227 39703 89261 39719
rect 1729 39417 1763 39433
rect 1729 39367 1763 39383
rect 89227 39417 89261 39433
rect 89227 39367 89261 39383
rect 1729 39081 1763 39097
rect 1729 39031 1763 39047
rect 89227 39081 89261 39097
rect 89227 39031 89261 39047
rect 1729 38745 1763 38761
rect 1729 38695 1763 38711
rect 89227 38745 89261 38761
rect 89227 38695 89261 38711
rect 1729 38409 1763 38425
rect 1729 38359 1763 38375
rect 89227 38409 89261 38425
rect 89227 38359 89261 38375
rect 1729 38073 1763 38089
rect 1729 38023 1763 38039
rect 89227 38073 89261 38089
rect 89227 38023 89261 38039
rect 1729 37737 1763 37753
rect 1729 37687 1763 37703
rect 89227 37737 89261 37753
rect 89227 37687 89261 37703
rect 1729 37401 1763 37417
rect 1729 37351 1763 37367
rect 89227 37401 89261 37417
rect 89227 37351 89261 37367
rect 1729 37065 1763 37081
rect 1729 37015 1763 37031
rect 89227 37065 89261 37081
rect 89227 37015 89261 37031
rect 1729 36729 1763 36745
rect 1729 36679 1763 36695
rect 89227 36729 89261 36745
rect 89227 36679 89261 36695
rect 1729 36393 1763 36409
rect 1729 36343 1763 36359
rect 89227 36393 89261 36409
rect 89227 36343 89261 36359
rect 1729 36057 1763 36073
rect 1729 36007 1763 36023
rect 89227 36057 89261 36073
rect 89227 36007 89261 36023
rect 1729 35721 1763 35737
rect 1729 35671 1763 35687
rect 89227 35721 89261 35737
rect 89227 35671 89261 35687
rect 1729 35385 1763 35401
rect 1729 35335 1763 35351
rect 89227 35385 89261 35401
rect 89227 35335 89261 35351
rect 1729 35049 1763 35065
rect 1729 34999 1763 35015
rect 89227 35049 89261 35065
rect 89227 34999 89261 35015
rect 1729 34713 1763 34729
rect 1729 34663 1763 34679
rect 89227 34713 89261 34729
rect 89227 34663 89261 34679
rect 1729 34377 1763 34393
rect 1729 34327 1763 34343
rect 89227 34377 89261 34393
rect 89227 34327 89261 34343
rect 1729 34041 1763 34057
rect 1729 33991 1763 34007
rect 89227 34041 89261 34057
rect 89227 33991 89261 34007
rect 1729 33705 1763 33721
rect 1729 33655 1763 33671
rect 89227 33705 89261 33721
rect 89227 33655 89261 33671
rect 1729 33369 1763 33385
rect 1729 33319 1763 33335
rect 89227 33369 89261 33385
rect 89227 33319 89261 33335
rect 1729 33033 1763 33049
rect 1729 32983 1763 32999
rect 89227 33033 89261 33049
rect 89227 32983 89261 32999
rect 1729 32697 1763 32713
rect 1729 32647 1763 32663
rect 89227 32697 89261 32713
rect 89227 32647 89261 32663
rect 1729 32361 1763 32377
rect 1729 32311 1763 32327
rect 89227 32361 89261 32377
rect 89227 32311 89261 32327
rect 1729 32025 1763 32041
rect 1729 31975 1763 31991
rect 89227 32025 89261 32041
rect 89227 31975 89261 31991
rect 1729 31689 1763 31705
rect 1729 31639 1763 31655
rect 89227 31689 89261 31705
rect 89227 31639 89261 31655
rect 1729 31353 1763 31369
rect 1729 31303 1763 31319
rect 89227 31353 89261 31369
rect 89227 31303 89261 31319
rect 1729 31017 1763 31033
rect 1729 30967 1763 30983
rect 89227 31017 89261 31033
rect 89227 30967 89261 30983
rect 1729 30681 1763 30697
rect 1729 30631 1763 30647
rect 89227 30681 89261 30697
rect 89227 30631 89261 30647
rect 1729 30345 1763 30361
rect 1729 30295 1763 30311
rect 89227 30345 89261 30361
rect 89227 30295 89261 30311
rect 1729 30009 1763 30025
rect 1729 29959 1763 29975
rect 89227 30009 89261 30025
rect 89227 29959 89261 29975
rect 1729 29673 1763 29689
rect 1729 29623 1763 29639
rect 89227 29673 89261 29689
rect 89227 29623 89261 29639
rect 1729 29337 1763 29353
rect 1729 29287 1763 29303
rect 89227 29337 89261 29353
rect 89227 29287 89261 29303
rect 1729 29001 1763 29017
rect 1729 28951 1763 28967
rect 89227 29001 89261 29017
rect 89227 28951 89261 28967
rect 1729 28665 1763 28681
rect 1729 28615 1763 28631
rect 89227 28665 89261 28681
rect 89227 28615 89261 28631
rect 1729 28329 1763 28345
rect 1729 28279 1763 28295
rect 89227 28329 89261 28345
rect 89227 28279 89261 28295
rect 1729 27993 1763 28009
rect 1729 27943 1763 27959
rect 89227 27993 89261 28009
rect 89227 27943 89261 27959
rect 1729 27657 1763 27673
rect 1729 27607 1763 27623
rect 89227 27657 89261 27673
rect 89227 27607 89261 27623
rect 1729 27321 1763 27337
rect 1729 27271 1763 27287
rect 89227 27321 89261 27337
rect 89227 27271 89261 27287
rect 1729 26985 1763 27001
rect 1729 26935 1763 26951
rect 89227 26985 89261 27001
rect 89227 26935 89261 26951
rect 1729 26649 1763 26665
rect 1729 26599 1763 26615
rect 89227 26649 89261 26665
rect 89227 26599 89261 26615
rect 1729 26313 1763 26329
rect 1729 26263 1763 26279
rect 89227 26313 89261 26329
rect 89227 26263 89261 26279
rect 1729 25977 1763 25993
rect 1729 25927 1763 25943
rect 89227 25977 89261 25993
rect 89227 25927 89261 25943
rect 1729 25641 1763 25657
rect 1729 25591 1763 25607
rect 89227 25641 89261 25657
rect 89227 25591 89261 25607
rect 1729 25305 1763 25321
rect 1729 25255 1763 25271
rect 89227 25305 89261 25321
rect 89227 25255 89261 25271
rect 1729 24969 1763 24985
rect 1729 24919 1763 24935
rect 89227 24969 89261 24985
rect 89227 24919 89261 24935
rect 1729 24633 1763 24649
rect 1729 24583 1763 24599
rect 89227 24633 89261 24649
rect 89227 24583 89261 24599
rect 1729 24297 1763 24313
rect 1729 24247 1763 24263
rect 89227 24297 89261 24313
rect 89227 24247 89261 24263
rect 1729 23961 1763 23977
rect 1729 23911 1763 23927
rect 89227 23961 89261 23977
rect 89227 23911 89261 23927
rect 1729 23625 1763 23641
rect 1729 23575 1763 23591
rect 89227 23625 89261 23641
rect 89227 23575 89261 23591
rect 1729 23289 1763 23305
rect 1729 23239 1763 23255
rect 89227 23289 89261 23305
rect 89227 23239 89261 23255
rect 1729 22953 1763 22969
rect 1729 22903 1763 22919
rect 89227 22953 89261 22969
rect 89227 22903 89261 22919
rect 1729 22617 1763 22633
rect 1729 22567 1763 22583
rect 89227 22617 89261 22633
rect 89227 22567 89261 22583
rect 1729 22281 1763 22297
rect 1729 22231 1763 22247
rect 89227 22281 89261 22297
rect 89227 22231 89261 22247
rect 1729 21945 1763 21961
rect 1729 21895 1763 21911
rect 89227 21945 89261 21961
rect 89227 21895 89261 21911
rect 1729 21609 1763 21625
rect 1729 21559 1763 21575
rect 89227 21609 89261 21625
rect 89227 21559 89261 21575
rect 1729 21273 1763 21289
rect 1729 21223 1763 21239
rect 89227 21273 89261 21289
rect 89227 21223 89261 21239
rect 1729 20937 1763 20953
rect 1729 20887 1763 20903
rect 89227 20937 89261 20953
rect 89227 20887 89261 20903
rect 1729 20601 1763 20617
rect 1729 20551 1763 20567
rect 89227 20601 89261 20617
rect 89227 20551 89261 20567
rect 1729 20265 1763 20281
rect 1729 20215 1763 20231
rect 89227 20265 89261 20281
rect 89227 20215 89261 20231
rect 1729 19929 1763 19945
rect 1729 19879 1763 19895
rect 89227 19929 89261 19945
rect 89227 19879 89261 19895
rect 1729 19593 1763 19609
rect 1729 19543 1763 19559
rect 89227 19593 89261 19609
rect 89227 19543 89261 19559
rect 1729 19257 1763 19273
rect 1729 19207 1763 19223
rect 89227 19257 89261 19273
rect 89227 19207 89261 19223
rect 1729 18921 1763 18937
rect 1729 18871 1763 18887
rect 89227 18921 89261 18937
rect 89227 18871 89261 18887
rect 1729 18585 1763 18601
rect 1729 18535 1763 18551
rect 89227 18585 89261 18601
rect 89227 18535 89261 18551
rect 1729 18249 1763 18265
rect 1729 18199 1763 18215
rect 89227 18249 89261 18265
rect 89227 18199 89261 18215
rect 1729 17913 1763 17929
rect 1729 17863 1763 17879
rect 89227 17913 89261 17929
rect 89227 17863 89261 17879
rect 1729 17577 1763 17593
rect 1729 17527 1763 17543
rect 89227 17577 89261 17593
rect 89227 17527 89261 17543
rect 1729 17241 1763 17257
rect 1729 17191 1763 17207
rect 89227 17241 89261 17257
rect 89227 17191 89261 17207
rect 1729 16905 1763 16921
rect 1729 16855 1763 16871
rect 89227 16905 89261 16921
rect 89227 16855 89261 16871
rect 1729 16569 1763 16585
rect 1729 16519 1763 16535
rect 89227 16569 89261 16585
rect 89227 16519 89261 16535
rect 1729 16233 1763 16249
rect 1729 16183 1763 16199
rect 89227 16233 89261 16249
rect 89227 16183 89261 16199
rect 1729 15897 1763 15913
rect 1729 15847 1763 15863
rect 89227 15897 89261 15913
rect 89227 15847 89261 15863
rect 1729 15561 1763 15577
rect 1729 15511 1763 15527
rect 89227 15561 89261 15577
rect 89227 15511 89261 15527
rect 1729 15225 1763 15241
rect 1729 15175 1763 15191
rect 89227 15225 89261 15241
rect 89227 15175 89261 15191
rect 1729 14889 1763 14905
rect 1729 14839 1763 14855
rect 89227 14889 89261 14905
rect 89227 14839 89261 14855
rect 1729 14553 1763 14569
rect 1729 14503 1763 14519
rect 89227 14553 89261 14569
rect 89227 14503 89261 14519
rect 1729 14217 1763 14233
rect 1729 14167 1763 14183
rect 89227 14217 89261 14233
rect 89227 14167 89261 14183
rect 1729 13881 1763 13897
rect 1729 13831 1763 13847
rect 89227 13881 89261 13897
rect 89227 13831 89261 13847
rect 1729 13545 1763 13561
rect 1729 13495 1763 13511
rect 89227 13545 89261 13561
rect 89227 13495 89261 13511
rect 1729 13209 1763 13225
rect 1729 13159 1763 13175
rect 89227 13209 89261 13225
rect 89227 13159 89261 13175
rect 1729 12873 1763 12889
rect 1729 12823 1763 12839
rect 89227 12873 89261 12889
rect 89227 12823 89261 12839
rect 1729 12537 1763 12553
rect 1729 12487 1763 12503
rect 89227 12537 89261 12553
rect 89227 12487 89261 12503
rect 1729 12201 1763 12217
rect 1729 12151 1763 12167
rect 89227 12201 89261 12217
rect 89227 12151 89261 12167
rect 1729 11865 1763 11881
rect 1729 11815 1763 11831
rect 89227 11865 89261 11881
rect 89227 11815 89261 11831
rect 1729 11529 1763 11545
rect 1729 11479 1763 11495
rect 89227 11529 89261 11545
rect 89227 11479 89261 11495
rect 1729 11193 1763 11209
rect 1729 11143 1763 11159
rect 89227 11193 89261 11209
rect 89227 11143 89261 11159
rect 1729 10857 1763 10873
rect 1729 10807 1763 10823
rect 89227 10857 89261 10873
rect 89227 10807 89261 10823
rect 1729 10521 1763 10537
rect 1729 10471 1763 10487
rect 89227 10521 89261 10537
rect 89227 10471 89261 10487
rect 1729 10185 1763 10201
rect 1729 10135 1763 10151
rect 89227 10185 89261 10201
rect 89227 10135 89261 10151
rect 1729 9849 1763 9865
rect 1729 9799 1763 9815
rect 89227 9849 89261 9865
rect 89227 9799 89261 9815
rect 1729 9513 1763 9529
rect 1729 9463 1763 9479
rect 89227 9513 89261 9529
rect 89227 9463 89261 9479
rect 1729 9177 1763 9193
rect 1729 9127 1763 9143
rect 89227 9177 89261 9193
rect 89227 9127 89261 9143
rect 1729 8841 1763 8857
rect 1729 8791 1763 8807
rect 89227 8841 89261 8857
rect 89227 8791 89261 8807
rect 1729 8505 1763 8521
rect 1729 8455 1763 8471
rect 89227 8505 89261 8521
rect 89227 8455 89261 8471
rect 1729 8169 1763 8185
rect 1729 8119 1763 8135
rect 89227 8169 89261 8185
rect 89227 8119 89261 8135
rect 1729 7833 1763 7849
rect 1729 7783 1763 7799
rect 89227 7833 89261 7849
rect 89227 7783 89261 7799
rect 1729 7497 1763 7513
rect 1729 7447 1763 7463
rect 89227 7497 89261 7513
rect 89227 7447 89261 7463
rect 1729 7161 1763 7177
rect 1729 7111 1763 7127
rect 89227 7161 89261 7177
rect 89227 7111 89261 7127
rect 1729 6825 1763 6841
rect 1729 6775 1763 6791
rect 89227 6825 89261 6841
rect 89227 6775 89261 6791
rect 1729 6489 1763 6505
rect 1729 6439 1763 6455
rect 89227 6489 89261 6505
rect 89227 6439 89261 6455
rect 1729 6153 1763 6169
rect 1729 6103 1763 6119
rect 89227 6153 89261 6169
rect 89227 6103 89261 6119
rect 1729 5817 1763 5833
rect 1729 5767 1763 5783
rect 89227 5817 89261 5833
rect 89227 5767 89261 5783
rect 1729 5481 1763 5497
rect 1729 5431 1763 5447
rect 89227 5481 89261 5497
rect 89227 5431 89261 5447
rect 1729 5145 1763 5161
rect 1729 5095 1763 5111
rect 89227 5145 89261 5161
rect 89227 5095 89261 5111
rect 1729 4809 1763 4825
rect 1729 4759 1763 4775
rect 89227 4809 89261 4825
rect 89227 4759 89261 4775
rect 1729 4473 1763 4489
rect 1729 4423 1763 4439
rect 89227 4473 89261 4489
rect 89227 4423 89261 4439
rect 1729 4137 1763 4153
rect 1729 4087 1763 4103
rect 89227 4137 89261 4153
rect 89227 4087 89261 4103
rect 1729 3801 1763 3817
rect 1729 3751 1763 3767
rect 89227 3801 89261 3817
rect 89227 3751 89261 3767
rect 1729 3465 1763 3481
rect 1729 3415 1763 3431
rect 89227 3465 89261 3481
rect 89227 3415 89261 3431
rect 1729 3129 1763 3145
rect 1729 3079 1763 3095
rect 89227 3129 89261 3145
rect 89227 3079 89261 3095
rect 1729 2793 1763 2809
rect 1729 2743 1763 2759
rect 89227 2793 89261 2809
rect 89227 2743 89261 2759
rect 1729 2457 1763 2473
rect 1729 2407 1763 2423
rect 89227 2457 89261 2473
rect 89227 2407 89261 2423
rect 1729 2121 1763 2137
rect 1729 2071 1763 2087
rect 89227 2121 89261 2137
rect 89227 2071 89261 2087
rect 2065 1785 2099 1801
rect 2065 1735 2099 1751
rect 2401 1785 2435 1801
rect 2401 1735 2435 1751
rect 2737 1785 2771 1801
rect 2737 1735 2771 1751
rect 3073 1785 3107 1801
rect 3073 1735 3107 1751
rect 3409 1785 3443 1801
rect 3409 1735 3443 1751
rect 3745 1785 3779 1801
rect 3745 1735 3779 1751
rect 4081 1785 4115 1801
rect 4081 1735 4115 1751
rect 4417 1785 4451 1801
rect 4417 1735 4451 1751
rect 4753 1785 4787 1801
rect 4753 1735 4787 1751
rect 5089 1785 5123 1801
rect 5089 1735 5123 1751
rect 5425 1785 5459 1801
rect 5425 1735 5459 1751
rect 5761 1785 5795 1801
rect 5761 1735 5795 1751
rect 6097 1785 6131 1801
rect 6097 1735 6131 1751
rect 6433 1785 6467 1801
rect 6433 1735 6467 1751
rect 6769 1785 6803 1801
rect 6769 1735 6803 1751
rect 7105 1785 7139 1801
rect 7105 1735 7139 1751
rect 7441 1785 7475 1801
rect 7441 1735 7475 1751
rect 7777 1785 7811 1801
rect 7777 1735 7811 1751
rect 8113 1785 8147 1801
rect 8113 1735 8147 1751
rect 8449 1785 8483 1801
rect 8449 1735 8483 1751
rect 8785 1785 8819 1801
rect 8785 1735 8819 1751
rect 9121 1785 9155 1801
rect 9121 1735 9155 1751
rect 9457 1785 9491 1801
rect 9457 1735 9491 1751
rect 9793 1785 9827 1801
rect 9793 1735 9827 1751
rect 10129 1785 10163 1801
rect 10129 1735 10163 1751
rect 10465 1785 10499 1801
rect 10465 1735 10499 1751
rect 10801 1785 10835 1801
rect 10801 1735 10835 1751
rect 11137 1785 11171 1801
rect 11137 1735 11171 1751
rect 11473 1785 11507 1801
rect 11473 1735 11507 1751
rect 11809 1785 11843 1801
rect 11809 1735 11843 1751
rect 12145 1785 12179 1801
rect 12145 1735 12179 1751
rect 12481 1785 12515 1801
rect 12481 1735 12515 1751
rect 12817 1785 12851 1801
rect 12817 1735 12851 1751
rect 13153 1785 13187 1801
rect 13153 1735 13187 1751
rect 13489 1785 13523 1801
rect 13489 1735 13523 1751
rect 13825 1785 13859 1801
rect 13825 1735 13859 1751
rect 14161 1785 14195 1801
rect 14161 1735 14195 1751
rect 14497 1785 14531 1801
rect 14497 1735 14531 1751
rect 14833 1785 14867 1801
rect 14833 1735 14867 1751
rect 15169 1785 15203 1801
rect 15169 1735 15203 1751
rect 15505 1785 15539 1801
rect 15505 1735 15539 1751
rect 15841 1785 15875 1801
rect 15841 1735 15875 1751
rect 16177 1785 16211 1801
rect 16177 1735 16211 1751
rect 16513 1785 16547 1801
rect 16513 1735 16547 1751
rect 16849 1785 16883 1801
rect 16849 1735 16883 1751
rect 17185 1785 17219 1801
rect 17185 1735 17219 1751
rect 17521 1785 17555 1801
rect 17521 1735 17555 1751
rect 17857 1785 17891 1801
rect 17857 1735 17891 1751
rect 18193 1785 18227 1801
rect 18193 1735 18227 1751
rect 18529 1785 18563 1801
rect 18529 1735 18563 1751
rect 18865 1785 18899 1801
rect 18865 1735 18899 1751
rect 19201 1785 19235 1801
rect 19201 1735 19235 1751
rect 19537 1785 19571 1801
rect 19537 1735 19571 1751
rect 19873 1785 19907 1801
rect 19873 1735 19907 1751
rect 20209 1785 20243 1801
rect 20209 1735 20243 1751
rect 20545 1785 20579 1801
rect 20545 1735 20579 1751
rect 20881 1785 20915 1801
rect 20881 1735 20915 1751
rect 21217 1785 21251 1801
rect 21217 1735 21251 1751
rect 21553 1785 21587 1801
rect 21553 1735 21587 1751
rect 21889 1785 21923 1801
rect 21889 1735 21923 1751
rect 22225 1785 22259 1801
rect 22225 1735 22259 1751
rect 22561 1785 22595 1801
rect 22561 1735 22595 1751
rect 22897 1785 22931 1801
rect 22897 1735 22931 1751
rect 23233 1785 23267 1801
rect 23233 1735 23267 1751
rect 23569 1785 23603 1801
rect 23569 1735 23603 1751
rect 23905 1785 23939 1801
rect 23905 1735 23939 1751
rect 24241 1785 24275 1801
rect 24241 1735 24275 1751
rect 24577 1785 24611 1801
rect 24577 1735 24611 1751
rect 24913 1785 24947 1801
rect 24913 1735 24947 1751
rect 25249 1785 25283 1801
rect 25249 1735 25283 1751
rect 25585 1785 25619 1801
rect 25585 1735 25619 1751
rect 25921 1785 25955 1801
rect 25921 1735 25955 1751
rect 26257 1785 26291 1801
rect 26257 1735 26291 1751
rect 26593 1785 26627 1801
rect 26593 1735 26627 1751
rect 26929 1785 26963 1801
rect 26929 1735 26963 1751
rect 27265 1785 27299 1801
rect 27265 1735 27299 1751
rect 27601 1785 27635 1801
rect 27601 1735 27635 1751
rect 27937 1785 27971 1801
rect 27937 1735 27971 1751
rect 28273 1785 28307 1801
rect 28273 1735 28307 1751
rect 28609 1785 28643 1801
rect 28609 1735 28643 1751
rect 28945 1785 28979 1801
rect 28945 1735 28979 1751
rect 29281 1785 29315 1801
rect 29281 1735 29315 1751
rect 29617 1785 29651 1801
rect 29617 1735 29651 1751
rect 29953 1785 29987 1801
rect 29953 1735 29987 1751
rect 30289 1785 30323 1801
rect 30289 1735 30323 1751
rect 30625 1785 30659 1801
rect 30625 1735 30659 1751
rect 30961 1785 30995 1801
rect 30961 1735 30995 1751
rect 31297 1785 31331 1801
rect 31297 1735 31331 1751
rect 31633 1785 31667 1801
rect 31633 1735 31667 1751
rect 31969 1785 32003 1801
rect 31969 1735 32003 1751
rect 32305 1785 32339 1801
rect 32305 1735 32339 1751
rect 32641 1785 32675 1801
rect 32641 1735 32675 1751
rect 32977 1785 33011 1801
rect 32977 1735 33011 1751
rect 33313 1785 33347 1801
rect 33313 1735 33347 1751
rect 33649 1785 33683 1801
rect 33649 1735 33683 1751
rect 33985 1785 34019 1801
rect 33985 1735 34019 1751
rect 34321 1785 34355 1801
rect 34321 1735 34355 1751
rect 34657 1785 34691 1801
rect 34657 1735 34691 1751
rect 34993 1785 35027 1801
rect 34993 1735 35027 1751
rect 35329 1785 35363 1801
rect 35329 1735 35363 1751
rect 35665 1785 35699 1801
rect 35665 1735 35699 1751
rect 36001 1785 36035 1801
rect 36001 1735 36035 1751
rect 36337 1785 36371 1801
rect 36337 1735 36371 1751
rect 36673 1785 36707 1801
rect 36673 1735 36707 1751
rect 37009 1785 37043 1801
rect 37009 1735 37043 1751
rect 37345 1785 37379 1801
rect 37345 1735 37379 1751
rect 37681 1785 37715 1801
rect 37681 1735 37715 1751
rect 38017 1785 38051 1801
rect 38017 1735 38051 1751
rect 38353 1785 38387 1801
rect 38353 1735 38387 1751
rect 38689 1785 38723 1801
rect 38689 1735 38723 1751
rect 39025 1785 39059 1801
rect 39025 1735 39059 1751
rect 39361 1785 39395 1801
rect 39361 1735 39395 1751
rect 39697 1785 39731 1801
rect 39697 1735 39731 1751
rect 40033 1785 40067 1801
rect 40033 1735 40067 1751
rect 40369 1785 40403 1801
rect 40369 1735 40403 1751
rect 40705 1785 40739 1801
rect 40705 1735 40739 1751
rect 41041 1785 41075 1801
rect 41041 1735 41075 1751
rect 41377 1785 41411 1801
rect 41377 1735 41411 1751
rect 41713 1785 41747 1801
rect 41713 1735 41747 1751
rect 42049 1785 42083 1801
rect 42049 1735 42083 1751
rect 42385 1785 42419 1801
rect 42385 1735 42419 1751
rect 42721 1785 42755 1801
rect 42721 1735 42755 1751
rect 43057 1785 43091 1801
rect 43057 1735 43091 1751
rect 43393 1785 43427 1801
rect 43393 1735 43427 1751
rect 43729 1785 43763 1801
rect 43729 1735 43763 1751
rect 44065 1785 44099 1801
rect 44065 1735 44099 1751
rect 44401 1785 44435 1801
rect 44401 1735 44435 1751
rect 44737 1785 44771 1801
rect 44737 1735 44771 1751
rect 45073 1785 45107 1801
rect 45073 1735 45107 1751
rect 45409 1785 45443 1801
rect 45409 1735 45443 1751
rect 45745 1785 45779 1801
rect 45745 1735 45779 1751
rect 46081 1785 46115 1801
rect 46081 1735 46115 1751
rect 46417 1785 46451 1801
rect 46417 1735 46451 1751
rect 46753 1785 46787 1801
rect 46753 1735 46787 1751
rect 47089 1785 47123 1801
rect 47089 1735 47123 1751
rect 47425 1785 47459 1801
rect 47425 1735 47459 1751
rect 47761 1785 47795 1801
rect 47761 1735 47795 1751
rect 48097 1785 48131 1801
rect 48097 1735 48131 1751
rect 48433 1785 48467 1801
rect 48433 1735 48467 1751
rect 48769 1785 48803 1801
rect 48769 1735 48803 1751
rect 49105 1785 49139 1801
rect 49105 1735 49139 1751
rect 49441 1785 49475 1801
rect 49441 1735 49475 1751
rect 49777 1785 49811 1801
rect 49777 1735 49811 1751
rect 50113 1785 50147 1801
rect 50113 1735 50147 1751
rect 50449 1785 50483 1801
rect 50449 1735 50483 1751
rect 50785 1785 50819 1801
rect 50785 1735 50819 1751
rect 51121 1785 51155 1801
rect 51121 1735 51155 1751
rect 51457 1785 51491 1801
rect 51457 1735 51491 1751
rect 51793 1785 51827 1801
rect 51793 1735 51827 1751
rect 52129 1785 52163 1801
rect 52129 1735 52163 1751
rect 52465 1785 52499 1801
rect 52465 1735 52499 1751
rect 52801 1785 52835 1801
rect 52801 1735 52835 1751
rect 53137 1785 53171 1801
rect 53137 1735 53171 1751
rect 53473 1785 53507 1801
rect 53473 1735 53507 1751
rect 53809 1785 53843 1801
rect 53809 1735 53843 1751
rect 54145 1785 54179 1801
rect 54145 1735 54179 1751
rect 54481 1785 54515 1801
rect 54481 1735 54515 1751
rect 54817 1785 54851 1801
rect 54817 1735 54851 1751
rect 55153 1785 55187 1801
rect 55153 1735 55187 1751
rect 55489 1785 55523 1801
rect 55489 1735 55523 1751
rect 55825 1785 55859 1801
rect 55825 1735 55859 1751
rect 56161 1785 56195 1801
rect 56161 1735 56195 1751
rect 56497 1785 56531 1801
rect 56497 1735 56531 1751
rect 56833 1785 56867 1801
rect 56833 1735 56867 1751
rect 57169 1785 57203 1801
rect 57169 1735 57203 1751
rect 57505 1785 57539 1801
rect 57505 1735 57539 1751
rect 57841 1785 57875 1801
rect 57841 1735 57875 1751
rect 58177 1785 58211 1801
rect 58177 1735 58211 1751
rect 58513 1785 58547 1801
rect 58513 1735 58547 1751
rect 58849 1785 58883 1801
rect 58849 1735 58883 1751
rect 59185 1785 59219 1801
rect 59185 1735 59219 1751
rect 59521 1785 59555 1801
rect 59521 1735 59555 1751
rect 59857 1785 59891 1801
rect 59857 1735 59891 1751
rect 60193 1785 60227 1801
rect 60193 1735 60227 1751
rect 60529 1785 60563 1801
rect 60529 1735 60563 1751
rect 60865 1785 60899 1801
rect 60865 1735 60899 1751
rect 61201 1785 61235 1801
rect 61201 1735 61235 1751
rect 61537 1785 61571 1801
rect 61537 1735 61571 1751
rect 61873 1785 61907 1801
rect 61873 1735 61907 1751
rect 62209 1785 62243 1801
rect 62209 1735 62243 1751
rect 62545 1785 62579 1801
rect 62545 1735 62579 1751
rect 62881 1785 62915 1801
rect 62881 1735 62915 1751
rect 63217 1785 63251 1801
rect 63217 1735 63251 1751
rect 63553 1785 63587 1801
rect 63553 1735 63587 1751
rect 63889 1785 63923 1801
rect 63889 1735 63923 1751
rect 64225 1785 64259 1801
rect 64225 1735 64259 1751
rect 64561 1785 64595 1801
rect 64561 1735 64595 1751
rect 64897 1785 64931 1801
rect 64897 1735 64931 1751
rect 65233 1785 65267 1801
rect 65233 1735 65267 1751
rect 65569 1785 65603 1801
rect 65569 1735 65603 1751
rect 65905 1785 65939 1801
rect 65905 1735 65939 1751
rect 66241 1785 66275 1801
rect 66241 1735 66275 1751
rect 66577 1785 66611 1801
rect 66577 1735 66611 1751
rect 66913 1785 66947 1801
rect 66913 1735 66947 1751
rect 67249 1785 67283 1801
rect 67249 1735 67283 1751
rect 67585 1785 67619 1801
rect 67585 1735 67619 1751
rect 67921 1785 67955 1801
rect 67921 1735 67955 1751
rect 68257 1785 68291 1801
rect 68257 1735 68291 1751
rect 68593 1785 68627 1801
rect 68593 1735 68627 1751
rect 68929 1785 68963 1801
rect 68929 1735 68963 1751
rect 69265 1785 69299 1801
rect 69265 1735 69299 1751
rect 69601 1785 69635 1801
rect 69601 1735 69635 1751
rect 69937 1785 69971 1801
rect 69937 1735 69971 1751
rect 70273 1785 70307 1801
rect 70273 1735 70307 1751
rect 70609 1785 70643 1801
rect 70609 1735 70643 1751
rect 70945 1785 70979 1801
rect 70945 1735 70979 1751
rect 71281 1785 71315 1801
rect 71281 1735 71315 1751
rect 71617 1785 71651 1801
rect 71617 1735 71651 1751
rect 71953 1785 71987 1801
rect 71953 1735 71987 1751
rect 72289 1785 72323 1801
rect 72289 1735 72323 1751
rect 72625 1785 72659 1801
rect 72625 1735 72659 1751
rect 72961 1785 72995 1801
rect 72961 1735 72995 1751
rect 73297 1785 73331 1801
rect 73297 1735 73331 1751
rect 73633 1785 73667 1801
rect 73633 1735 73667 1751
rect 73969 1785 74003 1801
rect 73969 1735 74003 1751
rect 74305 1785 74339 1801
rect 74305 1735 74339 1751
rect 74641 1785 74675 1801
rect 74641 1735 74675 1751
rect 74977 1785 75011 1801
rect 74977 1735 75011 1751
rect 75313 1785 75347 1801
rect 75313 1735 75347 1751
rect 75649 1785 75683 1801
rect 75649 1735 75683 1751
rect 75985 1785 76019 1801
rect 75985 1735 76019 1751
rect 76321 1785 76355 1801
rect 76321 1735 76355 1751
rect 76657 1785 76691 1801
rect 76657 1735 76691 1751
rect 76993 1785 77027 1801
rect 76993 1735 77027 1751
rect 77329 1785 77363 1801
rect 77329 1735 77363 1751
rect 77665 1785 77699 1801
rect 77665 1735 77699 1751
rect 78001 1785 78035 1801
rect 78001 1735 78035 1751
rect 78337 1785 78371 1801
rect 78337 1735 78371 1751
rect 78673 1785 78707 1801
rect 78673 1735 78707 1751
rect 79009 1785 79043 1801
rect 79009 1735 79043 1751
rect 79345 1785 79379 1801
rect 79345 1735 79379 1751
rect 79681 1785 79715 1801
rect 79681 1735 79715 1751
rect 80017 1785 80051 1801
rect 80017 1735 80051 1751
rect 80353 1785 80387 1801
rect 80353 1735 80387 1751
rect 80689 1785 80723 1801
rect 80689 1735 80723 1751
rect 81025 1785 81059 1801
rect 81025 1735 81059 1751
rect 81361 1785 81395 1801
rect 81361 1735 81395 1751
rect 81697 1785 81731 1801
rect 81697 1735 81731 1751
rect 82033 1785 82067 1801
rect 82033 1735 82067 1751
rect 82369 1785 82403 1801
rect 82369 1735 82403 1751
rect 82705 1785 82739 1801
rect 82705 1735 82739 1751
rect 83041 1785 83075 1801
rect 83041 1735 83075 1751
rect 83377 1785 83411 1801
rect 83377 1735 83411 1751
rect 83713 1785 83747 1801
rect 83713 1735 83747 1751
rect 84049 1785 84083 1801
rect 84049 1735 84083 1751
rect 84385 1785 84419 1801
rect 84385 1735 84419 1751
rect 84721 1785 84755 1801
rect 84721 1735 84755 1751
rect 85057 1785 85091 1801
rect 85057 1735 85091 1751
rect 85393 1785 85427 1801
rect 85393 1735 85427 1751
rect 85729 1785 85763 1801
rect 85729 1735 85763 1751
rect 86065 1785 86099 1801
rect 86065 1735 86099 1751
rect 86401 1785 86435 1801
rect 86401 1735 86435 1751
rect 86737 1785 86771 1801
rect 86737 1735 86771 1751
rect 87073 1785 87107 1801
rect 87073 1735 87107 1751
rect 87409 1785 87443 1801
rect 87409 1735 87443 1751
rect 87745 1785 87779 1801
rect 87745 1735 87779 1751
rect 88081 1785 88115 1801
rect 88081 1735 88115 1751
rect 88417 1785 88451 1801
rect 88417 1735 88451 1751
rect 88753 1785 88787 1801
rect 88753 1735 88787 1751
<< viali >>
rect 2065 87479 2099 87513
rect 2401 87479 2435 87513
rect 2737 87479 2771 87513
rect 3073 87479 3107 87513
rect 3409 87479 3443 87513
rect 3745 87479 3779 87513
rect 4081 87479 4115 87513
rect 4417 87479 4451 87513
rect 4753 87479 4787 87513
rect 5089 87479 5123 87513
rect 5425 87479 5459 87513
rect 5761 87479 5795 87513
rect 6097 87479 6131 87513
rect 6433 87479 6467 87513
rect 6769 87479 6803 87513
rect 7105 87479 7139 87513
rect 7441 87479 7475 87513
rect 7777 87479 7811 87513
rect 8113 87479 8147 87513
rect 8449 87479 8483 87513
rect 8785 87479 8819 87513
rect 9121 87479 9155 87513
rect 9457 87479 9491 87513
rect 9793 87479 9827 87513
rect 10129 87479 10163 87513
rect 10465 87479 10499 87513
rect 10801 87479 10835 87513
rect 11137 87479 11171 87513
rect 11473 87479 11507 87513
rect 11809 87479 11843 87513
rect 12145 87479 12179 87513
rect 12481 87479 12515 87513
rect 12817 87479 12851 87513
rect 13153 87479 13187 87513
rect 13489 87479 13523 87513
rect 13825 87479 13859 87513
rect 14161 87479 14195 87513
rect 14497 87479 14531 87513
rect 14833 87479 14867 87513
rect 15169 87479 15203 87513
rect 15505 87479 15539 87513
rect 15841 87479 15875 87513
rect 16177 87479 16211 87513
rect 16513 87479 16547 87513
rect 16849 87479 16883 87513
rect 17185 87479 17219 87513
rect 17521 87479 17555 87513
rect 17857 87479 17891 87513
rect 18193 87479 18227 87513
rect 18529 87479 18563 87513
rect 18865 87479 18899 87513
rect 19201 87479 19235 87513
rect 19537 87479 19571 87513
rect 19873 87479 19907 87513
rect 20209 87479 20243 87513
rect 20545 87479 20579 87513
rect 20881 87479 20915 87513
rect 21217 87479 21251 87513
rect 21553 87479 21587 87513
rect 21889 87479 21923 87513
rect 22225 87479 22259 87513
rect 22561 87479 22595 87513
rect 22897 87479 22931 87513
rect 23233 87479 23267 87513
rect 23569 87479 23603 87513
rect 23905 87479 23939 87513
rect 24241 87479 24275 87513
rect 24577 87479 24611 87513
rect 24913 87479 24947 87513
rect 25249 87479 25283 87513
rect 25585 87479 25619 87513
rect 25921 87479 25955 87513
rect 26257 87479 26291 87513
rect 26593 87479 26627 87513
rect 26929 87479 26963 87513
rect 27265 87479 27299 87513
rect 27601 87479 27635 87513
rect 27937 87479 27971 87513
rect 28273 87479 28307 87513
rect 28609 87479 28643 87513
rect 28945 87479 28979 87513
rect 29281 87479 29315 87513
rect 29617 87479 29651 87513
rect 29953 87479 29987 87513
rect 30289 87479 30323 87513
rect 30625 87479 30659 87513
rect 30961 87479 30995 87513
rect 31297 87479 31331 87513
rect 31633 87479 31667 87513
rect 31969 87479 32003 87513
rect 32305 87479 32339 87513
rect 32641 87479 32675 87513
rect 32977 87479 33011 87513
rect 33313 87479 33347 87513
rect 33649 87479 33683 87513
rect 33985 87479 34019 87513
rect 34321 87479 34355 87513
rect 34657 87479 34691 87513
rect 34993 87479 35027 87513
rect 35329 87479 35363 87513
rect 35665 87479 35699 87513
rect 36001 87479 36035 87513
rect 36337 87479 36371 87513
rect 36673 87479 36707 87513
rect 37009 87479 37043 87513
rect 37345 87479 37379 87513
rect 37681 87479 37715 87513
rect 38017 87479 38051 87513
rect 38353 87479 38387 87513
rect 38689 87479 38723 87513
rect 39025 87479 39059 87513
rect 39361 87479 39395 87513
rect 39697 87479 39731 87513
rect 40033 87479 40067 87513
rect 40369 87479 40403 87513
rect 40705 87479 40739 87513
rect 41041 87479 41075 87513
rect 41377 87479 41411 87513
rect 41713 87479 41747 87513
rect 42049 87479 42083 87513
rect 42385 87479 42419 87513
rect 42721 87479 42755 87513
rect 43057 87479 43091 87513
rect 43393 87479 43427 87513
rect 43729 87479 43763 87513
rect 44065 87479 44099 87513
rect 44401 87479 44435 87513
rect 44737 87479 44771 87513
rect 45073 87479 45107 87513
rect 45409 87479 45443 87513
rect 45745 87479 45779 87513
rect 46081 87479 46115 87513
rect 46417 87479 46451 87513
rect 46753 87479 46787 87513
rect 47089 87479 47123 87513
rect 47425 87479 47459 87513
rect 47761 87479 47795 87513
rect 48097 87479 48131 87513
rect 48433 87479 48467 87513
rect 48769 87479 48803 87513
rect 49105 87479 49139 87513
rect 49441 87479 49475 87513
rect 49777 87479 49811 87513
rect 50113 87479 50147 87513
rect 50449 87479 50483 87513
rect 50785 87479 50819 87513
rect 51121 87479 51155 87513
rect 51457 87479 51491 87513
rect 51793 87479 51827 87513
rect 52129 87479 52163 87513
rect 52465 87479 52499 87513
rect 52801 87479 52835 87513
rect 53137 87479 53171 87513
rect 53473 87479 53507 87513
rect 53809 87479 53843 87513
rect 54145 87479 54179 87513
rect 54481 87479 54515 87513
rect 54817 87479 54851 87513
rect 55153 87479 55187 87513
rect 55489 87479 55523 87513
rect 55825 87479 55859 87513
rect 56161 87479 56195 87513
rect 56497 87479 56531 87513
rect 56833 87479 56867 87513
rect 57169 87479 57203 87513
rect 57505 87479 57539 87513
rect 57841 87479 57875 87513
rect 58177 87479 58211 87513
rect 58513 87479 58547 87513
rect 58849 87479 58883 87513
rect 59185 87479 59219 87513
rect 59521 87479 59555 87513
rect 59857 87479 59891 87513
rect 60193 87479 60227 87513
rect 60529 87479 60563 87513
rect 60865 87479 60899 87513
rect 61201 87479 61235 87513
rect 61537 87479 61571 87513
rect 61873 87479 61907 87513
rect 62209 87479 62243 87513
rect 62545 87479 62579 87513
rect 62881 87479 62915 87513
rect 63217 87479 63251 87513
rect 63553 87479 63587 87513
rect 63889 87479 63923 87513
rect 64225 87479 64259 87513
rect 64561 87479 64595 87513
rect 64897 87479 64931 87513
rect 65233 87479 65267 87513
rect 65569 87479 65603 87513
rect 65905 87479 65939 87513
rect 66241 87479 66275 87513
rect 66577 87479 66611 87513
rect 66913 87479 66947 87513
rect 67249 87479 67283 87513
rect 67585 87479 67619 87513
rect 67921 87479 67955 87513
rect 68257 87479 68291 87513
rect 68593 87479 68627 87513
rect 68929 87479 68963 87513
rect 69265 87479 69299 87513
rect 69601 87479 69635 87513
rect 69937 87479 69971 87513
rect 70273 87479 70307 87513
rect 70609 87479 70643 87513
rect 70945 87479 70979 87513
rect 71281 87479 71315 87513
rect 71617 87479 71651 87513
rect 71953 87479 71987 87513
rect 72289 87479 72323 87513
rect 72625 87479 72659 87513
rect 72961 87479 72995 87513
rect 73297 87479 73331 87513
rect 73633 87479 73667 87513
rect 73969 87479 74003 87513
rect 74305 87479 74339 87513
rect 74641 87479 74675 87513
rect 74977 87479 75011 87513
rect 75313 87479 75347 87513
rect 75649 87479 75683 87513
rect 75985 87479 76019 87513
rect 76321 87479 76355 87513
rect 76657 87479 76691 87513
rect 76993 87479 77027 87513
rect 77329 87479 77363 87513
rect 77665 87479 77699 87513
rect 78001 87479 78035 87513
rect 78337 87479 78371 87513
rect 78673 87479 78707 87513
rect 79009 87479 79043 87513
rect 79345 87479 79379 87513
rect 79681 87479 79715 87513
rect 80017 87479 80051 87513
rect 80353 87479 80387 87513
rect 80689 87479 80723 87513
rect 81025 87479 81059 87513
rect 81361 87479 81395 87513
rect 81697 87479 81731 87513
rect 82033 87479 82067 87513
rect 82369 87479 82403 87513
rect 82705 87479 82739 87513
rect 83041 87479 83075 87513
rect 83377 87479 83411 87513
rect 83713 87479 83747 87513
rect 84049 87479 84083 87513
rect 84385 87479 84419 87513
rect 84721 87479 84755 87513
rect 85057 87479 85091 87513
rect 85393 87479 85427 87513
rect 85729 87479 85763 87513
rect 86065 87479 86099 87513
rect 86401 87479 86435 87513
rect 86737 87479 86771 87513
rect 87073 87479 87107 87513
rect 87409 87479 87443 87513
rect 87745 87479 87779 87513
rect 88081 87479 88115 87513
rect 88417 87479 88451 87513
rect 88753 87479 88787 87513
rect 1729 87095 1763 87129
rect 89227 87095 89261 87129
rect 1729 86759 1763 86793
rect 89227 86759 89261 86793
rect 1729 86423 1763 86457
rect 89227 86423 89261 86457
rect 1729 86087 1763 86121
rect 89227 86087 89261 86121
rect 1729 85751 1763 85785
rect 89227 85751 89261 85785
rect 1729 85415 1763 85449
rect 89227 85415 89261 85449
rect 1729 85079 1763 85113
rect 89227 85079 89261 85113
rect 1729 84743 1763 84777
rect 89227 84743 89261 84777
rect 1729 84407 1763 84441
rect 89227 84407 89261 84441
rect 1729 84071 1763 84105
rect 89227 84071 89261 84105
rect 1729 83735 1763 83769
rect 89227 83735 89261 83769
rect 1729 83399 1763 83433
rect 89227 83399 89261 83433
rect 1729 83063 1763 83097
rect 89227 83063 89261 83097
rect 1729 82727 1763 82761
rect 89227 82727 89261 82761
rect 1729 82391 1763 82425
rect 89227 82391 89261 82425
rect 1729 82055 1763 82089
rect 89227 82055 89261 82089
rect 1729 81719 1763 81753
rect 89227 81719 89261 81753
rect 1729 81383 1763 81417
rect 89227 81383 89261 81417
rect 1729 81047 1763 81081
rect 89227 81047 89261 81081
rect 1729 80711 1763 80745
rect 89227 80711 89261 80745
rect 1729 80375 1763 80409
rect 89227 80375 89261 80409
rect 1729 80039 1763 80073
rect 89227 80039 89261 80073
rect 1729 79703 1763 79737
rect 89227 79703 89261 79737
rect 1729 79367 1763 79401
rect 89227 79367 89261 79401
rect 1729 79031 1763 79065
rect 89227 79031 89261 79065
rect 1729 78695 1763 78729
rect 89227 78695 89261 78729
rect 1729 78359 1763 78393
rect 89227 78359 89261 78393
rect 1729 78023 1763 78057
rect 89227 78023 89261 78057
rect 1729 77687 1763 77721
rect 89227 77687 89261 77721
rect 1729 77351 1763 77385
rect 89227 77351 89261 77385
rect 1729 77015 1763 77049
rect 89227 77015 89261 77049
rect 1729 76679 1763 76713
rect 89227 76679 89261 76713
rect 1729 76343 1763 76377
rect 89227 76343 89261 76377
rect 1729 76007 1763 76041
rect 89227 76007 89261 76041
rect 1729 75671 1763 75705
rect 89227 75671 89261 75705
rect 1729 75335 1763 75369
rect 89227 75335 89261 75369
rect 1729 74999 1763 75033
rect 89227 74999 89261 75033
rect 1729 74663 1763 74697
rect 89227 74663 89261 74697
rect 1729 74327 1763 74361
rect 89227 74327 89261 74361
rect 1729 73991 1763 74025
rect 89227 73991 89261 74025
rect 1729 73655 1763 73689
rect 89227 73655 89261 73689
rect 1729 73319 1763 73353
rect 89227 73319 89261 73353
rect 1729 72983 1763 73017
rect 89227 72983 89261 73017
rect 1729 72647 1763 72681
rect 89227 72647 89261 72681
rect 1729 72311 1763 72345
rect 89227 72311 89261 72345
rect 1729 71975 1763 72009
rect 89227 71975 89261 72009
rect 1729 71639 1763 71673
rect 89227 71639 89261 71673
rect 1729 71303 1763 71337
rect 89227 71303 89261 71337
rect 1729 70967 1763 71001
rect 89227 70967 89261 71001
rect 1729 70631 1763 70665
rect 89227 70631 89261 70665
rect 1729 70295 1763 70329
rect 89227 70295 89261 70329
rect 1729 69959 1763 69993
rect 89227 69959 89261 69993
rect 1729 69623 1763 69657
rect 89227 69623 89261 69657
rect 1729 69287 1763 69321
rect 89227 69287 89261 69321
rect 1729 68951 1763 68985
rect 89227 68951 89261 68985
rect 1729 68615 1763 68649
rect 89227 68615 89261 68649
rect 1729 68279 1763 68313
rect 89227 68279 89261 68313
rect 1729 67943 1763 67977
rect 89227 67943 89261 67977
rect 1729 67607 1763 67641
rect 89227 67607 89261 67641
rect 1729 67271 1763 67305
rect 89227 67271 89261 67305
rect 1729 66935 1763 66969
rect 89227 66935 89261 66969
rect 1729 66599 1763 66633
rect 89227 66599 89261 66633
rect 1729 66263 1763 66297
rect 89227 66263 89261 66297
rect 1729 65927 1763 65961
rect 89227 65927 89261 65961
rect 1729 65591 1763 65625
rect 89227 65591 89261 65625
rect 1729 65255 1763 65289
rect 89227 65255 89261 65289
rect 1729 64919 1763 64953
rect 89227 64919 89261 64953
rect 1729 64583 1763 64617
rect 89227 64583 89261 64617
rect 1729 64247 1763 64281
rect 89227 64247 89261 64281
rect 1729 63911 1763 63945
rect 89227 63911 89261 63945
rect 1729 63575 1763 63609
rect 89227 63575 89261 63609
rect 1729 63239 1763 63273
rect 89227 63239 89261 63273
rect 1729 62903 1763 62937
rect 89227 62903 89261 62937
rect 1729 62567 1763 62601
rect 89227 62567 89261 62601
rect 1729 62231 1763 62265
rect 89227 62231 89261 62265
rect 1729 61895 1763 61929
rect 89227 61895 89261 61929
rect 1729 61559 1763 61593
rect 89227 61559 89261 61593
rect 1729 61223 1763 61257
rect 89227 61223 89261 61257
rect 1729 60887 1763 60921
rect 89227 60887 89261 60921
rect 1729 60551 1763 60585
rect 89227 60551 89261 60585
rect 1729 60215 1763 60249
rect 89227 60215 89261 60249
rect 1729 59879 1763 59913
rect 89227 59879 89261 59913
rect 1729 59543 1763 59577
rect 89227 59543 89261 59577
rect 1729 59207 1763 59241
rect 89227 59207 89261 59241
rect 1729 58871 1763 58905
rect 89227 58871 89261 58905
rect 1729 58535 1763 58569
rect 89227 58535 89261 58569
rect 1729 58199 1763 58233
rect 89227 58199 89261 58233
rect 1729 57863 1763 57897
rect 89227 57863 89261 57897
rect 1729 57527 1763 57561
rect 89227 57527 89261 57561
rect 1729 57191 1763 57225
rect 89227 57191 89261 57225
rect 1729 56855 1763 56889
rect 89227 56855 89261 56889
rect 1729 56519 1763 56553
rect 89227 56519 89261 56553
rect 1729 56183 1763 56217
rect 89227 56183 89261 56217
rect 1729 55847 1763 55881
rect 89227 55847 89261 55881
rect 1729 55511 1763 55545
rect 89227 55511 89261 55545
rect 1729 55175 1763 55209
rect 89227 55175 89261 55209
rect 1729 54839 1763 54873
rect 89227 54839 89261 54873
rect 1729 54503 1763 54537
rect 89227 54503 89261 54537
rect 1729 54167 1763 54201
rect 89227 54167 89261 54201
rect 1729 53831 1763 53865
rect 89227 53831 89261 53865
rect 1729 53495 1763 53529
rect 89227 53495 89261 53529
rect 1729 53159 1763 53193
rect 89227 53159 89261 53193
rect 1729 52823 1763 52857
rect 89227 52823 89261 52857
rect 1729 52487 1763 52521
rect 89227 52487 89261 52521
rect 1729 52151 1763 52185
rect 89227 52151 89261 52185
rect 1729 51815 1763 51849
rect 89227 51815 89261 51849
rect 1729 51479 1763 51513
rect 89227 51479 89261 51513
rect 1729 51143 1763 51177
rect 89227 51143 89261 51177
rect 1729 50807 1763 50841
rect 89227 50807 89261 50841
rect 1729 50471 1763 50505
rect 89227 50471 89261 50505
rect 1729 50135 1763 50169
rect 89227 50135 89261 50169
rect 1729 49799 1763 49833
rect 89227 49799 89261 49833
rect 1729 49463 1763 49497
rect 89227 49463 89261 49497
rect 1729 49127 1763 49161
rect 89227 49127 89261 49161
rect 1729 48791 1763 48825
rect 89227 48791 89261 48825
rect 1729 48455 1763 48489
rect 89227 48455 89261 48489
rect 1729 48119 1763 48153
rect 89227 48119 89261 48153
rect 1729 47783 1763 47817
rect 89227 47783 89261 47817
rect 1729 47447 1763 47481
rect 89227 47447 89261 47481
rect 1729 47111 1763 47145
rect 89227 47111 89261 47145
rect 1729 46775 1763 46809
rect 89227 46775 89261 46809
rect 1729 46439 1763 46473
rect 89227 46439 89261 46473
rect 1729 46103 1763 46137
rect 89227 46103 89261 46137
rect 1729 45767 1763 45801
rect 89227 45767 89261 45801
rect 1729 45431 1763 45465
rect 89227 45431 89261 45465
rect 1729 45095 1763 45129
rect 89227 45095 89261 45129
rect 1729 44759 1763 44793
rect 89227 44759 89261 44793
rect 1729 44423 1763 44457
rect 89227 44423 89261 44457
rect 1729 44087 1763 44121
rect 89227 44087 89261 44121
rect 1729 43751 1763 43785
rect 89227 43751 89261 43785
rect 1729 43415 1763 43449
rect 89227 43415 89261 43449
rect 1729 43079 1763 43113
rect 89227 43079 89261 43113
rect 1729 42743 1763 42777
rect 89227 42743 89261 42777
rect 1729 42407 1763 42441
rect 89227 42407 89261 42441
rect 1729 42071 1763 42105
rect 89227 42071 89261 42105
rect 1729 41735 1763 41769
rect 89227 41735 89261 41769
rect 1729 41399 1763 41433
rect 89227 41399 89261 41433
rect 1729 41063 1763 41097
rect 89227 41063 89261 41097
rect 1729 40727 1763 40761
rect 89227 40727 89261 40761
rect 1729 40391 1763 40425
rect 89227 40391 89261 40425
rect 1729 40055 1763 40089
rect 89227 40055 89261 40089
rect 1729 39719 1763 39753
rect 89227 39719 89261 39753
rect 1729 39383 1763 39417
rect 89227 39383 89261 39417
rect 1729 39047 1763 39081
rect 89227 39047 89261 39081
rect 1729 38711 1763 38745
rect 89227 38711 89261 38745
rect 1729 38375 1763 38409
rect 89227 38375 89261 38409
rect 1729 38039 1763 38073
rect 89227 38039 89261 38073
rect 1729 37703 1763 37737
rect 89227 37703 89261 37737
rect 1729 37367 1763 37401
rect 89227 37367 89261 37401
rect 1729 37031 1763 37065
rect 89227 37031 89261 37065
rect 1729 36695 1763 36729
rect 89227 36695 89261 36729
rect 1729 36359 1763 36393
rect 89227 36359 89261 36393
rect 1729 36023 1763 36057
rect 89227 36023 89261 36057
rect 1729 35687 1763 35721
rect 89227 35687 89261 35721
rect 1729 35351 1763 35385
rect 89227 35351 89261 35385
rect 1729 35015 1763 35049
rect 89227 35015 89261 35049
rect 1729 34679 1763 34713
rect 89227 34679 89261 34713
rect 1729 34343 1763 34377
rect 89227 34343 89261 34377
rect 1729 34007 1763 34041
rect 89227 34007 89261 34041
rect 1729 33671 1763 33705
rect 89227 33671 89261 33705
rect 1729 33335 1763 33369
rect 89227 33335 89261 33369
rect 1729 32999 1763 33033
rect 89227 32999 89261 33033
rect 1729 32663 1763 32697
rect 89227 32663 89261 32697
rect 1729 32327 1763 32361
rect 89227 32327 89261 32361
rect 1729 31991 1763 32025
rect 89227 31991 89261 32025
rect 1729 31655 1763 31689
rect 89227 31655 89261 31689
rect 1729 31319 1763 31353
rect 89227 31319 89261 31353
rect 1729 30983 1763 31017
rect 89227 30983 89261 31017
rect 1729 30647 1763 30681
rect 89227 30647 89261 30681
rect 1729 30311 1763 30345
rect 89227 30311 89261 30345
rect 1729 29975 1763 30009
rect 89227 29975 89261 30009
rect 1729 29639 1763 29673
rect 89227 29639 89261 29673
rect 1729 29303 1763 29337
rect 89227 29303 89261 29337
rect 1729 28967 1763 29001
rect 89227 28967 89261 29001
rect 1729 28631 1763 28665
rect 89227 28631 89261 28665
rect 1729 28295 1763 28329
rect 89227 28295 89261 28329
rect 1729 27959 1763 27993
rect 89227 27959 89261 27993
rect 1729 27623 1763 27657
rect 89227 27623 89261 27657
rect 1729 27287 1763 27321
rect 89227 27287 89261 27321
rect 1729 26951 1763 26985
rect 89227 26951 89261 26985
rect 1729 26615 1763 26649
rect 89227 26615 89261 26649
rect 1729 26279 1763 26313
rect 89227 26279 89261 26313
rect 1729 25943 1763 25977
rect 89227 25943 89261 25977
rect 1729 25607 1763 25641
rect 89227 25607 89261 25641
rect 1729 25271 1763 25305
rect 89227 25271 89261 25305
rect 1729 24935 1763 24969
rect 89227 24935 89261 24969
rect 1729 24599 1763 24633
rect 89227 24599 89261 24633
rect 1729 24263 1763 24297
rect 89227 24263 89261 24297
rect 1729 23927 1763 23961
rect 89227 23927 89261 23961
rect 1729 23591 1763 23625
rect 89227 23591 89261 23625
rect 1729 23255 1763 23289
rect 89227 23255 89261 23289
rect 1729 22919 1763 22953
rect 89227 22919 89261 22953
rect 1729 22583 1763 22617
rect 89227 22583 89261 22617
rect 1729 22247 1763 22281
rect 89227 22247 89261 22281
rect 1729 21911 1763 21945
rect 89227 21911 89261 21945
rect 1729 21575 1763 21609
rect 89227 21575 89261 21609
rect 1729 21239 1763 21273
rect 89227 21239 89261 21273
rect 1729 20903 1763 20937
rect 89227 20903 89261 20937
rect 1729 20567 1763 20601
rect 89227 20567 89261 20601
rect 1729 20231 1763 20265
rect 89227 20231 89261 20265
rect 1729 19895 1763 19929
rect 89227 19895 89261 19929
rect 1729 19559 1763 19593
rect 89227 19559 89261 19593
rect 1729 19223 1763 19257
rect 89227 19223 89261 19257
rect 1729 18887 1763 18921
rect 89227 18887 89261 18921
rect 1729 18551 1763 18585
rect 89227 18551 89261 18585
rect 1729 18215 1763 18249
rect 89227 18215 89261 18249
rect 1729 17879 1763 17913
rect 89227 17879 89261 17913
rect 1729 17543 1763 17577
rect 89227 17543 89261 17577
rect 1729 17207 1763 17241
rect 89227 17207 89261 17241
rect 1729 16871 1763 16905
rect 89227 16871 89261 16905
rect 1729 16535 1763 16569
rect 89227 16535 89261 16569
rect 1729 16199 1763 16233
rect 89227 16199 89261 16233
rect 1729 15863 1763 15897
rect 89227 15863 89261 15897
rect 1729 15527 1763 15561
rect 89227 15527 89261 15561
rect 1729 15191 1763 15225
rect 89227 15191 89261 15225
rect 1729 14855 1763 14889
rect 89227 14855 89261 14889
rect 1729 14519 1763 14553
rect 89227 14519 89261 14553
rect 1729 14183 1763 14217
rect 89227 14183 89261 14217
rect 1729 13847 1763 13881
rect 89227 13847 89261 13881
rect 1729 13511 1763 13545
rect 89227 13511 89261 13545
rect 1729 13175 1763 13209
rect 89227 13175 89261 13209
rect 1729 12839 1763 12873
rect 89227 12839 89261 12873
rect 1729 12503 1763 12537
rect 89227 12503 89261 12537
rect 1729 12167 1763 12201
rect 89227 12167 89261 12201
rect 1729 11831 1763 11865
rect 89227 11831 89261 11865
rect 1729 11495 1763 11529
rect 89227 11495 89261 11529
rect 1729 11159 1763 11193
rect 89227 11159 89261 11193
rect 1729 10823 1763 10857
rect 89227 10823 89261 10857
rect 1729 10487 1763 10521
rect 89227 10487 89261 10521
rect 1729 10151 1763 10185
rect 89227 10151 89261 10185
rect 1729 9815 1763 9849
rect 89227 9815 89261 9849
rect 1729 9479 1763 9513
rect 89227 9479 89261 9513
rect 1729 9143 1763 9177
rect 89227 9143 89261 9177
rect 1729 8807 1763 8841
rect 89227 8807 89261 8841
rect 1729 8471 1763 8505
rect 89227 8471 89261 8505
rect 1729 8135 1763 8169
rect 89227 8135 89261 8169
rect 1729 7799 1763 7833
rect 89227 7799 89261 7833
rect 1729 7463 1763 7497
rect 89227 7463 89261 7497
rect 1729 7127 1763 7161
rect 89227 7127 89261 7161
rect 1729 6791 1763 6825
rect 89227 6791 89261 6825
rect 1729 6455 1763 6489
rect 89227 6455 89261 6489
rect 1729 6119 1763 6153
rect 89227 6119 89261 6153
rect 1729 5783 1763 5817
rect 89227 5783 89261 5817
rect 1729 5447 1763 5481
rect 89227 5447 89261 5481
rect 1729 5111 1763 5145
rect 89227 5111 89261 5145
rect 1729 4775 1763 4809
rect 89227 4775 89261 4809
rect 1729 4439 1763 4473
rect 89227 4439 89261 4473
rect 1729 4103 1763 4137
rect 89227 4103 89261 4137
rect 1729 3767 1763 3801
rect 89227 3767 89261 3801
rect 1729 3431 1763 3465
rect 89227 3431 89261 3465
rect 1729 3095 1763 3129
rect 89227 3095 89261 3129
rect 1729 2759 1763 2793
rect 89227 2759 89261 2793
rect 1729 2423 1763 2457
rect 89227 2423 89261 2457
rect 1729 2087 1763 2121
rect 89227 2087 89261 2121
rect 2065 1751 2099 1785
rect 2401 1751 2435 1785
rect 2737 1751 2771 1785
rect 3073 1751 3107 1785
rect 3409 1751 3443 1785
rect 3745 1751 3779 1785
rect 4081 1751 4115 1785
rect 4417 1751 4451 1785
rect 4753 1751 4787 1785
rect 5089 1751 5123 1785
rect 5425 1751 5459 1785
rect 5761 1751 5795 1785
rect 6097 1751 6131 1785
rect 6433 1751 6467 1785
rect 6769 1751 6803 1785
rect 7105 1751 7139 1785
rect 7441 1751 7475 1785
rect 7777 1751 7811 1785
rect 8113 1751 8147 1785
rect 8449 1751 8483 1785
rect 8785 1751 8819 1785
rect 9121 1751 9155 1785
rect 9457 1751 9491 1785
rect 9793 1751 9827 1785
rect 10129 1751 10163 1785
rect 10465 1751 10499 1785
rect 10801 1751 10835 1785
rect 11137 1751 11171 1785
rect 11473 1751 11507 1785
rect 11809 1751 11843 1785
rect 12145 1751 12179 1785
rect 12481 1751 12515 1785
rect 12817 1751 12851 1785
rect 13153 1751 13187 1785
rect 13489 1751 13523 1785
rect 13825 1751 13859 1785
rect 14161 1751 14195 1785
rect 14497 1751 14531 1785
rect 14833 1751 14867 1785
rect 15169 1751 15203 1785
rect 15505 1751 15539 1785
rect 15841 1751 15875 1785
rect 16177 1751 16211 1785
rect 16513 1751 16547 1785
rect 16849 1751 16883 1785
rect 17185 1751 17219 1785
rect 17521 1751 17555 1785
rect 17857 1751 17891 1785
rect 18193 1751 18227 1785
rect 18529 1751 18563 1785
rect 18865 1751 18899 1785
rect 19201 1751 19235 1785
rect 19537 1751 19571 1785
rect 19873 1751 19907 1785
rect 20209 1751 20243 1785
rect 20545 1751 20579 1785
rect 20881 1751 20915 1785
rect 21217 1751 21251 1785
rect 21553 1751 21587 1785
rect 21889 1751 21923 1785
rect 22225 1751 22259 1785
rect 22561 1751 22595 1785
rect 22897 1751 22931 1785
rect 23233 1751 23267 1785
rect 23569 1751 23603 1785
rect 23905 1751 23939 1785
rect 24241 1751 24275 1785
rect 24577 1751 24611 1785
rect 24913 1751 24947 1785
rect 25249 1751 25283 1785
rect 25585 1751 25619 1785
rect 25921 1751 25955 1785
rect 26257 1751 26291 1785
rect 26593 1751 26627 1785
rect 26929 1751 26963 1785
rect 27265 1751 27299 1785
rect 27601 1751 27635 1785
rect 27937 1751 27971 1785
rect 28273 1751 28307 1785
rect 28609 1751 28643 1785
rect 28945 1751 28979 1785
rect 29281 1751 29315 1785
rect 29617 1751 29651 1785
rect 29953 1751 29987 1785
rect 30289 1751 30323 1785
rect 30625 1751 30659 1785
rect 30961 1751 30995 1785
rect 31297 1751 31331 1785
rect 31633 1751 31667 1785
rect 31969 1751 32003 1785
rect 32305 1751 32339 1785
rect 32641 1751 32675 1785
rect 32977 1751 33011 1785
rect 33313 1751 33347 1785
rect 33649 1751 33683 1785
rect 33985 1751 34019 1785
rect 34321 1751 34355 1785
rect 34657 1751 34691 1785
rect 34993 1751 35027 1785
rect 35329 1751 35363 1785
rect 35665 1751 35699 1785
rect 36001 1751 36035 1785
rect 36337 1751 36371 1785
rect 36673 1751 36707 1785
rect 37009 1751 37043 1785
rect 37345 1751 37379 1785
rect 37681 1751 37715 1785
rect 38017 1751 38051 1785
rect 38353 1751 38387 1785
rect 38689 1751 38723 1785
rect 39025 1751 39059 1785
rect 39361 1751 39395 1785
rect 39697 1751 39731 1785
rect 40033 1751 40067 1785
rect 40369 1751 40403 1785
rect 40705 1751 40739 1785
rect 41041 1751 41075 1785
rect 41377 1751 41411 1785
rect 41713 1751 41747 1785
rect 42049 1751 42083 1785
rect 42385 1751 42419 1785
rect 42721 1751 42755 1785
rect 43057 1751 43091 1785
rect 43393 1751 43427 1785
rect 43729 1751 43763 1785
rect 44065 1751 44099 1785
rect 44401 1751 44435 1785
rect 44737 1751 44771 1785
rect 45073 1751 45107 1785
rect 45409 1751 45443 1785
rect 45745 1751 45779 1785
rect 46081 1751 46115 1785
rect 46417 1751 46451 1785
rect 46753 1751 46787 1785
rect 47089 1751 47123 1785
rect 47425 1751 47459 1785
rect 47761 1751 47795 1785
rect 48097 1751 48131 1785
rect 48433 1751 48467 1785
rect 48769 1751 48803 1785
rect 49105 1751 49139 1785
rect 49441 1751 49475 1785
rect 49777 1751 49811 1785
rect 50113 1751 50147 1785
rect 50449 1751 50483 1785
rect 50785 1751 50819 1785
rect 51121 1751 51155 1785
rect 51457 1751 51491 1785
rect 51793 1751 51827 1785
rect 52129 1751 52163 1785
rect 52465 1751 52499 1785
rect 52801 1751 52835 1785
rect 53137 1751 53171 1785
rect 53473 1751 53507 1785
rect 53809 1751 53843 1785
rect 54145 1751 54179 1785
rect 54481 1751 54515 1785
rect 54817 1751 54851 1785
rect 55153 1751 55187 1785
rect 55489 1751 55523 1785
rect 55825 1751 55859 1785
rect 56161 1751 56195 1785
rect 56497 1751 56531 1785
rect 56833 1751 56867 1785
rect 57169 1751 57203 1785
rect 57505 1751 57539 1785
rect 57841 1751 57875 1785
rect 58177 1751 58211 1785
rect 58513 1751 58547 1785
rect 58849 1751 58883 1785
rect 59185 1751 59219 1785
rect 59521 1751 59555 1785
rect 59857 1751 59891 1785
rect 60193 1751 60227 1785
rect 60529 1751 60563 1785
rect 60865 1751 60899 1785
rect 61201 1751 61235 1785
rect 61537 1751 61571 1785
rect 61873 1751 61907 1785
rect 62209 1751 62243 1785
rect 62545 1751 62579 1785
rect 62881 1751 62915 1785
rect 63217 1751 63251 1785
rect 63553 1751 63587 1785
rect 63889 1751 63923 1785
rect 64225 1751 64259 1785
rect 64561 1751 64595 1785
rect 64897 1751 64931 1785
rect 65233 1751 65267 1785
rect 65569 1751 65603 1785
rect 65905 1751 65939 1785
rect 66241 1751 66275 1785
rect 66577 1751 66611 1785
rect 66913 1751 66947 1785
rect 67249 1751 67283 1785
rect 67585 1751 67619 1785
rect 67921 1751 67955 1785
rect 68257 1751 68291 1785
rect 68593 1751 68627 1785
rect 68929 1751 68963 1785
rect 69265 1751 69299 1785
rect 69601 1751 69635 1785
rect 69937 1751 69971 1785
rect 70273 1751 70307 1785
rect 70609 1751 70643 1785
rect 70945 1751 70979 1785
rect 71281 1751 71315 1785
rect 71617 1751 71651 1785
rect 71953 1751 71987 1785
rect 72289 1751 72323 1785
rect 72625 1751 72659 1785
rect 72961 1751 72995 1785
rect 73297 1751 73331 1785
rect 73633 1751 73667 1785
rect 73969 1751 74003 1785
rect 74305 1751 74339 1785
rect 74641 1751 74675 1785
rect 74977 1751 75011 1785
rect 75313 1751 75347 1785
rect 75649 1751 75683 1785
rect 75985 1751 76019 1785
rect 76321 1751 76355 1785
rect 76657 1751 76691 1785
rect 76993 1751 77027 1785
rect 77329 1751 77363 1785
rect 77665 1751 77699 1785
rect 78001 1751 78035 1785
rect 78337 1751 78371 1785
rect 78673 1751 78707 1785
rect 79009 1751 79043 1785
rect 79345 1751 79379 1785
rect 79681 1751 79715 1785
rect 80017 1751 80051 1785
rect 80353 1751 80387 1785
rect 80689 1751 80723 1785
rect 81025 1751 81059 1785
rect 81361 1751 81395 1785
rect 81697 1751 81731 1785
rect 82033 1751 82067 1785
rect 82369 1751 82403 1785
rect 82705 1751 82739 1785
rect 83041 1751 83075 1785
rect 83377 1751 83411 1785
rect 83713 1751 83747 1785
rect 84049 1751 84083 1785
rect 84385 1751 84419 1785
rect 84721 1751 84755 1785
rect 85057 1751 85091 1785
rect 85393 1751 85427 1785
rect 85729 1751 85763 1785
rect 86065 1751 86099 1785
rect 86401 1751 86435 1785
rect 86737 1751 86771 1785
rect 87073 1751 87107 1785
rect 87409 1751 87443 1785
rect 87745 1751 87779 1785
rect 88081 1751 88115 1785
rect 88417 1751 88451 1785
rect 88753 1751 88787 1785
<< metal1 >>
rect 1634 87522 89356 87608
rect 1634 87470 2056 87522
rect 2108 87513 3736 87522
rect 3788 87513 5416 87522
rect 5468 87513 7096 87522
rect 7148 87513 8776 87522
rect 8828 87513 10456 87522
rect 10508 87513 12136 87522
rect 12188 87513 13816 87522
rect 13868 87513 15496 87522
rect 15548 87513 17176 87522
rect 17228 87513 18856 87522
rect 18908 87513 20536 87522
rect 20588 87513 22216 87522
rect 22268 87513 23896 87522
rect 23948 87513 25576 87522
rect 25628 87513 27256 87522
rect 27308 87513 28936 87522
rect 28988 87513 30616 87522
rect 30668 87513 32296 87522
rect 32348 87513 33976 87522
rect 34028 87513 35656 87522
rect 35708 87513 37336 87522
rect 37388 87513 39016 87522
rect 39068 87513 40696 87522
rect 40748 87513 42376 87522
rect 42428 87513 44056 87522
rect 44108 87513 45736 87522
rect 45788 87513 47416 87522
rect 47468 87513 49096 87522
rect 49148 87513 50776 87522
rect 50828 87513 52456 87522
rect 52508 87513 54136 87522
rect 54188 87513 55816 87522
rect 55868 87513 57496 87522
rect 57548 87513 59176 87522
rect 59228 87513 60856 87522
rect 60908 87513 62536 87522
rect 62588 87513 64216 87522
rect 64268 87513 65896 87522
rect 65948 87513 67576 87522
rect 67628 87513 69256 87522
rect 69308 87513 70936 87522
rect 70988 87513 72616 87522
rect 72668 87513 74296 87522
rect 74348 87513 75976 87522
rect 76028 87513 77656 87522
rect 77708 87513 79336 87522
rect 79388 87513 81016 87522
rect 81068 87513 82696 87522
rect 82748 87513 84376 87522
rect 84428 87513 86056 87522
rect 86108 87513 87736 87522
rect 87788 87513 89356 87522
rect 2108 87479 2401 87513
rect 2435 87479 2737 87513
rect 2771 87479 3073 87513
rect 3107 87479 3409 87513
rect 3443 87479 3736 87513
rect 3788 87479 4081 87513
rect 4115 87479 4417 87513
rect 4451 87479 4753 87513
rect 4787 87479 5089 87513
rect 5123 87479 5416 87513
rect 5468 87479 5761 87513
rect 5795 87479 6097 87513
rect 6131 87479 6433 87513
rect 6467 87479 6769 87513
rect 6803 87479 7096 87513
rect 7148 87479 7441 87513
rect 7475 87479 7777 87513
rect 7811 87479 8113 87513
rect 8147 87479 8449 87513
rect 8483 87479 8776 87513
rect 8828 87479 9121 87513
rect 9155 87479 9457 87513
rect 9491 87479 9793 87513
rect 9827 87479 10129 87513
rect 10163 87479 10456 87513
rect 10508 87479 10801 87513
rect 10835 87479 11137 87513
rect 11171 87479 11473 87513
rect 11507 87479 11809 87513
rect 11843 87479 12136 87513
rect 12188 87479 12481 87513
rect 12515 87479 12817 87513
rect 12851 87479 13153 87513
rect 13187 87479 13489 87513
rect 13523 87479 13816 87513
rect 13868 87479 14161 87513
rect 14195 87479 14497 87513
rect 14531 87479 14833 87513
rect 14867 87479 15169 87513
rect 15203 87479 15496 87513
rect 15548 87479 15841 87513
rect 15875 87479 16177 87513
rect 16211 87479 16513 87513
rect 16547 87479 16849 87513
rect 16883 87479 17176 87513
rect 17228 87479 17521 87513
rect 17555 87479 17857 87513
rect 17891 87479 18193 87513
rect 18227 87479 18529 87513
rect 18563 87479 18856 87513
rect 18908 87479 19201 87513
rect 19235 87479 19537 87513
rect 19571 87479 19873 87513
rect 19907 87479 20209 87513
rect 20243 87479 20536 87513
rect 20588 87479 20881 87513
rect 20915 87479 21217 87513
rect 21251 87479 21553 87513
rect 21587 87479 21889 87513
rect 21923 87479 22216 87513
rect 22268 87479 22561 87513
rect 22595 87479 22897 87513
rect 22931 87479 23233 87513
rect 23267 87479 23569 87513
rect 23603 87479 23896 87513
rect 23948 87479 24241 87513
rect 24275 87479 24577 87513
rect 24611 87479 24913 87513
rect 24947 87479 25249 87513
rect 25283 87479 25576 87513
rect 25628 87479 25921 87513
rect 25955 87479 26257 87513
rect 26291 87479 26593 87513
rect 26627 87479 26929 87513
rect 26963 87479 27256 87513
rect 27308 87479 27601 87513
rect 27635 87479 27937 87513
rect 27971 87479 28273 87513
rect 28307 87479 28609 87513
rect 28643 87479 28936 87513
rect 28988 87479 29281 87513
rect 29315 87479 29617 87513
rect 29651 87479 29953 87513
rect 29987 87479 30289 87513
rect 30323 87479 30616 87513
rect 30668 87479 30961 87513
rect 30995 87479 31297 87513
rect 31331 87479 31633 87513
rect 31667 87479 31969 87513
rect 32003 87479 32296 87513
rect 32348 87479 32641 87513
rect 32675 87479 32977 87513
rect 33011 87479 33313 87513
rect 33347 87479 33649 87513
rect 33683 87479 33976 87513
rect 34028 87479 34321 87513
rect 34355 87479 34657 87513
rect 34691 87479 34993 87513
rect 35027 87479 35329 87513
rect 35363 87479 35656 87513
rect 35708 87479 36001 87513
rect 36035 87479 36337 87513
rect 36371 87479 36673 87513
rect 36707 87479 37009 87513
rect 37043 87479 37336 87513
rect 37388 87479 37681 87513
rect 37715 87479 38017 87513
rect 38051 87479 38353 87513
rect 38387 87479 38689 87513
rect 38723 87479 39016 87513
rect 39068 87479 39361 87513
rect 39395 87479 39697 87513
rect 39731 87479 40033 87513
rect 40067 87479 40369 87513
rect 40403 87479 40696 87513
rect 40748 87479 41041 87513
rect 41075 87479 41377 87513
rect 41411 87479 41713 87513
rect 41747 87479 42049 87513
rect 42083 87479 42376 87513
rect 42428 87479 42721 87513
rect 42755 87479 43057 87513
rect 43091 87479 43393 87513
rect 43427 87479 43729 87513
rect 43763 87479 44056 87513
rect 44108 87479 44401 87513
rect 44435 87479 44737 87513
rect 44771 87479 45073 87513
rect 45107 87479 45409 87513
rect 45443 87479 45736 87513
rect 45788 87479 46081 87513
rect 46115 87479 46417 87513
rect 46451 87479 46753 87513
rect 46787 87479 47089 87513
rect 47123 87479 47416 87513
rect 47468 87479 47761 87513
rect 47795 87479 48097 87513
rect 48131 87479 48433 87513
rect 48467 87479 48769 87513
rect 48803 87479 49096 87513
rect 49148 87479 49441 87513
rect 49475 87479 49777 87513
rect 49811 87479 50113 87513
rect 50147 87479 50449 87513
rect 50483 87479 50776 87513
rect 50828 87479 51121 87513
rect 51155 87479 51457 87513
rect 51491 87479 51793 87513
rect 51827 87479 52129 87513
rect 52163 87479 52456 87513
rect 52508 87479 52801 87513
rect 52835 87479 53137 87513
rect 53171 87479 53473 87513
rect 53507 87479 53809 87513
rect 53843 87479 54136 87513
rect 54188 87479 54481 87513
rect 54515 87479 54817 87513
rect 54851 87479 55153 87513
rect 55187 87479 55489 87513
rect 55523 87479 55816 87513
rect 55868 87479 56161 87513
rect 56195 87479 56497 87513
rect 56531 87479 56833 87513
rect 56867 87479 57169 87513
rect 57203 87479 57496 87513
rect 57548 87479 57841 87513
rect 57875 87479 58177 87513
rect 58211 87479 58513 87513
rect 58547 87479 58849 87513
rect 58883 87479 59176 87513
rect 59228 87479 59521 87513
rect 59555 87479 59857 87513
rect 59891 87479 60193 87513
rect 60227 87479 60529 87513
rect 60563 87479 60856 87513
rect 60908 87479 61201 87513
rect 61235 87479 61537 87513
rect 61571 87479 61873 87513
rect 61907 87479 62209 87513
rect 62243 87479 62536 87513
rect 62588 87479 62881 87513
rect 62915 87479 63217 87513
rect 63251 87479 63553 87513
rect 63587 87479 63889 87513
rect 63923 87479 64216 87513
rect 64268 87479 64561 87513
rect 64595 87479 64897 87513
rect 64931 87479 65233 87513
rect 65267 87479 65569 87513
rect 65603 87479 65896 87513
rect 65948 87479 66241 87513
rect 66275 87479 66577 87513
rect 66611 87479 66913 87513
rect 66947 87479 67249 87513
rect 67283 87479 67576 87513
rect 67628 87479 67921 87513
rect 67955 87479 68257 87513
rect 68291 87479 68593 87513
rect 68627 87479 68929 87513
rect 68963 87479 69256 87513
rect 69308 87479 69601 87513
rect 69635 87479 69937 87513
rect 69971 87479 70273 87513
rect 70307 87479 70609 87513
rect 70643 87479 70936 87513
rect 70988 87479 71281 87513
rect 71315 87479 71617 87513
rect 71651 87479 71953 87513
rect 71987 87479 72289 87513
rect 72323 87479 72616 87513
rect 72668 87479 72961 87513
rect 72995 87479 73297 87513
rect 73331 87479 73633 87513
rect 73667 87479 73969 87513
rect 74003 87479 74296 87513
rect 74348 87479 74641 87513
rect 74675 87479 74977 87513
rect 75011 87479 75313 87513
rect 75347 87479 75649 87513
rect 75683 87479 75976 87513
rect 76028 87479 76321 87513
rect 76355 87479 76657 87513
rect 76691 87479 76993 87513
rect 77027 87479 77329 87513
rect 77363 87479 77656 87513
rect 77708 87479 78001 87513
rect 78035 87479 78337 87513
rect 78371 87479 78673 87513
rect 78707 87479 79009 87513
rect 79043 87479 79336 87513
rect 79388 87479 79681 87513
rect 79715 87479 80017 87513
rect 80051 87479 80353 87513
rect 80387 87479 80689 87513
rect 80723 87479 81016 87513
rect 81068 87479 81361 87513
rect 81395 87479 81697 87513
rect 81731 87479 82033 87513
rect 82067 87479 82369 87513
rect 82403 87479 82696 87513
rect 82748 87479 83041 87513
rect 83075 87479 83377 87513
rect 83411 87479 83713 87513
rect 83747 87479 84049 87513
rect 84083 87479 84376 87513
rect 84428 87479 84721 87513
rect 84755 87479 85057 87513
rect 85091 87479 85393 87513
rect 85427 87479 85729 87513
rect 85763 87479 86056 87513
rect 86108 87479 86401 87513
rect 86435 87479 86737 87513
rect 86771 87479 87073 87513
rect 87107 87479 87409 87513
rect 87443 87479 87736 87513
rect 87788 87479 88081 87513
rect 88115 87479 88417 87513
rect 88451 87479 88753 87513
rect 88787 87479 89356 87513
rect 2108 87470 3736 87479
rect 3788 87470 5416 87479
rect 5468 87470 7096 87479
rect 7148 87470 8776 87479
rect 8828 87470 10456 87479
rect 10508 87470 12136 87479
rect 12188 87470 13816 87479
rect 13868 87470 15496 87479
rect 15548 87470 17176 87479
rect 17228 87470 18856 87479
rect 18908 87470 20536 87479
rect 20588 87470 22216 87479
rect 22268 87470 23896 87479
rect 23948 87470 25576 87479
rect 25628 87470 27256 87479
rect 27308 87470 28936 87479
rect 28988 87470 30616 87479
rect 30668 87470 32296 87479
rect 32348 87470 33976 87479
rect 34028 87470 35656 87479
rect 35708 87470 37336 87479
rect 37388 87470 39016 87479
rect 39068 87470 40696 87479
rect 40748 87470 42376 87479
rect 42428 87470 44056 87479
rect 44108 87470 45736 87479
rect 45788 87470 47416 87479
rect 47468 87470 49096 87479
rect 49148 87470 50776 87479
rect 50828 87470 52456 87479
rect 52508 87470 54136 87479
rect 54188 87470 55816 87479
rect 55868 87470 57496 87479
rect 57548 87470 59176 87479
rect 59228 87470 60856 87479
rect 60908 87470 62536 87479
rect 62588 87470 64216 87479
rect 64268 87470 65896 87479
rect 65948 87470 67576 87479
rect 67628 87470 69256 87479
rect 69308 87470 70936 87479
rect 70988 87470 72616 87479
rect 72668 87470 74296 87479
rect 74348 87470 75976 87479
rect 76028 87470 77656 87479
rect 77708 87470 79336 87479
rect 79388 87470 81016 87479
rect 81068 87470 82696 87479
rect 82748 87470 84376 87479
rect 84428 87470 86056 87479
rect 86108 87470 87736 87479
rect 87788 87470 89356 87479
rect 1634 87384 89356 87470
rect 1714 87086 1720 87138
rect 1772 87086 1778 87138
rect 89212 87086 89218 87138
rect 89270 87086 89276 87138
rect 1714 86750 1720 86802
rect 1772 86750 1778 86802
rect 89212 86750 89218 86802
rect 89270 86750 89276 86802
rect 1714 86414 1720 86466
rect 1772 86414 1778 86466
rect 89212 86414 89218 86466
rect 89270 86414 89276 86466
rect 1714 86078 1720 86130
rect 1772 86078 1778 86130
rect 89212 86078 89218 86130
rect 89270 86078 89276 86130
rect 1714 85742 1720 85794
rect 1772 85742 1778 85794
rect 89212 85742 89218 85794
rect 89270 85742 89276 85794
rect 1714 85406 1720 85458
rect 1772 85406 1778 85458
rect 89212 85406 89218 85458
rect 89270 85406 89276 85458
rect 1714 85070 1720 85122
rect 1772 85070 1778 85122
rect 89212 85070 89218 85122
rect 89270 85070 89276 85122
rect 1714 84734 1720 84786
rect 1772 84734 1778 84786
rect 89212 84734 89218 84786
rect 89270 84734 89276 84786
rect 1714 84398 1720 84450
rect 1772 84398 1778 84450
rect 89212 84398 89218 84450
rect 89270 84398 89276 84450
rect 1714 84062 1720 84114
rect 1772 84062 1778 84114
rect 89212 84062 89218 84114
rect 89270 84062 89276 84114
rect 1714 83726 1720 83778
rect 1772 83726 1778 83778
rect 89212 83726 89218 83778
rect 89270 83726 89276 83778
rect 1714 83390 1720 83442
rect 1772 83390 1778 83442
rect 89212 83390 89218 83442
rect 89270 83390 89276 83442
rect 1714 83054 1720 83106
rect 1772 83054 1778 83106
rect 89212 83054 89218 83106
rect 89270 83054 89276 83106
rect 1714 82718 1720 82770
rect 1772 82718 1778 82770
rect 89212 82718 89218 82770
rect 89270 82718 89276 82770
rect 1714 82382 1720 82434
rect 1772 82382 1778 82434
rect 89212 82382 89218 82434
rect 89270 82382 89276 82434
rect 1714 82046 1720 82098
rect 1772 82046 1778 82098
rect 89212 82046 89218 82098
rect 89270 82046 89276 82098
rect 1714 81710 1720 81762
rect 1772 81710 1778 81762
rect 89212 81710 89218 81762
rect 89270 81710 89276 81762
rect 1714 81374 1720 81426
rect 1772 81374 1778 81426
rect 89212 81374 89218 81426
rect 89270 81374 89276 81426
rect 1714 81038 1720 81090
rect 1772 81038 1778 81090
rect 89212 81038 89218 81090
rect 89270 81038 89276 81090
rect 1714 80702 1720 80754
rect 1772 80702 1778 80754
rect 89212 80702 89218 80754
rect 89270 80702 89276 80754
rect 1714 80366 1720 80418
rect 1772 80366 1778 80418
rect 89212 80366 89218 80418
rect 89270 80366 89276 80418
rect 1714 80030 1720 80082
rect 1772 80030 1778 80082
rect 89212 80030 89218 80082
rect 89270 80030 89276 80082
rect 1714 79694 1720 79746
rect 1772 79694 1778 79746
rect 89212 79694 89218 79746
rect 89270 79694 89276 79746
rect 1714 79358 1720 79410
rect 1772 79358 1778 79410
rect 89212 79358 89218 79410
rect 89270 79358 89276 79410
rect 1714 79022 1720 79074
rect 1772 79022 1778 79074
rect 89212 79022 89218 79074
rect 89270 79022 89276 79074
rect 1714 78686 1720 78738
rect 1772 78686 1778 78738
rect 89212 78686 89218 78738
rect 89270 78686 89276 78738
rect 1714 78350 1720 78402
rect 1772 78350 1778 78402
rect 89212 78350 89218 78402
rect 89270 78350 89276 78402
rect 1714 78014 1720 78066
rect 1772 78014 1778 78066
rect 89212 78014 89218 78066
rect 89270 78014 89276 78066
rect 25622 77856 25628 77908
rect 25680 77856 25686 77908
rect 30614 77856 30620 77908
rect 30672 77856 30678 77908
rect 35606 77856 35612 77908
rect 35664 77856 35670 77908
rect 40598 77856 40604 77908
rect 40656 77856 40662 77908
rect 45590 77856 45596 77908
rect 45648 77856 45654 77908
rect 50582 77856 50588 77908
rect 50640 77856 50646 77908
rect 55574 77856 55580 77908
rect 55632 77856 55638 77908
rect 60566 77856 60572 77908
rect 60624 77856 60630 77908
rect 1714 77678 1720 77730
rect 1772 77678 1778 77730
rect 89212 77678 89218 77730
rect 89270 77678 89276 77730
rect 1714 77342 1720 77394
rect 1772 77342 1778 77394
rect 89212 77342 89218 77394
rect 89270 77342 89276 77394
rect 1714 77006 1720 77058
rect 1772 77006 1778 77058
rect 89212 77006 89218 77058
rect 89270 77006 89276 77058
rect 1714 76670 1720 76722
rect 1772 76670 1778 76722
rect 89212 76670 89218 76722
rect 89270 76670 89276 76722
rect 1714 76334 1720 76386
rect 1772 76334 1778 76386
rect 89212 76334 89218 76386
rect 89270 76334 89276 76386
rect 1714 75998 1720 76050
rect 1772 75998 1778 76050
rect 89212 75998 89218 76050
rect 89270 75998 89276 76050
rect 1714 75662 1720 75714
rect 1772 75662 1778 75714
rect 89212 75662 89218 75714
rect 89270 75662 89276 75714
rect 1714 75326 1720 75378
rect 1772 75326 1778 75378
rect 89212 75326 89218 75378
rect 89270 75326 89276 75378
rect 1714 74990 1720 75042
rect 1772 74990 1778 75042
rect 89212 74990 89218 75042
rect 89270 74990 89276 75042
rect 1714 74654 1720 74706
rect 1772 74654 1778 74706
rect 89212 74654 89218 74706
rect 89270 74654 89276 74706
rect 1714 74318 1720 74370
rect 1772 74318 1778 74370
rect 89212 74318 89218 74370
rect 89270 74318 89276 74370
rect 1714 73982 1720 74034
rect 1772 73982 1778 74034
rect 89212 73982 89218 74034
rect 89270 73982 89276 74034
rect 1714 73646 1720 73698
rect 1772 73646 1778 73698
rect 89212 73646 89218 73698
rect 89270 73646 89276 73698
rect 1714 73310 1720 73362
rect 1772 73310 1778 73362
rect 89212 73310 89218 73362
rect 89270 73310 89276 73362
rect 1714 72974 1720 73026
rect 1772 72974 1778 73026
rect 89212 72974 89218 73026
rect 89270 72974 89276 73026
rect 1714 72638 1720 72690
rect 1772 72638 1778 72690
rect 89212 72638 89218 72690
rect 89270 72638 89276 72690
rect 1714 72302 1720 72354
rect 1772 72302 1778 72354
rect 89212 72302 89218 72354
rect 89270 72302 89276 72354
rect 1714 71966 1720 72018
rect 1772 71966 1778 72018
rect 89212 71966 89218 72018
rect 89270 71966 89276 72018
rect 1714 71630 1720 71682
rect 1772 71630 1778 71682
rect 89212 71630 89218 71682
rect 89270 71630 89276 71682
rect 1714 71294 1720 71346
rect 1772 71294 1778 71346
rect 89212 71294 89218 71346
rect 89270 71294 89276 71346
rect 1714 70958 1720 71010
rect 1772 70958 1778 71010
rect 89212 70958 89218 71010
rect 89270 70958 89276 71010
rect 1714 70622 1720 70674
rect 1772 70622 1778 70674
rect 89212 70622 89218 70674
rect 89270 70622 89276 70674
rect 1714 70286 1720 70338
rect 1772 70286 1778 70338
rect 89212 70286 89218 70338
rect 89270 70286 89276 70338
rect 1714 69950 1720 70002
rect 1772 69950 1778 70002
rect 89212 69950 89218 70002
rect 89270 69950 89276 70002
rect 1714 69614 1720 69666
rect 1772 69614 1778 69666
rect 89212 69614 89218 69666
rect 89270 69614 89276 69666
rect 1714 69278 1720 69330
rect 1772 69278 1778 69330
rect 89212 69278 89218 69330
rect 89270 69278 89276 69330
rect 1714 68942 1720 68994
rect 1772 68942 1778 68994
rect 89212 68942 89218 68994
rect 89270 68942 89276 68994
rect 1714 68606 1720 68658
rect 1772 68606 1778 68658
rect 89212 68606 89218 68658
rect 89270 68606 89276 68658
rect 1714 68270 1720 68322
rect 1772 68270 1778 68322
rect 89212 68270 89218 68322
rect 89270 68270 89276 68322
rect 1714 67934 1720 67986
rect 1772 67934 1778 67986
rect 89212 67934 89218 67986
rect 89270 67934 89276 67986
rect 1714 67598 1720 67650
rect 1772 67598 1778 67650
rect 89212 67598 89218 67650
rect 89270 67598 89276 67650
rect 1714 67262 1720 67314
rect 1772 67262 1778 67314
rect 89212 67262 89218 67314
rect 89270 67262 89276 67314
rect 1714 66926 1720 66978
rect 1772 66926 1778 66978
rect 89212 66926 89218 66978
rect 89270 66926 89276 66978
rect 1714 66590 1720 66642
rect 1772 66590 1778 66642
rect 89212 66590 89218 66642
rect 89270 66590 89276 66642
rect 1714 66254 1720 66306
rect 1772 66254 1778 66306
rect 89212 66254 89218 66306
rect 89270 66254 89276 66306
rect 1714 65918 1720 65970
rect 1772 65918 1778 65970
rect 89212 65918 89218 65970
rect 89270 65918 89276 65970
rect 1714 65582 1720 65634
rect 1772 65582 1778 65634
rect 89212 65582 89218 65634
rect 89270 65582 89276 65634
rect 1714 65246 1720 65298
rect 1772 65246 1778 65298
rect 89212 65246 89218 65298
rect 89270 65246 89276 65298
rect 1714 64910 1720 64962
rect 1772 64910 1778 64962
rect 89212 64910 89218 64962
rect 89270 64910 89276 64962
rect 1714 64574 1720 64626
rect 1772 64574 1778 64626
rect 89212 64574 89218 64626
rect 89270 64574 89276 64626
rect 1714 64238 1720 64290
rect 1772 64238 1778 64290
rect 89212 64238 89218 64290
rect 89270 64238 89276 64290
rect 1714 63902 1720 63954
rect 1772 63902 1778 63954
rect 89212 63902 89218 63954
rect 89270 63902 89276 63954
rect 1714 63566 1720 63618
rect 1772 63566 1778 63618
rect 89212 63566 89218 63618
rect 89270 63566 89276 63618
rect 1714 63230 1720 63282
rect 1772 63230 1778 63282
rect 89212 63230 89218 63282
rect 89270 63230 89276 63282
rect 1714 62894 1720 62946
rect 1772 62894 1778 62946
rect 89212 62894 89218 62946
rect 89270 62894 89276 62946
rect 1714 62558 1720 62610
rect 1772 62558 1778 62610
rect 89212 62558 89218 62610
rect 89270 62558 89276 62610
rect 1714 62222 1720 62274
rect 1772 62222 1778 62274
rect 89212 62222 89218 62274
rect 89270 62222 89276 62274
rect 1714 61886 1720 61938
rect 1772 61886 1778 61938
rect 89212 61886 89218 61938
rect 89270 61886 89276 61938
rect 1714 61550 1720 61602
rect 1772 61550 1778 61602
rect 89212 61550 89218 61602
rect 89270 61550 89276 61602
rect 1714 61214 1720 61266
rect 1772 61214 1778 61266
rect 89212 61214 89218 61266
rect 89270 61214 89276 61266
rect 1714 60878 1720 60930
rect 1772 60878 1778 60930
rect 89212 60878 89218 60930
rect 89270 60878 89276 60930
rect 1714 60542 1720 60594
rect 1772 60542 1778 60594
rect 89212 60542 89218 60594
rect 89270 60542 89276 60594
rect 1714 60206 1720 60258
rect 1772 60206 1778 60258
rect 89212 60206 89218 60258
rect 89270 60206 89276 60258
rect 1714 59870 1720 59922
rect 1772 59870 1778 59922
rect 89212 59870 89218 59922
rect 89270 59870 89276 59922
rect 1714 59534 1720 59586
rect 1772 59534 1778 59586
rect 89212 59534 89218 59586
rect 89270 59534 89276 59586
rect 1714 59198 1720 59250
rect 1772 59198 1778 59250
rect 89212 59198 89218 59250
rect 89270 59198 89276 59250
rect 1714 58862 1720 58914
rect 1772 58862 1778 58914
rect 89212 58862 89218 58914
rect 89270 58862 89276 58914
rect 1714 58526 1720 58578
rect 1772 58526 1778 58578
rect 89212 58526 89218 58578
rect 89270 58526 89276 58578
rect 1714 58190 1720 58242
rect 1772 58190 1778 58242
rect 89212 58190 89218 58242
rect 89270 58190 89276 58242
rect 1714 57854 1720 57906
rect 1772 57854 1778 57906
rect 89212 57854 89218 57906
rect 89270 57854 89276 57906
rect 1714 57518 1720 57570
rect 1772 57518 1778 57570
rect 89212 57518 89218 57570
rect 89270 57518 89276 57570
rect 1714 57182 1720 57234
rect 1772 57182 1778 57234
rect 89212 57182 89218 57234
rect 89270 57182 89276 57234
rect 1714 56846 1720 56898
rect 1772 56846 1778 56898
rect 89212 56846 89218 56898
rect 89270 56846 89276 56898
rect 1714 56510 1720 56562
rect 1772 56510 1778 56562
rect 89212 56510 89218 56562
rect 89270 56510 89276 56562
rect 1714 56174 1720 56226
rect 1772 56174 1778 56226
rect 89212 56174 89218 56226
rect 89270 56174 89276 56226
rect 1714 55838 1720 55890
rect 1772 55838 1778 55890
rect 89212 55838 89218 55890
rect 89270 55838 89276 55890
rect 1714 55502 1720 55554
rect 1772 55502 1778 55554
rect 89212 55502 89218 55554
rect 89270 55502 89276 55554
rect 1714 55166 1720 55218
rect 1772 55166 1778 55218
rect 89212 55166 89218 55218
rect 89270 55166 89276 55218
rect 1714 54830 1720 54882
rect 1772 54830 1778 54882
rect 89212 54830 89218 54882
rect 89270 54830 89276 54882
rect 1714 54494 1720 54546
rect 1772 54494 1778 54546
rect 89212 54494 89218 54546
rect 89270 54494 89276 54546
rect 1714 54158 1720 54210
rect 1772 54158 1778 54210
rect 89212 54158 89218 54210
rect 89270 54158 89276 54210
rect 1714 53822 1720 53874
rect 1772 53822 1778 53874
rect 89212 53822 89218 53874
rect 89270 53822 89276 53874
rect 1714 53486 1720 53538
rect 1772 53486 1778 53538
rect 89212 53486 89218 53538
rect 89270 53486 89276 53538
rect 1714 53150 1720 53202
rect 1772 53150 1778 53202
rect 89212 53150 89218 53202
rect 89270 53150 89276 53202
rect 1714 52814 1720 52866
rect 1772 52814 1778 52866
rect 89212 52814 89218 52866
rect 89270 52814 89276 52866
rect 1714 52478 1720 52530
rect 1772 52478 1778 52530
rect 89212 52478 89218 52530
rect 89270 52478 89276 52530
rect 1714 52142 1720 52194
rect 1772 52142 1778 52194
rect 89212 52142 89218 52194
rect 89270 52142 89276 52194
rect 1714 51806 1720 51858
rect 1772 51806 1778 51858
rect 89212 51806 89218 51858
rect 89270 51806 89276 51858
rect 1714 51470 1720 51522
rect 1772 51470 1778 51522
rect 89212 51470 89218 51522
rect 89270 51470 89276 51522
rect 1714 51134 1720 51186
rect 1772 51134 1778 51186
rect 89212 51134 89218 51186
rect 89270 51134 89276 51186
rect 1714 50798 1720 50850
rect 1772 50798 1778 50850
rect 89212 50798 89218 50850
rect 89270 50798 89276 50850
rect 1714 50462 1720 50514
rect 1772 50462 1778 50514
rect 89212 50462 89218 50514
rect 89270 50462 89276 50514
rect 1714 50126 1720 50178
rect 1772 50126 1778 50178
rect 89212 50126 89218 50178
rect 89270 50126 89276 50178
rect 1714 49790 1720 49842
rect 1772 49790 1778 49842
rect 89212 49790 89218 49842
rect 89270 49790 89276 49842
rect 1714 49454 1720 49506
rect 1772 49454 1778 49506
rect 89212 49454 89218 49506
rect 89270 49454 89276 49506
rect 1714 49118 1720 49170
rect 1772 49118 1778 49170
rect 89212 49118 89218 49170
rect 89270 49118 89276 49170
rect 1714 48782 1720 48834
rect 1772 48782 1778 48834
rect 89212 48782 89218 48834
rect 89270 48782 89276 48834
rect 1714 48446 1720 48498
rect 1772 48446 1778 48498
rect 89212 48446 89218 48498
rect 89270 48446 89276 48498
rect 1714 48110 1720 48162
rect 1772 48110 1778 48162
rect 89212 48110 89218 48162
rect 89270 48110 89276 48162
rect 1714 47774 1720 47826
rect 1772 47774 1778 47826
rect 89212 47774 89218 47826
rect 89270 47774 89276 47826
rect 1714 47438 1720 47490
rect 1772 47438 1778 47490
rect 89212 47438 89218 47490
rect 89270 47438 89276 47490
rect 1714 47102 1720 47154
rect 1772 47102 1778 47154
rect 89212 47102 89218 47154
rect 89270 47102 89276 47154
rect 1714 46766 1720 46818
rect 1772 46766 1778 46818
rect 89212 46766 89218 46818
rect 89270 46766 89276 46818
rect 1714 46430 1720 46482
rect 1772 46430 1778 46482
rect 89212 46430 89218 46482
rect 89270 46430 89276 46482
rect 1714 46094 1720 46146
rect 1772 46094 1778 46146
rect 89212 46094 89218 46146
rect 89270 46094 89276 46146
rect 1714 45758 1720 45810
rect 1772 45758 1778 45810
rect 89212 45758 89218 45810
rect 89270 45758 89276 45810
rect 1714 45422 1720 45474
rect 1772 45422 1778 45474
rect 89212 45422 89218 45474
rect 89270 45422 89276 45474
rect 1714 45086 1720 45138
rect 1772 45086 1778 45138
rect 89212 45086 89218 45138
rect 89270 45086 89276 45138
rect 1714 44750 1720 44802
rect 1772 44750 1778 44802
rect 89212 44750 89218 44802
rect 89270 44750 89276 44802
rect 1714 44414 1720 44466
rect 1772 44414 1778 44466
rect 89212 44414 89218 44466
rect 89270 44414 89276 44466
rect 1714 44078 1720 44130
rect 1772 44078 1778 44130
rect 89212 44078 89218 44130
rect 89270 44078 89276 44130
rect 1714 43742 1720 43794
rect 1772 43742 1778 43794
rect 89212 43742 89218 43794
rect 89270 43742 89276 43794
rect 1714 43406 1720 43458
rect 1772 43406 1778 43458
rect 89212 43406 89218 43458
rect 89270 43406 89276 43458
rect 1714 43070 1720 43122
rect 1772 43070 1778 43122
rect 89212 43070 89218 43122
rect 89270 43070 89276 43122
rect 1714 42734 1720 42786
rect 1772 42734 1778 42786
rect 89212 42734 89218 42786
rect 89270 42734 89276 42786
rect 1714 42398 1720 42450
rect 1772 42398 1778 42450
rect 89212 42398 89218 42450
rect 89270 42398 89276 42450
rect 1714 42062 1720 42114
rect 1772 42062 1778 42114
rect 89212 42062 89218 42114
rect 89270 42062 89276 42114
rect 1714 41726 1720 41778
rect 1772 41726 1778 41778
rect 89212 41726 89218 41778
rect 89270 41726 89276 41778
rect 1714 41390 1720 41442
rect 1772 41390 1778 41442
rect 89212 41390 89218 41442
rect 89270 41390 89276 41442
rect 1714 41054 1720 41106
rect 1772 41054 1778 41106
rect 89212 41054 89218 41106
rect 89270 41054 89276 41106
rect 1714 40718 1720 40770
rect 1772 40718 1778 40770
rect 89212 40718 89218 40770
rect 89270 40718 89276 40770
rect 1714 40382 1720 40434
rect 1772 40382 1778 40434
rect 89212 40382 89218 40434
rect 89270 40382 89276 40434
rect 1714 40046 1720 40098
rect 1772 40046 1778 40098
rect 89212 40046 89218 40098
rect 89270 40046 89276 40098
rect 1714 39710 1720 39762
rect 1772 39710 1778 39762
rect 89212 39710 89218 39762
rect 89270 39710 89276 39762
rect 1714 39374 1720 39426
rect 1772 39374 1778 39426
rect 89212 39374 89218 39426
rect 89270 39374 89276 39426
rect 1714 39038 1720 39090
rect 1772 39038 1778 39090
rect 89212 39038 89218 39090
rect 89270 39038 89276 39090
rect 1714 38702 1720 38754
rect 1772 38702 1778 38754
rect 89212 38702 89218 38754
rect 89270 38702 89276 38754
rect 1714 38366 1720 38418
rect 1772 38366 1778 38418
rect 89212 38366 89218 38418
rect 89270 38366 89276 38418
rect 1714 38030 1720 38082
rect 1772 38030 1778 38082
rect 89212 38030 89218 38082
rect 89270 38030 89276 38082
rect 1714 37694 1720 37746
rect 1772 37694 1778 37746
rect 89212 37694 89218 37746
rect 89270 37694 89276 37746
rect 1714 37358 1720 37410
rect 1772 37358 1778 37410
rect 89212 37358 89218 37410
rect 89270 37358 89276 37410
rect 12351 37206 12357 37258
rect 12409 37206 12415 37258
rect 1714 37022 1720 37074
rect 1772 37022 1778 37074
rect 1714 36686 1720 36738
rect 1772 36686 1778 36738
rect 1714 36350 1720 36402
rect 1772 36350 1778 36402
rect 1714 36014 1720 36066
rect 1772 36014 1778 36066
rect 12271 35936 12277 35988
rect 12329 35936 12335 35988
rect 1714 35678 1720 35730
rect 1772 35678 1778 35730
rect 1714 35342 1720 35394
rect 1772 35342 1778 35394
rect 1714 35006 1720 35058
rect 1772 35006 1778 35058
rect 1714 34670 1720 34722
rect 1772 34670 1778 34722
rect 1714 34334 1720 34386
rect 1772 34334 1778 34386
rect 12191 34378 12197 34430
rect 12249 34378 12255 34430
rect 1714 33998 1720 34050
rect 1772 33998 1778 34050
rect 1714 33662 1720 33714
rect 1772 33662 1778 33714
rect 1714 33326 1720 33378
rect 1772 33326 1778 33378
rect 12111 33108 12117 33160
rect 12169 33108 12175 33160
rect 1714 32990 1720 33042
rect 1772 32990 1778 33042
rect 1714 32654 1720 32706
rect 1772 32654 1778 32706
rect 1714 32318 1720 32370
rect 1772 32318 1778 32370
rect 1714 31982 1720 32034
rect 1772 31982 1778 32034
rect 1714 31646 1720 31698
rect 1772 31646 1778 31698
rect 12031 31550 12037 31602
rect 12089 31550 12095 31602
rect 1714 31310 1720 31362
rect 1772 31310 1778 31362
rect 1714 30974 1720 31026
rect 1772 30974 1778 31026
rect 1714 30638 1720 30690
rect 1772 30638 1778 30690
rect 1714 30302 1720 30354
rect 1772 30302 1778 30354
rect 11951 30280 11957 30332
rect 12009 30280 12015 30332
rect 1714 29966 1720 30018
rect 1772 29966 1778 30018
rect 1714 29630 1720 29682
rect 1772 29630 1778 29682
rect 1714 29294 1720 29346
rect 1772 29294 1778 29346
rect 1714 28958 1720 29010
rect 1772 28958 1778 29010
rect 11871 28722 11877 28774
rect 11929 28722 11935 28774
rect 1714 28622 1720 28674
rect 1772 28622 1778 28674
rect 1714 28286 1720 28338
rect 1772 28286 1778 28338
rect 1714 27950 1720 28002
rect 1772 27950 1778 28002
rect 1714 27614 1720 27666
rect 1772 27614 1778 27666
rect 1714 27278 1720 27330
rect 1772 27278 1778 27330
rect 1714 26942 1720 26994
rect 1772 26942 1778 26994
rect 1714 26606 1720 26658
rect 1772 26606 1778 26658
rect 1714 26270 1720 26322
rect 1772 26270 1778 26322
rect 1714 25934 1720 25986
rect 1772 25934 1778 25986
rect 1714 25598 1720 25650
rect 1772 25598 1778 25650
rect 1714 25262 1720 25314
rect 1772 25262 1778 25314
rect 1714 24926 1720 24978
rect 1772 24926 1778 24978
rect 1714 24590 1720 24642
rect 1772 24590 1778 24642
rect 1714 24254 1720 24306
rect 1772 24254 1778 24306
rect 11889 24163 11917 28722
rect 11969 24163 11997 30280
rect 12049 24163 12077 31550
rect 12129 24163 12157 33108
rect 12209 24163 12237 34378
rect 12289 24163 12317 35936
rect 12369 24163 12397 37206
rect 89212 37022 89218 37074
rect 89270 37022 89276 37074
rect 89212 36686 89218 36738
rect 89270 36686 89276 36738
rect 89212 36350 89218 36402
rect 89270 36350 89276 36402
rect 89212 36014 89218 36066
rect 89270 36014 89276 36066
rect 89212 35678 89218 35730
rect 89270 35678 89276 35730
rect 89212 35342 89218 35394
rect 89270 35342 89276 35394
rect 89212 35006 89218 35058
rect 89270 35006 89276 35058
rect 89212 34670 89218 34722
rect 89270 34670 89276 34722
rect 89212 34334 89218 34386
rect 89270 34334 89276 34386
rect 89212 33998 89218 34050
rect 89270 33998 89276 34050
rect 89212 33662 89218 33714
rect 89270 33662 89276 33714
rect 89212 33326 89218 33378
rect 89270 33326 89276 33378
rect 89212 32990 89218 33042
rect 89270 32990 89276 33042
rect 89212 32654 89218 32706
rect 89270 32654 89276 32706
rect 89212 32318 89218 32370
rect 89270 32318 89276 32370
rect 89212 31982 89218 32034
rect 89270 31982 89276 32034
rect 89212 31646 89218 31698
rect 89270 31646 89276 31698
rect 89212 31310 89218 31362
rect 89270 31310 89276 31362
rect 89212 30974 89218 31026
rect 89270 30974 89276 31026
rect 89212 30638 89218 30690
rect 89270 30638 89276 30690
rect 89212 30302 89218 30354
rect 89270 30302 89276 30354
rect 89212 29966 89218 30018
rect 89270 29966 89276 30018
rect 89212 29630 89218 29682
rect 89270 29630 89276 29682
rect 89212 29294 89218 29346
rect 89270 29294 89276 29346
rect 89212 28958 89218 29010
rect 89270 28958 89276 29010
rect 89212 28622 89218 28674
rect 89270 28622 89276 28674
rect 89212 28286 89218 28338
rect 89270 28286 89276 28338
rect 89212 27950 89218 28002
rect 89270 27950 89276 28002
rect 89212 27614 89218 27666
rect 89270 27614 89276 27666
rect 89212 27278 89218 27330
rect 89270 27278 89276 27330
rect 89212 26942 89218 26994
rect 89270 26942 89276 26994
rect 89212 26606 89218 26658
rect 89270 26606 89276 26658
rect 89212 26270 89218 26322
rect 89270 26270 89276 26322
rect 89212 25934 89218 25986
rect 89270 25934 89276 25986
rect 89212 25598 89218 25650
rect 89270 25598 89276 25650
rect 89212 25262 89218 25314
rect 89270 25262 89276 25314
rect 89212 24926 89218 24978
rect 89270 24926 89276 24978
rect 89212 24590 89218 24642
rect 89270 24590 89276 24642
rect 89212 24254 89218 24306
rect 89270 24254 89276 24306
rect 1714 23918 1720 23970
rect 1772 23918 1778 23970
rect 1714 23582 1720 23634
rect 1772 23582 1778 23634
rect 1714 23246 1720 23298
rect 1772 23246 1778 23298
rect 1714 22910 1720 22962
rect 1772 22910 1778 22962
rect 1714 22574 1720 22626
rect 1772 22574 1778 22626
rect 1714 22238 1720 22290
rect 1772 22238 1778 22290
rect 1714 21902 1720 21954
rect 1772 21902 1778 21954
rect 1714 21566 1720 21618
rect 1772 21566 1778 21618
rect 1714 21230 1720 21282
rect 1772 21230 1778 21282
rect 1714 20894 1720 20946
rect 1772 20894 1778 20946
rect 1714 20558 1720 20610
rect 1772 20558 1778 20610
rect 1714 20222 1720 20274
rect 1772 20222 1778 20274
rect 1714 19886 1720 19938
rect 1772 19886 1778 19938
rect 1714 19550 1720 19602
rect 1772 19550 1778 19602
rect 1714 19214 1720 19266
rect 1772 19214 1778 19266
rect 1714 18878 1720 18930
rect 1772 18878 1778 18930
rect 1714 18542 1720 18594
rect 1772 18542 1778 18594
rect 1714 18206 1720 18258
rect 1772 18206 1778 18258
rect 1714 17870 1720 17922
rect 1772 17870 1778 17922
rect 1714 17534 1720 17586
rect 1772 17534 1778 17586
rect 1714 17198 1720 17250
rect 1772 17198 1778 17250
rect 1714 16862 1720 16914
rect 1772 16862 1778 16914
rect 1714 16526 1720 16578
rect 1772 16526 1778 16578
rect 1714 16190 1720 16242
rect 1772 16190 1778 16242
rect 1714 15854 1720 15906
rect 1772 15854 1778 15906
rect 1714 15518 1720 15570
rect 1772 15518 1778 15570
rect 1714 15182 1720 15234
rect 1772 15182 1778 15234
rect 1714 14846 1720 14898
rect 1772 14846 1778 14898
rect 1714 14510 1720 14562
rect 1772 14510 1778 14562
rect 1714 14174 1720 14226
rect 1772 14174 1778 14226
rect 1714 13838 1720 13890
rect 1772 13838 1778 13890
rect 1714 13502 1720 13554
rect 1772 13502 1778 13554
rect 1714 13166 1720 13218
rect 1772 13166 1778 13218
rect 25622 13078 25628 13130
rect 25680 13078 25686 13130
rect 30614 13078 30620 13130
rect 30672 13078 30678 13130
rect 35606 13078 35612 13130
rect 35664 13078 35670 13130
rect 40598 13078 40604 13130
rect 40656 13078 40662 13130
rect 45590 13078 45596 13130
rect 45648 13078 45654 13130
rect 50582 13078 50588 13130
rect 50640 13078 50646 13130
rect 55574 13078 55580 13130
rect 55632 13078 55638 13130
rect 60566 13078 60572 13130
rect 60624 13078 60630 13130
rect 1714 12830 1720 12882
rect 1772 12830 1778 12882
rect 1714 12494 1720 12546
rect 1772 12494 1778 12546
rect 1714 12158 1720 12210
rect 1772 12158 1778 12210
rect 1714 11822 1720 11874
rect 1772 11822 1778 11874
rect 1714 11486 1720 11538
rect 1772 11486 1778 11538
rect 1714 11150 1720 11202
rect 1772 11150 1778 11202
rect 78593 11120 78621 24163
rect 78673 12390 78701 24163
rect 78753 13948 78781 24163
rect 78833 15218 78861 24163
rect 78913 16776 78941 24163
rect 78993 18046 79021 24163
rect 79073 19604 79101 24163
rect 89212 23918 89218 23970
rect 89270 23918 89276 23970
rect 89212 23582 89218 23634
rect 89270 23582 89276 23634
rect 89212 23246 89218 23298
rect 89270 23246 89276 23298
rect 89212 22910 89218 22962
rect 89270 22910 89276 22962
rect 89212 22574 89218 22626
rect 89270 22574 89276 22626
rect 89212 22238 89218 22290
rect 89270 22238 89276 22290
rect 89212 21902 89218 21954
rect 89270 21902 89276 21954
rect 89212 21566 89218 21618
rect 89270 21566 89276 21618
rect 89212 21230 89218 21282
rect 89270 21230 89276 21282
rect 89212 20894 89218 20946
rect 89270 20894 89276 20946
rect 89212 20558 89218 20610
rect 89270 20558 89276 20610
rect 89212 20222 89218 20274
rect 89270 20222 89276 20274
rect 89212 19886 89218 19938
rect 89270 19886 89276 19938
rect 79055 19552 79061 19604
rect 79113 19552 79119 19604
rect 89212 19550 89218 19602
rect 89270 19550 89276 19602
rect 89212 19214 89218 19266
rect 89270 19214 89276 19266
rect 89212 18878 89218 18930
rect 89270 18878 89276 18930
rect 89212 18542 89218 18594
rect 89270 18542 89276 18594
rect 89212 18206 89218 18258
rect 89270 18206 89276 18258
rect 78975 17994 78981 18046
rect 79033 17994 79039 18046
rect 89212 17870 89218 17922
rect 89270 17870 89276 17922
rect 89212 17534 89218 17586
rect 89270 17534 89276 17586
rect 89212 17198 89218 17250
rect 89270 17198 89276 17250
rect 89212 16862 89218 16914
rect 89270 16862 89276 16914
rect 78895 16724 78901 16776
rect 78953 16724 78959 16776
rect 89212 16526 89218 16578
rect 89270 16526 89276 16578
rect 89212 16190 89218 16242
rect 89270 16190 89276 16242
rect 89212 15854 89218 15906
rect 89270 15854 89276 15906
rect 89212 15518 89218 15570
rect 89270 15518 89276 15570
rect 78815 15166 78821 15218
rect 78873 15166 78879 15218
rect 89212 15182 89218 15234
rect 89270 15182 89276 15234
rect 89212 14846 89218 14898
rect 89270 14846 89276 14898
rect 89212 14510 89218 14562
rect 89270 14510 89276 14562
rect 89212 14174 89218 14226
rect 89270 14174 89276 14226
rect 78735 13896 78741 13948
rect 78793 13896 78799 13948
rect 89212 13838 89218 13890
rect 89270 13838 89276 13890
rect 89212 13502 89218 13554
rect 89270 13502 89276 13554
rect 89212 13166 89218 13218
rect 89270 13166 89276 13218
rect 89212 12830 89218 12882
rect 89270 12830 89276 12882
rect 89212 12494 89218 12546
rect 89270 12494 89276 12546
rect 78655 12338 78661 12390
rect 78713 12338 78719 12390
rect 89212 12158 89218 12210
rect 89270 12158 89276 12210
rect 89212 11822 89218 11874
rect 89270 11822 89276 11874
rect 89212 11486 89218 11538
rect 89270 11486 89276 11538
rect 89212 11150 89218 11202
rect 89270 11150 89276 11202
rect 78575 11068 78581 11120
rect 78633 11068 78639 11120
rect 1714 10814 1720 10866
rect 1772 10814 1778 10866
rect 89212 10814 89218 10866
rect 89270 10814 89276 10866
rect 1714 10478 1720 10530
rect 1772 10478 1778 10530
rect 89212 10478 89218 10530
rect 89270 10478 89276 10530
rect 1714 10142 1720 10194
rect 1772 10142 1778 10194
rect 89212 10142 89218 10194
rect 89270 10142 89276 10194
rect 1714 9806 1720 9858
rect 1772 9806 1778 9858
rect 89212 9806 89218 9858
rect 89270 9806 89276 9858
rect 1714 9470 1720 9522
rect 1772 9470 1778 9522
rect 89212 9470 89218 9522
rect 89270 9470 89276 9522
rect 1714 9134 1720 9186
rect 1772 9134 1778 9186
rect 89212 9134 89218 9186
rect 89270 9134 89276 9186
rect 1714 8798 1720 8850
rect 1772 8798 1778 8850
rect 89212 8798 89218 8850
rect 89270 8798 89276 8850
rect 1714 8462 1720 8514
rect 1772 8462 1778 8514
rect 89212 8462 89218 8514
rect 89270 8462 89276 8514
rect 1714 8126 1720 8178
rect 1772 8126 1778 8178
rect 89212 8126 89218 8178
rect 89270 8126 89276 8178
rect 1714 7790 1720 7842
rect 1772 7790 1778 7842
rect 89212 7790 89218 7842
rect 89270 7790 89276 7842
rect 1714 7454 1720 7506
rect 1772 7454 1778 7506
rect 89212 7454 89218 7506
rect 89270 7454 89276 7506
rect 1714 7118 1720 7170
rect 1772 7118 1778 7170
rect 89212 7118 89218 7170
rect 89270 7118 89276 7170
rect 1714 6782 1720 6834
rect 1772 6782 1778 6834
rect 89212 6782 89218 6834
rect 89270 6782 89276 6834
rect 1714 6446 1720 6498
rect 1772 6446 1778 6498
rect 89212 6446 89218 6498
rect 89270 6446 89276 6498
rect 1714 6110 1720 6162
rect 1772 6110 1778 6162
rect 89212 6110 89218 6162
rect 89270 6110 89276 6162
rect 1714 5774 1720 5826
rect 1772 5774 1778 5826
rect 89212 5774 89218 5826
rect 89270 5774 89276 5826
rect 1714 5438 1720 5490
rect 1772 5438 1778 5490
rect 89212 5438 89218 5490
rect 89270 5438 89276 5490
rect 1714 5102 1720 5154
rect 1772 5102 1778 5154
rect 89212 5102 89218 5154
rect 89270 5102 89276 5154
rect 1714 4766 1720 4818
rect 1772 4766 1778 4818
rect 89212 4766 89218 4818
rect 89270 4766 89276 4818
rect 1714 4430 1720 4482
rect 1772 4430 1778 4482
rect 89212 4430 89218 4482
rect 89270 4430 89276 4482
rect 1714 4094 1720 4146
rect 1772 4094 1778 4146
rect 89212 4094 89218 4146
rect 89270 4094 89276 4146
rect 1714 3758 1720 3810
rect 1772 3758 1778 3810
rect 89212 3758 89218 3810
rect 89270 3758 89276 3810
rect 1714 3422 1720 3474
rect 1772 3422 1778 3474
rect 89212 3422 89218 3474
rect 89270 3422 89276 3474
rect 1714 3086 1720 3138
rect 1772 3086 1778 3138
rect 89212 3086 89218 3138
rect 89270 3086 89276 3138
rect 1714 2750 1720 2802
rect 1772 2750 1778 2802
rect 89212 2750 89218 2802
rect 89270 2750 89276 2802
rect 1714 2414 1720 2466
rect 1772 2414 1778 2466
rect 89212 2414 89218 2466
rect 89270 2414 89276 2466
rect 1714 2078 1720 2130
rect 1772 2078 1778 2130
rect 89212 2078 89218 2130
rect 89270 2078 89276 2130
rect 1634 1794 89356 1880
rect 1634 1742 2056 1794
rect 2108 1785 3736 1794
rect 3788 1785 5416 1794
rect 5468 1785 7096 1794
rect 7148 1785 8776 1794
rect 8828 1785 10456 1794
rect 10508 1785 12136 1794
rect 12188 1785 13816 1794
rect 13868 1785 15496 1794
rect 15548 1785 17176 1794
rect 17228 1785 18856 1794
rect 18908 1785 20536 1794
rect 20588 1785 22216 1794
rect 22268 1785 23896 1794
rect 23948 1785 25576 1794
rect 25628 1785 27256 1794
rect 27308 1785 28936 1794
rect 28988 1785 30616 1794
rect 30668 1785 32296 1794
rect 32348 1785 33976 1794
rect 34028 1785 35656 1794
rect 35708 1785 37336 1794
rect 37388 1785 39016 1794
rect 39068 1785 40696 1794
rect 40748 1785 42376 1794
rect 42428 1785 44056 1794
rect 44108 1785 45736 1794
rect 45788 1785 47416 1794
rect 47468 1785 49096 1794
rect 49148 1785 50776 1794
rect 50828 1785 52456 1794
rect 52508 1785 54136 1794
rect 54188 1785 55816 1794
rect 55868 1785 57496 1794
rect 57548 1785 59176 1794
rect 59228 1785 60856 1794
rect 60908 1785 62536 1794
rect 62588 1785 64216 1794
rect 64268 1785 65896 1794
rect 65948 1785 67576 1794
rect 67628 1785 69256 1794
rect 69308 1785 70936 1794
rect 70988 1785 72616 1794
rect 72668 1785 74296 1794
rect 74348 1785 75976 1794
rect 76028 1785 77656 1794
rect 77708 1785 79336 1794
rect 79388 1785 81016 1794
rect 81068 1785 82696 1794
rect 82748 1785 84376 1794
rect 84428 1785 86056 1794
rect 86108 1785 87736 1794
rect 87788 1785 89356 1794
rect 2108 1751 2401 1785
rect 2435 1751 2737 1785
rect 2771 1751 3073 1785
rect 3107 1751 3409 1785
rect 3443 1751 3736 1785
rect 3788 1751 4081 1785
rect 4115 1751 4417 1785
rect 4451 1751 4753 1785
rect 4787 1751 5089 1785
rect 5123 1751 5416 1785
rect 5468 1751 5761 1785
rect 5795 1751 6097 1785
rect 6131 1751 6433 1785
rect 6467 1751 6769 1785
rect 6803 1751 7096 1785
rect 7148 1751 7441 1785
rect 7475 1751 7777 1785
rect 7811 1751 8113 1785
rect 8147 1751 8449 1785
rect 8483 1751 8776 1785
rect 8828 1751 9121 1785
rect 9155 1751 9457 1785
rect 9491 1751 9793 1785
rect 9827 1751 10129 1785
rect 10163 1751 10456 1785
rect 10508 1751 10801 1785
rect 10835 1751 11137 1785
rect 11171 1751 11473 1785
rect 11507 1751 11809 1785
rect 11843 1751 12136 1785
rect 12188 1751 12481 1785
rect 12515 1751 12817 1785
rect 12851 1751 13153 1785
rect 13187 1751 13489 1785
rect 13523 1751 13816 1785
rect 13868 1751 14161 1785
rect 14195 1751 14497 1785
rect 14531 1751 14833 1785
rect 14867 1751 15169 1785
rect 15203 1751 15496 1785
rect 15548 1751 15841 1785
rect 15875 1751 16177 1785
rect 16211 1751 16513 1785
rect 16547 1751 16849 1785
rect 16883 1751 17176 1785
rect 17228 1751 17521 1785
rect 17555 1751 17857 1785
rect 17891 1751 18193 1785
rect 18227 1751 18529 1785
rect 18563 1751 18856 1785
rect 18908 1751 19201 1785
rect 19235 1751 19537 1785
rect 19571 1751 19873 1785
rect 19907 1751 20209 1785
rect 20243 1751 20536 1785
rect 20588 1751 20881 1785
rect 20915 1751 21217 1785
rect 21251 1751 21553 1785
rect 21587 1751 21889 1785
rect 21923 1751 22216 1785
rect 22268 1751 22561 1785
rect 22595 1751 22897 1785
rect 22931 1751 23233 1785
rect 23267 1751 23569 1785
rect 23603 1751 23896 1785
rect 23948 1751 24241 1785
rect 24275 1751 24577 1785
rect 24611 1751 24913 1785
rect 24947 1751 25249 1785
rect 25283 1751 25576 1785
rect 25628 1751 25921 1785
rect 25955 1751 26257 1785
rect 26291 1751 26593 1785
rect 26627 1751 26929 1785
rect 26963 1751 27256 1785
rect 27308 1751 27601 1785
rect 27635 1751 27937 1785
rect 27971 1751 28273 1785
rect 28307 1751 28609 1785
rect 28643 1751 28936 1785
rect 28988 1751 29281 1785
rect 29315 1751 29617 1785
rect 29651 1751 29953 1785
rect 29987 1751 30289 1785
rect 30323 1751 30616 1785
rect 30668 1751 30961 1785
rect 30995 1751 31297 1785
rect 31331 1751 31633 1785
rect 31667 1751 31969 1785
rect 32003 1751 32296 1785
rect 32348 1751 32641 1785
rect 32675 1751 32977 1785
rect 33011 1751 33313 1785
rect 33347 1751 33649 1785
rect 33683 1751 33976 1785
rect 34028 1751 34321 1785
rect 34355 1751 34657 1785
rect 34691 1751 34993 1785
rect 35027 1751 35329 1785
rect 35363 1751 35656 1785
rect 35708 1751 36001 1785
rect 36035 1751 36337 1785
rect 36371 1751 36673 1785
rect 36707 1751 37009 1785
rect 37043 1751 37336 1785
rect 37388 1751 37681 1785
rect 37715 1751 38017 1785
rect 38051 1751 38353 1785
rect 38387 1751 38689 1785
rect 38723 1751 39016 1785
rect 39068 1751 39361 1785
rect 39395 1751 39697 1785
rect 39731 1751 40033 1785
rect 40067 1751 40369 1785
rect 40403 1751 40696 1785
rect 40748 1751 41041 1785
rect 41075 1751 41377 1785
rect 41411 1751 41713 1785
rect 41747 1751 42049 1785
rect 42083 1751 42376 1785
rect 42428 1751 42721 1785
rect 42755 1751 43057 1785
rect 43091 1751 43393 1785
rect 43427 1751 43729 1785
rect 43763 1751 44056 1785
rect 44108 1751 44401 1785
rect 44435 1751 44737 1785
rect 44771 1751 45073 1785
rect 45107 1751 45409 1785
rect 45443 1751 45736 1785
rect 45788 1751 46081 1785
rect 46115 1751 46417 1785
rect 46451 1751 46753 1785
rect 46787 1751 47089 1785
rect 47123 1751 47416 1785
rect 47468 1751 47761 1785
rect 47795 1751 48097 1785
rect 48131 1751 48433 1785
rect 48467 1751 48769 1785
rect 48803 1751 49096 1785
rect 49148 1751 49441 1785
rect 49475 1751 49777 1785
rect 49811 1751 50113 1785
rect 50147 1751 50449 1785
rect 50483 1751 50776 1785
rect 50828 1751 51121 1785
rect 51155 1751 51457 1785
rect 51491 1751 51793 1785
rect 51827 1751 52129 1785
rect 52163 1751 52456 1785
rect 52508 1751 52801 1785
rect 52835 1751 53137 1785
rect 53171 1751 53473 1785
rect 53507 1751 53809 1785
rect 53843 1751 54136 1785
rect 54188 1751 54481 1785
rect 54515 1751 54817 1785
rect 54851 1751 55153 1785
rect 55187 1751 55489 1785
rect 55523 1751 55816 1785
rect 55868 1751 56161 1785
rect 56195 1751 56497 1785
rect 56531 1751 56833 1785
rect 56867 1751 57169 1785
rect 57203 1751 57496 1785
rect 57548 1751 57841 1785
rect 57875 1751 58177 1785
rect 58211 1751 58513 1785
rect 58547 1751 58849 1785
rect 58883 1751 59176 1785
rect 59228 1751 59521 1785
rect 59555 1751 59857 1785
rect 59891 1751 60193 1785
rect 60227 1751 60529 1785
rect 60563 1751 60856 1785
rect 60908 1751 61201 1785
rect 61235 1751 61537 1785
rect 61571 1751 61873 1785
rect 61907 1751 62209 1785
rect 62243 1751 62536 1785
rect 62588 1751 62881 1785
rect 62915 1751 63217 1785
rect 63251 1751 63553 1785
rect 63587 1751 63889 1785
rect 63923 1751 64216 1785
rect 64268 1751 64561 1785
rect 64595 1751 64897 1785
rect 64931 1751 65233 1785
rect 65267 1751 65569 1785
rect 65603 1751 65896 1785
rect 65948 1751 66241 1785
rect 66275 1751 66577 1785
rect 66611 1751 66913 1785
rect 66947 1751 67249 1785
rect 67283 1751 67576 1785
rect 67628 1751 67921 1785
rect 67955 1751 68257 1785
rect 68291 1751 68593 1785
rect 68627 1751 68929 1785
rect 68963 1751 69256 1785
rect 69308 1751 69601 1785
rect 69635 1751 69937 1785
rect 69971 1751 70273 1785
rect 70307 1751 70609 1785
rect 70643 1751 70936 1785
rect 70988 1751 71281 1785
rect 71315 1751 71617 1785
rect 71651 1751 71953 1785
rect 71987 1751 72289 1785
rect 72323 1751 72616 1785
rect 72668 1751 72961 1785
rect 72995 1751 73297 1785
rect 73331 1751 73633 1785
rect 73667 1751 73969 1785
rect 74003 1751 74296 1785
rect 74348 1751 74641 1785
rect 74675 1751 74977 1785
rect 75011 1751 75313 1785
rect 75347 1751 75649 1785
rect 75683 1751 75976 1785
rect 76028 1751 76321 1785
rect 76355 1751 76657 1785
rect 76691 1751 76993 1785
rect 77027 1751 77329 1785
rect 77363 1751 77656 1785
rect 77708 1751 78001 1785
rect 78035 1751 78337 1785
rect 78371 1751 78673 1785
rect 78707 1751 79009 1785
rect 79043 1751 79336 1785
rect 79388 1751 79681 1785
rect 79715 1751 80017 1785
rect 80051 1751 80353 1785
rect 80387 1751 80689 1785
rect 80723 1751 81016 1785
rect 81068 1751 81361 1785
rect 81395 1751 81697 1785
rect 81731 1751 82033 1785
rect 82067 1751 82369 1785
rect 82403 1751 82696 1785
rect 82748 1751 83041 1785
rect 83075 1751 83377 1785
rect 83411 1751 83713 1785
rect 83747 1751 84049 1785
rect 84083 1751 84376 1785
rect 84428 1751 84721 1785
rect 84755 1751 85057 1785
rect 85091 1751 85393 1785
rect 85427 1751 85729 1785
rect 85763 1751 86056 1785
rect 86108 1751 86401 1785
rect 86435 1751 86737 1785
rect 86771 1751 87073 1785
rect 87107 1751 87409 1785
rect 87443 1751 87736 1785
rect 87788 1751 88081 1785
rect 88115 1751 88417 1785
rect 88451 1751 88753 1785
rect 88787 1751 89356 1785
rect 2108 1742 3736 1751
rect 3788 1742 5416 1751
rect 5468 1742 7096 1751
rect 7148 1742 8776 1751
rect 8828 1742 10456 1751
rect 10508 1742 12136 1751
rect 12188 1742 13816 1751
rect 13868 1742 15496 1751
rect 15548 1742 17176 1751
rect 17228 1742 18856 1751
rect 18908 1742 20536 1751
rect 20588 1742 22216 1751
rect 22268 1742 23896 1751
rect 23948 1742 25576 1751
rect 25628 1742 27256 1751
rect 27308 1742 28936 1751
rect 28988 1742 30616 1751
rect 30668 1742 32296 1751
rect 32348 1742 33976 1751
rect 34028 1742 35656 1751
rect 35708 1742 37336 1751
rect 37388 1742 39016 1751
rect 39068 1742 40696 1751
rect 40748 1742 42376 1751
rect 42428 1742 44056 1751
rect 44108 1742 45736 1751
rect 45788 1742 47416 1751
rect 47468 1742 49096 1751
rect 49148 1742 50776 1751
rect 50828 1742 52456 1751
rect 52508 1742 54136 1751
rect 54188 1742 55816 1751
rect 55868 1742 57496 1751
rect 57548 1742 59176 1751
rect 59228 1742 60856 1751
rect 60908 1742 62536 1751
rect 62588 1742 64216 1751
rect 64268 1742 65896 1751
rect 65948 1742 67576 1751
rect 67628 1742 69256 1751
rect 69308 1742 70936 1751
rect 70988 1742 72616 1751
rect 72668 1742 74296 1751
rect 74348 1742 75976 1751
rect 76028 1742 77656 1751
rect 77708 1742 79336 1751
rect 79388 1742 81016 1751
rect 81068 1742 82696 1751
rect 82748 1742 84376 1751
rect 84428 1742 86056 1751
rect 86108 1742 87736 1751
rect 87788 1742 89356 1751
rect 1634 1656 89356 1742
<< via1 >>
rect 2056 87513 2108 87522
rect 3736 87513 3788 87522
rect 5416 87513 5468 87522
rect 7096 87513 7148 87522
rect 8776 87513 8828 87522
rect 10456 87513 10508 87522
rect 12136 87513 12188 87522
rect 13816 87513 13868 87522
rect 15496 87513 15548 87522
rect 17176 87513 17228 87522
rect 18856 87513 18908 87522
rect 20536 87513 20588 87522
rect 22216 87513 22268 87522
rect 23896 87513 23948 87522
rect 25576 87513 25628 87522
rect 27256 87513 27308 87522
rect 28936 87513 28988 87522
rect 30616 87513 30668 87522
rect 32296 87513 32348 87522
rect 33976 87513 34028 87522
rect 35656 87513 35708 87522
rect 37336 87513 37388 87522
rect 39016 87513 39068 87522
rect 40696 87513 40748 87522
rect 42376 87513 42428 87522
rect 44056 87513 44108 87522
rect 45736 87513 45788 87522
rect 47416 87513 47468 87522
rect 49096 87513 49148 87522
rect 50776 87513 50828 87522
rect 52456 87513 52508 87522
rect 54136 87513 54188 87522
rect 55816 87513 55868 87522
rect 57496 87513 57548 87522
rect 59176 87513 59228 87522
rect 60856 87513 60908 87522
rect 62536 87513 62588 87522
rect 64216 87513 64268 87522
rect 65896 87513 65948 87522
rect 67576 87513 67628 87522
rect 69256 87513 69308 87522
rect 70936 87513 70988 87522
rect 72616 87513 72668 87522
rect 74296 87513 74348 87522
rect 75976 87513 76028 87522
rect 77656 87513 77708 87522
rect 79336 87513 79388 87522
rect 81016 87513 81068 87522
rect 82696 87513 82748 87522
rect 84376 87513 84428 87522
rect 86056 87513 86108 87522
rect 87736 87513 87788 87522
rect 2056 87479 2065 87513
rect 2065 87479 2099 87513
rect 2099 87479 2108 87513
rect 3736 87479 3745 87513
rect 3745 87479 3779 87513
rect 3779 87479 3788 87513
rect 5416 87479 5425 87513
rect 5425 87479 5459 87513
rect 5459 87479 5468 87513
rect 7096 87479 7105 87513
rect 7105 87479 7139 87513
rect 7139 87479 7148 87513
rect 8776 87479 8785 87513
rect 8785 87479 8819 87513
rect 8819 87479 8828 87513
rect 10456 87479 10465 87513
rect 10465 87479 10499 87513
rect 10499 87479 10508 87513
rect 12136 87479 12145 87513
rect 12145 87479 12179 87513
rect 12179 87479 12188 87513
rect 13816 87479 13825 87513
rect 13825 87479 13859 87513
rect 13859 87479 13868 87513
rect 15496 87479 15505 87513
rect 15505 87479 15539 87513
rect 15539 87479 15548 87513
rect 17176 87479 17185 87513
rect 17185 87479 17219 87513
rect 17219 87479 17228 87513
rect 18856 87479 18865 87513
rect 18865 87479 18899 87513
rect 18899 87479 18908 87513
rect 20536 87479 20545 87513
rect 20545 87479 20579 87513
rect 20579 87479 20588 87513
rect 22216 87479 22225 87513
rect 22225 87479 22259 87513
rect 22259 87479 22268 87513
rect 23896 87479 23905 87513
rect 23905 87479 23939 87513
rect 23939 87479 23948 87513
rect 25576 87479 25585 87513
rect 25585 87479 25619 87513
rect 25619 87479 25628 87513
rect 27256 87479 27265 87513
rect 27265 87479 27299 87513
rect 27299 87479 27308 87513
rect 28936 87479 28945 87513
rect 28945 87479 28979 87513
rect 28979 87479 28988 87513
rect 30616 87479 30625 87513
rect 30625 87479 30659 87513
rect 30659 87479 30668 87513
rect 32296 87479 32305 87513
rect 32305 87479 32339 87513
rect 32339 87479 32348 87513
rect 33976 87479 33985 87513
rect 33985 87479 34019 87513
rect 34019 87479 34028 87513
rect 35656 87479 35665 87513
rect 35665 87479 35699 87513
rect 35699 87479 35708 87513
rect 37336 87479 37345 87513
rect 37345 87479 37379 87513
rect 37379 87479 37388 87513
rect 39016 87479 39025 87513
rect 39025 87479 39059 87513
rect 39059 87479 39068 87513
rect 40696 87479 40705 87513
rect 40705 87479 40739 87513
rect 40739 87479 40748 87513
rect 42376 87479 42385 87513
rect 42385 87479 42419 87513
rect 42419 87479 42428 87513
rect 44056 87479 44065 87513
rect 44065 87479 44099 87513
rect 44099 87479 44108 87513
rect 45736 87479 45745 87513
rect 45745 87479 45779 87513
rect 45779 87479 45788 87513
rect 47416 87479 47425 87513
rect 47425 87479 47459 87513
rect 47459 87479 47468 87513
rect 49096 87479 49105 87513
rect 49105 87479 49139 87513
rect 49139 87479 49148 87513
rect 50776 87479 50785 87513
rect 50785 87479 50819 87513
rect 50819 87479 50828 87513
rect 52456 87479 52465 87513
rect 52465 87479 52499 87513
rect 52499 87479 52508 87513
rect 54136 87479 54145 87513
rect 54145 87479 54179 87513
rect 54179 87479 54188 87513
rect 55816 87479 55825 87513
rect 55825 87479 55859 87513
rect 55859 87479 55868 87513
rect 57496 87479 57505 87513
rect 57505 87479 57539 87513
rect 57539 87479 57548 87513
rect 59176 87479 59185 87513
rect 59185 87479 59219 87513
rect 59219 87479 59228 87513
rect 60856 87479 60865 87513
rect 60865 87479 60899 87513
rect 60899 87479 60908 87513
rect 62536 87479 62545 87513
rect 62545 87479 62579 87513
rect 62579 87479 62588 87513
rect 64216 87479 64225 87513
rect 64225 87479 64259 87513
rect 64259 87479 64268 87513
rect 65896 87479 65905 87513
rect 65905 87479 65939 87513
rect 65939 87479 65948 87513
rect 67576 87479 67585 87513
rect 67585 87479 67619 87513
rect 67619 87479 67628 87513
rect 69256 87479 69265 87513
rect 69265 87479 69299 87513
rect 69299 87479 69308 87513
rect 70936 87479 70945 87513
rect 70945 87479 70979 87513
rect 70979 87479 70988 87513
rect 72616 87479 72625 87513
rect 72625 87479 72659 87513
rect 72659 87479 72668 87513
rect 74296 87479 74305 87513
rect 74305 87479 74339 87513
rect 74339 87479 74348 87513
rect 75976 87479 75985 87513
rect 75985 87479 76019 87513
rect 76019 87479 76028 87513
rect 77656 87479 77665 87513
rect 77665 87479 77699 87513
rect 77699 87479 77708 87513
rect 79336 87479 79345 87513
rect 79345 87479 79379 87513
rect 79379 87479 79388 87513
rect 81016 87479 81025 87513
rect 81025 87479 81059 87513
rect 81059 87479 81068 87513
rect 82696 87479 82705 87513
rect 82705 87479 82739 87513
rect 82739 87479 82748 87513
rect 84376 87479 84385 87513
rect 84385 87479 84419 87513
rect 84419 87479 84428 87513
rect 86056 87479 86065 87513
rect 86065 87479 86099 87513
rect 86099 87479 86108 87513
rect 87736 87479 87745 87513
rect 87745 87479 87779 87513
rect 87779 87479 87788 87513
rect 2056 87470 2108 87479
rect 3736 87470 3788 87479
rect 5416 87470 5468 87479
rect 7096 87470 7148 87479
rect 8776 87470 8828 87479
rect 10456 87470 10508 87479
rect 12136 87470 12188 87479
rect 13816 87470 13868 87479
rect 15496 87470 15548 87479
rect 17176 87470 17228 87479
rect 18856 87470 18908 87479
rect 20536 87470 20588 87479
rect 22216 87470 22268 87479
rect 23896 87470 23948 87479
rect 25576 87470 25628 87479
rect 27256 87470 27308 87479
rect 28936 87470 28988 87479
rect 30616 87470 30668 87479
rect 32296 87470 32348 87479
rect 33976 87470 34028 87479
rect 35656 87470 35708 87479
rect 37336 87470 37388 87479
rect 39016 87470 39068 87479
rect 40696 87470 40748 87479
rect 42376 87470 42428 87479
rect 44056 87470 44108 87479
rect 45736 87470 45788 87479
rect 47416 87470 47468 87479
rect 49096 87470 49148 87479
rect 50776 87470 50828 87479
rect 52456 87470 52508 87479
rect 54136 87470 54188 87479
rect 55816 87470 55868 87479
rect 57496 87470 57548 87479
rect 59176 87470 59228 87479
rect 60856 87470 60908 87479
rect 62536 87470 62588 87479
rect 64216 87470 64268 87479
rect 65896 87470 65948 87479
rect 67576 87470 67628 87479
rect 69256 87470 69308 87479
rect 70936 87470 70988 87479
rect 72616 87470 72668 87479
rect 74296 87470 74348 87479
rect 75976 87470 76028 87479
rect 77656 87470 77708 87479
rect 79336 87470 79388 87479
rect 81016 87470 81068 87479
rect 82696 87470 82748 87479
rect 84376 87470 84428 87479
rect 86056 87470 86108 87479
rect 87736 87470 87788 87479
rect 1720 87129 1772 87138
rect 1720 87095 1729 87129
rect 1729 87095 1763 87129
rect 1763 87095 1772 87129
rect 1720 87086 1772 87095
rect 89218 87129 89270 87138
rect 89218 87095 89227 87129
rect 89227 87095 89261 87129
rect 89261 87095 89270 87129
rect 89218 87086 89270 87095
rect 1720 86793 1772 86802
rect 1720 86759 1729 86793
rect 1729 86759 1763 86793
rect 1763 86759 1772 86793
rect 1720 86750 1772 86759
rect 89218 86793 89270 86802
rect 89218 86759 89227 86793
rect 89227 86759 89261 86793
rect 89261 86759 89270 86793
rect 89218 86750 89270 86759
rect 1720 86457 1772 86466
rect 1720 86423 1729 86457
rect 1729 86423 1763 86457
rect 1763 86423 1772 86457
rect 1720 86414 1772 86423
rect 89218 86457 89270 86466
rect 89218 86423 89227 86457
rect 89227 86423 89261 86457
rect 89261 86423 89270 86457
rect 89218 86414 89270 86423
rect 1720 86121 1772 86130
rect 1720 86087 1729 86121
rect 1729 86087 1763 86121
rect 1763 86087 1772 86121
rect 1720 86078 1772 86087
rect 89218 86121 89270 86130
rect 89218 86087 89227 86121
rect 89227 86087 89261 86121
rect 89261 86087 89270 86121
rect 89218 86078 89270 86087
rect 1720 85785 1772 85794
rect 1720 85751 1729 85785
rect 1729 85751 1763 85785
rect 1763 85751 1772 85785
rect 1720 85742 1772 85751
rect 89218 85785 89270 85794
rect 89218 85751 89227 85785
rect 89227 85751 89261 85785
rect 89261 85751 89270 85785
rect 89218 85742 89270 85751
rect 1720 85449 1772 85458
rect 1720 85415 1729 85449
rect 1729 85415 1763 85449
rect 1763 85415 1772 85449
rect 1720 85406 1772 85415
rect 89218 85449 89270 85458
rect 89218 85415 89227 85449
rect 89227 85415 89261 85449
rect 89261 85415 89270 85449
rect 89218 85406 89270 85415
rect 1720 85113 1772 85122
rect 1720 85079 1729 85113
rect 1729 85079 1763 85113
rect 1763 85079 1772 85113
rect 1720 85070 1772 85079
rect 89218 85113 89270 85122
rect 89218 85079 89227 85113
rect 89227 85079 89261 85113
rect 89261 85079 89270 85113
rect 89218 85070 89270 85079
rect 1720 84777 1772 84786
rect 1720 84743 1729 84777
rect 1729 84743 1763 84777
rect 1763 84743 1772 84777
rect 1720 84734 1772 84743
rect 89218 84777 89270 84786
rect 89218 84743 89227 84777
rect 89227 84743 89261 84777
rect 89261 84743 89270 84777
rect 89218 84734 89270 84743
rect 1720 84441 1772 84450
rect 1720 84407 1729 84441
rect 1729 84407 1763 84441
rect 1763 84407 1772 84441
rect 1720 84398 1772 84407
rect 89218 84441 89270 84450
rect 89218 84407 89227 84441
rect 89227 84407 89261 84441
rect 89261 84407 89270 84441
rect 89218 84398 89270 84407
rect 1720 84105 1772 84114
rect 1720 84071 1729 84105
rect 1729 84071 1763 84105
rect 1763 84071 1772 84105
rect 1720 84062 1772 84071
rect 89218 84105 89270 84114
rect 89218 84071 89227 84105
rect 89227 84071 89261 84105
rect 89261 84071 89270 84105
rect 89218 84062 89270 84071
rect 1720 83769 1772 83778
rect 1720 83735 1729 83769
rect 1729 83735 1763 83769
rect 1763 83735 1772 83769
rect 1720 83726 1772 83735
rect 89218 83769 89270 83778
rect 89218 83735 89227 83769
rect 89227 83735 89261 83769
rect 89261 83735 89270 83769
rect 89218 83726 89270 83735
rect 1720 83433 1772 83442
rect 1720 83399 1729 83433
rect 1729 83399 1763 83433
rect 1763 83399 1772 83433
rect 1720 83390 1772 83399
rect 89218 83433 89270 83442
rect 89218 83399 89227 83433
rect 89227 83399 89261 83433
rect 89261 83399 89270 83433
rect 89218 83390 89270 83399
rect 1720 83097 1772 83106
rect 1720 83063 1729 83097
rect 1729 83063 1763 83097
rect 1763 83063 1772 83097
rect 1720 83054 1772 83063
rect 89218 83097 89270 83106
rect 89218 83063 89227 83097
rect 89227 83063 89261 83097
rect 89261 83063 89270 83097
rect 89218 83054 89270 83063
rect 1720 82761 1772 82770
rect 1720 82727 1729 82761
rect 1729 82727 1763 82761
rect 1763 82727 1772 82761
rect 1720 82718 1772 82727
rect 89218 82761 89270 82770
rect 89218 82727 89227 82761
rect 89227 82727 89261 82761
rect 89261 82727 89270 82761
rect 89218 82718 89270 82727
rect 1720 82425 1772 82434
rect 1720 82391 1729 82425
rect 1729 82391 1763 82425
rect 1763 82391 1772 82425
rect 1720 82382 1772 82391
rect 89218 82425 89270 82434
rect 89218 82391 89227 82425
rect 89227 82391 89261 82425
rect 89261 82391 89270 82425
rect 89218 82382 89270 82391
rect 1720 82089 1772 82098
rect 1720 82055 1729 82089
rect 1729 82055 1763 82089
rect 1763 82055 1772 82089
rect 1720 82046 1772 82055
rect 89218 82089 89270 82098
rect 89218 82055 89227 82089
rect 89227 82055 89261 82089
rect 89261 82055 89270 82089
rect 89218 82046 89270 82055
rect 1720 81753 1772 81762
rect 1720 81719 1729 81753
rect 1729 81719 1763 81753
rect 1763 81719 1772 81753
rect 1720 81710 1772 81719
rect 89218 81753 89270 81762
rect 89218 81719 89227 81753
rect 89227 81719 89261 81753
rect 89261 81719 89270 81753
rect 89218 81710 89270 81719
rect 1720 81417 1772 81426
rect 1720 81383 1729 81417
rect 1729 81383 1763 81417
rect 1763 81383 1772 81417
rect 1720 81374 1772 81383
rect 89218 81417 89270 81426
rect 89218 81383 89227 81417
rect 89227 81383 89261 81417
rect 89261 81383 89270 81417
rect 89218 81374 89270 81383
rect 1720 81081 1772 81090
rect 1720 81047 1729 81081
rect 1729 81047 1763 81081
rect 1763 81047 1772 81081
rect 1720 81038 1772 81047
rect 89218 81081 89270 81090
rect 89218 81047 89227 81081
rect 89227 81047 89261 81081
rect 89261 81047 89270 81081
rect 89218 81038 89270 81047
rect 1720 80745 1772 80754
rect 1720 80711 1729 80745
rect 1729 80711 1763 80745
rect 1763 80711 1772 80745
rect 1720 80702 1772 80711
rect 89218 80745 89270 80754
rect 89218 80711 89227 80745
rect 89227 80711 89261 80745
rect 89261 80711 89270 80745
rect 89218 80702 89270 80711
rect 1720 80409 1772 80418
rect 1720 80375 1729 80409
rect 1729 80375 1763 80409
rect 1763 80375 1772 80409
rect 1720 80366 1772 80375
rect 89218 80409 89270 80418
rect 89218 80375 89227 80409
rect 89227 80375 89261 80409
rect 89261 80375 89270 80409
rect 89218 80366 89270 80375
rect 1720 80073 1772 80082
rect 1720 80039 1729 80073
rect 1729 80039 1763 80073
rect 1763 80039 1772 80073
rect 1720 80030 1772 80039
rect 89218 80073 89270 80082
rect 89218 80039 89227 80073
rect 89227 80039 89261 80073
rect 89261 80039 89270 80073
rect 89218 80030 89270 80039
rect 1720 79737 1772 79746
rect 1720 79703 1729 79737
rect 1729 79703 1763 79737
rect 1763 79703 1772 79737
rect 1720 79694 1772 79703
rect 89218 79737 89270 79746
rect 89218 79703 89227 79737
rect 89227 79703 89261 79737
rect 89261 79703 89270 79737
rect 89218 79694 89270 79703
rect 1720 79401 1772 79410
rect 1720 79367 1729 79401
rect 1729 79367 1763 79401
rect 1763 79367 1772 79401
rect 1720 79358 1772 79367
rect 89218 79401 89270 79410
rect 89218 79367 89227 79401
rect 89227 79367 89261 79401
rect 89261 79367 89270 79401
rect 89218 79358 89270 79367
rect 1720 79065 1772 79074
rect 1720 79031 1729 79065
rect 1729 79031 1763 79065
rect 1763 79031 1772 79065
rect 1720 79022 1772 79031
rect 89218 79065 89270 79074
rect 89218 79031 89227 79065
rect 89227 79031 89261 79065
rect 89261 79031 89270 79065
rect 89218 79022 89270 79031
rect 1720 78729 1772 78738
rect 1720 78695 1729 78729
rect 1729 78695 1763 78729
rect 1763 78695 1772 78729
rect 1720 78686 1772 78695
rect 89218 78729 89270 78738
rect 89218 78695 89227 78729
rect 89227 78695 89261 78729
rect 89261 78695 89270 78729
rect 89218 78686 89270 78695
rect 1720 78393 1772 78402
rect 1720 78359 1729 78393
rect 1729 78359 1763 78393
rect 1763 78359 1772 78393
rect 1720 78350 1772 78359
rect 89218 78393 89270 78402
rect 89218 78359 89227 78393
rect 89227 78359 89261 78393
rect 89261 78359 89270 78393
rect 89218 78350 89270 78359
rect 1720 78057 1772 78066
rect 1720 78023 1729 78057
rect 1729 78023 1763 78057
rect 1763 78023 1772 78057
rect 1720 78014 1772 78023
rect 89218 78057 89270 78066
rect 89218 78023 89227 78057
rect 89227 78023 89261 78057
rect 89261 78023 89270 78057
rect 89218 78014 89270 78023
rect 25628 77856 25680 77908
rect 30620 77856 30672 77908
rect 35612 77856 35664 77908
rect 40604 77856 40656 77908
rect 45596 77856 45648 77908
rect 50588 77856 50640 77908
rect 55580 77856 55632 77908
rect 60572 77856 60624 77908
rect 1720 77721 1772 77730
rect 1720 77687 1729 77721
rect 1729 77687 1763 77721
rect 1763 77687 1772 77721
rect 1720 77678 1772 77687
rect 89218 77721 89270 77730
rect 89218 77687 89227 77721
rect 89227 77687 89261 77721
rect 89261 77687 89270 77721
rect 89218 77678 89270 77687
rect 1720 77385 1772 77394
rect 1720 77351 1729 77385
rect 1729 77351 1763 77385
rect 1763 77351 1772 77385
rect 1720 77342 1772 77351
rect 89218 77385 89270 77394
rect 89218 77351 89227 77385
rect 89227 77351 89261 77385
rect 89261 77351 89270 77385
rect 89218 77342 89270 77351
rect 1720 77049 1772 77058
rect 1720 77015 1729 77049
rect 1729 77015 1763 77049
rect 1763 77015 1772 77049
rect 1720 77006 1772 77015
rect 89218 77049 89270 77058
rect 89218 77015 89227 77049
rect 89227 77015 89261 77049
rect 89261 77015 89270 77049
rect 89218 77006 89270 77015
rect 1720 76713 1772 76722
rect 1720 76679 1729 76713
rect 1729 76679 1763 76713
rect 1763 76679 1772 76713
rect 1720 76670 1772 76679
rect 89218 76713 89270 76722
rect 89218 76679 89227 76713
rect 89227 76679 89261 76713
rect 89261 76679 89270 76713
rect 89218 76670 89270 76679
rect 1720 76377 1772 76386
rect 1720 76343 1729 76377
rect 1729 76343 1763 76377
rect 1763 76343 1772 76377
rect 1720 76334 1772 76343
rect 89218 76377 89270 76386
rect 89218 76343 89227 76377
rect 89227 76343 89261 76377
rect 89261 76343 89270 76377
rect 89218 76334 89270 76343
rect 1720 76041 1772 76050
rect 1720 76007 1729 76041
rect 1729 76007 1763 76041
rect 1763 76007 1772 76041
rect 1720 75998 1772 76007
rect 89218 76041 89270 76050
rect 89218 76007 89227 76041
rect 89227 76007 89261 76041
rect 89261 76007 89270 76041
rect 89218 75998 89270 76007
rect 1720 75705 1772 75714
rect 1720 75671 1729 75705
rect 1729 75671 1763 75705
rect 1763 75671 1772 75705
rect 1720 75662 1772 75671
rect 89218 75705 89270 75714
rect 89218 75671 89227 75705
rect 89227 75671 89261 75705
rect 89261 75671 89270 75705
rect 89218 75662 89270 75671
rect 1720 75369 1772 75378
rect 1720 75335 1729 75369
rect 1729 75335 1763 75369
rect 1763 75335 1772 75369
rect 1720 75326 1772 75335
rect 89218 75369 89270 75378
rect 89218 75335 89227 75369
rect 89227 75335 89261 75369
rect 89261 75335 89270 75369
rect 89218 75326 89270 75335
rect 1720 75033 1772 75042
rect 1720 74999 1729 75033
rect 1729 74999 1763 75033
rect 1763 74999 1772 75033
rect 1720 74990 1772 74999
rect 89218 75033 89270 75042
rect 89218 74999 89227 75033
rect 89227 74999 89261 75033
rect 89261 74999 89270 75033
rect 89218 74990 89270 74999
rect 1720 74697 1772 74706
rect 1720 74663 1729 74697
rect 1729 74663 1763 74697
rect 1763 74663 1772 74697
rect 1720 74654 1772 74663
rect 89218 74697 89270 74706
rect 89218 74663 89227 74697
rect 89227 74663 89261 74697
rect 89261 74663 89270 74697
rect 89218 74654 89270 74663
rect 1720 74361 1772 74370
rect 1720 74327 1729 74361
rect 1729 74327 1763 74361
rect 1763 74327 1772 74361
rect 1720 74318 1772 74327
rect 89218 74361 89270 74370
rect 89218 74327 89227 74361
rect 89227 74327 89261 74361
rect 89261 74327 89270 74361
rect 89218 74318 89270 74327
rect 1720 74025 1772 74034
rect 1720 73991 1729 74025
rect 1729 73991 1763 74025
rect 1763 73991 1772 74025
rect 1720 73982 1772 73991
rect 89218 74025 89270 74034
rect 89218 73991 89227 74025
rect 89227 73991 89261 74025
rect 89261 73991 89270 74025
rect 89218 73982 89270 73991
rect 1720 73689 1772 73698
rect 1720 73655 1729 73689
rect 1729 73655 1763 73689
rect 1763 73655 1772 73689
rect 1720 73646 1772 73655
rect 89218 73689 89270 73698
rect 89218 73655 89227 73689
rect 89227 73655 89261 73689
rect 89261 73655 89270 73689
rect 89218 73646 89270 73655
rect 1720 73353 1772 73362
rect 1720 73319 1729 73353
rect 1729 73319 1763 73353
rect 1763 73319 1772 73353
rect 1720 73310 1772 73319
rect 89218 73353 89270 73362
rect 89218 73319 89227 73353
rect 89227 73319 89261 73353
rect 89261 73319 89270 73353
rect 89218 73310 89270 73319
rect 1720 73017 1772 73026
rect 1720 72983 1729 73017
rect 1729 72983 1763 73017
rect 1763 72983 1772 73017
rect 1720 72974 1772 72983
rect 89218 73017 89270 73026
rect 89218 72983 89227 73017
rect 89227 72983 89261 73017
rect 89261 72983 89270 73017
rect 89218 72974 89270 72983
rect 1720 72681 1772 72690
rect 1720 72647 1729 72681
rect 1729 72647 1763 72681
rect 1763 72647 1772 72681
rect 1720 72638 1772 72647
rect 89218 72681 89270 72690
rect 89218 72647 89227 72681
rect 89227 72647 89261 72681
rect 89261 72647 89270 72681
rect 89218 72638 89270 72647
rect 1720 72345 1772 72354
rect 1720 72311 1729 72345
rect 1729 72311 1763 72345
rect 1763 72311 1772 72345
rect 1720 72302 1772 72311
rect 89218 72345 89270 72354
rect 89218 72311 89227 72345
rect 89227 72311 89261 72345
rect 89261 72311 89270 72345
rect 89218 72302 89270 72311
rect 1720 72009 1772 72018
rect 1720 71975 1729 72009
rect 1729 71975 1763 72009
rect 1763 71975 1772 72009
rect 1720 71966 1772 71975
rect 89218 72009 89270 72018
rect 89218 71975 89227 72009
rect 89227 71975 89261 72009
rect 89261 71975 89270 72009
rect 89218 71966 89270 71975
rect 1720 71673 1772 71682
rect 1720 71639 1729 71673
rect 1729 71639 1763 71673
rect 1763 71639 1772 71673
rect 1720 71630 1772 71639
rect 89218 71673 89270 71682
rect 89218 71639 89227 71673
rect 89227 71639 89261 71673
rect 89261 71639 89270 71673
rect 89218 71630 89270 71639
rect 1720 71337 1772 71346
rect 1720 71303 1729 71337
rect 1729 71303 1763 71337
rect 1763 71303 1772 71337
rect 1720 71294 1772 71303
rect 89218 71337 89270 71346
rect 89218 71303 89227 71337
rect 89227 71303 89261 71337
rect 89261 71303 89270 71337
rect 89218 71294 89270 71303
rect 1720 71001 1772 71010
rect 1720 70967 1729 71001
rect 1729 70967 1763 71001
rect 1763 70967 1772 71001
rect 1720 70958 1772 70967
rect 89218 71001 89270 71010
rect 89218 70967 89227 71001
rect 89227 70967 89261 71001
rect 89261 70967 89270 71001
rect 89218 70958 89270 70967
rect 1720 70665 1772 70674
rect 1720 70631 1729 70665
rect 1729 70631 1763 70665
rect 1763 70631 1772 70665
rect 1720 70622 1772 70631
rect 89218 70665 89270 70674
rect 89218 70631 89227 70665
rect 89227 70631 89261 70665
rect 89261 70631 89270 70665
rect 89218 70622 89270 70631
rect 1720 70329 1772 70338
rect 1720 70295 1729 70329
rect 1729 70295 1763 70329
rect 1763 70295 1772 70329
rect 1720 70286 1772 70295
rect 89218 70329 89270 70338
rect 89218 70295 89227 70329
rect 89227 70295 89261 70329
rect 89261 70295 89270 70329
rect 89218 70286 89270 70295
rect 1720 69993 1772 70002
rect 1720 69959 1729 69993
rect 1729 69959 1763 69993
rect 1763 69959 1772 69993
rect 1720 69950 1772 69959
rect 89218 69993 89270 70002
rect 89218 69959 89227 69993
rect 89227 69959 89261 69993
rect 89261 69959 89270 69993
rect 89218 69950 89270 69959
rect 1720 69657 1772 69666
rect 1720 69623 1729 69657
rect 1729 69623 1763 69657
rect 1763 69623 1772 69657
rect 1720 69614 1772 69623
rect 89218 69657 89270 69666
rect 89218 69623 89227 69657
rect 89227 69623 89261 69657
rect 89261 69623 89270 69657
rect 89218 69614 89270 69623
rect 1720 69321 1772 69330
rect 1720 69287 1729 69321
rect 1729 69287 1763 69321
rect 1763 69287 1772 69321
rect 1720 69278 1772 69287
rect 89218 69321 89270 69330
rect 89218 69287 89227 69321
rect 89227 69287 89261 69321
rect 89261 69287 89270 69321
rect 89218 69278 89270 69287
rect 1720 68985 1772 68994
rect 1720 68951 1729 68985
rect 1729 68951 1763 68985
rect 1763 68951 1772 68985
rect 1720 68942 1772 68951
rect 89218 68985 89270 68994
rect 89218 68951 89227 68985
rect 89227 68951 89261 68985
rect 89261 68951 89270 68985
rect 89218 68942 89270 68951
rect 1720 68649 1772 68658
rect 1720 68615 1729 68649
rect 1729 68615 1763 68649
rect 1763 68615 1772 68649
rect 1720 68606 1772 68615
rect 89218 68649 89270 68658
rect 89218 68615 89227 68649
rect 89227 68615 89261 68649
rect 89261 68615 89270 68649
rect 89218 68606 89270 68615
rect 1720 68313 1772 68322
rect 1720 68279 1729 68313
rect 1729 68279 1763 68313
rect 1763 68279 1772 68313
rect 1720 68270 1772 68279
rect 89218 68313 89270 68322
rect 89218 68279 89227 68313
rect 89227 68279 89261 68313
rect 89261 68279 89270 68313
rect 89218 68270 89270 68279
rect 1720 67977 1772 67986
rect 1720 67943 1729 67977
rect 1729 67943 1763 67977
rect 1763 67943 1772 67977
rect 1720 67934 1772 67943
rect 89218 67977 89270 67986
rect 89218 67943 89227 67977
rect 89227 67943 89261 67977
rect 89261 67943 89270 67977
rect 89218 67934 89270 67943
rect 1720 67641 1772 67650
rect 1720 67607 1729 67641
rect 1729 67607 1763 67641
rect 1763 67607 1772 67641
rect 1720 67598 1772 67607
rect 89218 67641 89270 67650
rect 89218 67607 89227 67641
rect 89227 67607 89261 67641
rect 89261 67607 89270 67641
rect 89218 67598 89270 67607
rect 1720 67305 1772 67314
rect 1720 67271 1729 67305
rect 1729 67271 1763 67305
rect 1763 67271 1772 67305
rect 1720 67262 1772 67271
rect 89218 67305 89270 67314
rect 89218 67271 89227 67305
rect 89227 67271 89261 67305
rect 89261 67271 89270 67305
rect 89218 67262 89270 67271
rect 1720 66969 1772 66978
rect 1720 66935 1729 66969
rect 1729 66935 1763 66969
rect 1763 66935 1772 66969
rect 1720 66926 1772 66935
rect 89218 66969 89270 66978
rect 89218 66935 89227 66969
rect 89227 66935 89261 66969
rect 89261 66935 89270 66969
rect 89218 66926 89270 66935
rect 1720 66633 1772 66642
rect 1720 66599 1729 66633
rect 1729 66599 1763 66633
rect 1763 66599 1772 66633
rect 1720 66590 1772 66599
rect 89218 66633 89270 66642
rect 89218 66599 89227 66633
rect 89227 66599 89261 66633
rect 89261 66599 89270 66633
rect 89218 66590 89270 66599
rect 1720 66297 1772 66306
rect 1720 66263 1729 66297
rect 1729 66263 1763 66297
rect 1763 66263 1772 66297
rect 1720 66254 1772 66263
rect 89218 66297 89270 66306
rect 89218 66263 89227 66297
rect 89227 66263 89261 66297
rect 89261 66263 89270 66297
rect 89218 66254 89270 66263
rect 1720 65961 1772 65970
rect 1720 65927 1729 65961
rect 1729 65927 1763 65961
rect 1763 65927 1772 65961
rect 1720 65918 1772 65927
rect 89218 65961 89270 65970
rect 89218 65927 89227 65961
rect 89227 65927 89261 65961
rect 89261 65927 89270 65961
rect 89218 65918 89270 65927
rect 1720 65625 1772 65634
rect 1720 65591 1729 65625
rect 1729 65591 1763 65625
rect 1763 65591 1772 65625
rect 1720 65582 1772 65591
rect 89218 65625 89270 65634
rect 89218 65591 89227 65625
rect 89227 65591 89261 65625
rect 89261 65591 89270 65625
rect 89218 65582 89270 65591
rect 1720 65289 1772 65298
rect 1720 65255 1729 65289
rect 1729 65255 1763 65289
rect 1763 65255 1772 65289
rect 1720 65246 1772 65255
rect 89218 65289 89270 65298
rect 89218 65255 89227 65289
rect 89227 65255 89261 65289
rect 89261 65255 89270 65289
rect 89218 65246 89270 65255
rect 1720 64953 1772 64962
rect 1720 64919 1729 64953
rect 1729 64919 1763 64953
rect 1763 64919 1772 64953
rect 1720 64910 1772 64919
rect 89218 64953 89270 64962
rect 89218 64919 89227 64953
rect 89227 64919 89261 64953
rect 89261 64919 89270 64953
rect 89218 64910 89270 64919
rect 1720 64617 1772 64626
rect 1720 64583 1729 64617
rect 1729 64583 1763 64617
rect 1763 64583 1772 64617
rect 1720 64574 1772 64583
rect 89218 64617 89270 64626
rect 89218 64583 89227 64617
rect 89227 64583 89261 64617
rect 89261 64583 89270 64617
rect 89218 64574 89270 64583
rect 1720 64281 1772 64290
rect 1720 64247 1729 64281
rect 1729 64247 1763 64281
rect 1763 64247 1772 64281
rect 1720 64238 1772 64247
rect 89218 64281 89270 64290
rect 89218 64247 89227 64281
rect 89227 64247 89261 64281
rect 89261 64247 89270 64281
rect 89218 64238 89270 64247
rect 1720 63945 1772 63954
rect 1720 63911 1729 63945
rect 1729 63911 1763 63945
rect 1763 63911 1772 63945
rect 1720 63902 1772 63911
rect 89218 63945 89270 63954
rect 89218 63911 89227 63945
rect 89227 63911 89261 63945
rect 89261 63911 89270 63945
rect 89218 63902 89270 63911
rect 1720 63609 1772 63618
rect 1720 63575 1729 63609
rect 1729 63575 1763 63609
rect 1763 63575 1772 63609
rect 1720 63566 1772 63575
rect 89218 63609 89270 63618
rect 89218 63575 89227 63609
rect 89227 63575 89261 63609
rect 89261 63575 89270 63609
rect 89218 63566 89270 63575
rect 1720 63273 1772 63282
rect 1720 63239 1729 63273
rect 1729 63239 1763 63273
rect 1763 63239 1772 63273
rect 1720 63230 1772 63239
rect 89218 63273 89270 63282
rect 89218 63239 89227 63273
rect 89227 63239 89261 63273
rect 89261 63239 89270 63273
rect 89218 63230 89270 63239
rect 1720 62937 1772 62946
rect 1720 62903 1729 62937
rect 1729 62903 1763 62937
rect 1763 62903 1772 62937
rect 1720 62894 1772 62903
rect 89218 62937 89270 62946
rect 89218 62903 89227 62937
rect 89227 62903 89261 62937
rect 89261 62903 89270 62937
rect 89218 62894 89270 62903
rect 1720 62601 1772 62610
rect 1720 62567 1729 62601
rect 1729 62567 1763 62601
rect 1763 62567 1772 62601
rect 1720 62558 1772 62567
rect 89218 62601 89270 62610
rect 89218 62567 89227 62601
rect 89227 62567 89261 62601
rect 89261 62567 89270 62601
rect 89218 62558 89270 62567
rect 1720 62265 1772 62274
rect 1720 62231 1729 62265
rect 1729 62231 1763 62265
rect 1763 62231 1772 62265
rect 1720 62222 1772 62231
rect 89218 62265 89270 62274
rect 89218 62231 89227 62265
rect 89227 62231 89261 62265
rect 89261 62231 89270 62265
rect 89218 62222 89270 62231
rect 1720 61929 1772 61938
rect 1720 61895 1729 61929
rect 1729 61895 1763 61929
rect 1763 61895 1772 61929
rect 1720 61886 1772 61895
rect 89218 61929 89270 61938
rect 89218 61895 89227 61929
rect 89227 61895 89261 61929
rect 89261 61895 89270 61929
rect 89218 61886 89270 61895
rect 1720 61593 1772 61602
rect 1720 61559 1729 61593
rect 1729 61559 1763 61593
rect 1763 61559 1772 61593
rect 1720 61550 1772 61559
rect 89218 61593 89270 61602
rect 89218 61559 89227 61593
rect 89227 61559 89261 61593
rect 89261 61559 89270 61593
rect 89218 61550 89270 61559
rect 1720 61257 1772 61266
rect 1720 61223 1729 61257
rect 1729 61223 1763 61257
rect 1763 61223 1772 61257
rect 1720 61214 1772 61223
rect 89218 61257 89270 61266
rect 89218 61223 89227 61257
rect 89227 61223 89261 61257
rect 89261 61223 89270 61257
rect 89218 61214 89270 61223
rect 1720 60921 1772 60930
rect 1720 60887 1729 60921
rect 1729 60887 1763 60921
rect 1763 60887 1772 60921
rect 1720 60878 1772 60887
rect 89218 60921 89270 60930
rect 89218 60887 89227 60921
rect 89227 60887 89261 60921
rect 89261 60887 89270 60921
rect 89218 60878 89270 60887
rect 1720 60585 1772 60594
rect 1720 60551 1729 60585
rect 1729 60551 1763 60585
rect 1763 60551 1772 60585
rect 1720 60542 1772 60551
rect 89218 60585 89270 60594
rect 89218 60551 89227 60585
rect 89227 60551 89261 60585
rect 89261 60551 89270 60585
rect 89218 60542 89270 60551
rect 1720 60249 1772 60258
rect 1720 60215 1729 60249
rect 1729 60215 1763 60249
rect 1763 60215 1772 60249
rect 1720 60206 1772 60215
rect 89218 60249 89270 60258
rect 89218 60215 89227 60249
rect 89227 60215 89261 60249
rect 89261 60215 89270 60249
rect 89218 60206 89270 60215
rect 1720 59913 1772 59922
rect 1720 59879 1729 59913
rect 1729 59879 1763 59913
rect 1763 59879 1772 59913
rect 1720 59870 1772 59879
rect 89218 59913 89270 59922
rect 89218 59879 89227 59913
rect 89227 59879 89261 59913
rect 89261 59879 89270 59913
rect 89218 59870 89270 59879
rect 1720 59577 1772 59586
rect 1720 59543 1729 59577
rect 1729 59543 1763 59577
rect 1763 59543 1772 59577
rect 1720 59534 1772 59543
rect 89218 59577 89270 59586
rect 89218 59543 89227 59577
rect 89227 59543 89261 59577
rect 89261 59543 89270 59577
rect 89218 59534 89270 59543
rect 1720 59241 1772 59250
rect 1720 59207 1729 59241
rect 1729 59207 1763 59241
rect 1763 59207 1772 59241
rect 1720 59198 1772 59207
rect 89218 59241 89270 59250
rect 89218 59207 89227 59241
rect 89227 59207 89261 59241
rect 89261 59207 89270 59241
rect 89218 59198 89270 59207
rect 1720 58905 1772 58914
rect 1720 58871 1729 58905
rect 1729 58871 1763 58905
rect 1763 58871 1772 58905
rect 1720 58862 1772 58871
rect 89218 58905 89270 58914
rect 89218 58871 89227 58905
rect 89227 58871 89261 58905
rect 89261 58871 89270 58905
rect 89218 58862 89270 58871
rect 1720 58569 1772 58578
rect 1720 58535 1729 58569
rect 1729 58535 1763 58569
rect 1763 58535 1772 58569
rect 1720 58526 1772 58535
rect 89218 58569 89270 58578
rect 89218 58535 89227 58569
rect 89227 58535 89261 58569
rect 89261 58535 89270 58569
rect 89218 58526 89270 58535
rect 1720 58233 1772 58242
rect 1720 58199 1729 58233
rect 1729 58199 1763 58233
rect 1763 58199 1772 58233
rect 1720 58190 1772 58199
rect 89218 58233 89270 58242
rect 89218 58199 89227 58233
rect 89227 58199 89261 58233
rect 89261 58199 89270 58233
rect 89218 58190 89270 58199
rect 1720 57897 1772 57906
rect 1720 57863 1729 57897
rect 1729 57863 1763 57897
rect 1763 57863 1772 57897
rect 1720 57854 1772 57863
rect 89218 57897 89270 57906
rect 89218 57863 89227 57897
rect 89227 57863 89261 57897
rect 89261 57863 89270 57897
rect 89218 57854 89270 57863
rect 1720 57561 1772 57570
rect 1720 57527 1729 57561
rect 1729 57527 1763 57561
rect 1763 57527 1772 57561
rect 1720 57518 1772 57527
rect 89218 57561 89270 57570
rect 89218 57527 89227 57561
rect 89227 57527 89261 57561
rect 89261 57527 89270 57561
rect 89218 57518 89270 57527
rect 1720 57225 1772 57234
rect 1720 57191 1729 57225
rect 1729 57191 1763 57225
rect 1763 57191 1772 57225
rect 1720 57182 1772 57191
rect 89218 57225 89270 57234
rect 89218 57191 89227 57225
rect 89227 57191 89261 57225
rect 89261 57191 89270 57225
rect 89218 57182 89270 57191
rect 1720 56889 1772 56898
rect 1720 56855 1729 56889
rect 1729 56855 1763 56889
rect 1763 56855 1772 56889
rect 1720 56846 1772 56855
rect 89218 56889 89270 56898
rect 89218 56855 89227 56889
rect 89227 56855 89261 56889
rect 89261 56855 89270 56889
rect 89218 56846 89270 56855
rect 1720 56553 1772 56562
rect 1720 56519 1729 56553
rect 1729 56519 1763 56553
rect 1763 56519 1772 56553
rect 1720 56510 1772 56519
rect 89218 56553 89270 56562
rect 89218 56519 89227 56553
rect 89227 56519 89261 56553
rect 89261 56519 89270 56553
rect 89218 56510 89270 56519
rect 1720 56217 1772 56226
rect 1720 56183 1729 56217
rect 1729 56183 1763 56217
rect 1763 56183 1772 56217
rect 1720 56174 1772 56183
rect 89218 56217 89270 56226
rect 89218 56183 89227 56217
rect 89227 56183 89261 56217
rect 89261 56183 89270 56217
rect 89218 56174 89270 56183
rect 1720 55881 1772 55890
rect 1720 55847 1729 55881
rect 1729 55847 1763 55881
rect 1763 55847 1772 55881
rect 1720 55838 1772 55847
rect 89218 55881 89270 55890
rect 89218 55847 89227 55881
rect 89227 55847 89261 55881
rect 89261 55847 89270 55881
rect 89218 55838 89270 55847
rect 1720 55545 1772 55554
rect 1720 55511 1729 55545
rect 1729 55511 1763 55545
rect 1763 55511 1772 55545
rect 1720 55502 1772 55511
rect 89218 55545 89270 55554
rect 89218 55511 89227 55545
rect 89227 55511 89261 55545
rect 89261 55511 89270 55545
rect 89218 55502 89270 55511
rect 1720 55209 1772 55218
rect 1720 55175 1729 55209
rect 1729 55175 1763 55209
rect 1763 55175 1772 55209
rect 1720 55166 1772 55175
rect 89218 55209 89270 55218
rect 89218 55175 89227 55209
rect 89227 55175 89261 55209
rect 89261 55175 89270 55209
rect 89218 55166 89270 55175
rect 1720 54873 1772 54882
rect 1720 54839 1729 54873
rect 1729 54839 1763 54873
rect 1763 54839 1772 54873
rect 1720 54830 1772 54839
rect 89218 54873 89270 54882
rect 89218 54839 89227 54873
rect 89227 54839 89261 54873
rect 89261 54839 89270 54873
rect 89218 54830 89270 54839
rect 1720 54537 1772 54546
rect 1720 54503 1729 54537
rect 1729 54503 1763 54537
rect 1763 54503 1772 54537
rect 1720 54494 1772 54503
rect 89218 54537 89270 54546
rect 89218 54503 89227 54537
rect 89227 54503 89261 54537
rect 89261 54503 89270 54537
rect 89218 54494 89270 54503
rect 1720 54201 1772 54210
rect 1720 54167 1729 54201
rect 1729 54167 1763 54201
rect 1763 54167 1772 54201
rect 1720 54158 1772 54167
rect 89218 54201 89270 54210
rect 89218 54167 89227 54201
rect 89227 54167 89261 54201
rect 89261 54167 89270 54201
rect 89218 54158 89270 54167
rect 1720 53865 1772 53874
rect 1720 53831 1729 53865
rect 1729 53831 1763 53865
rect 1763 53831 1772 53865
rect 1720 53822 1772 53831
rect 89218 53865 89270 53874
rect 89218 53831 89227 53865
rect 89227 53831 89261 53865
rect 89261 53831 89270 53865
rect 89218 53822 89270 53831
rect 1720 53529 1772 53538
rect 1720 53495 1729 53529
rect 1729 53495 1763 53529
rect 1763 53495 1772 53529
rect 1720 53486 1772 53495
rect 89218 53529 89270 53538
rect 89218 53495 89227 53529
rect 89227 53495 89261 53529
rect 89261 53495 89270 53529
rect 89218 53486 89270 53495
rect 1720 53193 1772 53202
rect 1720 53159 1729 53193
rect 1729 53159 1763 53193
rect 1763 53159 1772 53193
rect 1720 53150 1772 53159
rect 89218 53193 89270 53202
rect 89218 53159 89227 53193
rect 89227 53159 89261 53193
rect 89261 53159 89270 53193
rect 89218 53150 89270 53159
rect 1720 52857 1772 52866
rect 1720 52823 1729 52857
rect 1729 52823 1763 52857
rect 1763 52823 1772 52857
rect 1720 52814 1772 52823
rect 89218 52857 89270 52866
rect 89218 52823 89227 52857
rect 89227 52823 89261 52857
rect 89261 52823 89270 52857
rect 89218 52814 89270 52823
rect 1720 52521 1772 52530
rect 1720 52487 1729 52521
rect 1729 52487 1763 52521
rect 1763 52487 1772 52521
rect 1720 52478 1772 52487
rect 89218 52521 89270 52530
rect 89218 52487 89227 52521
rect 89227 52487 89261 52521
rect 89261 52487 89270 52521
rect 89218 52478 89270 52487
rect 1720 52185 1772 52194
rect 1720 52151 1729 52185
rect 1729 52151 1763 52185
rect 1763 52151 1772 52185
rect 1720 52142 1772 52151
rect 89218 52185 89270 52194
rect 89218 52151 89227 52185
rect 89227 52151 89261 52185
rect 89261 52151 89270 52185
rect 89218 52142 89270 52151
rect 1720 51849 1772 51858
rect 1720 51815 1729 51849
rect 1729 51815 1763 51849
rect 1763 51815 1772 51849
rect 1720 51806 1772 51815
rect 89218 51849 89270 51858
rect 89218 51815 89227 51849
rect 89227 51815 89261 51849
rect 89261 51815 89270 51849
rect 89218 51806 89270 51815
rect 1720 51513 1772 51522
rect 1720 51479 1729 51513
rect 1729 51479 1763 51513
rect 1763 51479 1772 51513
rect 1720 51470 1772 51479
rect 89218 51513 89270 51522
rect 89218 51479 89227 51513
rect 89227 51479 89261 51513
rect 89261 51479 89270 51513
rect 89218 51470 89270 51479
rect 1720 51177 1772 51186
rect 1720 51143 1729 51177
rect 1729 51143 1763 51177
rect 1763 51143 1772 51177
rect 1720 51134 1772 51143
rect 89218 51177 89270 51186
rect 89218 51143 89227 51177
rect 89227 51143 89261 51177
rect 89261 51143 89270 51177
rect 89218 51134 89270 51143
rect 1720 50841 1772 50850
rect 1720 50807 1729 50841
rect 1729 50807 1763 50841
rect 1763 50807 1772 50841
rect 1720 50798 1772 50807
rect 89218 50841 89270 50850
rect 89218 50807 89227 50841
rect 89227 50807 89261 50841
rect 89261 50807 89270 50841
rect 89218 50798 89270 50807
rect 1720 50505 1772 50514
rect 1720 50471 1729 50505
rect 1729 50471 1763 50505
rect 1763 50471 1772 50505
rect 1720 50462 1772 50471
rect 89218 50505 89270 50514
rect 89218 50471 89227 50505
rect 89227 50471 89261 50505
rect 89261 50471 89270 50505
rect 89218 50462 89270 50471
rect 1720 50169 1772 50178
rect 1720 50135 1729 50169
rect 1729 50135 1763 50169
rect 1763 50135 1772 50169
rect 1720 50126 1772 50135
rect 89218 50169 89270 50178
rect 89218 50135 89227 50169
rect 89227 50135 89261 50169
rect 89261 50135 89270 50169
rect 89218 50126 89270 50135
rect 1720 49833 1772 49842
rect 1720 49799 1729 49833
rect 1729 49799 1763 49833
rect 1763 49799 1772 49833
rect 1720 49790 1772 49799
rect 89218 49833 89270 49842
rect 89218 49799 89227 49833
rect 89227 49799 89261 49833
rect 89261 49799 89270 49833
rect 89218 49790 89270 49799
rect 1720 49497 1772 49506
rect 1720 49463 1729 49497
rect 1729 49463 1763 49497
rect 1763 49463 1772 49497
rect 1720 49454 1772 49463
rect 89218 49497 89270 49506
rect 89218 49463 89227 49497
rect 89227 49463 89261 49497
rect 89261 49463 89270 49497
rect 89218 49454 89270 49463
rect 1720 49161 1772 49170
rect 1720 49127 1729 49161
rect 1729 49127 1763 49161
rect 1763 49127 1772 49161
rect 1720 49118 1772 49127
rect 89218 49161 89270 49170
rect 89218 49127 89227 49161
rect 89227 49127 89261 49161
rect 89261 49127 89270 49161
rect 89218 49118 89270 49127
rect 1720 48825 1772 48834
rect 1720 48791 1729 48825
rect 1729 48791 1763 48825
rect 1763 48791 1772 48825
rect 1720 48782 1772 48791
rect 89218 48825 89270 48834
rect 89218 48791 89227 48825
rect 89227 48791 89261 48825
rect 89261 48791 89270 48825
rect 89218 48782 89270 48791
rect 1720 48489 1772 48498
rect 1720 48455 1729 48489
rect 1729 48455 1763 48489
rect 1763 48455 1772 48489
rect 1720 48446 1772 48455
rect 89218 48489 89270 48498
rect 89218 48455 89227 48489
rect 89227 48455 89261 48489
rect 89261 48455 89270 48489
rect 89218 48446 89270 48455
rect 1720 48153 1772 48162
rect 1720 48119 1729 48153
rect 1729 48119 1763 48153
rect 1763 48119 1772 48153
rect 1720 48110 1772 48119
rect 89218 48153 89270 48162
rect 89218 48119 89227 48153
rect 89227 48119 89261 48153
rect 89261 48119 89270 48153
rect 89218 48110 89270 48119
rect 1720 47817 1772 47826
rect 1720 47783 1729 47817
rect 1729 47783 1763 47817
rect 1763 47783 1772 47817
rect 1720 47774 1772 47783
rect 89218 47817 89270 47826
rect 89218 47783 89227 47817
rect 89227 47783 89261 47817
rect 89261 47783 89270 47817
rect 89218 47774 89270 47783
rect 1720 47481 1772 47490
rect 1720 47447 1729 47481
rect 1729 47447 1763 47481
rect 1763 47447 1772 47481
rect 1720 47438 1772 47447
rect 89218 47481 89270 47490
rect 89218 47447 89227 47481
rect 89227 47447 89261 47481
rect 89261 47447 89270 47481
rect 89218 47438 89270 47447
rect 1720 47145 1772 47154
rect 1720 47111 1729 47145
rect 1729 47111 1763 47145
rect 1763 47111 1772 47145
rect 1720 47102 1772 47111
rect 89218 47145 89270 47154
rect 89218 47111 89227 47145
rect 89227 47111 89261 47145
rect 89261 47111 89270 47145
rect 89218 47102 89270 47111
rect 1720 46809 1772 46818
rect 1720 46775 1729 46809
rect 1729 46775 1763 46809
rect 1763 46775 1772 46809
rect 1720 46766 1772 46775
rect 89218 46809 89270 46818
rect 89218 46775 89227 46809
rect 89227 46775 89261 46809
rect 89261 46775 89270 46809
rect 89218 46766 89270 46775
rect 1720 46473 1772 46482
rect 1720 46439 1729 46473
rect 1729 46439 1763 46473
rect 1763 46439 1772 46473
rect 1720 46430 1772 46439
rect 89218 46473 89270 46482
rect 89218 46439 89227 46473
rect 89227 46439 89261 46473
rect 89261 46439 89270 46473
rect 89218 46430 89270 46439
rect 1720 46137 1772 46146
rect 1720 46103 1729 46137
rect 1729 46103 1763 46137
rect 1763 46103 1772 46137
rect 1720 46094 1772 46103
rect 89218 46137 89270 46146
rect 89218 46103 89227 46137
rect 89227 46103 89261 46137
rect 89261 46103 89270 46137
rect 89218 46094 89270 46103
rect 1720 45801 1772 45810
rect 1720 45767 1729 45801
rect 1729 45767 1763 45801
rect 1763 45767 1772 45801
rect 1720 45758 1772 45767
rect 89218 45801 89270 45810
rect 89218 45767 89227 45801
rect 89227 45767 89261 45801
rect 89261 45767 89270 45801
rect 89218 45758 89270 45767
rect 1720 45465 1772 45474
rect 1720 45431 1729 45465
rect 1729 45431 1763 45465
rect 1763 45431 1772 45465
rect 1720 45422 1772 45431
rect 89218 45465 89270 45474
rect 89218 45431 89227 45465
rect 89227 45431 89261 45465
rect 89261 45431 89270 45465
rect 89218 45422 89270 45431
rect 1720 45129 1772 45138
rect 1720 45095 1729 45129
rect 1729 45095 1763 45129
rect 1763 45095 1772 45129
rect 1720 45086 1772 45095
rect 89218 45129 89270 45138
rect 89218 45095 89227 45129
rect 89227 45095 89261 45129
rect 89261 45095 89270 45129
rect 89218 45086 89270 45095
rect 1720 44793 1772 44802
rect 1720 44759 1729 44793
rect 1729 44759 1763 44793
rect 1763 44759 1772 44793
rect 1720 44750 1772 44759
rect 89218 44793 89270 44802
rect 89218 44759 89227 44793
rect 89227 44759 89261 44793
rect 89261 44759 89270 44793
rect 89218 44750 89270 44759
rect 1720 44457 1772 44466
rect 1720 44423 1729 44457
rect 1729 44423 1763 44457
rect 1763 44423 1772 44457
rect 1720 44414 1772 44423
rect 89218 44457 89270 44466
rect 89218 44423 89227 44457
rect 89227 44423 89261 44457
rect 89261 44423 89270 44457
rect 89218 44414 89270 44423
rect 1720 44121 1772 44130
rect 1720 44087 1729 44121
rect 1729 44087 1763 44121
rect 1763 44087 1772 44121
rect 1720 44078 1772 44087
rect 89218 44121 89270 44130
rect 89218 44087 89227 44121
rect 89227 44087 89261 44121
rect 89261 44087 89270 44121
rect 89218 44078 89270 44087
rect 1720 43785 1772 43794
rect 1720 43751 1729 43785
rect 1729 43751 1763 43785
rect 1763 43751 1772 43785
rect 1720 43742 1772 43751
rect 89218 43785 89270 43794
rect 89218 43751 89227 43785
rect 89227 43751 89261 43785
rect 89261 43751 89270 43785
rect 89218 43742 89270 43751
rect 1720 43449 1772 43458
rect 1720 43415 1729 43449
rect 1729 43415 1763 43449
rect 1763 43415 1772 43449
rect 1720 43406 1772 43415
rect 89218 43449 89270 43458
rect 89218 43415 89227 43449
rect 89227 43415 89261 43449
rect 89261 43415 89270 43449
rect 89218 43406 89270 43415
rect 1720 43113 1772 43122
rect 1720 43079 1729 43113
rect 1729 43079 1763 43113
rect 1763 43079 1772 43113
rect 1720 43070 1772 43079
rect 89218 43113 89270 43122
rect 89218 43079 89227 43113
rect 89227 43079 89261 43113
rect 89261 43079 89270 43113
rect 89218 43070 89270 43079
rect 1720 42777 1772 42786
rect 1720 42743 1729 42777
rect 1729 42743 1763 42777
rect 1763 42743 1772 42777
rect 1720 42734 1772 42743
rect 89218 42777 89270 42786
rect 89218 42743 89227 42777
rect 89227 42743 89261 42777
rect 89261 42743 89270 42777
rect 89218 42734 89270 42743
rect 1720 42441 1772 42450
rect 1720 42407 1729 42441
rect 1729 42407 1763 42441
rect 1763 42407 1772 42441
rect 1720 42398 1772 42407
rect 89218 42441 89270 42450
rect 89218 42407 89227 42441
rect 89227 42407 89261 42441
rect 89261 42407 89270 42441
rect 89218 42398 89270 42407
rect 1720 42105 1772 42114
rect 1720 42071 1729 42105
rect 1729 42071 1763 42105
rect 1763 42071 1772 42105
rect 1720 42062 1772 42071
rect 89218 42105 89270 42114
rect 89218 42071 89227 42105
rect 89227 42071 89261 42105
rect 89261 42071 89270 42105
rect 89218 42062 89270 42071
rect 1720 41769 1772 41778
rect 1720 41735 1729 41769
rect 1729 41735 1763 41769
rect 1763 41735 1772 41769
rect 1720 41726 1772 41735
rect 89218 41769 89270 41778
rect 89218 41735 89227 41769
rect 89227 41735 89261 41769
rect 89261 41735 89270 41769
rect 89218 41726 89270 41735
rect 1720 41433 1772 41442
rect 1720 41399 1729 41433
rect 1729 41399 1763 41433
rect 1763 41399 1772 41433
rect 1720 41390 1772 41399
rect 89218 41433 89270 41442
rect 89218 41399 89227 41433
rect 89227 41399 89261 41433
rect 89261 41399 89270 41433
rect 89218 41390 89270 41399
rect 1720 41097 1772 41106
rect 1720 41063 1729 41097
rect 1729 41063 1763 41097
rect 1763 41063 1772 41097
rect 1720 41054 1772 41063
rect 89218 41097 89270 41106
rect 89218 41063 89227 41097
rect 89227 41063 89261 41097
rect 89261 41063 89270 41097
rect 89218 41054 89270 41063
rect 1720 40761 1772 40770
rect 1720 40727 1729 40761
rect 1729 40727 1763 40761
rect 1763 40727 1772 40761
rect 1720 40718 1772 40727
rect 89218 40761 89270 40770
rect 89218 40727 89227 40761
rect 89227 40727 89261 40761
rect 89261 40727 89270 40761
rect 89218 40718 89270 40727
rect 1720 40425 1772 40434
rect 1720 40391 1729 40425
rect 1729 40391 1763 40425
rect 1763 40391 1772 40425
rect 1720 40382 1772 40391
rect 89218 40425 89270 40434
rect 89218 40391 89227 40425
rect 89227 40391 89261 40425
rect 89261 40391 89270 40425
rect 89218 40382 89270 40391
rect 1720 40089 1772 40098
rect 1720 40055 1729 40089
rect 1729 40055 1763 40089
rect 1763 40055 1772 40089
rect 1720 40046 1772 40055
rect 89218 40089 89270 40098
rect 89218 40055 89227 40089
rect 89227 40055 89261 40089
rect 89261 40055 89270 40089
rect 89218 40046 89270 40055
rect 1720 39753 1772 39762
rect 1720 39719 1729 39753
rect 1729 39719 1763 39753
rect 1763 39719 1772 39753
rect 1720 39710 1772 39719
rect 89218 39753 89270 39762
rect 89218 39719 89227 39753
rect 89227 39719 89261 39753
rect 89261 39719 89270 39753
rect 89218 39710 89270 39719
rect 1720 39417 1772 39426
rect 1720 39383 1729 39417
rect 1729 39383 1763 39417
rect 1763 39383 1772 39417
rect 1720 39374 1772 39383
rect 89218 39417 89270 39426
rect 89218 39383 89227 39417
rect 89227 39383 89261 39417
rect 89261 39383 89270 39417
rect 89218 39374 89270 39383
rect 1720 39081 1772 39090
rect 1720 39047 1729 39081
rect 1729 39047 1763 39081
rect 1763 39047 1772 39081
rect 1720 39038 1772 39047
rect 89218 39081 89270 39090
rect 89218 39047 89227 39081
rect 89227 39047 89261 39081
rect 89261 39047 89270 39081
rect 89218 39038 89270 39047
rect 1720 38745 1772 38754
rect 1720 38711 1729 38745
rect 1729 38711 1763 38745
rect 1763 38711 1772 38745
rect 1720 38702 1772 38711
rect 89218 38745 89270 38754
rect 89218 38711 89227 38745
rect 89227 38711 89261 38745
rect 89261 38711 89270 38745
rect 89218 38702 89270 38711
rect 1720 38409 1772 38418
rect 1720 38375 1729 38409
rect 1729 38375 1763 38409
rect 1763 38375 1772 38409
rect 1720 38366 1772 38375
rect 89218 38409 89270 38418
rect 89218 38375 89227 38409
rect 89227 38375 89261 38409
rect 89261 38375 89270 38409
rect 89218 38366 89270 38375
rect 1720 38073 1772 38082
rect 1720 38039 1729 38073
rect 1729 38039 1763 38073
rect 1763 38039 1772 38073
rect 1720 38030 1772 38039
rect 89218 38073 89270 38082
rect 89218 38039 89227 38073
rect 89227 38039 89261 38073
rect 89261 38039 89270 38073
rect 89218 38030 89270 38039
rect 1720 37737 1772 37746
rect 1720 37703 1729 37737
rect 1729 37703 1763 37737
rect 1763 37703 1772 37737
rect 1720 37694 1772 37703
rect 89218 37737 89270 37746
rect 89218 37703 89227 37737
rect 89227 37703 89261 37737
rect 89261 37703 89270 37737
rect 89218 37694 89270 37703
rect 1720 37401 1772 37410
rect 1720 37367 1729 37401
rect 1729 37367 1763 37401
rect 1763 37367 1772 37401
rect 1720 37358 1772 37367
rect 89218 37401 89270 37410
rect 89218 37367 89227 37401
rect 89227 37367 89261 37401
rect 89261 37367 89270 37401
rect 89218 37358 89270 37367
rect 12357 37206 12409 37258
rect 1720 37065 1772 37074
rect 1720 37031 1729 37065
rect 1729 37031 1763 37065
rect 1763 37031 1772 37065
rect 1720 37022 1772 37031
rect 1720 36729 1772 36738
rect 1720 36695 1729 36729
rect 1729 36695 1763 36729
rect 1763 36695 1772 36729
rect 1720 36686 1772 36695
rect 1720 36393 1772 36402
rect 1720 36359 1729 36393
rect 1729 36359 1763 36393
rect 1763 36359 1772 36393
rect 1720 36350 1772 36359
rect 1720 36057 1772 36066
rect 1720 36023 1729 36057
rect 1729 36023 1763 36057
rect 1763 36023 1772 36057
rect 1720 36014 1772 36023
rect 12277 35936 12329 35988
rect 1720 35721 1772 35730
rect 1720 35687 1729 35721
rect 1729 35687 1763 35721
rect 1763 35687 1772 35721
rect 1720 35678 1772 35687
rect 1720 35385 1772 35394
rect 1720 35351 1729 35385
rect 1729 35351 1763 35385
rect 1763 35351 1772 35385
rect 1720 35342 1772 35351
rect 1720 35049 1772 35058
rect 1720 35015 1729 35049
rect 1729 35015 1763 35049
rect 1763 35015 1772 35049
rect 1720 35006 1772 35015
rect 1720 34713 1772 34722
rect 1720 34679 1729 34713
rect 1729 34679 1763 34713
rect 1763 34679 1772 34713
rect 1720 34670 1772 34679
rect 1720 34377 1772 34386
rect 1720 34343 1729 34377
rect 1729 34343 1763 34377
rect 1763 34343 1772 34377
rect 1720 34334 1772 34343
rect 12197 34378 12249 34430
rect 1720 34041 1772 34050
rect 1720 34007 1729 34041
rect 1729 34007 1763 34041
rect 1763 34007 1772 34041
rect 1720 33998 1772 34007
rect 1720 33705 1772 33714
rect 1720 33671 1729 33705
rect 1729 33671 1763 33705
rect 1763 33671 1772 33705
rect 1720 33662 1772 33671
rect 1720 33369 1772 33378
rect 1720 33335 1729 33369
rect 1729 33335 1763 33369
rect 1763 33335 1772 33369
rect 1720 33326 1772 33335
rect 12117 33108 12169 33160
rect 1720 33033 1772 33042
rect 1720 32999 1729 33033
rect 1729 32999 1763 33033
rect 1763 32999 1772 33033
rect 1720 32990 1772 32999
rect 1720 32697 1772 32706
rect 1720 32663 1729 32697
rect 1729 32663 1763 32697
rect 1763 32663 1772 32697
rect 1720 32654 1772 32663
rect 1720 32361 1772 32370
rect 1720 32327 1729 32361
rect 1729 32327 1763 32361
rect 1763 32327 1772 32361
rect 1720 32318 1772 32327
rect 1720 32025 1772 32034
rect 1720 31991 1729 32025
rect 1729 31991 1763 32025
rect 1763 31991 1772 32025
rect 1720 31982 1772 31991
rect 1720 31689 1772 31698
rect 1720 31655 1729 31689
rect 1729 31655 1763 31689
rect 1763 31655 1772 31689
rect 1720 31646 1772 31655
rect 12037 31550 12089 31602
rect 1720 31353 1772 31362
rect 1720 31319 1729 31353
rect 1729 31319 1763 31353
rect 1763 31319 1772 31353
rect 1720 31310 1772 31319
rect 1720 31017 1772 31026
rect 1720 30983 1729 31017
rect 1729 30983 1763 31017
rect 1763 30983 1772 31017
rect 1720 30974 1772 30983
rect 1720 30681 1772 30690
rect 1720 30647 1729 30681
rect 1729 30647 1763 30681
rect 1763 30647 1772 30681
rect 1720 30638 1772 30647
rect 1720 30345 1772 30354
rect 1720 30311 1729 30345
rect 1729 30311 1763 30345
rect 1763 30311 1772 30345
rect 1720 30302 1772 30311
rect 11957 30280 12009 30332
rect 1720 30009 1772 30018
rect 1720 29975 1729 30009
rect 1729 29975 1763 30009
rect 1763 29975 1772 30009
rect 1720 29966 1772 29975
rect 1720 29673 1772 29682
rect 1720 29639 1729 29673
rect 1729 29639 1763 29673
rect 1763 29639 1772 29673
rect 1720 29630 1772 29639
rect 1720 29337 1772 29346
rect 1720 29303 1729 29337
rect 1729 29303 1763 29337
rect 1763 29303 1772 29337
rect 1720 29294 1772 29303
rect 1720 29001 1772 29010
rect 1720 28967 1729 29001
rect 1729 28967 1763 29001
rect 1763 28967 1772 29001
rect 1720 28958 1772 28967
rect 11877 28722 11929 28774
rect 1720 28665 1772 28674
rect 1720 28631 1729 28665
rect 1729 28631 1763 28665
rect 1763 28631 1772 28665
rect 1720 28622 1772 28631
rect 1720 28329 1772 28338
rect 1720 28295 1729 28329
rect 1729 28295 1763 28329
rect 1763 28295 1772 28329
rect 1720 28286 1772 28295
rect 1720 27993 1772 28002
rect 1720 27959 1729 27993
rect 1729 27959 1763 27993
rect 1763 27959 1772 27993
rect 1720 27950 1772 27959
rect 1720 27657 1772 27666
rect 1720 27623 1729 27657
rect 1729 27623 1763 27657
rect 1763 27623 1772 27657
rect 1720 27614 1772 27623
rect 1720 27321 1772 27330
rect 1720 27287 1729 27321
rect 1729 27287 1763 27321
rect 1763 27287 1772 27321
rect 1720 27278 1772 27287
rect 1720 26985 1772 26994
rect 1720 26951 1729 26985
rect 1729 26951 1763 26985
rect 1763 26951 1772 26985
rect 1720 26942 1772 26951
rect 1720 26649 1772 26658
rect 1720 26615 1729 26649
rect 1729 26615 1763 26649
rect 1763 26615 1772 26649
rect 1720 26606 1772 26615
rect 1720 26313 1772 26322
rect 1720 26279 1729 26313
rect 1729 26279 1763 26313
rect 1763 26279 1772 26313
rect 1720 26270 1772 26279
rect 1720 25977 1772 25986
rect 1720 25943 1729 25977
rect 1729 25943 1763 25977
rect 1763 25943 1772 25977
rect 1720 25934 1772 25943
rect 1720 25641 1772 25650
rect 1720 25607 1729 25641
rect 1729 25607 1763 25641
rect 1763 25607 1772 25641
rect 1720 25598 1772 25607
rect 1720 25305 1772 25314
rect 1720 25271 1729 25305
rect 1729 25271 1763 25305
rect 1763 25271 1772 25305
rect 1720 25262 1772 25271
rect 1720 24969 1772 24978
rect 1720 24935 1729 24969
rect 1729 24935 1763 24969
rect 1763 24935 1772 24969
rect 1720 24926 1772 24935
rect 1720 24633 1772 24642
rect 1720 24599 1729 24633
rect 1729 24599 1763 24633
rect 1763 24599 1772 24633
rect 1720 24590 1772 24599
rect 1720 24297 1772 24306
rect 1720 24263 1729 24297
rect 1729 24263 1763 24297
rect 1763 24263 1772 24297
rect 1720 24254 1772 24263
rect 89218 37065 89270 37074
rect 89218 37031 89227 37065
rect 89227 37031 89261 37065
rect 89261 37031 89270 37065
rect 89218 37022 89270 37031
rect 89218 36729 89270 36738
rect 89218 36695 89227 36729
rect 89227 36695 89261 36729
rect 89261 36695 89270 36729
rect 89218 36686 89270 36695
rect 89218 36393 89270 36402
rect 89218 36359 89227 36393
rect 89227 36359 89261 36393
rect 89261 36359 89270 36393
rect 89218 36350 89270 36359
rect 89218 36057 89270 36066
rect 89218 36023 89227 36057
rect 89227 36023 89261 36057
rect 89261 36023 89270 36057
rect 89218 36014 89270 36023
rect 89218 35721 89270 35730
rect 89218 35687 89227 35721
rect 89227 35687 89261 35721
rect 89261 35687 89270 35721
rect 89218 35678 89270 35687
rect 89218 35385 89270 35394
rect 89218 35351 89227 35385
rect 89227 35351 89261 35385
rect 89261 35351 89270 35385
rect 89218 35342 89270 35351
rect 89218 35049 89270 35058
rect 89218 35015 89227 35049
rect 89227 35015 89261 35049
rect 89261 35015 89270 35049
rect 89218 35006 89270 35015
rect 89218 34713 89270 34722
rect 89218 34679 89227 34713
rect 89227 34679 89261 34713
rect 89261 34679 89270 34713
rect 89218 34670 89270 34679
rect 89218 34377 89270 34386
rect 89218 34343 89227 34377
rect 89227 34343 89261 34377
rect 89261 34343 89270 34377
rect 89218 34334 89270 34343
rect 89218 34041 89270 34050
rect 89218 34007 89227 34041
rect 89227 34007 89261 34041
rect 89261 34007 89270 34041
rect 89218 33998 89270 34007
rect 89218 33705 89270 33714
rect 89218 33671 89227 33705
rect 89227 33671 89261 33705
rect 89261 33671 89270 33705
rect 89218 33662 89270 33671
rect 89218 33369 89270 33378
rect 89218 33335 89227 33369
rect 89227 33335 89261 33369
rect 89261 33335 89270 33369
rect 89218 33326 89270 33335
rect 89218 33033 89270 33042
rect 89218 32999 89227 33033
rect 89227 32999 89261 33033
rect 89261 32999 89270 33033
rect 89218 32990 89270 32999
rect 89218 32697 89270 32706
rect 89218 32663 89227 32697
rect 89227 32663 89261 32697
rect 89261 32663 89270 32697
rect 89218 32654 89270 32663
rect 89218 32361 89270 32370
rect 89218 32327 89227 32361
rect 89227 32327 89261 32361
rect 89261 32327 89270 32361
rect 89218 32318 89270 32327
rect 89218 32025 89270 32034
rect 89218 31991 89227 32025
rect 89227 31991 89261 32025
rect 89261 31991 89270 32025
rect 89218 31982 89270 31991
rect 89218 31689 89270 31698
rect 89218 31655 89227 31689
rect 89227 31655 89261 31689
rect 89261 31655 89270 31689
rect 89218 31646 89270 31655
rect 89218 31353 89270 31362
rect 89218 31319 89227 31353
rect 89227 31319 89261 31353
rect 89261 31319 89270 31353
rect 89218 31310 89270 31319
rect 89218 31017 89270 31026
rect 89218 30983 89227 31017
rect 89227 30983 89261 31017
rect 89261 30983 89270 31017
rect 89218 30974 89270 30983
rect 89218 30681 89270 30690
rect 89218 30647 89227 30681
rect 89227 30647 89261 30681
rect 89261 30647 89270 30681
rect 89218 30638 89270 30647
rect 89218 30345 89270 30354
rect 89218 30311 89227 30345
rect 89227 30311 89261 30345
rect 89261 30311 89270 30345
rect 89218 30302 89270 30311
rect 89218 30009 89270 30018
rect 89218 29975 89227 30009
rect 89227 29975 89261 30009
rect 89261 29975 89270 30009
rect 89218 29966 89270 29975
rect 89218 29673 89270 29682
rect 89218 29639 89227 29673
rect 89227 29639 89261 29673
rect 89261 29639 89270 29673
rect 89218 29630 89270 29639
rect 89218 29337 89270 29346
rect 89218 29303 89227 29337
rect 89227 29303 89261 29337
rect 89261 29303 89270 29337
rect 89218 29294 89270 29303
rect 89218 29001 89270 29010
rect 89218 28967 89227 29001
rect 89227 28967 89261 29001
rect 89261 28967 89270 29001
rect 89218 28958 89270 28967
rect 89218 28665 89270 28674
rect 89218 28631 89227 28665
rect 89227 28631 89261 28665
rect 89261 28631 89270 28665
rect 89218 28622 89270 28631
rect 89218 28329 89270 28338
rect 89218 28295 89227 28329
rect 89227 28295 89261 28329
rect 89261 28295 89270 28329
rect 89218 28286 89270 28295
rect 89218 27993 89270 28002
rect 89218 27959 89227 27993
rect 89227 27959 89261 27993
rect 89261 27959 89270 27993
rect 89218 27950 89270 27959
rect 89218 27657 89270 27666
rect 89218 27623 89227 27657
rect 89227 27623 89261 27657
rect 89261 27623 89270 27657
rect 89218 27614 89270 27623
rect 89218 27321 89270 27330
rect 89218 27287 89227 27321
rect 89227 27287 89261 27321
rect 89261 27287 89270 27321
rect 89218 27278 89270 27287
rect 89218 26985 89270 26994
rect 89218 26951 89227 26985
rect 89227 26951 89261 26985
rect 89261 26951 89270 26985
rect 89218 26942 89270 26951
rect 89218 26649 89270 26658
rect 89218 26615 89227 26649
rect 89227 26615 89261 26649
rect 89261 26615 89270 26649
rect 89218 26606 89270 26615
rect 89218 26313 89270 26322
rect 89218 26279 89227 26313
rect 89227 26279 89261 26313
rect 89261 26279 89270 26313
rect 89218 26270 89270 26279
rect 89218 25977 89270 25986
rect 89218 25943 89227 25977
rect 89227 25943 89261 25977
rect 89261 25943 89270 25977
rect 89218 25934 89270 25943
rect 89218 25641 89270 25650
rect 89218 25607 89227 25641
rect 89227 25607 89261 25641
rect 89261 25607 89270 25641
rect 89218 25598 89270 25607
rect 89218 25305 89270 25314
rect 89218 25271 89227 25305
rect 89227 25271 89261 25305
rect 89261 25271 89270 25305
rect 89218 25262 89270 25271
rect 89218 24969 89270 24978
rect 89218 24935 89227 24969
rect 89227 24935 89261 24969
rect 89261 24935 89270 24969
rect 89218 24926 89270 24935
rect 89218 24633 89270 24642
rect 89218 24599 89227 24633
rect 89227 24599 89261 24633
rect 89261 24599 89270 24633
rect 89218 24590 89270 24599
rect 89218 24297 89270 24306
rect 89218 24263 89227 24297
rect 89227 24263 89261 24297
rect 89261 24263 89270 24297
rect 89218 24254 89270 24263
rect 1720 23961 1772 23970
rect 1720 23927 1729 23961
rect 1729 23927 1763 23961
rect 1763 23927 1772 23961
rect 1720 23918 1772 23927
rect 1720 23625 1772 23634
rect 1720 23591 1729 23625
rect 1729 23591 1763 23625
rect 1763 23591 1772 23625
rect 1720 23582 1772 23591
rect 1720 23289 1772 23298
rect 1720 23255 1729 23289
rect 1729 23255 1763 23289
rect 1763 23255 1772 23289
rect 1720 23246 1772 23255
rect 1720 22953 1772 22962
rect 1720 22919 1729 22953
rect 1729 22919 1763 22953
rect 1763 22919 1772 22953
rect 1720 22910 1772 22919
rect 1720 22617 1772 22626
rect 1720 22583 1729 22617
rect 1729 22583 1763 22617
rect 1763 22583 1772 22617
rect 1720 22574 1772 22583
rect 1720 22281 1772 22290
rect 1720 22247 1729 22281
rect 1729 22247 1763 22281
rect 1763 22247 1772 22281
rect 1720 22238 1772 22247
rect 1720 21945 1772 21954
rect 1720 21911 1729 21945
rect 1729 21911 1763 21945
rect 1763 21911 1772 21945
rect 1720 21902 1772 21911
rect 1720 21609 1772 21618
rect 1720 21575 1729 21609
rect 1729 21575 1763 21609
rect 1763 21575 1772 21609
rect 1720 21566 1772 21575
rect 1720 21273 1772 21282
rect 1720 21239 1729 21273
rect 1729 21239 1763 21273
rect 1763 21239 1772 21273
rect 1720 21230 1772 21239
rect 1720 20937 1772 20946
rect 1720 20903 1729 20937
rect 1729 20903 1763 20937
rect 1763 20903 1772 20937
rect 1720 20894 1772 20903
rect 1720 20601 1772 20610
rect 1720 20567 1729 20601
rect 1729 20567 1763 20601
rect 1763 20567 1772 20601
rect 1720 20558 1772 20567
rect 1720 20265 1772 20274
rect 1720 20231 1729 20265
rect 1729 20231 1763 20265
rect 1763 20231 1772 20265
rect 1720 20222 1772 20231
rect 1720 19929 1772 19938
rect 1720 19895 1729 19929
rect 1729 19895 1763 19929
rect 1763 19895 1772 19929
rect 1720 19886 1772 19895
rect 1720 19593 1772 19602
rect 1720 19559 1729 19593
rect 1729 19559 1763 19593
rect 1763 19559 1772 19593
rect 1720 19550 1772 19559
rect 1720 19257 1772 19266
rect 1720 19223 1729 19257
rect 1729 19223 1763 19257
rect 1763 19223 1772 19257
rect 1720 19214 1772 19223
rect 1720 18921 1772 18930
rect 1720 18887 1729 18921
rect 1729 18887 1763 18921
rect 1763 18887 1772 18921
rect 1720 18878 1772 18887
rect 1720 18585 1772 18594
rect 1720 18551 1729 18585
rect 1729 18551 1763 18585
rect 1763 18551 1772 18585
rect 1720 18542 1772 18551
rect 1720 18249 1772 18258
rect 1720 18215 1729 18249
rect 1729 18215 1763 18249
rect 1763 18215 1772 18249
rect 1720 18206 1772 18215
rect 1720 17913 1772 17922
rect 1720 17879 1729 17913
rect 1729 17879 1763 17913
rect 1763 17879 1772 17913
rect 1720 17870 1772 17879
rect 1720 17577 1772 17586
rect 1720 17543 1729 17577
rect 1729 17543 1763 17577
rect 1763 17543 1772 17577
rect 1720 17534 1772 17543
rect 1720 17241 1772 17250
rect 1720 17207 1729 17241
rect 1729 17207 1763 17241
rect 1763 17207 1772 17241
rect 1720 17198 1772 17207
rect 1720 16905 1772 16914
rect 1720 16871 1729 16905
rect 1729 16871 1763 16905
rect 1763 16871 1772 16905
rect 1720 16862 1772 16871
rect 1720 16569 1772 16578
rect 1720 16535 1729 16569
rect 1729 16535 1763 16569
rect 1763 16535 1772 16569
rect 1720 16526 1772 16535
rect 1720 16233 1772 16242
rect 1720 16199 1729 16233
rect 1729 16199 1763 16233
rect 1763 16199 1772 16233
rect 1720 16190 1772 16199
rect 1720 15897 1772 15906
rect 1720 15863 1729 15897
rect 1729 15863 1763 15897
rect 1763 15863 1772 15897
rect 1720 15854 1772 15863
rect 1720 15561 1772 15570
rect 1720 15527 1729 15561
rect 1729 15527 1763 15561
rect 1763 15527 1772 15561
rect 1720 15518 1772 15527
rect 1720 15225 1772 15234
rect 1720 15191 1729 15225
rect 1729 15191 1763 15225
rect 1763 15191 1772 15225
rect 1720 15182 1772 15191
rect 1720 14889 1772 14898
rect 1720 14855 1729 14889
rect 1729 14855 1763 14889
rect 1763 14855 1772 14889
rect 1720 14846 1772 14855
rect 1720 14553 1772 14562
rect 1720 14519 1729 14553
rect 1729 14519 1763 14553
rect 1763 14519 1772 14553
rect 1720 14510 1772 14519
rect 1720 14217 1772 14226
rect 1720 14183 1729 14217
rect 1729 14183 1763 14217
rect 1763 14183 1772 14217
rect 1720 14174 1772 14183
rect 1720 13881 1772 13890
rect 1720 13847 1729 13881
rect 1729 13847 1763 13881
rect 1763 13847 1772 13881
rect 1720 13838 1772 13847
rect 1720 13545 1772 13554
rect 1720 13511 1729 13545
rect 1729 13511 1763 13545
rect 1763 13511 1772 13545
rect 1720 13502 1772 13511
rect 1720 13209 1772 13218
rect 1720 13175 1729 13209
rect 1729 13175 1763 13209
rect 1763 13175 1772 13209
rect 1720 13166 1772 13175
rect 25628 13078 25680 13130
rect 30620 13078 30672 13130
rect 35612 13078 35664 13130
rect 40604 13078 40656 13130
rect 45596 13078 45648 13130
rect 50588 13078 50640 13130
rect 55580 13078 55632 13130
rect 60572 13078 60624 13130
rect 1720 12873 1772 12882
rect 1720 12839 1729 12873
rect 1729 12839 1763 12873
rect 1763 12839 1772 12873
rect 1720 12830 1772 12839
rect 1720 12537 1772 12546
rect 1720 12503 1729 12537
rect 1729 12503 1763 12537
rect 1763 12503 1772 12537
rect 1720 12494 1772 12503
rect 1720 12201 1772 12210
rect 1720 12167 1729 12201
rect 1729 12167 1763 12201
rect 1763 12167 1772 12201
rect 1720 12158 1772 12167
rect 1720 11865 1772 11874
rect 1720 11831 1729 11865
rect 1729 11831 1763 11865
rect 1763 11831 1772 11865
rect 1720 11822 1772 11831
rect 1720 11529 1772 11538
rect 1720 11495 1729 11529
rect 1729 11495 1763 11529
rect 1763 11495 1772 11529
rect 1720 11486 1772 11495
rect 1720 11193 1772 11202
rect 1720 11159 1729 11193
rect 1729 11159 1763 11193
rect 1763 11159 1772 11193
rect 1720 11150 1772 11159
rect 89218 23961 89270 23970
rect 89218 23927 89227 23961
rect 89227 23927 89261 23961
rect 89261 23927 89270 23961
rect 89218 23918 89270 23927
rect 89218 23625 89270 23634
rect 89218 23591 89227 23625
rect 89227 23591 89261 23625
rect 89261 23591 89270 23625
rect 89218 23582 89270 23591
rect 89218 23289 89270 23298
rect 89218 23255 89227 23289
rect 89227 23255 89261 23289
rect 89261 23255 89270 23289
rect 89218 23246 89270 23255
rect 89218 22953 89270 22962
rect 89218 22919 89227 22953
rect 89227 22919 89261 22953
rect 89261 22919 89270 22953
rect 89218 22910 89270 22919
rect 89218 22617 89270 22626
rect 89218 22583 89227 22617
rect 89227 22583 89261 22617
rect 89261 22583 89270 22617
rect 89218 22574 89270 22583
rect 89218 22281 89270 22290
rect 89218 22247 89227 22281
rect 89227 22247 89261 22281
rect 89261 22247 89270 22281
rect 89218 22238 89270 22247
rect 89218 21945 89270 21954
rect 89218 21911 89227 21945
rect 89227 21911 89261 21945
rect 89261 21911 89270 21945
rect 89218 21902 89270 21911
rect 89218 21609 89270 21618
rect 89218 21575 89227 21609
rect 89227 21575 89261 21609
rect 89261 21575 89270 21609
rect 89218 21566 89270 21575
rect 89218 21273 89270 21282
rect 89218 21239 89227 21273
rect 89227 21239 89261 21273
rect 89261 21239 89270 21273
rect 89218 21230 89270 21239
rect 89218 20937 89270 20946
rect 89218 20903 89227 20937
rect 89227 20903 89261 20937
rect 89261 20903 89270 20937
rect 89218 20894 89270 20903
rect 89218 20601 89270 20610
rect 89218 20567 89227 20601
rect 89227 20567 89261 20601
rect 89261 20567 89270 20601
rect 89218 20558 89270 20567
rect 89218 20265 89270 20274
rect 89218 20231 89227 20265
rect 89227 20231 89261 20265
rect 89261 20231 89270 20265
rect 89218 20222 89270 20231
rect 89218 19929 89270 19938
rect 89218 19895 89227 19929
rect 89227 19895 89261 19929
rect 89261 19895 89270 19929
rect 89218 19886 89270 19895
rect 79061 19552 79113 19604
rect 89218 19593 89270 19602
rect 89218 19559 89227 19593
rect 89227 19559 89261 19593
rect 89261 19559 89270 19593
rect 89218 19550 89270 19559
rect 89218 19257 89270 19266
rect 89218 19223 89227 19257
rect 89227 19223 89261 19257
rect 89261 19223 89270 19257
rect 89218 19214 89270 19223
rect 89218 18921 89270 18930
rect 89218 18887 89227 18921
rect 89227 18887 89261 18921
rect 89261 18887 89270 18921
rect 89218 18878 89270 18887
rect 89218 18585 89270 18594
rect 89218 18551 89227 18585
rect 89227 18551 89261 18585
rect 89261 18551 89270 18585
rect 89218 18542 89270 18551
rect 89218 18249 89270 18258
rect 89218 18215 89227 18249
rect 89227 18215 89261 18249
rect 89261 18215 89270 18249
rect 89218 18206 89270 18215
rect 78981 17994 79033 18046
rect 89218 17913 89270 17922
rect 89218 17879 89227 17913
rect 89227 17879 89261 17913
rect 89261 17879 89270 17913
rect 89218 17870 89270 17879
rect 89218 17577 89270 17586
rect 89218 17543 89227 17577
rect 89227 17543 89261 17577
rect 89261 17543 89270 17577
rect 89218 17534 89270 17543
rect 89218 17241 89270 17250
rect 89218 17207 89227 17241
rect 89227 17207 89261 17241
rect 89261 17207 89270 17241
rect 89218 17198 89270 17207
rect 89218 16905 89270 16914
rect 89218 16871 89227 16905
rect 89227 16871 89261 16905
rect 89261 16871 89270 16905
rect 89218 16862 89270 16871
rect 78901 16724 78953 16776
rect 89218 16569 89270 16578
rect 89218 16535 89227 16569
rect 89227 16535 89261 16569
rect 89261 16535 89270 16569
rect 89218 16526 89270 16535
rect 89218 16233 89270 16242
rect 89218 16199 89227 16233
rect 89227 16199 89261 16233
rect 89261 16199 89270 16233
rect 89218 16190 89270 16199
rect 89218 15897 89270 15906
rect 89218 15863 89227 15897
rect 89227 15863 89261 15897
rect 89261 15863 89270 15897
rect 89218 15854 89270 15863
rect 89218 15561 89270 15570
rect 89218 15527 89227 15561
rect 89227 15527 89261 15561
rect 89261 15527 89270 15561
rect 89218 15518 89270 15527
rect 78821 15166 78873 15218
rect 89218 15225 89270 15234
rect 89218 15191 89227 15225
rect 89227 15191 89261 15225
rect 89261 15191 89270 15225
rect 89218 15182 89270 15191
rect 89218 14889 89270 14898
rect 89218 14855 89227 14889
rect 89227 14855 89261 14889
rect 89261 14855 89270 14889
rect 89218 14846 89270 14855
rect 89218 14553 89270 14562
rect 89218 14519 89227 14553
rect 89227 14519 89261 14553
rect 89261 14519 89270 14553
rect 89218 14510 89270 14519
rect 89218 14217 89270 14226
rect 89218 14183 89227 14217
rect 89227 14183 89261 14217
rect 89261 14183 89270 14217
rect 89218 14174 89270 14183
rect 78741 13896 78793 13948
rect 89218 13881 89270 13890
rect 89218 13847 89227 13881
rect 89227 13847 89261 13881
rect 89261 13847 89270 13881
rect 89218 13838 89270 13847
rect 89218 13545 89270 13554
rect 89218 13511 89227 13545
rect 89227 13511 89261 13545
rect 89261 13511 89270 13545
rect 89218 13502 89270 13511
rect 89218 13209 89270 13218
rect 89218 13175 89227 13209
rect 89227 13175 89261 13209
rect 89261 13175 89270 13209
rect 89218 13166 89270 13175
rect 89218 12873 89270 12882
rect 89218 12839 89227 12873
rect 89227 12839 89261 12873
rect 89261 12839 89270 12873
rect 89218 12830 89270 12839
rect 89218 12537 89270 12546
rect 89218 12503 89227 12537
rect 89227 12503 89261 12537
rect 89261 12503 89270 12537
rect 89218 12494 89270 12503
rect 78661 12338 78713 12390
rect 89218 12201 89270 12210
rect 89218 12167 89227 12201
rect 89227 12167 89261 12201
rect 89261 12167 89270 12201
rect 89218 12158 89270 12167
rect 89218 11865 89270 11874
rect 89218 11831 89227 11865
rect 89227 11831 89261 11865
rect 89261 11831 89270 11865
rect 89218 11822 89270 11831
rect 89218 11529 89270 11538
rect 89218 11495 89227 11529
rect 89227 11495 89261 11529
rect 89261 11495 89270 11529
rect 89218 11486 89270 11495
rect 89218 11193 89270 11202
rect 89218 11159 89227 11193
rect 89227 11159 89261 11193
rect 89261 11159 89270 11193
rect 89218 11150 89270 11159
rect 78581 11068 78633 11120
rect 1720 10857 1772 10866
rect 1720 10823 1729 10857
rect 1729 10823 1763 10857
rect 1763 10823 1772 10857
rect 1720 10814 1772 10823
rect 89218 10857 89270 10866
rect 89218 10823 89227 10857
rect 89227 10823 89261 10857
rect 89261 10823 89270 10857
rect 89218 10814 89270 10823
rect 1720 10521 1772 10530
rect 1720 10487 1729 10521
rect 1729 10487 1763 10521
rect 1763 10487 1772 10521
rect 1720 10478 1772 10487
rect 89218 10521 89270 10530
rect 89218 10487 89227 10521
rect 89227 10487 89261 10521
rect 89261 10487 89270 10521
rect 89218 10478 89270 10487
rect 1720 10185 1772 10194
rect 1720 10151 1729 10185
rect 1729 10151 1763 10185
rect 1763 10151 1772 10185
rect 1720 10142 1772 10151
rect 89218 10185 89270 10194
rect 89218 10151 89227 10185
rect 89227 10151 89261 10185
rect 89261 10151 89270 10185
rect 89218 10142 89270 10151
rect 1720 9849 1772 9858
rect 1720 9815 1729 9849
rect 1729 9815 1763 9849
rect 1763 9815 1772 9849
rect 1720 9806 1772 9815
rect 89218 9849 89270 9858
rect 89218 9815 89227 9849
rect 89227 9815 89261 9849
rect 89261 9815 89270 9849
rect 89218 9806 89270 9815
rect 1720 9513 1772 9522
rect 1720 9479 1729 9513
rect 1729 9479 1763 9513
rect 1763 9479 1772 9513
rect 1720 9470 1772 9479
rect 89218 9513 89270 9522
rect 89218 9479 89227 9513
rect 89227 9479 89261 9513
rect 89261 9479 89270 9513
rect 89218 9470 89270 9479
rect 1720 9177 1772 9186
rect 1720 9143 1729 9177
rect 1729 9143 1763 9177
rect 1763 9143 1772 9177
rect 1720 9134 1772 9143
rect 89218 9177 89270 9186
rect 89218 9143 89227 9177
rect 89227 9143 89261 9177
rect 89261 9143 89270 9177
rect 89218 9134 89270 9143
rect 1720 8841 1772 8850
rect 1720 8807 1729 8841
rect 1729 8807 1763 8841
rect 1763 8807 1772 8841
rect 1720 8798 1772 8807
rect 89218 8841 89270 8850
rect 89218 8807 89227 8841
rect 89227 8807 89261 8841
rect 89261 8807 89270 8841
rect 89218 8798 89270 8807
rect 1720 8505 1772 8514
rect 1720 8471 1729 8505
rect 1729 8471 1763 8505
rect 1763 8471 1772 8505
rect 1720 8462 1772 8471
rect 89218 8505 89270 8514
rect 89218 8471 89227 8505
rect 89227 8471 89261 8505
rect 89261 8471 89270 8505
rect 89218 8462 89270 8471
rect 1720 8169 1772 8178
rect 1720 8135 1729 8169
rect 1729 8135 1763 8169
rect 1763 8135 1772 8169
rect 1720 8126 1772 8135
rect 89218 8169 89270 8178
rect 89218 8135 89227 8169
rect 89227 8135 89261 8169
rect 89261 8135 89270 8169
rect 89218 8126 89270 8135
rect 1720 7833 1772 7842
rect 1720 7799 1729 7833
rect 1729 7799 1763 7833
rect 1763 7799 1772 7833
rect 1720 7790 1772 7799
rect 89218 7833 89270 7842
rect 89218 7799 89227 7833
rect 89227 7799 89261 7833
rect 89261 7799 89270 7833
rect 89218 7790 89270 7799
rect 1720 7497 1772 7506
rect 1720 7463 1729 7497
rect 1729 7463 1763 7497
rect 1763 7463 1772 7497
rect 1720 7454 1772 7463
rect 89218 7497 89270 7506
rect 89218 7463 89227 7497
rect 89227 7463 89261 7497
rect 89261 7463 89270 7497
rect 89218 7454 89270 7463
rect 1720 7161 1772 7170
rect 1720 7127 1729 7161
rect 1729 7127 1763 7161
rect 1763 7127 1772 7161
rect 1720 7118 1772 7127
rect 89218 7161 89270 7170
rect 89218 7127 89227 7161
rect 89227 7127 89261 7161
rect 89261 7127 89270 7161
rect 89218 7118 89270 7127
rect 1720 6825 1772 6834
rect 1720 6791 1729 6825
rect 1729 6791 1763 6825
rect 1763 6791 1772 6825
rect 1720 6782 1772 6791
rect 89218 6825 89270 6834
rect 89218 6791 89227 6825
rect 89227 6791 89261 6825
rect 89261 6791 89270 6825
rect 89218 6782 89270 6791
rect 1720 6489 1772 6498
rect 1720 6455 1729 6489
rect 1729 6455 1763 6489
rect 1763 6455 1772 6489
rect 1720 6446 1772 6455
rect 89218 6489 89270 6498
rect 89218 6455 89227 6489
rect 89227 6455 89261 6489
rect 89261 6455 89270 6489
rect 89218 6446 89270 6455
rect 1720 6153 1772 6162
rect 1720 6119 1729 6153
rect 1729 6119 1763 6153
rect 1763 6119 1772 6153
rect 1720 6110 1772 6119
rect 89218 6153 89270 6162
rect 89218 6119 89227 6153
rect 89227 6119 89261 6153
rect 89261 6119 89270 6153
rect 89218 6110 89270 6119
rect 1720 5817 1772 5826
rect 1720 5783 1729 5817
rect 1729 5783 1763 5817
rect 1763 5783 1772 5817
rect 1720 5774 1772 5783
rect 89218 5817 89270 5826
rect 89218 5783 89227 5817
rect 89227 5783 89261 5817
rect 89261 5783 89270 5817
rect 89218 5774 89270 5783
rect 1720 5481 1772 5490
rect 1720 5447 1729 5481
rect 1729 5447 1763 5481
rect 1763 5447 1772 5481
rect 1720 5438 1772 5447
rect 89218 5481 89270 5490
rect 89218 5447 89227 5481
rect 89227 5447 89261 5481
rect 89261 5447 89270 5481
rect 89218 5438 89270 5447
rect 1720 5145 1772 5154
rect 1720 5111 1729 5145
rect 1729 5111 1763 5145
rect 1763 5111 1772 5145
rect 1720 5102 1772 5111
rect 89218 5145 89270 5154
rect 89218 5111 89227 5145
rect 89227 5111 89261 5145
rect 89261 5111 89270 5145
rect 89218 5102 89270 5111
rect 1720 4809 1772 4818
rect 1720 4775 1729 4809
rect 1729 4775 1763 4809
rect 1763 4775 1772 4809
rect 1720 4766 1772 4775
rect 89218 4809 89270 4818
rect 89218 4775 89227 4809
rect 89227 4775 89261 4809
rect 89261 4775 89270 4809
rect 89218 4766 89270 4775
rect 1720 4473 1772 4482
rect 1720 4439 1729 4473
rect 1729 4439 1763 4473
rect 1763 4439 1772 4473
rect 1720 4430 1772 4439
rect 89218 4473 89270 4482
rect 89218 4439 89227 4473
rect 89227 4439 89261 4473
rect 89261 4439 89270 4473
rect 89218 4430 89270 4439
rect 1720 4137 1772 4146
rect 1720 4103 1729 4137
rect 1729 4103 1763 4137
rect 1763 4103 1772 4137
rect 1720 4094 1772 4103
rect 89218 4137 89270 4146
rect 89218 4103 89227 4137
rect 89227 4103 89261 4137
rect 89261 4103 89270 4137
rect 89218 4094 89270 4103
rect 1720 3801 1772 3810
rect 1720 3767 1729 3801
rect 1729 3767 1763 3801
rect 1763 3767 1772 3801
rect 1720 3758 1772 3767
rect 89218 3801 89270 3810
rect 89218 3767 89227 3801
rect 89227 3767 89261 3801
rect 89261 3767 89270 3801
rect 89218 3758 89270 3767
rect 1720 3465 1772 3474
rect 1720 3431 1729 3465
rect 1729 3431 1763 3465
rect 1763 3431 1772 3465
rect 1720 3422 1772 3431
rect 89218 3465 89270 3474
rect 89218 3431 89227 3465
rect 89227 3431 89261 3465
rect 89261 3431 89270 3465
rect 89218 3422 89270 3431
rect 1720 3129 1772 3138
rect 1720 3095 1729 3129
rect 1729 3095 1763 3129
rect 1763 3095 1772 3129
rect 1720 3086 1772 3095
rect 89218 3129 89270 3138
rect 89218 3095 89227 3129
rect 89227 3095 89261 3129
rect 89261 3095 89270 3129
rect 89218 3086 89270 3095
rect 1720 2793 1772 2802
rect 1720 2759 1729 2793
rect 1729 2759 1763 2793
rect 1763 2759 1772 2793
rect 1720 2750 1772 2759
rect 89218 2793 89270 2802
rect 89218 2759 89227 2793
rect 89227 2759 89261 2793
rect 89261 2759 89270 2793
rect 89218 2750 89270 2759
rect 1720 2457 1772 2466
rect 1720 2423 1729 2457
rect 1729 2423 1763 2457
rect 1763 2423 1772 2457
rect 1720 2414 1772 2423
rect 89218 2457 89270 2466
rect 89218 2423 89227 2457
rect 89227 2423 89261 2457
rect 89261 2423 89270 2457
rect 89218 2414 89270 2423
rect 1720 2121 1772 2130
rect 1720 2087 1729 2121
rect 1729 2087 1763 2121
rect 1763 2087 1772 2121
rect 1720 2078 1772 2087
rect 89218 2121 89270 2130
rect 89218 2087 89227 2121
rect 89227 2087 89261 2121
rect 89261 2087 89270 2121
rect 89218 2078 89270 2087
rect 2056 1785 2108 1794
rect 3736 1785 3788 1794
rect 5416 1785 5468 1794
rect 7096 1785 7148 1794
rect 8776 1785 8828 1794
rect 10456 1785 10508 1794
rect 12136 1785 12188 1794
rect 13816 1785 13868 1794
rect 15496 1785 15548 1794
rect 17176 1785 17228 1794
rect 18856 1785 18908 1794
rect 20536 1785 20588 1794
rect 22216 1785 22268 1794
rect 23896 1785 23948 1794
rect 25576 1785 25628 1794
rect 27256 1785 27308 1794
rect 28936 1785 28988 1794
rect 30616 1785 30668 1794
rect 32296 1785 32348 1794
rect 33976 1785 34028 1794
rect 35656 1785 35708 1794
rect 37336 1785 37388 1794
rect 39016 1785 39068 1794
rect 40696 1785 40748 1794
rect 42376 1785 42428 1794
rect 44056 1785 44108 1794
rect 45736 1785 45788 1794
rect 47416 1785 47468 1794
rect 49096 1785 49148 1794
rect 50776 1785 50828 1794
rect 52456 1785 52508 1794
rect 54136 1785 54188 1794
rect 55816 1785 55868 1794
rect 57496 1785 57548 1794
rect 59176 1785 59228 1794
rect 60856 1785 60908 1794
rect 62536 1785 62588 1794
rect 64216 1785 64268 1794
rect 65896 1785 65948 1794
rect 67576 1785 67628 1794
rect 69256 1785 69308 1794
rect 70936 1785 70988 1794
rect 72616 1785 72668 1794
rect 74296 1785 74348 1794
rect 75976 1785 76028 1794
rect 77656 1785 77708 1794
rect 79336 1785 79388 1794
rect 81016 1785 81068 1794
rect 82696 1785 82748 1794
rect 84376 1785 84428 1794
rect 86056 1785 86108 1794
rect 87736 1785 87788 1794
rect 2056 1751 2065 1785
rect 2065 1751 2099 1785
rect 2099 1751 2108 1785
rect 3736 1751 3745 1785
rect 3745 1751 3779 1785
rect 3779 1751 3788 1785
rect 5416 1751 5425 1785
rect 5425 1751 5459 1785
rect 5459 1751 5468 1785
rect 7096 1751 7105 1785
rect 7105 1751 7139 1785
rect 7139 1751 7148 1785
rect 8776 1751 8785 1785
rect 8785 1751 8819 1785
rect 8819 1751 8828 1785
rect 10456 1751 10465 1785
rect 10465 1751 10499 1785
rect 10499 1751 10508 1785
rect 12136 1751 12145 1785
rect 12145 1751 12179 1785
rect 12179 1751 12188 1785
rect 13816 1751 13825 1785
rect 13825 1751 13859 1785
rect 13859 1751 13868 1785
rect 15496 1751 15505 1785
rect 15505 1751 15539 1785
rect 15539 1751 15548 1785
rect 17176 1751 17185 1785
rect 17185 1751 17219 1785
rect 17219 1751 17228 1785
rect 18856 1751 18865 1785
rect 18865 1751 18899 1785
rect 18899 1751 18908 1785
rect 20536 1751 20545 1785
rect 20545 1751 20579 1785
rect 20579 1751 20588 1785
rect 22216 1751 22225 1785
rect 22225 1751 22259 1785
rect 22259 1751 22268 1785
rect 23896 1751 23905 1785
rect 23905 1751 23939 1785
rect 23939 1751 23948 1785
rect 25576 1751 25585 1785
rect 25585 1751 25619 1785
rect 25619 1751 25628 1785
rect 27256 1751 27265 1785
rect 27265 1751 27299 1785
rect 27299 1751 27308 1785
rect 28936 1751 28945 1785
rect 28945 1751 28979 1785
rect 28979 1751 28988 1785
rect 30616 1751 30625 1785
rect 30625 1751 30659 1785
rect 30659 1751 30668 1785
rect 32296 1751 32305 1785
rect 32305 1751 32339 1785
rect 32339 1751 32348 1785
rect 33976 1751 33985 1785
rect 33985 1751 34019 1785
rect 34019 1751 34028 1785
rect 35656 1751 35665 1785
rect 35665 1751 35699 1785
rect 35699 1751 35708 1785
rect 37336 1751 37345 1785
rect 37345 1751 37379 1785
rect 37379 1751 37388 1785
rect 39016 1751 39025 1785
rect 39025 1751 39059 1785
rect 39059 1751 39068 1785
rect 40696 1751 40705 1785
rect 40705 1751 40739 1785
rect 40739 1751 40748 1785
rect 42376 1751 42385 1785
rect 42385 1751 42419 1785
rect 42419 1751 42428 1785
rect 44056 1751 44065 1785
rect 44065 1751 44099 1785
rect 44099 1751 44108 1785
rect 45736 1751 45745 1785
rect 45745 1751 45779 1785
rect 45779 1751 45788 1785
rect 47416 1751 47425 1785
rect 47425 1751 47459 1785
rect 47459 1751 47468 1785
rect 49096 1751 49105 1785
rect 49105 1751 49139 1785
rect 49139 1751 49148 1785
rect 50776 1751 50785 1785
rect 50785 1751 50819 1785
rect 50819 1751 50828 1785
rect 52456 1751 52465 1785
rect 52465 1751 52499 1785
rect 52499 1751 52508 1785
rect 54136 1751 54145 1785
rect 54145 1751 54179 1785
rect 54179 1751 54188 1785
rect 55816 1751 55825 1785
rect 55825 1751 55859 1785
rect 55859 1751 55868 1785
rect 57496 1751 57505 1785
rect 57505 1751 57539 1785
rect 57539 1751 57548 1785
rect 59176 1751 59185 1785
rect 59185 1751 59219 1785
rect 59219 1751 59228 1785
rect 60856 1751 60865 1785
rect 60865 1751 60899 1785
rect 60899 1751 60908 1785
rect 62536 1751 62545 1785
rect 62545 1751 62579 1785
rect 62579 1751 62588 1785
rect 64216 1751 64225 1785
rect 64225 1751 64259 1785
rect 64259 1751 64268 1785
rect 65896 1751 65905 1785
rect 65905 1751 65939 1785
rect 65939 1751 65948 1785
rect 67576 1751 67585 1785
rect 67585 1751 67619 1785
rect 67619 1751 67628 1785
rect 69256 1751 69265 1785
rect 69265 1751 69299 1785
rect 69299 1751 69308 1785
rect 70936 1751 70945 1785
rect 70945 1751 70979 1785
rect 70979 1751 70988 1785
rect 72616 1751 72625 1785
rect 72625 1751 72659 1785
rect 72659 1751 72668 1785
rect 74296 1751 74305 1785
rect 74305 1751 74339 1785
rect 74339 1751 74348 1785
rect 75976 1751 75985 1785
rect 75985 1751 76019 1785
rect 76019 1751 76028 1785
rect 77656 1751 77665 1785
rect 77665 1751 77699 1785
rect 77699 1751 77708 1785
rect 79336 1751 79345 1785
rect 79345 1751 79379 1785
rect 79379 1751 79388 1785
rect 81016 1751 81025 1785
rect 81025 1751 81059 1785
rect 81059 1751 81068 1785
rect 82696 1751 82705 1785
rect 82705 1751 82739 1785
rect 82739 1751 82748 1785
rect 84376 1751 84385 1785
rect 84385 1751 84419 1785
rect 84419 1751 84428 1785
rect 86056 1751 86065 1785
rect 86065 1751 86099 1785
rect 86099 1751 86108 1785
rect 87736 1751 87745 1785
rect 87745 1751 87779 1785
rect 87779 1751 87788 1785
rect 2056 1742 2108 1751
rect 3736 1742 3788 1751
rect 5416 1742 5468 1751
rect 7096 1742 7148 1751
rect 8776 1742 8828 1751
rect 10456 1742 10508 1751
rect 12136 1742 12188 1751
rect 13816 1742 13868 1751
rect 15496 1742 15548 1751
rect 17176 1742 17228 1751
rect 18856 1742 18908 1751
rect 20536 1742 20588 1751
rect 22216 1742 22268 1751
rect 23896 1742 23948 1751
rect 25576 1742 25628 1751
rect 27256 1742 27308 1751
rect 28936 1742 28988 1751
rect 30616 1742 30668 1751
rect 32296 1742 32348 1751
rect 33976 1742 34028 1751
rect 35656 1742 35708 1751
rect 37336 1742 37388 1751
rect 39016 1742 39068 1751
rect 40696 1742 40748 1751
rect 42376 1742 42428 1751
rect 44056 1742 44108 1751
rect 45736 1742 45788 1751
rect 47416 1742 47468 1751
rect 49096 1742 49148 1751
rect 50776 1742 50828 1751
rect 52456 1742 52508 1751
rect 54136 1742 54188 1751
rect 55816 1742 55868 1751
rect 57496 1742 57548 1751
rect 59176 1742 59228 1751
rect 60856 1742 60908 1751
rect 62536 1742 62588 1751
rect 64216 1742 64268 1751
rect 65896 1742 65948 1751
rect 67576 1742 67628 1751
rect 69256 1742 69308 1751
rect 70936 1742 70988 1751
rect 72616 1742 72668 1751
rect 74296 1742 74348 1751
rect 75976 1742 76028 1751
rect 77656 1742 77708 1751
rect 79336 1742 79388 1751
rect 81016 1742 81068 1751
rect 82696 1742 82748 1751
rect 84376 1742 84428 1751
rect 86056 1742 86108 1751
rect 87736 1742 87788 1751
<< metal2 >>
rect 1634 87138 1858 87608
rect 2054 87524 2110 87533
rect 2054 87459 2110 87468
rect 3734 87524 3790 87533
rect 3734 87459 3790 87468
rect 5414 87524 5470 87533
rect 5414 87459 5470 87468
rect 7094 87524 7150 87533
rect 7094 87459 7150 87468
rect 8774 87524 8830 87533
rect 8774 87459 8830 87468
rect 10454 87524 10510 87533
rect 10454 87459 10510 87468
rect 12134 87524 12190 87533
rect 12134 87459 12190 87468
rect 13814 87524 13870 87533
rect 13814 87459 13870 87468
rect 15494 87524 15550 87533
rect 15494 87459 15550 87468
rect 17174 87524 17230 87533
rect 17174 87459 17230 87468
rect 18854 87524 18910 87533
rect 18854 87459 18910 87468
rect 20534 87524 20590 87533
rect 20534 87459 20590 87468
rect 22214 87524 22270 87533
rect 22214 87459 22270 87468
rect 23894 87524 23950 87533
rect 23894 87459 23950 87468
rect 25574 87524 25630 87533
rect 25574 87459 25630 87468
rect 27254 87524 27310 87533
rect 27254 87459 27310 87468
rect 28934 87524 28990 87533
rect 28934 87459 28990 87468
rect 30614 87524 30670 87533
rect 30614 87459 30670 87468
rect 32294 87524 32350 87533
rect 32294 87459 32350 87468
rect 33974 87524 34030 87533
rect 33974 87459 34030 87468
rect 35654 87524 35710 87533
rect 35654 87459 35710 87468
rect 37334 87524 37390 87533
rect 37334 87459 37390 87468
rect 39014 87524 39070 87533
rect 39014 87459 39070 87468
rect 40694 87524 40750 87533
rect 40694 87459 40750 87468
rect 42374 87524 42430 87533
rect 42374 87459 42430 87468
rect 44054 87524 44110 87533
rect 44054 87459 44110 87468
rect 45734 87524 45790 87533
rect 45734 87459 45790 87468
rect 47414 87524 47470 87533
rect 47414 87459 47470 87468
rect 49094 87524 49150 87533
rect 49094 87459 49150 87468
rect 50774 87524 50830 87533
rect 50774 87459 50830 87468
rect 52454 87524 52510 87533
rect 52454 87459 52510 87468
rect 54134 87524 54190 87533
rect 54134 87459 54190 87468
rect 55814 87524 55870 87533
rect 55814 87459 55870 87468
rect 57494 87524 57550 87533
rect 57494 87459 57550 87468
rect 59174 87524 59230 87533
rect 59174 87459 59230 87468
rect 60854 87524 60910 87533
rect 60854 87459 60910 87468
rect 62534 87524 62590 87533
rect 62534 87459 62590 87468
rect 64214 87524 64270 87533
rect 64214 87459 64270 87468
rect 65894 87524 65950 87533
rect 65894 87459 65950 87468
rect 67574 87524 67630 87533
rect 67574 87459 67630 87468
rect 69254 87524 69310 87533
rect 69254 87459 69310 87468
rect 70934 87524 70990 87533
rect 70934 87459 70990 87468
rect 72614 87524 72670 87533
rect 72614 87459 72670 87468
rect 74294 87524 74350 87533
rect 74294 87459 74350 87468
rect 75974 87524 76030 87533
rect 75974 87459 76030 87468
rect 77654 87524 77710 87533
rect 77654 87459 77710 87468
rect 79334 87524 79390 87533
rect 79334 87459 79390 87468
rect 81014 87524 81070 87533
rect 81014 87459 81070 87468
rect 82694 87524 82750 87533
rect 82694 87459 82750 87468
rect 84374 87524 84430 87533
rect 84374 87459 84430 87468
rect 86054 87524 86110 87533
rect 86054 87459 86110 87468
rect 87734 87524 87790 87533
rect 87734 87459 87790 87468
rect 1634 87086 1720 87138
rect 1772 87086 1858 87138
rect 1634 86802 1858 87086
rect 1634 86750 1720 86802
rect 1772 86750 1858 86802
rect 1634 86466 1858 86750
rect 89132 87138 89356 87608
rect 89132 87086 89218 87138
rect 89270 87086 89356 87138
rect 89132 86802 89356 87086
rect 89132 86750 89218 86802
rect 89270 86750 89356 86802
rect 79260 86544 79316 86553
rect 79260 86479 79316 86488
rect 1634 86414 1720 86466
rect 1772 86414 1858 86466
rect 1634 86132 1858 86414
rect 74502 86288 74558 86297
rect 74502 86223 74558 86232
rect 75670 86288 75726 86297
rect 75670 86223 75726 86232
rect 76838 86288 76894 86297
rect 76838 86223 76894 86232
rect 1634 86076 1718 86132
rect 1774 86076 1858 86132
rect 1634 85794 1858 86076
rect 1634 85742 1720 85794
rect 1772 85742 1858 85794
rect 1634 85458 1858 85742
rect 1634 85406 1720 85458
rect 1772 85406 1858 85458
rect 1634 85122 1858 85406
rect 1634 85070 1720 85122
rect 1772 85070 1858 85122
rect 1634 84786 1858 85070
rect 1634 84734 1720 84786
rect 1772 84734 1858 84786
rect 1634 84452 1858 84734
rect 1634 84396 1718 84452
rect 1774 84396 1858 84452
rect 1634 84114 1858 84396
rect 1634 84062 1720 84114
rect 1772 84062 1858 84114
rect 1634 83778 1858 84062
rect 1634 83726 1720 83778
rect 1772 83726 1858 83778
rect 1634 83442 1858 83726
rect 1634 83390 1720 83442
rect 1772 83390 1858 83442
rect 1634 83106 1858 83390
rect 1634 83054 1720 83106
rect 1772 83054 1858 83106
rect 1634 82772 1858 83054
rect 1634 82716 1718 82772
rect 1774 82716 1858 82772
rect 1634 82434 1858 82716
rect 1634 82382 1720 82434
rect 1772 82382 1858 82434
rect 1634 82098 1858 82382
rect 1634 82046 1720 82098
rect 1772 82046 1858 82098
rect 1634 81762 1858 82046
rect 1634 81710 1720 81762
rect 1772 81710 1858 81762
rect 1634 81426 1858 81710
rect 1634 81374 1720 81426
rect 1772 81374 1858 81426
rect 1634 81092 1858 81374
rect 1634 81036 1718 81092
rect 1774 81036 1858 81092
rect 1634 80754 1858 81036
rect 1634 80702 1720 80754
rect 1772 80702 1858 80754
rect 1634 80418 1858 80702
rect 1634 80366 1720 80418
rect 1772 80366 1858 80418
rect 1634 80082 1858 80366
rect 1634 80030 1720 80082
rect 1772 80030 1858 80082
rect 1634 79746 1858 80030
rect 1634 79694 1720 79746
rect 1772 79694 1858 79746
rect 1634 79412 1858 79694
rect 1634 79356 1718 79412
rect 1774 79356 1858 79412
rect 1634 79074 1858 79356
rect 1634 79022 1720 79074
rect 1772 79022 1858 79074
rect 1634 78738 1858 79022
rect 1634 78686 1720 78738
rect 1772 78686 1858 78738
rect 1634 78402 1858 78686
rect 1634 78350 1720 78402
rect 1772 78350 1858 78402
rect 1634 78066 1858 78350
rect 1634 78014 1720 78066
rect 1772 78014 1858 78066
rect 1634 77732 1858 78014
rect 79274 79478 79302 86479
rect 89132 86466 89356 86750
rect 89132 86414 89218 86466
rect 89270 86414 89356 86466
rect 89132 86132 89356 86414
rect 89132 86076 89216 86132
rect 89272 86076 89356 86132
rect 89132 85794 89356 86076
rect 89132 85742 89218 85794
rect 89270 85742 89356 85794
rect 89132 85458 89356 85742
rect 89132 85406 89218 85458
rect 89270 85406 89356 85458
rect 89132 85122 89356 85406
rect 89132 85070 89218 85122
rect 89270 85070 89356 85122
rect 89132 84786 89356 85070
rect 89132 84734 89218 84786
rect 89270 84734 89356 84786
rect 89132 84452 89356 84734
rect 89132 84396 89216 84452
rect 89272 84396 89356 84452
rect 89132 84114 89356 84396
rect 89132 84062 89218 84114
rect 89270 84062 89356 84114
rect 89132 83778 89356 84062
rect 89132 83726 89218 83778
rect 89270 83726 89356 83778
rect 89132 83442 89356 83726
rect 89132 83390 89218 83442
rect 89270 83390 89356 83442
rect 89132 83106 89356 83390
rect 89132 83054 89218 83106
rect 89270 83054 89356 83106
rect 89132 82772 89356 83054
rect 89132 82716 89216 82772
rect 89272 82716 89356 82772
rect 89132 82434 89356 82716
rect 89132 82382 89218 82434
rect 89270 82382 89356 82434
rect 89132 82098 89356 82382
rect 89132 82046 89218 82098
rect 89270 82046 89356 82098
rect 89132 81762 89356 82046
rect 89132 81710 89218 81762
rect 89270 81710 89356 81762
rect 89132 81426 89356 81710
rect 89132 81374 89218 81426
rect 89270 81374 89356 81426
rect 89132 81092 89356 81374
rect 89132 81036 89216 81092
rect 89272 81036 89356 81092
rect 89132 80754 89356 81036
rect 89132 80702 89218 80754
rect 89270 80702 89356 80754
rect 89132 80418 89356 80702
rect 89132 80366 89218 80418
rect 89270 80366 89356 80418
rect 89132 80082 89356 80366
rect 89132 80030 89218 80082
rect 89270 80030 89356 80082
rect 89132 79746 89356 80030
rect 89132 79694 89218 79746
rect 89270 79694 89356 79746
rect 88256 79635 88312 79644
rect 88256 79570 88312 79579
rect 85119 79530 85175 79539
rect 79274 79450 79372 79478
rect 85119 79465 85175 79474
rect 25626 77910 25682 77919
rect 25626 77845 25682 77854
rect 30618 77910 30674 77919
rect 30618 77845 30674 77854
rect 35610 77910 35666 77919
rect 35610 77845 35666 77854
rect 40602 77910 40658 77919
rect 40602 77845 40658 77854
rect 45594 77910 45650 77919
rect 45594 77845 45650 77854
rect 50586 77910 50642 77919
rect 50586 77845 50642 77854
rect 55578 77910 55634 77919
rect 55578 77845 55634 77854
rect 60570 77910 60626 77919
rect 60570 77845 60626 77854
rect 1634 77676 1718 77732
rect 1774 77676 1858 77732
rect 1634 77394 1858 77676
rect 1634 77342 1720 77394
rect 1772 77342 1858 77394
rect 1634 77058 1858 77342
rect 1634 77006 1720 77058
rect 1772 77006 1858 77058
rect 1634 76722 1858 77006
rect 1634 76670 1720 76722
rect 1772 76670 1858 76722
rect 1634 76386 1858 76670
rect 1634 76334 1720 76386
rect 1772 76334 1858 76386
rect 1634 76052 1858 76334
rect 1634 75996 1718 76052
rect 1774 75996 1858 76052
rect 1634 75714 1858 75996
rect 1634 75662 1720 75714
rect 1772 75662 1858 75714
rect 1634 75378 1858 75662
rect 1634 75326 1720 75378
rect 1772 75326 1858 75378
rect 1634 75042 1858 75326
rect 67133 75254 67189 75263
rect 67133 75189 67189 75198
rect 1634 74990 1720 75042
rect 1772 74990 1858 75042
rect 1634 74706 1858 74990
rect 1634 74654 1720 74706
rect 1772 74654 1858 74706
rect 1634 74372 1858 74654
rect 1634 74316 1718 74372
rect 1774 74316 1858 74372
rect 1634 74034 1858 74316
rect 1634 73982 1720 74034
rect 1772 73982 1858 74034
rect 1634 73698 1858 73982
rect 1634 73646 1720 73698
rect 1772 73646 1858 73698
rect 1634 73362 1858 73646
rect 1634 73310 1720 73362
rect 1772 73310 1858 73362
rect 1634 73026 1858 73310
rect 1634 72974 1720 73026
rect 1772 72974 1858 73026
rect 1634 72692 1858 72974
rect 1634 72636 1718 72692
rect 1774 72636 1858 72692
rect 1634 72354 1858 72636
rect 1634 72302 1720 72354
rect 1772 72302 1858 72354
rect 1634 72018 1858 72302
rect 1634 71966 1720 72018
rect 1772 71966 1858 72018
rect 1634 71682 1858 71966
rect 1634 71630 1720 71682
rect 1772 71630 1858 71682
rect 1634 71346 1858 71630
rect 67147 71549 67175 75189
rect 67257 73836 67313 73845
rect 67257 73771 67313 73780
rect 67271 71549 67299 73771
rect 71118 72422 71174 72431
rect 71118 72357 71174 72366
rect 1634 71294 1720 71346
rect 1772 71294 1858 71346
rect 1634 71012 1858 71294
rect 71132 71072 71160 72357
rect 1634 70956 1718 71012
rect 1774 70956 1858 71012
rect 1634 70674 1858 70956
rect 1634 70622 1720 70674
rect 1772 70622 1858 70674
rect 1634 70338 1858 70622
rect 1634 70286 1720 70338
rect 1772 70286 1858 70338
rect 1634 70002 1858 70286
rect 1634 69950 1720 70002
rect 1772 69950 1858 70002
rect 1634 69666 1858 69950
rect 1634 69614 1720 69666
rect 1772 69614 1858 69666
rect 1634 69332 1858 69614
rect 1634 69276 1718 69332
rect 1774 69276 1858 69332
rect 1634 68994 1858 69276
rect 1634 68942 1720 68994
rect 1772 68942 1858 68994
rect 1634 68658 1858 68942
rect 1634 68606 1720 68658
rect 1772 68606 1858 68658
rect 1634 68322 1858 68606
rect 1634 68270 1720 68322
rect 1772 68270 1858 68322
rect 1634 67986 1858 68270
rect 1634 67934 1720 67986
rect 1772 67934 1858 67986
rect 1634 67652 1858 67934
rect 1634 67596 1718 67652
rect 1774 67596 1858 67652
rect 1634 67314 1858 67596
rect 1634 67262 1720 67314
rect 1772 67262 1858 67314
rect 1634 66978 1858 67262
rect 1634 66926 1720 66978
rect 1772 66926 1858 66978
rect 1634 66642 1858 66926
rect 1634 66590 1720 66642
rect 1772 66590 1858 66642
rect 1634 66306 1858 66590
rect 1634 66254 1720 66306
rect 1772 66254 1858 66306
rect 1634 65972 1858 66254
rect 1634 65916 1718 65972
rect 1774 65916 1858 65972
rect 1634 65634 1858 65916
rect 1634 65582 1720 65634
rect 1772 65582 1858 65634
rect 1634 65298 1858 65582
rect 1634 65246 1720 65298
rect 1772 65246 1858 65298
rect 1634 64962 1858 65246
rect 1634 64910 1720 64962
rect 1772 64910 1858 64962
rect 1634 64626 1858 64910
rect 1634 64574 1720 64626
rect 1772 64574 1858 64626
rect 1634 64292 1858 64574
rect 1634 64236 1718 64292
rect 1774 64236 1858 64292
rect 1634 63954 1858 64236
rect 1634 63902 1720 63954
rect 1772 63902 1858 63954
rect 1634 63618 1858 63902
rect 1634 63566 1720 63618
rect 1772 63566 1858 63618
rect 1634 63282 1858 63566
rect 1634 63230 1720 63282
rect 1772 63230 1858 63282
rect 1634 62946 1858 63230
rect 1634 62894 1720 62946
rect 1772 62894 1858 62946
rect 1634 62612 1858 62894
rect 1634 62556 1718 62612
rect 1774 62556 1858 62612
rect 1634 62274 1858 62556
rect 1634 62222 1720 62274
rect 1772 62222 1858 62274
rect 1634 61938 1858 62222
rect 1634 61886 1720 61938
rect 1772 61886 1858 61938
rect 1634 61602 1858 61886
rect 1634 61550 1720 61602
rect 1772 61550 1858 61602
rect 1634 61266 1858 61550
rect 1634 61214 1720 61266
rect 1772 61214 1858 61266
rect 1634 60932 1858 61214
rect 1634 60876 1718 60932
rect 1774 60876 1858 60932
rect 1634 60594 1858 60876
rect 1634 60542 1720 60594
rect 1772 60542 1858 60594
rect 1634 60258 1858 60542
rect 1634 60206 1720 60258
rect 1772 60206 1858 60258
rect 1634 59922 1858 60206
rect 1634 59870 1720 59922
rect 1772 59870 1858 59922
rect 1634 59586 1858 59870
rect 1634 59534 1720 59586
rect 1772 59534 1858 59586
rect 1634 59252 1858 59534
rect 1634 59196 1718 59252
rect 1774 59196 1858 59252
rect 1634 58914 1858 59196
rect 1634 58862 1720 58914
rect 1772 58862 1858 58914
rect 1634 58578 1858 58862
rect 1634 58526 1720 58578
rect 1772 58526 1858 58578
rect 1634 58242 1858 58526
rect 1634 58190 1720 58242
rect 1772 58190 1858 58242
rect 1634 57906 1858 58190
rect 1634 57854 1720 57906
rect 1772 57854 1858 57906
rect 1634 57572 1858 57854
rect 1634 57516 1718 57572
rect 1774 57516 1858 57572
rect 1634 57234 1858 57516
rect 1634 57182 1720 57234
rect 1772 57182 1858 57234
rect 1634 56898 1858 57182
rect 1634 56846 1720 56898
rect 1772 56846 1858 56898
rect 1634 56562 1858 56846
rect 1634 56510 1720 56562
rect 1772 56510 1858 56562
rect 1634 56226 1858 56510
rect 1634 56174 1720 56226
rect 1772 56174 1858 56226
rect 1634 55892 1858 56174
rect 1634 55836 1718 55892
rect 1774 55836 1858 55892
rect 1634 55554 1858 55836
rect 1634 55502 1720 55554
rect 1772 55502 1858 55554
rect 1634 55218 1858 55502
rect 1634 55166 1720 55218
rect 1772 55166 1858 55218
rect 1634 54882 1858 55166
rect 1634 54830 1720 54882
rect 1772 54830 1858 54882
rect 1634 54546 1858 54830
rect 1634 54494 1720 54546
rect 1772 54494 1858 54546
rect 1634 54212 1858 54494
rect 1634 54156 1718 54212
rect 1774 54156 1858 54212
rect 1634 53874 1858 54156
rect 1634 53822 1720 53874
rect 1772 53822 1858 53874
rect 1634 53538 1858 53822
rect 1634 53486 1720 53538
rect 1772 53486 1858 53538
rect 1634 53202 1858 53486
rect 1634 53150 1720 53202
rect 1772 53150 1858 53202
rect 1634 52866 1858 53150
rect 1634 52814 1720 52866
rect 1772 52814 1858 52866
rect 1634 52532 1858 52814
rect 1634 52476 1718 52532
rect 1774 52476 1858 52532
rect 1634 52194 1858 52476
rect 1634 52142 1720 52194
rect 1772 52142 1858 52194
rect 1634 51858 1858 52142
rect 1634 51806 1720 51858
rect 1772 51806 1858 51858
rect 1634 51522 1858 51806
rect 1634 51470 1720 51522
rect 1772 51470 1858 51522
rect 1634 51186 1858 51470
rect 1634 51134 1720 51186
rect 1772 51134 1858 51186
rect 1634 50852 1858 51134
rect 1634 50796 1718 50852
rect 1774 50796 1858 50852
rect 1634 50514 1858 50796
rect 1634 50462 1720 50514
rect 1772 50462 1858 50514
rect 1634 50178 1858 50462
rect 1634 50126 1720 50178
rect 1772 50126 1858 50178
rect 1634 49842 1858 50126
rect 1634 49790 1720 49842
rect 1772 49790 1858 49842
rect 1634 49506 1858 49790
rect 1634 49454 1720 49506
rect 1772 49454 1858 49506
rect 1634 49172 1858 49454
rect 1634 49116 1718 49172
rect 1774 49116 1858 49172
rect 1634 48834 1858 49116
rect 1634 48782 1720 48834
rect 1772 48782 1858 48834
rect 1634 48498 1858 48782
rect 1634 48446 1720 48498
rect 1772 48446 1858 48498
rect 1634 48162 1858 48446
rect 1634 48110 1720 48162
rect 1772 48110 1858 48162
rect 1634 47826 1858 48110
rect 1634 47774 1720 47826
rect 1772 47774 1858 47826
rect 1634 47492 1858 47774
rect 1634 47436 1718 47492
rect 1774 47436 1858 47492
rect 1634 47154 1858 47436
rect 1634 47102 1720 47154
rect 1772 47102 1858 47154
rect 1634 46818 1858 47102
rect 1634 46766 1720 46818
rect 1772 46766 1858 46818
rect 1634 46482 1858 46766
rect 1634 46430 1720 46482
rect 1772 46430 1858 46482
rect 1634 46146 1858 46430
rect 1634 46094 1720 46146
rect 1772 46094 1858 46146
rect 1634 45812 1858 46094
rect 1634 45756 1718 45812
rect 1774 45756 1858 45812
rect 1634 45474 1858 45756
rect 1634 45422 1720 45474
rect 1772 45422 1858 45474
rect 1634 45138 1858 45422
rect 1634 45086 1720 45138
rect 1772 45086 1858 45138
rect 1634 44802 1858 45086
rect 1634 44750 1720 44802
rect 1772 44750 1858 44802
rect 1634 44466 1858 44750
rect 1634 44414 1720 44466
rect 1772 44414 1858 44466
rect 1634 44132 1858 44414
rect 1634 44076 1718 44132
rect 1774 44076 1858 44132
rect 1634 43794 1858 44076
rect 1634 43742 1720 43794
rect 1772 43742 1858 43794
rect 1634 43458 1858 43742
rect 1634 43406 1720 43458
rect 1772 43406 1858 43458
rect 1634 43122 1858 43406
rect 1634 43070 1720 43122
rect 1772 43070 1858 43122
rect 1634 42786 1858 43070
rect 1634 42734 1720 42786
rect 1772 42734 1858 42786
rect 1634 42452 1858 42734
rect 1634 42396 1718 42452
rect 1774 42396 1858 42452
rect 1634 42114 1858 42396
rect 1634 42062 1720 42114
rect 1772 42062 1858 42114
rect 1634 41778 1858 42062
rect 1634 41726 1720 41778
rect 1772 41726 1858 41778
rect 1634 41442 1858 41726
rect 1634 41390 1720 41442
rect 1772 41390 1858 41442
rect 1634 41106 1858 41390
rect 1634 41054 1720 41106
rect 1772 41054 1858 41106
rect 1634 40772 1858 41054
rect 1634 40716 1718 40772
rect 1774 40716 1858 40772
rect 1634 40434 1858 40716
rect 1634 40382 1720 40434
rect 1772 40382 1858 40434
rect 1634 40098 1858 40382
rect 1634 40046 1720 40098
rect 1772 40046 1858 40098
rect 1634 39762 1858 40046
rect 1634 39710 1720 39762
rect 1772 39710 1858 39762
rect 1634 39426 1858 39710
rect 1634 39374 1720 39426
rect 1772 39374 1858 39426
rect 1634 39092 1858 39374
rect 1634 39036 1718 39092
rect 1774 39036 1858 39092
rect 1634 38754 1858 39036
rect 1634 38702 1720 38754
rect 1772 38702 1858 38754
rect 1634 38418 1858 38702
rect 1634 38366 1720 38418
rect 1772 38366 1858 38418
rect 1634 38082 1858 38366
rect 1634 38030 1720 38082
rect 1772 38030 1858 38082
rect 1634 37746 1858 38030
rect 1634 37694 1720 37746
rect 1772 37694 1858 37746
rect 1634 37412 1858 37694
rect 1634 37356 1718 37412
rect 1774 37356 1858 37412
rect 1634 37074 1858 37356
rect 11621 37260 11677 37269
rect 10676 37189 10732 37198
rect 11621 37195 11677 37204
rect 12355 37260 12411 37269
rect 12355 37195 12411 37204
rect 10676 37124 10732 37133
rect 1634 37022 1720 37074
rect 1772 37022 1858 37074
rect 1634 36738 1858 37022
rect 1634 36686 1720 36738
rect 1772 36686 1858 36738
rect 1634 36402 1858 36686
rect 1634 36350 1720 36402
rect 1772 36350 1858 36402
rect 1634 36066 1858 36350
rect 1634 36014 1720 36066
rect 1772 36014 1858 36066
rect 1634 35732 1858 36014
rect 10676 36061 10732 36070
rect 10676 35996 10732 36005
rect 11621 35990 11677 35999
rect 11621 35925 11677 35934
rect 12275 35990 12331 35999
rect 12275 35925 12331 35934
rect 1634 35676 1718 35732
rect 1774 35676 1858 35732
rect 1634 35394 1858 35676
rect 1634 35342 1720 35394
rect 1772 35342 1858 35394
rect 1634 35058 1858 35342
rect 1634 35006 1720 35058
rect 1772 35006 1858 35058
rect 1634 34722 1858 35006
rect 1634 34670 1720 34722
rect 1772 34670 1858 34722
rect 1634 34386 1858 34670
rect 1634 34334 1720 34386
rect 1772 34334 1858 34386
rect 11621 34432 11677 34441
rect 1634 34052 1858 34334
rect 10676 34361 10732 34370
rect 11621 34367 11677 34376
rect 12195 34432 12251 34441
rect 12195 34367 12251 34376
rect 10676 34296 10732 34305
rect 1634 33996 1718 34052
rect 1774 33996 1858 34052
rect 1634 33714 1858 33996
rect 1634 33662 1720 33714
rect 1772 33662 1858 33714
rect 1634 33378 1858 33662
rect 1634 33326 1720 33378
rect 1772 33326 1858 33378
rect 1634 33042 1858 33326
rect 10676 33233 10732 33242
rect 10676 33168 10732 33177
rect 11621 33162 11677 33171
rect 11621 33097 11677 33106
rect 12115 33162 12171 33171
rect 12115 33097 12171 33106
rect 1634 32990 1720 33042
rect 1772 32990 1858 33042
rect 1634 32706 1858 32990
rect 1634 32654 1720 32706
rect 1772 32654 1858 32706
rect 1634 32372 1858 32654
rect 1634 32316 1718 32372
rect 1774 32316 1858 32372
rect 1634 32034 1858 32316
rect 1634 31982 1720 32034
rect 1772 31982 1858 32034
rect 1634 31698 1858 31982
rect 1634 31646 1720 31698
rect 1772 31646 1858 31698
rect 1634 31362 1858 31646
rect 11621 31604 11677 31613
rect 10676 31533 10732 31542
rect 11621 31539 11677 31548
rect 12035 31604 12091 31613
rect 12035 31539 12091 31548
rect 10676 31468 10732 31477
rect 1634 31310 1720 31362
rect 1772 31310 1858 31362
rect 1634 31026 1858 31310
rect 1634 30974 1720 31026
rect 1772 30974 1858 31026
rect 1634 30692 1858 30974
rect 1634 30636 1718 30692
rect 1774 30636 1858 30692
rect 1634 30354 1858 30636
rect 1634 30302 1720 30354
rect 1772 30302 1858 30354
rect 10676 30405 10732 30414
rect 10676 30340 10732 30349
rect 1634 30018 1858 30302
rect 11621 30334 11677 30343
rect 11621 30269 11677 30278
rect 11955 30334 12011 30343
rect 11955 30269 12011 30278
rect 1634 29966 1720 30018
rect 1772 29966 1858 30018
rect 1634 29682 1858 29966
rect 1634 29630 1720 29682
rect 1772 29630 1858 29682
rect 1634 29346 1858 29630
rect 1634 29294 1720 29346
rect 1772 29294 1858 29346
rect 1634 29012 1858 29294
rect 1634 28956 1718 29012
rect 1774 28956 1858 29012
rect 1634 28674 1858 28956
rect 11621 28776 11677 28785
rect 1634 28622 1720 28674
rect 1772 28622 1858 28674
rect 10676 28705 10732 28714
rect 11621 28711 11677 28720
rect 11875 28776 11931 28785
rect 11875 28711 11931 28720
rect 10676 28640 10732 28649
rect 1634 28338 1858 28622
rect 11758 28449 11814 28458
rect 11758 28384 11814 28393
rect 1634 28286 1720 28338
rect 1772 28286 1858 28338
rect 1634 28002 1858 28286
rect 1634 27950 1720 28002
rect 1772 27950 1858 28002
rect 1634 27666 1858 27950
rect 1634 27614 1720 27666
rect 1772 27614 1858 27666
rect 1634 27332 1858 27614
rect 1634 27276 1718 27332
rect 1774 27276 1858 27332
rect 1634 26994 1858 27276
rect 1634 26942 1720 26994
rect 1772 26942 1858 26994
rect 1634 26658 1858 26942
rect 1634 26606 1720 26658
rect 1772 26606 1858 26658
rect 1634 26322 1858 26606
rect 1634 26270 1720 26322
rect 1772 26270 1858 26322
rect 1634 25986 1858 26270
rect 1634 25934 1720 25986
rect 1772 25934 1858 25986
rect 1634 25652 1858 25934
rect 2465 25728 2521 25737
rect 2465 25663 2521 25672
rect 1634 25596 1718 25652
rect 1774 25596 1858 25652
rect 1634 25314 1858 25596
rect 1634 25262 1720 25314
rect 1772 25262 1858 25314
rect 1634 24978 1858 25262
rect 1634 24926 1720 24978
rect 1772 24926 1858 24978
rect 1634 24642 1858 24926
rect 1634 24590 1720 24642
rect 1772 24590 1858 24642
rect 1634 24306 1858 24590
rect 1634 24254 1720 24306
rect 1772 24254 1858 24306
rect 1634 23972 1858 24254
rect 1634 23916 1718 23972
rect 1774 23916 1858 23972
rect 1634 23634 1858 23916
rect 1634 23582 1720 23634
rect 1772 23582 1858 23634
rect 1634 23298 1858 23582
rect 1634 23246 1720 23298
rect 1772 23246 1858 23298
rect 1634 22962 1858 23246
rect 1634 22910 1720 22962
rect 1772 22910 1858 22962
rect 1634 22626 1858 22910
rect 1634 22574 1720 22626
rect 1772 22574 1858 22626
rect 1634 22292 1858 22574
rect 1634 22236 1718 22292
rect 1774 22236 1858 22292
rect 1634 21954 1858 22236
rect 1634 21902 1720 21954
rect 1772 21902 1858 21954
rect 1634 21618 1858 21902
rect 1634 21566 1720 21618
rect 1772 21566 1858 21618
rect 1634 21282 1858 21566
rect 1634 21230 1720 21282
rect 1772 21230 1858 21282
rect 1634 20946 1858 21230
rect 1634 20894 1720 20946
rect 1772 20894 1858 20946
rect 1634 20612 1858 20894
rect 1634 20556 1718 20612
rect 1774 20556 1858 20612
rect 1634 20274 1858 20556
rect 1634 20222 1720 20274
rect 1772 20222 1858 20274
rect 1634 19938 1858 20222
rect 1634 19886 1720 19938
rect 1772 19886 1858 19938
rect 1634 19602 1858 19886
rect 1634 19550 1720 19602
rect 1772 19550 1858 19602
rect 1634 19266 1858 19550
rect 1634 19214 1720 19266
rect 1772 19214 1858 19266
rect 1634 18932 1858 19214
rect 1634 18876 1718 18932
rect 1774 18876 1858 18932
rect 1634 18594 1858 18876
rect 1634 18542 1720 18594
rect 1772 18542 1858 18594
rect 11674 18620 11730 18629
rect 11674 18555 11730 18564
rect 1634 18258 1858 18542
rect 1634 18206 1720 18258
rect 1772 18206 1858 18258
rect 1634 17922 1858 18206
rect 1634 17870 1720 17922
rect 1772 17870 1858 17922
rect 1634 17586 1858 17870
rect 1634 17534 1720 17586
rect 1772 17534 1858 17586
rect 1634 17252 1858 17534
rect 1634 17196 1718 17252
rect 1774 17196 1858 17252
rect 1634 16914 1858 17196
rect 1634 16862 1720 16914
rect 1772 16862 1858 16914
rect 1634 16578 1858 16862
rect 1634 16526 1720 16578
rect 1772 16526 1858 16578
rect 1634 16242 1858 16526
rect 1634 16190 1720 16242
rect 1772 16190 1858 16242
rect 1634 15906 1858 16190
rect 1634 15854 1720 15906
rect 1772 15854 1858 15906
rect 1634 15572 1858 15854
rect 11674 15792 11730 15801
rect 11674 15727 11730 15736
rect 1634 15516 1718 15572
rect 1774 15516 1858 15572
rect 1634 15234 1858 15516
rect 1634 15182 1720 15234
rect 1772 15182 1858 15234
rect 1634 14898 1858 15182
rect 1634 14846 1720 14898
rect 1772 14846 1858 14898
rect 1634 14562 1858 14846
rect 1634 14510 1720 14562
rect 1772 14510 1858 14562
rect 1634 14226 1858 14510
rect 11674 14378 11730 14387
rect 11674 14313 11730 14322
rect 1634 14174 1720 14226
rect 1772 14174 1858 14226
rect 1634 13892 1858 14174
rect 1634 13836 1718 13892
rect 1774 13836 1858 13892
rect 1634 13554 1858 13836
rect 1634 13502 1720 13554
rect 1772 13502 1858 13554
rect 1634 13218 1858 13502
rect 1634 13166 1720 13218
rect 1772 13166 1858 13218
rect 1634 12882 1858 13166
rect 11674 12980 11730 12989
rect 11674 12915 11730 12924
rect 1634 12830 1720 12882
rect 1772 12830 1858 12882
rect 1634 12546 1858 12830
rect 1634 12494 1720 12546
rect 1772 12494 1858 12546
rect 1634 12212 1858 12494
rect 1634 12156 1718 12212
rect 1774 12156 1858 12212
rect 1634 11874 1858 12156
rect 1634 11822 1720 11874
rect 1772 11822 1858 11874
rect 1634 11538 1858 11822
rect 1634 11486 1720 11538
rect 1772 11486 1858 11538
rect 1634 11202 1858 11486
rect 1634 11150 1720 11202
rect 1772 11150 1858 11202
rect 1634 10866 1858 11150
rect 1634 10814 1720 10866
rect 1772 10814 1858 10866
rect 1634 10532 1858 10814
rect 1634 10476 1718 10532
rect 1774 10476 1858 10532
rect 1634 10194 1858 10476
rect 2678 10279 2734 10288
rect 2678 10214 2734 10223
rect 1634 10142 1720 10194
rect 1772 10142 1858 10194
rect 1634 9858 1858 10142
rect 1634 9806 1720 9858
rect 1772 9806 1858 9858
rect 1634 9522 1858 9806
rect 1634 9470 1720 9522
rect 1772 9470 1858 9522
rect 1634 9186 1858 9470
rect 1634 9134 1720 9186
rect 1772 9134 1858 9186
rect 1634 8852 1858 9134
rect 1634 8796 1718 8852
rect 1774 8796 1858 8852
rect 1634 8514 1858 8796
rect 11772 8708 11800 28384
rect 79274 19942 79302 79450
rect 89132 79412 89356 79694
rect 89132 79356 89216 79412
rect 89272 79356 89356 79412
rect 89132 79074 89356 79356
rect 89132 79022 89218 79074
rect 89270 79022 89356 79074
rect 89132 78738 89356 79022
rect 89132 78686 89218 78738
rect 89270 78686 89356 78738
rect 89132 78402 89356 78686
rect 89132 78350 89218 78402
rect 89270 78350 89356 78402
rect 89132 78066 89356 78350
rect 89132 78014 89218 78066
rect 89270 78014 89356 78066
rect 89132 77732 89356 78014
rect 89132 77676 89216 77732
rect 89272 77676 89356 77732
rect 89132 77394 89356 77676
rect 89132 77342 89218 77394
rect 89270 77342 89356 77394
rect 89132 77058 89356 77342
rect 89132 77006 89218 77058
rect 89270 77006 89356 77058
rect 89132 76722 89356 77006
rect 89132 76670 89218 76722
rect 89270 76670 89356 76722
rect 89132 76386 89356 76670
rect 89132 76334 89218 76386
rect 89270 76334 89356 76386
rect 89132 76052 89356 76334
rect 89132 75996 89216 76052
rect 89272 75996 89356 76052
rect 89132 75714 89356 75996
rect 89132 75662 89218 75714
rect 89270 75662 89356 75714
rect 89132 75378 89356 75662
rect 89132 75326 89218 75378
rect 89270 75326 89356 75378
rect 79344 75234 79400 75243
rect 79344 75169 79400 75178
rect 89132 75042 89356 75326
rect 89132 74990 89218 75042
rect 89270 74990 89356 75042
rect 89132 74706 89356 74990
rect 89132 74654 89218 74706
rect 89270 74654 89356 74706
rect 89132 74372 89356 74654
rect 89132 74316 89216 74372
rect 89272 74316 89356 74372
rect 89132 74034 89356 74316
rect 89132 73982 89218 74034
rect 89270 73982 89356 74034
rect 79344 73836 79400 73845
rect 79344 73771 79400 73780
rect 89132 73698 89356 73982
rect 89132 73646 89218 73698
rect 89270 73646 89356 73698
rect 89132 73362 89356 73646
rect 89132 73310 89218 73362
rect 89270 73310 89356 73362
rect 89132 73026 89356 73310
rect 89132 72974 89218 73026
rect 89270 72974 89356 73026
rect 89132 72692 89356 72974
rect 89132 72636 89216 72692
rect 89272 72636 89356 72692
rect 79344 72422 79400 72431
rect 79344 72357 79400 72366
rect 89132 72354 89356 72636
rect 89132 72302 89218 72354
rect 89270 72302 89356 72354
rect 89132 72018 89356 72302
rect 89132 71966 89218 72018
rect 89270 71966 89356 72018
rect 89132 71682 89356 71966
rect 89132 71630 89218 71682
rect 89270 71630 89356 71682
rect 89132 71346 89356 71630
rect 89132 71294 89218 71346
rect 89270 71294 89356 71346
rect 89132 71012 89356 71294
rect 89132 70956 89216 71012
rect 89272 70956 89356 71012
rect 89132 70674 89356 70956
rect 89132 70622 89218 70674
rect 89270 70622 89356 70674
rect 89132 70338 89356 70622
rect 89132 70286 89218 70338
rect 89270 70286 89356 70338
rect 89132 70002 89356 70286
rect 89132 69950 89218 70002
rect 89270 69950 89356 70002
rect 89132 69666 89356 69950
rect 89132 69614 89218 69666
rect 89270 69614 89356 69666
rect 89132 69332 89356 69614
rect 89132 69276 89216 69332
rect 89272 69276 89356 69332
rect 89132 68994 89356 69276
rect 89132 68942 89218 68994
rect 89270 68942 89356 68994
rect 89132 68658 89356 68942
rect 89132 68606 89218 68658
rect 89270 68606 89356 68658
rect 89132 68322 89356 68606
rect 89132 68270 89218 68322
rect 89270 68270 89356 68322
rect 89132 67986 89356 68270
rect 89132 67934 89218 67986
rect 89270 67934 89356 67986
rect 89132 67652 89356 67934
rect 89132 67596 89216 67652
rect 89272 67596 89356 67652
rect 89132 67314 89356 67596
rect 89132 67262 89218 67314
rect 89270 67262 89356 67314
rect 89132 66978 89356 67262
rect 89132 66926 89218 66978
rect 89270 66926 89356 66978
rect 89132 66642 89356 66926
rect 89132 66590 89218 66642
rect 89270 66590 89356 66642
rect 89132 66306 89356 66590
rect 89132 66254 89218 66306
rect 89270 66254 89356 66306
rect 89132 65972 89356 66254
rect 89132 65916 89216 65972
rect 89272 65916 89356 65972
rect 89132 65634 89356 65916
rect 89132 65582 89218 65634
rect 89270 65582 89356 65634
rect 89132 65298 89356 65582
rect 89132 65246 89218 65298
rect 89270 65246 89356 65298
rect 89132 64962 89356 65246
rect 89132 64910 89218 64962
rect 89270 64910 89356 64962
rect 89132 64626 89356 64910
rect 89132 64574 89218 64626
rect 89270 64574 89356 64626
rect 89132 64292 89356 64574
rect 89132 64236 89216 64292
rect 89272 64236 89356 64292
rect 89132 63954 89356 64236
rect 89132 63902 89218 63954
rect 89270 63902 89356 63954
rect 89132 63618 89356 63902
rect 89132 63566 89218 63618
rect 89270 63566 89356 63618
rect 89132 63282 89356 63566
rect 89132 63230 89218 63282
rect 89270 63230 89356 63282
rect 89132 62946 89356 63230
rect 89132 62894 89218 62946
rect 89270 62894 89356 62946
rect 89132 62612 89356 62894
rect 89132 62556 89216 62612
rect 89272 62556 89356 62612
rect 88469 62486 88525 62495
rect 88469 62421 88525 62430
rect 89132 62274 89356 62556
rect 89132 62222 89218 62274
rect 89270 62222 89356 62274
rect 89132 61938 89356 62222
rect 89132 61886 89218 61938
rect 89270 61886 89356 61938
rect 89132 61602 89356 61886
rect 89132 61550 89218 61602
rect 89270 61550 89356 61602
rect 89132 61266 89356 61550
rect 89132 61214 89218 61266
rect 89270 61214 89356 61266
rect 89132 60932 89356 61214
rect 89132 60876 89216 60932
rect 89272 60876 89356 60932
rect 89132 60594 89356 60876
rect 89132 60542 89218 60594
rect 89270 60542 89356 60594
rect 89132 60258 89356 60542
rect 89132 60206 89218 60258
rect 89270 60206 89356 60258
rect 89132 59922 89356 60206
rect 89132 59870 89218 59922
rect 89270 59870 89356 59922
rect 89132 59586 89356 59870
rect 89132 59534 89218 59586
rect 89270 59534 89356 59586
rect 89132 59252 89356 59534
rect 89132 59196 89216 59252
rect 89272 59196 89356 59252
rect 89132 58914 89356 59196
rect 89132 58862 89218 58914
rect 89270 58862 89356 58914
rect 89132 58578 89356 58862
rect 89132 58526 89218 58578
rect 89270 58526 89356 58578
rect 89132 58242 89356 58526
rect 89132 58190 89218 58242
rect 89270 58190 89356 58242
rect 89132 57906 89356 58190
rect 89132 57854 89218 57906
rect 89270 57854 89356 57906
rect 89132 57572 89356 57854
rect 89132 57516 89216 57572
rect 89272 57516 89356 57572
rect 89132 57234 89356 57516
rect 89132 57182 89218 57234
rect 89270 57182 89356 57234
rect 89132 56898 89356 57182
rect 89132 56846 89218 56898
rect 89270 56846 89356 56898
rect 89132 56562 89356 56846
rect 89132 56510 89218 56562
rect 89270 56510 89356 56562
rect 89132 56226 89356 56510
rect 89132 56174 89218 56226
rect 89270 56174 89356 56226
rect 89132 55892 89356 56174
rect 89132 55836 89216 55892
rect 89272 55836 89356 55892
rect 89132 55554 89356 55836
rect 89132 55502 89218 55554
rect 89270 55502 89356 55554
rect 89132 55218 89356 55502
rect 89132 55166 89218 55218
rect 89270 55166 89356 55218
rect 89132 54882 89356 55166
rect 89132 54830 89218 54882
rect 89270 54830 89356 54882
rect 89132 54546 89356 54830
rect 89132 54494 89218 54546
rect 89270 54494 89356 54546
rect 89132 54212 89356 54494
rect 89132 54156 89216 54212
rect 89272 54156 89356 54212
rect 89132 53874 89356 54156
rect 89132 53822 89218 53874
rect 89270 53822 89356 53874
rect 89132 53538 89356 53822
rect 89132 53486 89218 53538
rect 89270 53486 89356 53538
rect 89132 53202 89356 53486
rect 89132 53150 89218 53202
rect 89270 53150 89356 53202
rect 89132 52866 89356 53150
rect 89132 52814 89218 52866
rect 89270 52814 89356 52866
rect 89132 52532 89356 52814
rect 89132 52476 89216 52532
rect 89272 52476 89356 52532
rect 89132 52194 89356 52476
rect 89132 52142 89218 52194
rect 89270 52142 89356 52194
rect 89132 51858 89356 52142
rect 89132 51806 89218 51858
rect 89270 51806 89356 51858
rect 89132 51522 89356 51806
rect 89132 51470 89218 51522
rect 89270 51470 89356 51522
rect 89132 51186 89356 51470
rect 89132 51134 89218 51186
rect 89270 51134 89356 51186
rect 89132 50852 89356 51134
rect 89132 50796 89216 50852
rect 89272 50796 89356 50852
rect 89132 50514 89356 50796
rect 89132 50462 89218 50514
rect 89270 50462 89356 50514
rect 89132 50178 89356 50462
rect 89132 50126 89218 50178
rect 89270 50126 89356 50178
rect 89132 49842 89356 50126
rect 89132 49790 89218 49842
rect 89270 49790 89356 49842
rect 89132 49506 89356 49790
rect 89132 49454 89218 49506
rect 89270 49454 89356 49506
rect 89132 49172 89356 49454
rect 89132 49116 89216 49172
rect 89272 49116 89356 49172
rect 89132 48834 89356 49116
rect 89132 48782 89218 48834
rect 89270 48782 89356 48834
rect 89132 48498 89356 48782
rect 89132 48446 89218 48498
rect 89270 48446 89356 48498
rect 89132 48162 89356 48446
rect 89132 48110 89218 48162
rect 89270 48110 89356 48162
rect 89132 47826 89356 48110
rect 89132 47774 89218 47826
rect 89270 47774 89356 47826
rect 89132 47492 89356 47774
rect 89132 47436 89216 47492
rect 89272 47436 89356 47492
rect 89132 47154 89356 47436
rect 89132 47102 89218 47154
rect 89270 47102 89356 47154
rect 89132 46818 89356 47102
rect 89132 46766 89218 46818
rect 89270 46766 89356 46818
rect 89132 46482 89356 46766
rect 89132 46430 89218 46482
rect 89270 46430 89356 46482
rect 89132 46146 89356 46430
rect 89132 46094 89218 46146
rect 89270 46094 89356 46146
rect 89132 45812 89356 46094
rect 89132 45756 89216 45812
rect 89272 45756 89356 45812
rect 89132 45474 89356 45756
rect 89132 45422 89218 45474
rect 89270 45422 89356 45474
rect 89132 45138 89356 45422
rect 89132 45086 89218 45138
rect 89270 45086 89356 45138
rect 89132 44802 89356 45086
rect 89132 44750 89218 44802
rect 89270 44750 89356 44802
rect 89132 44466 89356 44750
rect 89132 44414 89218 44466
rect 89270 44414 89356 44466
rect 89132 44132 89356 44414
rect 89132 44076 89216 44132
rect 89272 44076 89356 44132
rect 89132 43794 89356 44076
rect 89132 43742 89218 43794
rect 89270 43742 89356 43794
rect 89132 43458 89356 43742
rect 89132 43406 89218 43458
rect 89270 43406 89356 43458
rect 89132 43122 89356 43406
rect 89132 43070 89218 43122
rect 89270 43070 89356 43122
rect 89132 42786 89356 43070
rect 89132 42734 89218 42786
rect 89270 42734 89356 42786
rect 89132 42452 89356 42734
rect 89132 42396 89216 42452
rect 89272 42396 89356 42452
rect 89132 42114 89356 42396
rect 89132 42062 89218 42114
rect 89270 42062 89356 42114
rect 89132 41778 89356 42062
rect 89132 41726 89218 41778
rect 89270 41726 89356 41778
rect 89132 41442 89356 41726
rect 89132 41390 89218 41442
rect 89270 41390 89356 41442
rect 89132 41106 89356 41390
rect 89132 41054 89218 41106
rect 89270 41054 89356 41106
rect 89132 40772 89356 41054
rect 89132 40716 89216 40772
rect 89272 40716 89356 40772
rect 89132 40434 89356 40716
rect 89132 40382 89218 40434
rect 89270 40382 89356 40434
rect 89132 40098 89356 40382
rect 89132 40046 89218 40098
rect 89270 40046 89356 40098
rect 89132 39762 89356 40046
rect 89132 39710 89218 39762
rect 89270 39710 89356 39762
rect 89132 39426 89356 39710
rect 89132 39374 89218 39426
rect 89270 39374 89356 39426
rect 89132 39092 89356 39374
rect 89132 39036 89216 39092
rect 89272 39036 89356 39092
rect 89132 38754 89356 39036
rect 89132 38702 89218 38754
rect 89270 38702 89356 38754
rect 89132 38418 89356 38702
rect 89132 38366 89218 38418
rect 89270 38366 89356 38418
rect 89132 38082 89356 38366
rect 89132 38030 89218 38082
rect 89270 38030 89356 38082
rect 89132 37746 89356 38030
rect 89132 37694 89218 37746
rect 89270 37694 89356 37746
rect 89132 37412 89356 37694
rect 89132 37356 89216 37412
rect 89272 37356 89356 37412
rect 89132 37074 89356 37356
rect 89132 37022 89218 37074
rect 89270 37022 89356 37074
rect 89132 36738 89356 37022
rect 89132 36686 89218 36738
rect 89270 36686 89356 36738
rect 89132 36402 89356 36686
rect 89132 36350 89218 36402
rect 89270 36350 89356 36402
rect 89132 36066 89356 36350
rect 89132 36014 89218 36066
rect 89270 36014 89356 36066
rect 89132 35732 89356 36014
rect 89132 35676 89216 35732
rect 89272 35676 89356 35732
rect 89132 35394 89356 35676
rect 89132 35342 89218 35394
rect 89270 35342 89356 35394
rect 89132 35058 89356 35342
rect 89132 35006 89218 35058
rect 89270 35006 89356 35058
rect 89132 34722 89356 35006
rect 89132 34670 89218 34722
rect 89270 34670 89356 34722
rect 89132 34386 89356 34670
rect 89132 34334 89218 34386
rect 89270 34334 89356 34386
rect 89132 34052 89356 34334
rect 89132 33996 89216 34052
rect 89272 33996 89356 34052
rect 89132 33714 89356 33996
rect 89132 33662 89218 33714
rect 89270 33662 89356 33714
rect 89132 33378 89356 33662
rect 89132 33326 89218 33378
rect 89270 33326 89356 33378
rect 89132 33042 89356 33326
rect 89132 32990 89218 33042
rect 89270 32990 89356 33042
rect 89132 32706 89356 32990
rect 89132 32654 89218 32706
rect 89270 32654 89356 32706
rect 89132 32372 89356 32654
rect 89132 32316 89216 32372
rect 89272 32316 89356 32372
rect 89132 32034 89356 32316
rect 89132 31982 89218 32034
rect 89270 31982 89356 32034
rect 89132 31698 89356 31982
rect 89132 31646 89218 31698
rect 89270 31646 89356 31698
rect 89132 31362 89356 31646
rect 89132 31310 89218 31362
rect 89270 31310 89356 31362
rect 89132 31026 89356 31310
rect 89132 30974 89218 31026
rect 89270 30974 89356 31026
rect 89132 30692 89356 30974
rect 89132 30636 89216 30692
rect 89272 30636 89356 30692
rect 89132 30354 89356 30636
rect 89132 30302 89218 30354
rect 89270 30302 89356 30354
rect 89132 30018 89356 30302
rect 89132 29966 89218 30018
rect 89270 29966 89356 30018
rect 89132 29682 89356 29966
rect 89132 29630 89218 29682
rect 89270 29630 89356 29682
rect 89132 29346 89356 29630
rect 89132 29294 89218 29346
rect 89270 29294 89356 29346
rect 89132 29012 89356 29294
rect 89132 28956 89216 29012
rect 89272 28956 89356 29012
rect 89132 28674 89356 28956
rect 89132 28622 89218 28674
rect 89270 28622 89356 28674
rect 89132 28338 89356 28622
rect 89132 28286 89218 28338
rect 89270 28286 89356 28338
rect 89132 28002 89356 28286
rect 89132 27950 89218 28002
rect 89270 27950 89356 28002
rect 89132 27666 89356 27950
rect 89132 27614 89218 27666
rect 89270 27614 89356 27666
rect 89132 27332 89356 27614
rect 89132 27276 89216 27332
rect 89272 27276 89356 27332
rect 89132 26994 89356 27276
rect 89132 26942 89218 26994
rect 89270 26942 89356 26994
rect 89132 26658 89356 26942
rect 89132 26606 89218 26658
rect 89270 26606 89356 26658
rect 89132 26322 89356 26606
rect 89132 26270 89218 26322
rect 89270 26270 89356 26322
rect 89132 25986 89356 26270
rect 89132 25934 89218 25986
rect 89270 25934 89356 25986
rect 89132 25652 89356 25934
rect 89132 25596 89216 25652
rect 89272 25596 89356 25652
rect 89132 25314 89356 25596
rect 89132 25262 89218 25314
rect 89270 25262 89356 25314
rect 89132 24978 89356 25262
rect 89132 24926 89218 24978
rect 89270 24926 89356 24978
rect 89132 24642 89356 24926
rect 89132 24590 89218 24642
rect 89270 24590 89356 24642
rect 89132 24306 89356 24590
rect 89132 24254 89218 24306
rect 89270 24254 89356 24306
rect 89132 23972 89356 24254
rect 89132 23916 89216 23972
rect 89272 23916 89356 23972
rect 89132 23634 89356 23916
rect 89132 23582 89218 23634
rect 89270 23582 89356 23634
rect 89132 23298 89356 23582
rect 89132 23246 89218 23298
rect 89270 23246 89356 23298
rect 89132 22962 89356 23246
rect 89132 22910 89218 22962
rect 89270 22910 89356 22962
rect 89132 22626 89356 22910
rect 89132 22574 89218 22626
rect 89270 22574 89356 22626
rect 89132 22292 89356 22574
rect 89132 22236 89216 22292
rect 89272 22236 89356 22292
rect 89132 21954 89356 22236
rect 89132 21902 89218 21954
rect 89270 21902 89356 21954
rect 89132 21618 89356 21902
rect 89132 21566 89218 21618
rect 89270 21566 89356 21618
rect 89132 21282 89356 21566
rect 89132 21230 89218 21282
rect 89270 21230 89356 21282
rect 89132 20946 89356 21230
rect 89132 20894 89218 20946
rect 89270 20894 89356 20946
rect 89132 20612 89356 20894
rect 89132 20556 89216 20612
rect 89272 20556 89356 20612
rect 89132 20274 89356 20556
rect 89132 20222 89218 20274
rect 89270 20222 89356 20274
rect 79260 19933 79316 19942
rect 19830 18629 19858 19914
rect 79260 19868 79316 19877
rect 89132 19938 89356 20222
rect 89132 19886 89218 19938
rect 89270 19886 89356 19938
rect 80342 19677 80398 19686
rect 79059 19606 79115 19615
rect 79059 19541 79115 19550
rect 79397 19606 79453 19615
rect 80342 19612 80398 19621
rect 79397 19541 79453 19550
rect 89132 19602 89356 19886
rect 89132 19550 89218 19602
rect 89270 19550 89356 19602
rect 19816 18620 19872 18629
rect 19816 18555 19872 18564
rect 23533 15781 23561 19437
rect 23519 15772 23575 15781
rect 23519 15707 23575 15716
rect 23657 12989 23685 19437
rect 23781 14387 23809 19437
rect 89132 19266 89356 19550
rect 89132 19214 89218 19266
rect 89270 19214 89356 19266
rect 89132 18932 89356 19214
rect 89132 18876 89216 18932
rect 89272 18876 89356 18932
rect 89132 18594 89356 18876
rect 89132 18542 89218 18594
rect 89270 18542 89356 18594
rect 89132 18258 89356 18542
rect 89132 18206 89218 18258
rect 89270 18206 89356 18258
rect 78979 18048 79035 18057
rect 78979 17983 79035 17992
rect 79397 18048 79453 18057
rect 79397 17983 79453 17992
rect 80342 17977 80398 17986
rect 80342 17912 80398 17921
rect 89132 17922 89356 18206
rect 89132 17870 89218 17922
rect 89270 17870 89356 17922
rect 89132 17586 89356 17870
rect 89132 17534 89218 17586
rect 89270 17534 89356 17586
rect 89132 17252 89356 17534
rect 89132 17196 89216 17252
rect 89272 17196 89356 17252
rect 89132 16914 89356 17196
rect 89132 16862 89218 16914
rect 89270 16862 89356 16914
rect 80342 16849 80398 16858
rect 78899 16778 78955 16787
rect 78899 16713 78955 16722
rect 79397 16778 79453 16787
rect 80342 16784 80398 16793
rect 79397 16713 79453 16722
rect 89132 16578 89356 16862
rect 89132 16526 89218 16578
rect 89270 16526 89356 16578
rect 89132 16242 89356 16526
rect 89132 16190 89218 16242
rect 89270 16190 89356 16242
rect 89132 15906 89356 16190
rect 89132 15854 89218 15906
rect 89270 15854 89356 15906
rect 89132 15572 89356 15854
rect 89132 15516 89216 15572
rect 89272 15516 89356 15572
rect 89132 15234 89356 15516
rect 78819 15220 78875 15229
rect 78819 15155 78875 15164
rect 79397 15220 79453 15229
rect 79397 15155 79453 15164
rect 89132 15182 89218 15234
rect 89270 15182 89356 15234
rect 80342 15149 80398 15158
rect 80342 15084 80398 15093
rect 89132 14898 89356 15182
rect 89132 14846 89218 14898
rect 89270 14846 89356 14898
rect 89132 14562 89356 14846
rect 89132 14510 89218 14562
rect 89270 14510 89356 14562
rect 23767 14378 23823 14387
rect 23767 14313 23823 14322
rect 89132 14226 89356 14510
rect 89132 14174 89218 14226
rect 89270 14174 89356 14226
rect 80342 14021 80398 14030
rect 78739 13950 78795 13959
rect 78739 13885 78795 13894
rect 79397 13950 79453 13959
rect 80342 13956 80398 13965
rect 79397 13885 79453 13894
rect 89132 13892 89356 14174
rect 89132 13836 89216 13892
rect 89272 13836 89356 13892
rect 89132 13554 89356 13836
rect 89132 13502 89218 13554
rect 89270 13502 89356 13554
rect 89132 13218 89356 13502
rect 89132 13166 89218 13218
rect 89270 13166 89356 13218
rect 25626 13132 25682 13141
rect 25626 13067 25682 13076
rect 30618 13132 30674 13141
rect 30618 13067 30674 13076
rect 35610 13132 35666 13141
rect 35610 13067 35666 13076
rect 40602 13132 40658 13141
rect 40602 13067 40658 13076
rect 45594 13132 45650 13141
rect 45594 13067 45650 13076
rect 50586 13132 50642 13141
rect 50586 13067 50642 13076
rect 55578 13132 55634 13141
rect 55578 13067 55634 13076
rect 60570 13132 60626 13141
rect 60570 13067 60626 13076
rect 23643 12980 23699 12989
rect 23643 12915 23699 12924
rect 89132 12882 89356 13166
rect 89132 12830 89218 12882
rect 89270 12830 89356 12882
rect 89132 12546 89356 12830
rect 89132 12494 89218 12546
rect 89270 12494 89356 12546
rect 78659 12392 78715 12401
rect 78659 12327 78715 12336
rect 79397 12392 79453 12401
rect 79397 12327 79453 12336
rect 80342 12321 80398 12330
rect 80342 12256 80398 12265
rect 89132 12212 89356 12494
rect 89132 12156 89216 12212
rect 89272 12156 89356 12212
rect 89132 11874 89356 12156
rect 89132 11822 89218 11874
rect 89270 11822 89356 11874
rect 89132 11538 89356 11822
rect 89132 11486 89218 11538
rect 89270 11486 89356 11538
rect 89132 11202 89356 11486
rect 80342 11193 80398 11202
rect 78579 11122 78635 11131
rect 78579 11057 78635 11066
rect 79397 11122 79453 11131
rect 80342 11128 80398 11137
rect 89132 11150 89218 11202
rect 89270 11150 89356 11202
rect 79397 11057 79453 11066
rect 5899 8684 5955 8693
rect 11702 8680 11800 8708
rect 5899 8619 5955 8628
rect 2678 8579 2734 8588
rect 2678 8514 2734 8523
rect 1634 8462 1720 8514
rect 1772 8462 1858 8514
rect 1634 8178 1858 8462
rect 1634 8126 1720 8178
rect 1772 8126 1858 8178
rect 1634 7842 1858 8126
rect 1634 7790 1720 7842
rect 1772 7790 1858 7842
rect 1634 7506 1858 7790
rect 1634 7454 1720 7506
rect 1772 7454 1858 7506
rect 1634 7172 1858 7454
rect 1634 7116 1718 7172
rect 1774 7116 1858 7172
rect 1634 6834 1858 7116
rect 1634 6782 1720 6834
rect 1772 6782 1858 6834
rect 1634 6498 1858 6782
rect 1634 6446 1720 6498
rect 1772 6446 1858 6498
rect 1634 6162 1858 6446
rect 1634 6110 1720 6162
rect 1772 6110 1858 6162
rect 1634 5826 1858 6110
rect 1634 5774 1720 5826
rect 1772 5774 1858 5826
rect 1634 5492 1858 5774
rect 1634 5436 1718 5492
rect 1774 5436 1858 5492
rect 1634 5154 1858 5436
rect 1634 5102 1720 5154
rect 1772 5102 1858 5154
rect 1634 4818 1858 5102
rect 1634 4766 1720 4818
rect 1772 4766 1858 4818
rect 1634 4482 1858 4766
rect 1634 4430 1720 4482
rect 1772 4430 1858 4482
rect 1634 4146 1858 4430
rect 1634 4094 1720 4146
rect 1772 4094 1858 4146
rect 1634 3812 1858 4094
rect 1634 3756 1718 3812
rect 1774 3756 1858 3812
rect 1634 3474 1858 3756
rect 1634 3422 1720 3474
rect 1772 3422 1858 3474
rect 1634 3138 1858 3422
rect 1634 3086 1720 3138
rect 1772 3086 1858 3138
rect 1634 2802 1858 3086
rect 1634 2750 1720 2802
rect 1772 2750 1858 2802
rect 11772 2785 11800 8680
rect 89132 10866 89356 11150
rect 89132 10814 89218 10866
rect 89270 10814 89356 10866
rect 89132 10532 89356 10814
rect 89132 10476 89216 10532
rect 89272 10476 89356 10532
rect 89132 10194 89356 10476
rect 89132 10142 89218 10194
rect 89270 10142 89356 10194
rect 89132 9858 89356 10142
rect 89132 9806 89218 9858
rect 89270 9806 89356 9858
rect 89132 9522 89356 9806
rect 89132 9470 89218 9522
rect 89270 9470 89356 9522
rect 89132 9186 89356 9470
rect 89132 9134 89218 9186
rect 89270 9134 89356 9186
rect 89132 8852 89356 9134
rect 89132 8796 89216 8852
rect 89272 8796 89356 8852
rect 89132 8514 89356 8796
rect 89132 8462 89218 8514
rect 89270 8462 89356 8514
rect 89132 8178 89356 8462
rect 89132 8126 89218 8178
rect 89270 8126 89356 8178
rect 89132 7842 89356 8126
rect 89132 7790 89218 7842
rect 89270 7790 89356 7842
rect 89132 7506 89356 7790
rect 89132 7454 89218 7506
rect 89270 7454 89356 7506
rect 89132 7172 89356 7454
rect 89132 7116 89216 7172
rect 89272 7116 89356 7172
rect 89132 6834 89356 7116
rect 89132 6782 89218 6834
rect 89270 6782 89356 6834
rect 89132 6498 89356 6782
rect 89132 6446 89218 6498
rect 89270 6446 89356 6498
rect 89132 6162 89356 6446
rect 89132 6110 89218 6162
rect 89270 6110 89356 6162
rect 89132 5826 89356 6110
rect 89132 5774 89218 5826
rect 89270 5774 89356 5826
rect 89132 5492 89356 5774
rect 89132 5436 89216 5492
rect 89272 5436 89356 5492
rect 89132 5154 89356 5436
rect 89132 5102 89218 5154
rect 89270 5102 89356 5154
rect 89132 4818 89356 5102
rect 89132 4766 89218 4818
rect 89270 4766 89356 4818
rect 89132 4482 89356 4766
rect 89132 4430 89218 4482
rect 89270 4430 89356 4482
rect 89132 4146 89356 4430
rect 89132 4094 89218 4146
rect 89270 4094 89356 4146
rect 89132 3812 89356 4094
rect 89132 3756 89216 3812
rect 89272 3756 89356 3812
rect 89132 3474 89356 3756
rect 89132 3422 89218 3474
rect 89270 3422 89356 3474
rect 89132 3138 89356 3422
rect 89132 3086 89218 3138
rect 89270 3086 89356 3138
rect 13012 3032 13068 3041
rect 13012 2967 13068 2976
rect 14180 3032 14236 3041
rect 14180 2967 14236 2976
rect 15348 3032 15404 3041
rect 15348 2967 15404 2976
rect 16516 3032 16572 3041
rect 16516 2967 16572 2976
rect 17684 3032 17740 3041
rect 17684 2967 17740 2976
rect 18852 3032 18908 3041
rect 18852 2967 18908 2976
rect 20020 3032 20076 3041
rect 20020 2967 20076 2976
rect 21188 3032 21244 3041
rect 21188 2967 21244 2976
rect 22356 3032 22412 3041
rect 22356 2967 22412 2976
rect 23524 3032 23580 3041
rect 23524 2967 23580 2976
rect 24692 3032 24748 3041
rect 24692 2967 24748 2976
rect 25860 3032 25916 3041
rect 25860 2967 25916 2976
rect 89132 2802 89356 3086
rect 1634 2466 1858 2750
rect 11758 2776 11814 2785
rect 11758 2711 11814 2720
rect 89132 2750 89218 2802
rect 89270 2750 89356 2802
rect 1634 2414 1720 2466
rect 1772 2414 1858 2466
rect 1634 2132 1858 2414
rect 1634 2076 1718 2132
rect 1774 2076 1858 2132
rect 1634 1656 1858 2076
rect 89132 2466 89356 2750
rect 89132 2414 89218 2466
rect 89270 2414 89356 2466
rect 89132 2132 89356 2414
rect 89132 2076 89216 2132
rect 89272 2076 89356 2132
rect 2054 1796 2110 1805
rect 2054 1731 2110 1740
rect 3734 1796 3790 1805
rect 3734 1731 3790 1740
rect 5414 1796 5470 1805
rect 5414 1731 5470 1740
rect 7094 1796 7150 1805
rect 7094 1731 7150 1740
rect 8774 1796 8830 1805
rect 8774 1731 8830 1740
rect 10454 1796 10510 1805
rect 10454 1731 10510 1740
rect 12134 1796 12190 1805
rect 12134 1731 12190 1740
rect 13814 1796 13870 1805
rect 13814 1731 13870 1740
rect 15494 1796 15550 1805
rect 15494 1731 15550 1740
rect 17174 1796 17230 1805
rect 17174 1731 17230 1740
rect 18854 1796 18910 1805
rect 18854 1731 18910 1740
rect 20534 1796 20590 1805
rect 20534 1731 20590 1740
rect 22214 1796 22270 1805
rect 22214 1731 22270 1740
rect 23894 1796 23950 1805
rect 23894 1731 23950 1740
rect 25574 1796 25630 1805
rect 25574 1731 25630 1740
rect 27254 1796 27310 1805
rect 27254 1731 27310 1740
rect 28934 1796 28990 1805
rect 28934 1731 28990 1740
rect 30614 1796 30670 1805
rect 30614 1731 30670 1740
rect 32294 1796 32350 1805
rect 32294 1731 32350 1740
rect 33974 1796 34030 1805
rect 33974 1731 34030 1740
rect 35654 1796 35710 1805
rect 35654 1731 35710 1740
rect 37334 1796 37390 1805
rect 37334 1731 37390 1740
rect 39014 1796 39070 1805
rect 39014 1731 39070 1740
rect 40694 1796 40750 1805
rect 40694 1731 40750 1740
rect 42374 1796 42430 1805
rect 42374 1731 42430 1740
rect 44054 1796 44110 1805
rect 44054 1731 44110 1740
rect 45734 1796 45790 1805
rect 45734 1731 45790 1740
rect 47414 1796 47470 1805
rect 47414 1731 47470 1740
rect 49094 1796 49150 1805
rect 49094 1731 49150 1740
rect 50774 1796 50830 1805
rect 50774 1731 50830 1740
rect 52454 1796 52510 1805
rect 52454 1731 52510 1740
rect 54134 1796 54190 1805
rect 54134 1731 54190 1740
rect 55814 1796 55870 1805
rect 55814 1731 55870 1740
rect 57494 1796 57550 1805
rect 57494 1731 57550 1740
rect 59174 1796 59230 1805
rect 59174 1731 59230 1740
rect 60854 1796 60910 1805
rect 60854 1731 60910 1740
rect 62534 1796 62590 1805
rect 62534 1731 62590 1740
rect 64214 1796 64270 1805
rect 64214 1731 64270 1740
rect 65894 1796 65950 1805
rect 65894 1731 65950 1740
rect 67574 1796 67630 1805
rect 67574 1731 67630 1740
rect 69254 1796 69310 1805
rect 69254 1731 69310 1740
rect 70934 1796 70990 1805
rect 70934 1731 70990 1740
rect 72614 1796 72670 1805
rect 72614 1731 72670 1740
rect 74294 1796 74350 1805
rect 74294 1731 74350 1740
rect 75974 1796 76030 1805
rect 75974 1731 76030 1740
rect 77654 1796 77710 1805
rect 77654 1731 77710 1740
rect 79334 1796 79390 1805
rect 79334 1731 79390 1740
rect 81014 1796 81070 1805
rect 81014 1731 81070 1740
rect 82694 1796 82750 1805
rect 82694 1731 82750 1740
rect 84374 1796 84430 1805
rect 84374 1731 84430 1740
rect 86054 1796 86110 1805
rect 86054 1731 86110 1740
rect 87734 1796 87790 1805
rect 87734 1731 87790 1740
rect 89132 1656 89356 2076
<< via2 >>
rect 2054 87522 2110 87524
rect 2054 87470 2056 87522
rect 2056 87470 2108 87522
rect 2108 87470 2110 87522
rect 2054 87468 2110 87470
rect 3734 87522 3790 87524
rect 3734 87470 3736 87522
rect 3736 87470 3788 87522
rect 3788 87470 3790 87522
rect 3734 87468 3790 87470
rect 5414 87522 5470 87524
rect 5414 87470 5416 87522
rect 5416 87470 5468 87522
rect 5468 87470 5470 87522
rect 5414 87468 5470 87470
rect 7094 87522 7150 87524
rect 7094 87470 7096 87522
rect 7096 87470 7148 87522
rect 7148 87470 7150 87522
rect 7094 87468 7150 87470
rect 8774 87522 8830 87524
rect 8774 87470 8776 87522
rect 8776 87470 8828 87522
rect 8828 87470 8830 87522
rect 8774 87468 8830 87470
rect 10454 87522 10510 87524
rect 10454 87470 10456 87522
rect 10456 87470 10508 87522
rect 10508 87470 10510 87522
rect 10454 87468 10510 87470
rect 12134 87522 12190 87524
rect 12134 87470 12136 87522
rect 12136 87470 12188 87522
rect 12188 87470 12190 87522
rect 12134 87468 12190 87470
rect 13814 87522 13870 87524
rect 13814 87470 13816 87522
rect 13816 87470 13868 87522
rect 13868 87470 13870 87522
rect 13814 87468 13870 87470
rect 15494 87522 15550 87524
rect 15494 87470 15496 87522
rect 15496 87470 15548 87522
rect 15548 87470 15550 87522
rect 15494 87468 15550 87470
rect 17174 87522 17230 87524
rect 17174 87470 17176 87522
rect 17176 87470 17228 87522
rect 17228 87470 17230 87522
rect 17174 87468 17230 87470
rect 18854 87522 18910 87524
rect 18854 87470 18856 87522
rect 18856 87470 18908 87522
rect 18908 87470 18910 87522
rect 18854 87468 18910 87470
rect 20534 87522 20590 87524
rect 20534 87470 20536 87522
rect 20536 87470 20588 87522
rect 20588 87470 20590 87522
rect 20534 87468 20590 87470
rect 22214 87522 22270 87524
rect 22214 87470 22216 87522
rect 22216 87470 22268 87522
rect 22268 87470 22270 87522
rect 22214 87468 22270 87470
rect 23894 87522 23950 87524
rect 23894 87470 23896 87522
rect 23896 87470 23948 87522
rect 23948 87470 23950 87522
rect 23894 87468 23950 87470
rect 25574 87522 25630 87524
rect 25574 87470 25576 87522
rect 25576 87470 25628 87522
rect 25628 87470 25630 87522
rect 25574 87468 25630 87470
rect 27254 87522 27310 87524
rect 27254 87470 27256 87522
rect 27256 87470 27308 87522
rect 27308 87470 27310 87522
rect 27254 87468 27310 87470
rect 28934 87522 28990 87524
rect 28934 87470 28936 87522
rect 28936 87470 28988 87522
rect 28988 87470 28990 87522
rect 28934 87468 28990 87470
rect 30614 87522 30670 87524
rect 30614 87470 30616 87522
rect 30616 87470 30668 87522
rect 30668 87470 30670 87522
rect 30614 87468 30670 87470
rect 32294 87522 32350 87524
rect 32294 87470 32296 87522
rect 32296 87470 32348 87522
rect 32348 87470 32350 87522
rect 32294 87468 32350 87470
rect 33974 87522 34030 87524
rect 33974 87470 33976 87522
rect 33976 87470 34028 87522
rect 34028 87470 34030 87522
rect 33974 87468 34030 87470
rect 35654 87522 35710 87524
rect 35654 87470 35656 87522
rect 35656 87470 35708 87522
rect 35708 87470 35710 87522
rect 35654 87468 35710 87470
rect 37334 87522 37390 87524
rect 37334 87470 37336 87522
rect 37336 87470 37388 87522
rect 37388 87470 37390 87522
rect 37334 87468 37390 87470
rect 39014 87522 39070 87524
rect 39014 87470 39016 87522
rect 39016 87470 39068 87522
rect 39068 87470 39070 87522
rect 39014 87468 39070 87470
rect 40694 87522 40750 87524
rect 40694 87470 40696 87522
rect 40696 87470 40748 87522
rect 40748 87470 40750 87522
rect 40694 87468 40750 87470
rect 42374 87522 42430 87524
rect 42374 87470 42376 87522
rect 42376 87470 42428 87522
rect 42428 87470 42430 87522
rect 42374 87468 42430 87470
rect 44054 87522 44110 87524
rect 44054 87470 44056 87522
rect 44056 87470 44108 87522
rect 44108 87470 44110 87522
rect 44054 87468 44110 87470
rect 45734 87522 45790 87524
rect 45734 87470 45736 87522
rect 45736 87470 45788 87522
rect 45788 87470 45790 87522
rect 45734 87468 45790 87470
rect 47414 87522 47470 87524
rect 47414 87470 47416 87522
rect 47416 87470 47468 87522
rect 47468 87470 47470 87522
rect 47414 87468 47470 87470
rect 49094 87522 49150 87524
rect 49094 87470 49096 87522
rect 49096 87470 49148 87522
rect 49148 87470 49150 87522
rect 49094 87468 49150 87470
rect 50774 87522 50830 87524
rect 50774 87470 50776 87522
rect 50776 87470 50828 87522
rect 50828 87470 50830 87522
rect 50774 87468 50830 87470
rect 52454 87522 52510 87524
rect 52454 87470 52456 87522
rect 52456 87470 52508 87522
rect 52508 87470 52510 87522
rect 52454 87468 52510 87470
rect 54134 87522 54190 87524
rect 54134 87470 54136 87522
rect 54136 87470 54188 87522
rect 54188 87470 54190 87522
rect 54134 87468 54190 87470
rect 55814 87522 55870 87524
rect 55814 87470 55816 87522
rect 55816 87470 55868 87522
rect 55868 87470 55870 87522
rect 55814 87468 55870 87470
rect 57494 87522 57550 87524
rect 57494 87470 57496 87522
rect 57496 87470 57548 87522
rect 57548 87470 57550 87522
rect 57494 87468 57550 87470
rect 59174 87522 59230 87524
rect 59174 87470 59176 87522
rect 59176 87470 59228 87522
rect 59228 87470 59230 87522
rect 59174 87468 59230 87470
rect 60854 87522 60910 87524
rect 60854 87470 60856 87522
rect 60856 87470 60908 87522
rect 60908 87470 60910 87522
rect 60854 87468 60910 87470
rect 62534 87522 62590 87524
rect 62534 87470 62536 87522
rect 62536 87470 62588 87522
rect 62588 87470 62590 87522
rect 62534 87468 62590 87470
rect 64214 87522 64270 87524
rect 64214 87470 64216 87522
rect 64216 87470 64268 87522
rect 64268 87470 64270 87522
rect 64214 87468 64270 87470
rect 65894 87522 65950 87524
rect 65894 87470 65896 87522
rect 65896 87470 65948 87522
rect 65948 87470 65950 87522
rect 65894 87468 65950 87470
rect 67574 87522 67630 87524
rect 67574 87470 67576 87522
rect 67576 87470 67628 87522
rect 67628 87470 67630 87522
rect 67574 87468 67630 87470
rect 69254 87522 69310 87524
rect 69254 87470 69256 87522
rect 69256 87470 69308 87522
rect 69308 87470 69310 87522
rect 69254 87468 69310 87470
rect 70934 87522 70990 87524
rect 70934 87470 70936 87522
rect 70936 87470 70988 87522
rect 70988 87470 70990 87522
rect 70934 87468 70990 87470
rect 72614 87522 72670 87524
rect 72614 87470 72616 87522
rect 72616 87470 72668 87522
rect 72668 87470 72670 87522
rect 72614 87468 72670 87470
rect 74294 87522 74350 87524
rect 74294 87470 74296 87522
rect 74296 87470 74348 87522
rect 74348 87470 74350 87522
rect 74294 87468 74350 87470
rect 75974 87522 76030 87524
rect 75974 87470 75976 87522
rect 75976 87470 76028 87522
rect 76028 87470 76030 87522
rect 75974 87468 76030 87470
rect 77654 87522 77710 87524
rect 77654 87470 77656 87522
rect 77656 87470 77708 87522
rect 77708 87470 77710 87522
rect 77654 87468 77710 87470
rect 79334 87522 79390 87524
rect 79334 87470 79336 87522
rect 79336 87470 79388 87522
rect 79388 87470 79390 87522
rect 79334 87468 79390 87470
rect 81014 87522 81070 87524
rect 81014 87470 81016 87522
rect 81016 87470 81068 87522
rect 81068 87470 81070 87522
rect 81014 87468 81070 87470
rect 82694 87522 82750 87524
rect 82694 87470 82696 87522
rect 82696 87470 82748 87522
rect 82748 87470 82750 87522
rect 82694 87468 82750 87470
rect 84374 87522 84430 87524
rect 84374 87470 84376 87522
rect 84376 87470 84428 87522
rect 84428 87470 84430 87522
rect 84374 87468 84430 87470
rect 86054 87522 86110 87524
rect 86054 87470 86056 87522
rect 86056 87470 86108 87522
rect 86108 87470 86110 87522
rect 86054 87468 86110 87470
rect 87734 87522 87790 87524
rect 87734 87470 87736 87522
rect 87736 87470 87788 87522
rect 87788 87470 87790 87522
rect 87734 87468 87790 87470
rect 79260 86488 79316 86544
rect 74502 86232 74558 86288
rect 75670 86232 75726 86288
rect 76838 86232 76894 86288
rect 1718 86130 1774 86132
rect 1718 86078 1720 86130
rect 1720 86078 1772 86130
rect 1772 86078 1774 86130
rect 1718 86076 1774 86078
rect 1718 84450 1774 84452
rect 1718 84398 1720 84450
rect 1720 84398 1772 84450
rect 1772 84398 1774 84450
rect 1718 84396 1774 84398
rect 1718 82770 1774 82772
rect 1718 82718 1720 82770
rect 1720 82718 1772 82770
rect 1772 82718 1774 82770
rect 1718 82716 1774 82718
rect 1718 81090 1774 81092
rect 1718 81038 1720 81090
rect 1720 81038 1772 81090
rect 1772 81038 1774 81090
rect 1718 81036 1774 81038
rect 1718 79410 1774 79412
rect 1718 79358 1720 79410
rect 1720 79358 1772 79410
rect 1772 79358 1774 79410
rect 1718 79356 1774 79358
rect 89216 86130 89272 86132
rect 89216 86078 89218 86130
rect 89218 86078 89270 86130
rect 89270 86078 89272 86130
rect 89216 86076 89272 86078
rect 89216 84450 89272 84452
rect 89216 84398 89218 84450
rect 89218 84398 89270 84450
rect 89270 84398 89272 84450
rect 89216 84396 89272 84398
rect 89216 82770 89272 82772
rect 89216 82718 89218 82770
rect 89218 82718 89270 82770
rect 89270 82718 89272 82770
rect 89216 82716 89272 82718
rect 89216 81090 89272 81092
rect 89216 81038 89218 81090
rect 89218 81038 89270 81090
rect 89270 81038 89272 81090
rect 89216 81036 89272 81038
rect 88256 79579 88312 79635
rect 85119 79474 85175 79530
rect 25626 77908 25682 77910
rect 25626 77856 25628 77908
rect 25628 77856 25680 77908
rect 25680 77856 25682 77908
rect 25626 77854 25682 77856
rect 30618 77908 30674 77910
rect 30618 77856 30620 77908
rect 30620 77856 30672 77908
rect 30672 77856 30674 77908
rect 30618 77854 30674 77856
rect 35610 77908 35666 77910
rect 35610 77856 35612 77908
rect 35612 77856 35664 77908
rect 35664 77856 35666 77908
rect 35610 77854 35666 77856
rect 40602 77908 40658 77910
rect 40602 77856 40604 77908
rect 40604 77856 40656 77908
rect 40656 77856 40658 77908
rect 40602 77854 40658 77856
rect 45594 77908 45650 77910
rect 45594 77856 45596 77908
rect 45596 77856 45648 77908
rect 45648 77856 45650 77908
rect 45594 77854 45650 77856
rect 50586 77908 50642 77910
rect 50586 77856 50588 77908
rect 50588 77856 50640 77908
rect 50640 77856 50642 77908
rect 50586 77854 50642 77856
rect 55578 77908 55634 77910
rect 55578 77856 55580 77908
rect 55580 77856 55632 77908
rect 55632 77856 55634 77908
rect 55578 77854 55634 77856
rect 60570 77908 60626 77910
rect 60570 77856 60572 77908
rect 60572 77856 60624 77908
rect 60624 77856 60626 77908
rect 60570 77854 60626 77856
rect 1718 77730 1774 77732
rect 1718 77678 1720 77730
rect 1720 77678 1772 77730
rect 1772 77678 1774 77730
rect 1718 77676 1774 77678
rect 1718 76050 1774 76052
rect 1718 75998 1720 76050
rect 1720 75998 1772 76050
rect 1772 75998 1774 76050
rect 1718 75996 1774 75998
rect 67133 75198 67189 75254
rect 1718 74370 1774 74372
rect 1718 74318 1720 74370
rect 1720 74318 1772 74370
rect 1772 74318 1774 74370
rect 1718 74316 1774 74318
rect 1718 72690 1774 72692
rect 1718 72638 1720 72690
rect 1720 72638 1772 72690
rect 1772 72638 1774 72690
rect 1718 72636 1774 72638
rect 67257 73780 67313 73836
rect 71118 72366 71174 72422
rect 1718 71010 1774 71012
rect 1718 70958 1720 71010
rect 1720 70958 1772 71010
rect 1772 70958 1774 71010
rect 1718 70956 1774 70958
rect 1718 69330 1774 69332
rect 1718 69278 1720 69330
rect 1720 69278 1772 69330
rect 1772 69278 1774 69330
rect 1718 69276 1774 69278
rect 1718 67650 1774 67652
rect 1718 67598 1720 67650
rect 1720 67598 1772 67650
rect 1772 67598 1774 67650
rect 1718 67596 1774 67598
rect 1718 65970 1774 65972
rect 1718 65918 1720 65970
rect 1720 65918 1772 65970
rect 1772 65918 1774 65970
rect 1718 65916 1774 65918
rect 1718 64290 1774 64292
rect 1718 64238 1720 64290
rect 1720 64238 1772 64290
rect 1772 64238 1774 64290
rect 1718 64236 1774 64238
rect 1718 62610 1774 62612
rect 1718 62558 1720 62610
rect 1720 62558 1772 62610
rect 1772 62558 1774 62610
rect 1718 62556 1774 62558
rect 1718 60930 1774 60932
rect 1718 60878 1720 60930
rect 1720 60878 1772 60930
rect 1772 60878 1774 60930
rect 1718 60876 1774 60878
rect 1718 59250 1774 59252
rect 1718 59198 1720 59250
rect 1720 59198 1772 59250
rect 1772 59198 1774 59250
rect 1718 59196 1774 59198
rect 1718 57570 1774 57572
rect 1718 57518 1720 57570
rect 1720 57518 1772 57570
rect 1772 57518 1774 57570
rect 1718 57516 1774 57518
rect 1718 55890 1774 55892
rect 1718 55838 1720 55890
rect 1720 55838 1772 55890
rect 1772 55838 1774 55890
rect 1718 55836 1774 55838
rect 1718 54210 1774 54212
rect 1718 54158 1720 54210
rect 1720 54158 1772 54210
rect 1772 54158 1774 54210
rect 1718 54156 1774 54158
rect 1718 52530 1774 52532
rect 1718 52478 1720 52530
rect 1720 52478 1772 52530
rect 1772 52478 1774 52530
rect 1718 52476 1774 52478
rect 1718 50850 1774 50852
rect 1718 50798 1720 50850
rect 1720 50798 1772 50850
rect 1772 50798 1774 50850
rect 1718 50796 1774 50798
rect 1718 49170 1774 49172
rect 1718 49118 1720 49170
rect 1720 49118 1772 49170
rect 1772 49118 1774 49170
rect 1718 49116 1774 49118
rect 1718 47490 1774 47492
rect 1718 47438 1720 47490
rect 1720 47438 1772 47490
rect 1772 47438 1774 47490
rect 1718 47436 1774 47438
rect 1718 45810 1774 45812
rect 1718 45758 1720 45810
rect 1720 45758 1772 45810
rect 1772 45758 1774 45810
rect 1718 45756 1774 45758
rect 1718 44130 1774 44132
rect 1718 44078 1720 44130
rect 1720 44078 1772 44130
rect 1772 44078 1774 44130
rect 1718 44076 1774 44078
rect 1718 42450 1774 42452
rect 1718 42398 1720 42450
rect 1720 42398 1772 42450
rect 1772 42398 1774 42450
rect 1718 42396 1774 42398
rect 1718 40770 1774 40772
rect 1718 40718 1720 40770
rect 1720 40718 1772 40770
rect 1772 40718 1774 40770
rect 1718 40716 1774 40718
rect 1718 39090 1774 39092
rect 1718 39038 1720 39090
rect 1720 39038 1772 39090
rect 1772 39038 1774 39090
rect 1718 39036 1774 39038
rect 1718 37410 1774 37412
rect 1718 37358 1720 37410
rect 1720 37358 1772 37410
rect 1772 37358 1774 37410
rect 1718 37356 1774 37358
rect 11621 37204 11677 37260
rect 12355 37258 12411 37260
rect 12355 37206 12357 37258
rect 12357 37206 12409 37258
rect 12409 37206 12411 37258
rect 12355 37204 12411 37206
rect 10676 37133 10732 37189
rect 10676 36005 10732 36061
rect 11621 35934 11677 35990
rect 12275 35988 12331 35990
rect 12275 35936 12277 35988
rect 12277 35936 12329 35988
rect 12329 35936 12331 35988
rect 12275 35934 12331 35936
rect 1718 35730 1774 35732
rect 1718 35678 1720 35730
rect 1720 35678 1772 35730
rect 1772 35678 1774 35730
rect 1718 35676 1774 35678
rect 11621 34376 11677 34432
rect 12195 34430 12251 34432
rect 12195 34378 12197 34430
rect 12197 34378 12249 34430
rect 12249 34378 12251 34430
rect 12195 34376 12251 34378
rect 10676 34305 10732 34361
rect 1718 34050 1774 34052
rect 1718 33998 1720 34050
rect 1720 33998 1772 34050
rect 1772 33998 1774 34050
rect 1718 33996 1774 33998
rect 10676 33177 10732 33233
rect 11621 33106 11677 33162
rect 12115 33160 12171 33162
rect 12115 33108 12117 33160
rect 12117 33108 12169 33160
rect 12169 33108 12171 33160
rect 12115 33106 12171 33108
rect 1718 32370 1774 32372
rect 1718 32318 1720 32370
rect 1720 32318 1772 32370
rect 1772 32318 1774 32370
rect 1718 32316 1774 32318
rect 11621 31548 11677 31604
rect 12035 31602 12091 31604
rect 12035 31550 12037 31602
rect 12037 31550 12089 31602
rect 12089 31550 12091 31602
rect 12035 31548 12091 31550
rect 10676 31477 10732 31533
rect 1718 30690 1774 30692
rect 1718 30638 1720 30690
rect 1720 30638 1772 30690
rect 1772 30638 1774 30690
rect 1718 30636 1774 30638
rect 10676 30349 10732 30405
rect 11621 30278 11677 30334
rect 11955 30332 12011 30334
rect 11955 30280 11957 30332
rect 11957 30280 12009 30332
rect 12009 30280 12011 30332
rect 11955 30278 12011 30280
rect 1718 29010 1774 29012
rect 1718 28958 1720 29010
rect 1720 28958 1772 29010
rect 1772 28958 1774 29010
rect 1718 28956 1774 28958
rect 11621 28720 11677 28776
rect 11875 28774 11931 28776
rect 11875 28722 11877 28774
rect 11877 28722 11929 28774
rect 11929 28722 11931 28774
rect 11875 28720 11931 28722
rect 10676 28649 10732 28705
rect 11758 28393 11814 28449
rect 1718 27330 1774 27332
rect 1718 27278 1720 27330
rect 1720 27278 1772 27330
rect 1772 27278 1774 27330
rect 1718 27276 1774 27278
rect 2465 25672 2521 25728
rect 1718 25650 1774 25652
rect 1718 25598 1720 25650
rect 1720 25598 1772 25650
rect 1772 25598 1774 25650
rect 1718 25596 1774 25598
rect 1718 23970 1774 23972
rect 1718 23918 1720 23970
rect 1720 23918 1772 23970
rect 1772 23918 1774 23970
rect 1718 23916 1774 23918
rect 1718 22290 1774 22292
rect 1718 22238 1720 22290
rect 1720 22238 1772 22290
rect 1772 22238 1774 22290
rect 1718 22236 1774 22238
rect 1718 20610 1774 20612
rect 1718 20558 1720 20610
rect 1720 20558 1772 20610
rect 1772 20558 1774 20610
rect 1718 20556 1774 20558
rect 1718 18930 1774 18932
rect 1718 18878 1720 18930
rect 1720 18878 1772 18930
rect 1772 18878 1774 18930
rect 1718 18876 1774 18878
rect 11674 18564 11730 18620
rect 1718 17250 1774 17252
rect 1718 17198 1720 17250
rect 1720 17198 1772 17250
rect 1772 17198 1774 17250
rect 1718 17196 1774 17198
rect 11674 15736 11730 15792
rect 1718 15570 1774 15572
rect 1718 15518 1720 15570
rect 1720 15518 1772 15570
rect 1772 15518 1774 15570
rect 1718 15516 1774 15518
rect 11674 14322 11730 14378
rect 1718 13890 1774 13892
rect 1718 13838 1720 13890
rect 1720 13838 1772 13890
rect 1772 13838 1774 13890
rect 1718 13836 1774 13838
rect 11674 12924 11730 12980
rect 1718 12210 1774 12212
rect 1718 12158 1720 12210
rect 1720 12158 1772 12210
rect 1772 12158 1774 12210
rect 1718 12156 1774 12158
rect 1718 10530 1774 10532
rect 1718 10478 1720 10530
rect 1720 10478 1772 10530
rect 1772 10478 1774 10530
rect 1718 10476 1774 10478
rect 2678 10223 2734 10279
rect 1718 8850 1774 8852
rect 1718 8798 1720 8850
rect 1720 8798 1772 8850
rect 1772 8798 1774 8850
rect 1718 8796 1774 8798
rect 89216 79410 89272 79412
rect 89216 79358 89218 79410
rect 89218 79358 89270 79410
rect 89270 79358 89272 79410
rect 89216 79356 89272 79358
rect 89216 77730 89272 77732
rect 89216 77678 89218 77730
rect 89218 77678 89270 77730
rect 89270 77678 89272 77730
rect 89216 77676 89272 77678
rect 89216 76050 89272 76052
rect 89216 75998 89218 76050
rect 89218 75998 89270 76050
rect 89270 75998 89272 76050
rect 89216 75996 89272 75998
rect 79344 75178 79400 75234
rect 89216 74370 89272 74372
rect 89216 74318 89218 74370
rect 89218 74318 89270 74370
rect 89270 74318 89272 74370
rect 89216 74316 89272 74318
rect 79344 73780 79400 73836
rect 89216 72690 89272 72692
rect 89216 72638 89218 72690
rect 89218 72638 89270 72690
rect 89270 72638 89272 72690
rect 89216 72636 89272 72638
rect 79344 72366 79400 72422
rect 89216 71010 89272 71012
rect 89216 70958 89218 71010
rect 89218 70958 89270 71010
rect 89270 70958 89272 71010
rect 89216 70956 89272 70958
rect 89216 69330 89272 69332
rect 89216 69278 89218 69330
rect 89218 69278 89270 69330
rect 89270 69278 89272 69330
rect 89216 69276 89272 69278
rect 89216 67650 89272 67652
rect 89216 67598 89218 67650
rect 89218 67598 89270 67650
rect 89270 67598 89272 67650
rect 89216 67596 89272 67598
rect 89216 65970 89272 65972
rect 89216 65918 89218 65970
rect 89218 65918 89270 65970
rect 89270 65918 89272 65970
rect 89216 65916 89272 65918
rect 89216 64290 89272 64292
rect 89216 64238 89218 64290
rect 89218 64238 89270 64290
rect 89270 64238 89272 64290
rect 89216 64236 89272 64238
rect 89216 62610 89272 62612
rect 89216 62558 89218 62610
rect 89218 62558 89270 62610
rect 89270 62558 89272 62610
rect 89216 62556 89272 62558
rect 88469 62430 88525 62486
rect 89216 60930 89272 60932
rect 89216 60878 89218 60930
rect 89218 60878 89270 60930
rect 89270 60878 89272 60930
rect 89216 60876 89272 60878
rect 89216 59250 89272 59252
rect 89216 59198 89218 59250
rect 89218 59198 89270 59250
rect 89270 59198 89272 59250
rect 89216 59196 89272 59198
rect 89216 57570 89272 57572
rect 89216 57518 89218 57570
rect 89218 57518 89270 57570
rect 89270 57518 89272 57570
rect 89216 57516 89272 57518
rect 89216 55890 89272 55892
rect 89216 55838 89218 55890
rect 89218 55838 89270 55890
rect 89270 55838 89272 55890
rect 89216 55836 89272 55838
rect 89216 54210 89272 54212
rect 89216 54158 89218 54210
rect 89218 54158 89270 54210
rect 89270 54158 89272 54210
rect 89216 54156 89272 54158
rect 89216 52530 89272 52532
rect 89216 52478 89218 52530
rect 89218 52478 89270 52530
rect 89270 52478 89272 52530
rect 89216 52476 89272 52478
rect 89216 50850 89272 50852
rect 89216 50798 89218 50850
rect 89218 50798 89270 50850
rect 89270 50798 89272 50850
rect 89216 50796 89272 50798
rect 89216 49170 89272 49172
rect 89216 49118 89218 49170
rect 89218 49118 89270 49170
rect 89270 49118 89272 49170
rect 89216 49116 89272 49118
rect 89216 47490 89272 47492
rect 89216 47438 89218 47490
rect 89218 47438 89270 47490
rect 89270 47438 89272 47490
rect 89216 47436 89272 47438
rect 89216 45810 89272 45812
rect 89216 45758 89218 45810
rect 89218 45758 89270 45810
rect 89270 45758 89272 45810
rect 89216 45756 89272 45758
rect 89216 44130 89272 44132
rect 89216 44078 89218 44130
rect 89218 44078 89270 44130
rect 89270 44078 89272 44130
rect 89216 44076 89272 44078
rect 89216 42450 89272 42452
rect 89216 42398 89218 42450
rect 89218 42398 89270 42450
rect 89270 42398 89272 42450
rect 89216 42396 89272 42398
rect 89216 40770 89272 40772
rect 89216 40718 89218 40770
rect 89218 40718 89270 40770
rect 89270 40718 89272 40770
rect 89216 40716 89272 40718
rect 89216 39090 89272 39092
rect 89216 39038 89218 39090
rect 89218 39038 89270 39090
rect 89270 39038 89272 39090
rect 89216 39036 89272 39038
rect 89216 37410 89272 37412
rect 89216 37358 89218 37410
rect 89218 37358 89270 37410
rect 89270 37358 89272 37410
rect 89216 37356 89272 37358
rect 89216 35730 89272 35732
rect 89216 35678 89218 35730
rect 89218 35678 89270 35730
rect 89270 35678 89272 35730
rect 89216 35676 89272 35678
rect 89216 34050 89272 34052
rect 89216 33998 89218 34050
rect 89218 33998 89270 34050
rect 89270 33998 89272 34050
rect 89216 33996 89272 33998
rect 89216 32370 89272 32372
rect 89216 32318 89218 32370
rect 89218 32318 89270 32370
rect 89270 32318 89272 32370
rect 89216 32316 89272 32318
rect 89216 30690 89272 30692
rect 89216 30638 89218 30690
rect 89218 30638 89270 30690
rect 89270 30638 89272 30690
rect 89216 30636 89272 30638
rect 89216 29010 89272 29012
rect 89216 28958 89218 29010
rect 89218 28958 89270 29010
rect 89270 28958 89272 29010
rect 89216 28956 89272 28958
rect 89216 27330 89272 27332
rect 89216 27278 89218 27330
rect 89218 27278 89270 27330
rect 89270 27278 89272 27330
rect 89216 27276 89272 27278
rect 89216 25650 89272 25652
rect 89216 25598 89218 25650
rect 89218 25598 89270 25650
rect 89270 25598 89272 25650
rect 89216 25596 89272 25598
rect 89216 23970 89272 23972
rect 89216 23918 89218 23970
rect 89218 23918 89270 23970
rect 89270 23918 89272 23970
rect 89216 23916 89272 23918
rect 89216 22290 89272 22292
rect 89216 22238 89218 22290
rect 89218 22238 89270 22290
rect 89270 22238 89272 22290
rect 89216 22236 89272 22238
rect 89216 20610 89272 20612
rect 89216 20558 89218 20610
rect 89218 20558 89270 20610
rect 89270 20558 89272 20610
rect 89216 20556 89272 20558
rect 79260 19877 79316 19933
rect 80342 19621 80398 19677
rect 79059 19604 79115 19606
rect 79059 19552 79061 19604
rect 79061 19552 79113 19604
rect 79113 19552 79115 19604
rect 79059 19550 79115 19552
rect 79397 19550 79453 19606
rect 19816 18564 19872 18620
rect 23519 15716 23575 15772
rect 89216 18930 89272 18932
rect 89216 18878 89218 18930
rect 89218 18878 89270 18930
rect 89270 18878 89272 18930
rect 89216 18876 89272 18878
rect 78979 18046 79035 18048
rect 78979 17994 78981 18046
rect 78981 17994 79033 18046
rect 79033 17994 79035 18046
rect 78979 17992 79035 17994
rect 79397 17992 79453 18048
rect 80342 17921 80398 17977
rect 89216 17250 89272 17252
rect 89216 17198 89218 17250
rect 89218 17198 89270 17250
rect 89270 17198 89272 17250
rect 89216 17196 89272 17198
rect 80342 16793 80398 16849
rect 78899 16776 78955 16778
rect 78899 16724 78901 16776
rect 78901 16724 78953 16776
rect 78953 16724 78955 16776
rect 78899 16722 78955 16724
rect 79397 16722 79453 16778
rect 89216 15570 89272 15572
rect 89216 15518 89218 15570
rect 89218 15518 89270 15570
rect 89270 15518 89272 15570
rect 89216 15516 89272 15518
rect 78819 15218 78875 15220
rect 78819 15166 78821 15218
rect 78821 15166 78873 15218
rect 78873 15166 78875 15218
rect 78819 15164 78875 15166
rect 79397 15164 79453 15220
rect 80342 15093 80398 15149
rect 23767 14322 23823 14378
rect 80342 13965 80398 14021
rect 78739 13948 78795 13950
rect 78739 13896 78741 13948
rect 78741 13896 78793 13948
rect 78793 13896 78795 13948
rect 78739 13894 78795 13896
rect 79397 13894 79453 13950
rect 89216 13890 89272 13892
rect 89216 13838 89218 13890
rect 89218 13838 89270 13890
rect 89270 13838 89272 13890
rect 89216 13836 89272 13838
rect 25626 13130 25682 13132
rect 25626 13078 25628 13130
rect 25628 13078 25680 13130
rect 25680 13078 25682 13130
rect 25626 13076 25682 13078
rect 30618 13130 30674 13132
rect 30618 13078 30620 13130
rect 30620 13078 30672 13130
rect 30672 13078 30674 13130
rect 30618 13076 30674 13078
rect 35610 13130 35666 13132
rect 35610 13078 35612 13130
rect 35612 13078 35664 13130
rect 35664 13078 35666 13130
rect 35610 13076 35666 13078
rect 40602 13130 40658 13132
rect 40602 13078 40604 13130
rect 40604 13078 40656 13130
rect 40656 13078 40658 13130
rect 40602 13076 40658 13078
rect 45594 13130 45650 13132
rect 45594 13078 45596 13130
rect 45596 13078 45648 13130
rect 45648 13078 45650 13130
rect 45594 13076 45650 13078
rect 50586 13130 50642 13132
rect 50586 13078 50588 13130
rect 50588 13078 50640 13130
rect 50640 13078 50642 13130
rect 50586 13076 50642 13078
rect 55578 13130 55634 13132
rect 55578 13078 55580 13130
rect 55580 13078 55632 13130
rect 55632 13078 55634 13130
rect 55578 13076 55634 13078
rect 60570 13130 60626 13132
rect 60570 13078 60572 13130
rect 60572 13078 60624 13130
rect 60624 13078 60626 13130
rect 60570 13076 60626 13078
rect 23643 12924 23699 12980
rect 78659 12390 78715 12392
rect 78659 12338 78661 12390
rect 78661 12338 78713 12390
rect 78713 12338 78715 12390
rect 78659 12336 78715 12338
rect 79397 12336 79453 12392
rect 80342 12265 80398 12321
rect 89216 12210 89272 12212
rect 89216 12158 89218 12210
rect 89218 12158 89270 12210
rect 89270 12158 89272 12210
rect 89216 12156 89272 12158
rect 80342 11137 80398 11193
rect 78579 11120 78635 11122
rect 78579 11068 78581 11120
rect 78581 11068 78633 11120
rect 78633 11068 78635 11120
rect 78579 11066 78635 11068
rect 79397 11066 79453 11122
rect 5899 8628 5955 8684
rect 2678 8523 2734 8579
rect 1718 7170 1774 7172
rect 1718 7118 1720 7170
rect 1720 7118 1772 7170
rect 1772 7118 1774 7170
rect 1718 7116 1774 7118
rect 1718 5490 1774 5492
rect 1718 5438 1720 5490
rect 1720 5438 1772 5490
rect 1772 5438 1774 5490
rect 1718 5436 1774 5438
rect 1718 3810 1774 3812
rect 1718 3758 1720 3810
rect 1720 3758 1772 3810
rect 1772 3758 1774 3810
rect 1718 3756 1774 3758
rect 89216 10530 89272 10532
rect 89216 10478 89218 10530
rect 89218 10478 89270 10530
rect 89270 10478 89272 10530
rect 89216 10476 89272 10478
rect 89216 8850 89272 8852
rect 89216 8798 89218 8850
rect 89218 8798 89270 8850
rect 89270 8798 89272 8850
rect 89216 8796 89272 8798
rect 89216 7170 89272 7172
rect 89216 7118 89218 7170
rect 89218 7118 89270 7170
rect 89270 7118 89272 7170
rect 89216 7116 89272 7118
rect 89216 5490 89272 5492
rect 89216 5438 89218 5490
rect 89218 5438 89270 5490
rect 89270 5438 89272 5490
rect 89216 5436 89272 5438
rect 89216 3810 89272 3812
rect 89216 3758 89218 3810
rect 89218 3758 89270 3810
rect 89270 3758 89272 3810
rect 89216 3756 89272 3758
rect 13012 2976 13068 3032
rect 14180 2976 14236 3032
rect 15348 2976 15404 3032
rect 16516 2976 16572 3032
rect 17684 2976 17740 3032
rect 18852 2976 18908 3032
rect 20020 2976 20076 3032
rect 21188 2976 21244 3032
rect 22356 2976 22412 3032
rect 23524 2976 23580 3032
rect 24692 2976 24748 3032
rect 25860 2976 25916 3032
rect 11758 2720 11814 2776
rect 1718 2130 1774 2132
rect 1718 2078 1720 2130
rect 1720 2078 1772 2130
rect 1772 2078 1774 2130
rect 1718 2076 1774 2078
rect 89216 2130 89272 2132
rect 89216 2078 89218 2130
rect 89218 2078 89270 2130
rect 89270 2078 89272 2130
rect 89216 2076 89272 2078
rect 2054 1794 2110 1796
rect 2054 1742 2056 1794
rect 2056 1742 2108 1794
rect 2108 1742 2110 1794
rect 2054 1740 2110 1742
rect 3734 1794 3790 1796
rect 3734 1742 3736 1794
rect 3736 1742 3788 1794
rect 3788 1742 3790 1794
rect 3734 1740 3790 1742
rect 5414 1794 5470 1796
rect 5414 1742 5416 1794
rect 5416 1742 5468 1794
rect 5468 1742 5470 1794
rect 5414 1740 5470 1742
rect 7094 1794 7150 1796
rect 7094 1742 7096 1794
rect 7096 1742 7148 1794
rect 7148 1742 7150 1794
rect 7094 1740 7150 1742
rect 8774 1794 8830 1796
rect 8774 1742 8776 1794
rect 8776 1742 8828 1794
rect 8828 1742 8830 1794
rect 8774 1740 8830 1742
rect 10454 1794 10510 1796
rect 10454 1742 10456 1794
rect 10456 1742 10508 1794
rect 10508 1742 10510 1794
rect 10454 1740 10510 1742
rect 12134 1794 12190 1796
rect 12134 1742 12136 1794
rect 12136 1742 12188 1794
rect 12188 1742 12190 1794
rect 12134 1740 12190 1742
rect 13814 1794 13870 1796
rect 13814 1742 13816 1794
rect 13816 1742 13868 1794
rect 13868 1742 13870 1794
rect 13814 1740 13870 1742
rect 15494 1794 15550 1796
rect 15494 1742 15496 1794
rect 15496 1742 15548 1794
rect 15548 1742 15550 1794
rect 15494 1740 15550 1742
rect 17174 1794 17230 1796
rect 17174 1742 17176 1794
rect 17176 1742 17228 1794
rect 17228 1742 17230 1794
rect 17174 1740 17230 1742
rect 18854 1794 18910 1796
rect 18854 1742 18856 1794
rect 18856 1742 18908 1794
rect 18908 1742 18910 1794
rect 18854 1740 18910 1742
rect 20534 1794 20590 1796
rect 20534 1742 20536 1794
rect 20536 1742 20588 1794
rect 20588 1742 20590 1794
rect 20534 1740 20590 1742
rect 22214 1794 22270 1796
rect 22214 1742 22216 1794
rect 22216 1742 22268 1794
rect 22268 1742 22270 1794
rect 22214 1740 22270 1742
rect 23894 1794 23950 1796
rect 23894 1742 23896 1794
rect 23896 1742 23948 1794
rect 23948 1742 23950 1794
rect 23894 1740 23950 1742
rect 25574 1794 25630 1796
rect 25574 1742 25576 1794
rect 25576 1742 25628 1794
rect 25628 1742 25630 1794
rect 25574 1740 25630 1742
rect 27254 1794 27310 1796
rect 27254 1742 27256 1794
rect 27256 1742 27308 1794
rect 27308 1742 27310 1794
rect 27254 1740 27310 1742
rect 28934 1794 28990 1796
rect 28934 1742 28936 1794
rect 28936 1742 28988 1794
rect 28988 1742 28990 1794
rect 28934 1740 28990 1742
rect 30614 1794 30670 1796
rect 30614 1742 30616 1794
rect 30616 1742 30668 1794
rect 30668 1742 30670 1794
rect 30614 1740 30670 1742
rect 32294 1794 32350 1796
rect 32294 1742 32296 1794
rect 32296 1742 32348 1794
rect 32348 1742 32350 1794
rect 32294 1740 32350 1742
rect 33974 1794 34030 1796
rect 33974 1742 33976 1794
rect 33976 1742 34028 1794
rect 34028 1742 34030 1794
rect 33974 1740 34030 1742
rect 35654 1794 35710 1796
rect 35654 1742 35656 1794
rect 35656 1742 35708 1794
rect 35708 1742 35710 1794
rect 35654 1740 35710 1742
rect 37334 1794 37390 1796
rect 37334 1742 37336 1794
rect 37336 1742 37388 1794
rect 37388 1742 37390 1794
rect 37334 1740 37390 1742
rect 39014 1794 39070 1796
rect 39014 1742 39016 1794
rect 39016 1742 39068 1794
rect 39068 1742 39070 1794
rect 39014 1740 39070 1742
rect 40694 1794 40750 1796
rect 40694 1742 40696 1794
rect 40696 1742 40748 1794
rect 40748 1742 40750 1794
rect 40694 1740 40750 1742
rect 42374 1794 42430 1796
rect 42374 1742 42376 1794
rect 42376 1742 42428 1794
rect 42428 1742 42430 1794
rect 42374 1740 42430 1742
rect 44054 1794 44110 1796
rect 44054 1742 44056 1794
rect 44056 1742 44108 1794
rect 44108 1742 44110 1794
rect 44054 1740 44110 1742
rect 45734 1794 45790 1796
rect 45734 1742 45736 1794
rect 45736 1742 45788 1794
rect 45788 1742 45790 1794
rect 45734 1740 45790 1742
rect 47414 1794 47470 1796
rect 47414 1742 47416 1794
rect 47416 1742 47468 1794
rect 47468 1742 47470 1794
rect 47414 1740 47470 1742
rect 49094 1794 49150 1796
rect 49094 1742 49096 1794
rect 49096 1742 49148 1794
rect 49148 1742 49150 1794
rect 49094 1740 49150 1742
rect 50774 1794 50830 1796
rect 50774 1742 50776 1794
rect 50776 1742 50828 1794
rect 50828 1742 50830 1794
rect 50774 1740 50830 1742
rect 52454 1794 52510 1796
rect 52454 1742 52456 1794
rect 52456 1742 52508 1794
rect 52508 1742 52510 1794
rect 52454 1740 52510 1742
rect 54134 1794 54190 1796
rect 54134 1742 54136 1794
rect 54136 1742 54188 1794
rect 54188 1742 54190 1794
rect 54134 1740 54190 1742
rect 55814 1794 55870 1796
rect 55814 1742 55816 1794
rect 55816 1742 55868 1794
rect 55868 1742 55870 1794
rect 55814 1740 55870 1742
rect 57494 1794 57550 1796
rect 57494 1742 57496 1794
rect 57496 1742 57548 1794
rect 57548 1742 57550 1794
rect 57494 1740 57550 1742
rect 59174 1794 59230 1796
rect 59174 1742 59176 1794
rect 59176 1742 59228 1794
rect 59228 1742 59230 1794
rect 59174 1740 59230 1742
rect 60854 1794 60910 1796
rect 60854 1742 60856 1794
rect 60856 1742 60908 1794
rect 60908 1742 60910 1794
rect 60854 1740 60910 1742
rect 62534 1794 62590 1796
rect 62534 1742 62536 1794
rect 62536 1742 62588 1794
rect 62588 1742 62590 1794
rect 62534 1740 62590 1742
rect 64214 1794 64270 1796
rect 64214 1742 64216 1794
rect 64216 1742 64268 1794
rect 64268 1742 64270 1794
rect 64214 1740 64270 1742
rect 65894 1794 65950 1796
rect 65894 1742 65896 1794
rect 65896 1742 65948 1794
rect 65948 1742 65950 1794
rect 65894 1740 65950 1742
rect 67574 1794 67630 1796
rect 67574 1742 67576 1794
rect 67576 1742 67628 1794
rect 67628 1742 67630 1794
rect 67574 1740 67630 1742
rect 69254 1794 69310 1796
rect 69254 1742 69256 1794
rect 69256 1742 69308 1794
rect 69308 1742 69310 1794
rect 69254 1740 69310 1742
rect 70934 1794 70990 1796
rect 70934 1742 70936 1794
rect 70936 1742 70988 1794
rect 70988 1742 70990 1794
rect 70934 1740 70990 1742
rect 72614 1794 72670 1796
rect 72614 1742 72616 1794
rect 72616 1742 72668 1794
rect 72668 1742 72670 1794
rect 72614 1740 72670 1742
rect 74294 1794 74350 1796
rect 74294 1742 74296 1794
rect 74296 1742 74348 1794
rect 74348 1742 74350 1794
rect 74294 1740 74350 1742
rect 75974 1794 76030 1796
rect 75974 1742 75976 1794
rect 75976 1742 76028 1794
rect 76028 1742 76030 1794
rect 75974 1740 76030 1742
rect 77654 1794 77710 1796
rect 77654 1742 77656 1794
rect 77656 1742 77708 1794
rect 77708 1742 77710 1794
rect 77654 1740 77710 1742
rect 79334 1794 79390 1796
rect 79334 1742 79336 1794
rect 79336 1742 79388 1794
rect 79388 1742 79390 1794
rect 79334 1740 79390 1742
rect 81014 1794 81070 1796
rect 81014 1742 81016 1794
rect 81016 1742 81068 1794
rect 81068 1742 81070 1794
rect 81014 1740 81070 1742
rect 82694 1794 82750 1796
rect 82694 1742 82696 1794
rect 82696 1742 82748 1794
rect 82748 1742 82750 1794
rect 82694 1740 82750 1742
rect 84374 1794 84430 1796
rect 84374 1742 84376 1794
rect 84376 1742 84428 1794
rect 84428 1742 84430 1794
rect 84374 1740 84430 1742
rect 86054 1794 86110 1796
rect 86054 1742 86056 1794
rect 86056 1742 86108 1794
rect 86108 1742 86110 1794
rect 86054 1740 86110 1742
rect 87734 1794 87790 1796
rect 87734 1742 87736 1794
rect 87736 1742 87788 1794
rect 87788 1742 87790 1794
rect 87734 1740 87790 1742
<< metal3 >>
rect 272 89014 90788 89020
rect 272 88950 278 89014
rect 342 88950 414 89014
rect 478 88950 550 89014
rect 614 88950 90446 89014
rect 90510 88950 90582 89014
rect 90646 88950 90718 89014
rect 90782 88950 90788 89014
rect 272 88878 90788 88950
rect 272 88814 278 88878
rect 342 88814 414 88878
rect 478 88814 550 88878
rect 614 88814 90446 88878
rect 90510 88814 90582 88878
rect 90646 88814 90718 88878
rect 90782 88814 90788 88878
rect 272 88742 90788 88814
rect 272 88678 278 88742
rect 342 88678 414 88742
rect 478 88678 550 88742
rect 614 88678 73990 88742
rect 74054 88678 90446 88742
rect 90510 88678 90582 88742
rect 90646 88678 90718 88742
rect 90782 88678 90788 88742
rect 272 88672 90788 88678
rect 952 88334 90108 88340
rect 952 88270 958 88334
rect 1022 88270 1094 88334
rect 1158 88270 1230 88334
rect 1294 88270 89766 88334
rect 89830 88270 89902 88334
rect 89966 88270 90038 88334
rect 90102 88270 90108 88334
rect 952 88198 90108 88270
rect 952 88134 958 88198
rect 1022 88134 1094 88198
rect 1158 88134 1230 88198
rect 1294 88134 89766 88198
rect 89830 88134 89902 88198
rect 89966 88134 90038 88198
rect 90102 88134 90108 88198
rect 952 88062 90108 88134
rect 952 87998 958 88062
rect 1022 87998 1094 88062
rect 1158 87998 1230 88062
rect 1294 87998 2182 88062
rect 2246 87998 3814 88062
rect 3878 87998 5310 88062
rect 5374 87998 7078 88062
rect 7142 87998 8846 88062
rect 8910 87998 10342 88062
rect 10406 87998 12110 88062
rect 12174 87998 13878 88062
rect 13942 87998 15374 88062
rect 15438 87998 17278 88062
rect 17342 87998 18910 88062
rect 18974 87998 20542 88062
rect 20606 87998 22174 88062
rect 22238 87998 23942 88062
rect 24006 87998 25438 88062
rect 25502 87998 27342 88062
rect 27406 87998 28838 88062
rect 28902 87998 30470 88062
rect 30534 87998 32374 88062
rect 32438 87998 33870 88062
rect 33934 87998 35910 88062
rect 35974 87998 37406 88062
rect 37470 87998 39038 88062
rect 39102 87998 40942 88062
rect 41006 87998 42438 88062
rect 42502 87998 43934 88062
rect 43998 87998 45838 88062
rect 45902 87998 47334 88062
rect 47398 87998 49102 88062
rect 49166 87998 50870 88062
rect 50934 87998 52502 88062
rect 52566 87998 54270 88062
rect 54334 87998 55902 88062
rect 55966 87998 57398 88062
rect 57462 87998 59302 88062
rect 59366 87998 60934 88062
rect 60998 87998 62566 88062
rect 62630 87998 64334 88062
rect 64398 87998 65966 88062
rect 66030 87998 67598 88062
rect 67662 87998 69366 88062
rect 69430 87998 70862 88062
rect 70926 87998 72630 88062
rect 72694 87998 74262 88062
rect 74326 87998 76030 88062
rect 76094 87998 77662 88062
rect 77726 87998 79430 88062
rect 79494 87998 81062 88062
rect 81126 87998 82558 88062
rect 82622 87998 84326 88062
rect 84390 87998 86094 88062
rect 86158 87998 87862 88062
rect 87926 87998 89766 88062
rect 89830 87998 89902 88062
rect 89966 87998 90038 88062
rect 90102 87998 90108 88062
rect 952 87992 90108 87998
rect 1904 87654 2252 87660
rect 1904 87590 2182 87654
rect 2246 87590 2252 87654
rect 1904 87524 2252 87590
rect 1904 87468 2054 87524
rect 2110 87468 2252 87524
rect 1904 87312 2252 87468
rect 3672 87654 3884 87660
rect 3672 87590 3814 87654
rect 3878 87590 3884 87654
rect 3672 87524 3884 87590
rect 3672 87468 3734 87524
rect 3790 87468 3884 87524
rect 3672 87312 3884 87468
rect 5304 87654 5516 87660
rect 5304 87590 5310 87654
rect 5374 87590 5516 87654
rect 5304 87524 5516 87590
rect 5304 87468 5414 87524
rect 5470 87468 5516 87524
rect 5304 87312 5516 87468
rect 7072 87654 7284 87660
rect 7072 87590 7078 87654
rect 7142 87590 7284 87654
rect 7072 87524 7284 87590
rect 7072 87468 7094 87524
rect 7150 87468 7284 87524
rect 7072 87312 7284 87468
rect 8704 87654 8916 87660
rect 8704 87590 8846 87654
rect 8910 87590 8916 87654
rect 8704 87524 8916 87590
rect 8704 87468 8774 87524
rect 8830 87468 8916 87524
rect 8704 87312 8916 87468
rect 10336 87654 10548 87660
rect 10336 87590 10342 87654
rect 10406 87590 10548 87654
rect 10336 87524 10548 87590
rect 10336 87468 10454 87524
rect 10510 87468 10548 87524
rect 10336 87312 10548 87468
rect 12104 87654 12316 87660
rect 12104 87590 12110 87654
rect 12174 87590 12316 87654
rect 12104 87524 12316 87590
rect 12104 87468 12134 87524
rect 12190 87468 12316 87524
rect 12104 87312 12316 87468
rect 13736 87654 13948 87660
rect 13736 87590 13878 87654
rect 13942 87590 13948 87654
rect 13736 87524 13948 87590
rect 13736 87468 13814 87524
rect 13870 87468 13948 87524
rect 13736 87312 13948 87468
rect 15368 87654 15580 87660
rect 15368 87590 15374 87654
rect 15438 87590 15580 87654
rect 15368 87524 15580 87590
rect 15368 87468 15494 87524
rect 15550 87468 15580 87524
rect 15368 87312 15580 87468
rect 17136 87654 17348 87660
rect 17136 87590 17278 87654
rect 17342 87590 17348 87654
rect 17136 87524 17348 87590
rect 17136 87468 17174 87524
rect 17230 87468 17348 87524
rect 17136 87312 17348 87468
rect 18768 87654 18980 87660
rect 18768 87590 18910 87654
rect 18974 87590 18980 87654
rect 18768 87524 18980 87590
rect 18768 87468 18854 87524
rect 18910 87468 18980 87524
rect 18768 87312 18980 87468
rect 20400 87654 20612 87660
rect 20400 87590 20542 87654
rect 20606 87590 20612 87654
rect 20400 87524 20612 87590
rect 20400 87468 20534 87524
rect 20590 87468 20612 87524
rect 20400 87312 20612 87468
rect 22168 87654 22380 87660
rect 22168 87590 22174 87654
rect 22238 87590 22380 87654
rect 22168 87524 22380 87590
rect 22168 87468 22214 87524
rect 22270 87468 22380 87524
rect 22168 87312 22380 87468
rect 23800 87654 24012 87660
rect 23800 87590 23942 87654
rect 24006 87590 24012 87654
rect 23800 87524 24012 87590
rect 23800 87468 23894 87524
rect 23950 87468 24012 87524
rect 23800 87312 24012 87468
rect 25432 87654 25780 87660
rect 25432 87590 25438 87654
rect 25502 87590 25780 87654
rect 25432 87524 25780 87590
rect 25432 87468 25574 87524
rect 25630 87468 25780 87524
rect 25432 87312 25780 87468
rect 27200 87654 27412 87660
rect 27200 87590 27342 87654
rect 27406 87590 27412 87654
rect 27200 87524 27412 87590
rect 27200 87468 27254 87524
rect 27310 87468 27412 87524
rect 27200 87312 27412 87468
rect 28832 87654 29044 87660
rect 28832 87590 28838 87654
rect 28902 87590 29044 87654
rect 28832 87524 29044 87590
rect 28832 87468 28934 87524
rect 28990 87468 29044 87524
rect 28832 87312 29044 87468
rect 30464 87654 30812 87660
rect 30464 87590 30470 87654
rect 30534 87590 30812 87654
rect 30464 87524 30812 87590
rect 30464 87468 30614 87524
rect 30670 87468 30812 87524
rect 30464 87312 30812 87468
rect 32232 87654 32444 87660
rect 32232 87590 32374 87654
rect 32438 87590 32444 87654
rect 32232 87524 32444 87590
rect 32232 87468 32294 87524
rect 32350 87468 32444 87524
rect 32232 87312 32444 87468
rect 33864 87654 34076 87660
rect 33864 87590 33870 87654
rect 33934 87590 34076 87654
rect 33864 87524 34076 87590
rect 33864 87468 33974 87524
rect 34030 87468 34076 87524
rect 33864 87312 34076 87468
rect 35632 87654 35980 87660
rect 35632 87590 35910 87654
rect 35974 87590 35980 87654
rect 35632 87584 35980 87590
rect 37264 87654 37476 87660
rect 37264 87590 37406 87654
rect 37470 87590 37476 87654
rect 35632 87524 35844 87584
rect 35632 87468 35654 87524
rect 35710 87468 35844 87524
rect 35632 87312 35844 87468
rect 37264 87524 37476 87590
rect 37264 87468 37334 87524
rect 37390 87468 37476 87524
rect 37264 87312 37476 87468
rect 38896 87654 39108 87660
rect 38896 87590 39038 87654
rect 39102 87590 39108 87654
rect 38896 87524 39108 87590
rect 38896 87468 39014 87524
rect 39070 87468 39108 87524
rect 38896 87312 39108 87468
rect 40664 87654 41012 87660
rect 40664 87590 40942 87654
rect 41006 87590 41012 87654
rect 40664 87584 41012 87590
rect 42296 87654 42508 87660
rect 42296 87590 42438 87654
rect 42502 87590 42508 87654
rect 40664 87524 40876 87584
rect 40664 87468 40694 87524
rect 40750 87468 40876 87524
rect 40664 87312 40876 87468
rect 42296 87524 42508 87590
rect 42296 87468 42374 87524
rect 42430 87468 42508 87524
rect 42296 87312 42508 87468
rect 43928 87654 44140 87660
rect 43928 87590 43934 87654
rect 43998 87590 44140 87654
rect 43928 87524 44140 87590
rect 43928 87468 44054 87524
rect 44110 87468 44140 87524
rect 43928 87312 44140 87468
rect 45696 87654 45908 87660
rect 45696 87590 45838 87654
rect 45902 87590 45908 87654
rect 45696 87524 45908 87590
rect 45696 87468 45734 87524
rect 45790 87468 45908 87524
rect 45696 87312 45908 87468
rect 47328 87654 47540 87660
rect 47328 87590 47334 87654
rect 47398 87590 47540 87654
rect 47328 87524 47540 87590
rect 47328 87468 47414 87524
rect 47470 87468 47540 87524
rect 47328 87312 47540 87468
rect 48960 87654 49172 87660
rect 48960 87590 49102 87654
rect 49166 87590 49172 87654
rect 48960 87524 49172 87590
rect 48960 87468 49094 87524
rect 49150 87468 49172 87524
rect 48960 87312 49172 87468
rect 50728 87654 50940 87660
rect 50728 87590 50870 87654
rect 50934 87590 50940 87654
rect 50728 87524 50940 87590
rect 50728 87468 50774 87524
rect 50830 87468 50940 87524
rect 50728 87312 50940 87468
rect 52360 87654 52572 87660
rect 52360 87590 52502 87654
rect 52566 87590 52572 87654
rect 52360 87524 52572 87590
rect 52360 87468 52454 87524
rect 52510 87468 52572 87524
rect 52360 87312 52572 87468
rect 53992 87654 54340 87660
rect 53992 87590 54270 87654
rect 54334 87590 54340 87654
rect 53992 87524 54340 87590
rect 53992 87468 54134 87524
rect 54190 87468 54340 87524
rect 53992 87312 54340 87468
rect 55760 87654 55972 87660
rect 55760 87590 55902 87654
rect 55966 87590 55972 87654
rect 55760 87524 55972 87590
rect 55760 87468 55814 87524
rect 55870 87468 55972 87524
rect 55760 87312 55972 87468
rect 57392 87654 57604 87660
rect 57392 87590 57398 87654
rect 57462 87590 57604 87654
rect 57392 87524 57604 87590
rect 57392 87468 57494 87524
rect 57550 87468 57604 87524
rect 57392 87312 57604 87468
rect 59024 87654 59372 87660
rect 59024 87590 59302 87654
rect 59366 87590 59372 87654
rect 59024 87524 59372 87590
rect 59024 87468 59174 87524
rect 59230 87468 59372 87524
rect 59024 87312 59372 87468
rect 60792 87654 61004 87660
rect 60792 87590 60934 87654
rect 60998 87590 61004 87654
rect 60792 87524 61004 87590
rect 60792 87468 60854 87524
rect 60910 87468 61004 87524
rect 60792 87312 61004 87468
rect 62424 87654 62636 87660
rect 62424 87590 62566 87654
rect 62630 87590 62636 87654
rect 62424 87524 62636 87590
rect 62424 87468 62534 87524
rect 62590 87468 62636 87524
rect 62424 87312 62636 87468
rect 64192 87654 64404 87660
rect 64192 87590 64334 87654
rect 64398 87590 64404 87654
rect 64192 87524 64404 87590
rect 64192 87468 64214 87524
rect 64270 87468 64404 87524
rect 64192 87312 64404 87468
rect 65824 87654 66036 87660
rect 65824 87590 65966 87654
rect 66030 87590 66036 87654
rect 65824 87524 66036 87590
rect 65824 87468 65894 87524
rect 65950 87468 66036 87524
rect 65824 87312 66036 87468
rect 67456 87654 67668 87660
rect 67456 87590 67598 87654
rect 67662 87590 67668 87654
rect 67456 87524 67668 87590
rect 67456 87468 67574 87524
rect 67630 87468 67668 87524
rect 67456 87312 67668 87468
rect 69224 87654 69436 87660
rect 69224 87590 69366 87654
rect 69430 87590 69436 87654
rect 69224 87524 69436 87590
rect 69224 87468 69254 87524
rect 69310 87468 69436 87524
rect 69224 87312 69436 87468
rect 70856 87654 71068 87660
rect 70856 87590 70862 87654
rect 70926 87590 71068 87654
rect 70856 87524 71068 87590
rect 70856 87468 70934 87524
rect 70990 87468 71068 87524
rect 70856 87312 71068 87468
rect 72488 87654 72700 87660
rect 72488 87590 72630 87654
rect 72694 87590 72700 87654
rect 72488 87524 72700 87590
rect 72488 87468 72614 87524
rect 72670 87468 72700 87524
rect 72488 87312 72700 87468
rect 74256 87654 74468 87660
rect 74256 87590 74262 87654
rect 74326 87590 74468 87654
rect 74256 87524 74468 87590
rect 74256 87468 74294 87524
rect 74350 87468 74468 87524
rect 74256 87312 74468 87468
rect 75888 87654 76100 87660
rect 75888 87590 76030 87654
rect 76094 87590 76100 87654
rect 75888 87524 76100 87590
rect 75888 87468 75974 87524
rect 76030 87468 76100 87524
rect 75888 87388 76100 87468
rect 77520 87654 77732 87660
rect 77520 87590 77662 87654
rect 77726 87590 77732 87654
rect 77520 87524 77732 87590
rect 77520 87468 77654 87524
rect 77710 87468 77732 87524
rect 75888 87382 76372 87388
rect 75888 87318 76302 87382
rect 76366 87318 76372 87382
rect 75888 87312 76372 87318
rect 77520 87312 77732 87468
rect 79288 87654 79500 87660
rect 79288 87590 79430 87654
rect 79494 87590 79500 87654
rect 79288 87524 79500 87590
rect 79288 87468 79334 87524
rect 79390 87468 79500 87524
rect 79288 87312 79500 87468
rect 80920 87654 81132 87660
rect 80920 87590 81062 87654
rect 81126 87590 81132 87654
rect 80920 87524 81132 87590
rect 80920 87468 81014 87524
rect 81070 87468 81132 87524
rect 80920 87312 81132 87468
rect 82552 87654 82900 87660
rect 82552 87590 82558 87654
rect 82622 87590 82900 87654
rect 82552 87524 82900 87590
rect 82552 87468 82694 87524
rect 82750 87468 82900 87524
rect 82552 87312 82900 87468
rect 84320 87654 84532 87660
rect 84320 87590 84326 87654
rect 84390 87590 84532 87654
rect 84320 87524 84532 87590
rect 84320 87468 84374 87524
rect 84430 87468 84532 87524
rect 84320 87312 84532 87468
rect 85952 87654 86164 87660
rect 85952 87590 86094 87654
rect 86158 87590 86164 87654
rect 85952 87524 86164 87590
rect 85952 87468 86054 87524
rect 86110 87468 86164 87524
rect 85952 87312 86164 87468
rect 87584 87654 87932 87660
rect 87584 87590 87862 87654
rect 87926 87590 87932 87654
rect 87584 87524 87932 87590
rect 87584 87468 87734 87524
rect 87790 87468 87932 87524
rect 87584 87312 87932 87468
rect 73984 86974 75420 86980
rect 73984 86910 73990 86974
rect 74054 86910 75420 86974
rect 73984 86904 75420 86910
rect 73984 86844 74196 86904
rect 75208 86844 75420 86904
rect 76296 86844 76508 86980
rect 73984 86838 74332 86844
rect 73984 86774 74262 86838
rect 74326 86774 74332 86838
rect 73984 86768 74332 86774
rect 75208 86768 76508 86844
rect 79255 86546 79321 86549
rect 75284 86544 79321 86546
rect 75284 86488 79260 86544
rect 79316 86488 79321 86544
rect 75284 86486 79321 86488
rect 79255 86483 79321 86486
rect 74481 86300 74579 86309
rect 75649 86300 75747 86309
rect 76817 86300 76915 86309
rect 74392 86294 74604 86300
rect 74392 86288 74534 86294
rect 74392 86232 74502 86288
rect 74392 86230 74534 86232
rect 74598 86230 74604 86294
rect 1632 86132 1844 86164
rect 1632 86076 1718 86132
rect 1774 86076 1844 86132
rect 74392 86088 74604 86230
rect 75616 86294 75828 86300
rect 75616 86230 75622 86294
rect 75686 86288 75828 86294
rect 75726 86232 75828 86288
rect 75686 86230 75828 86232
rect 75616 86088 75828 86230
rect 76704 86294 76916 86300
rect 76704 86230 76710 86294
rect 76774 86288 76916 86294
rect 76774 86232 76838 86288
rect 76894 86232 76916 86288
rect 76774 86230 76916 86232
rect 76704 86088 76916 86230
rect 89080 86132 89428 86164
rect 1632 86028 1844 86076
rect 1224 86022 1844 86028
rect 1224 85958 1230 86022
rect 1294 85958 1844 86022
rect 1224 85952 1844 85958
rect 89080 86076 89216 86132
rect 89272 86076 89428 86132
rect 89080 86028 89428 86076
rect 89080 86022 89836 86028
rect 89080 85958 89766 86022
rect 89830 85958 89836 86022
rect 89080 85952 89836 85958
rect 73984 85348 74196 85484
rect 75208 85478 76508 85484
rect 75208 85414 76302 85478
rect 76366 85414 76508 85478
rect 75208 85408 76508 85414
rect 75208 85348 75420 85408
rect 73984 85342 75420 85348
rect 73984 85278 74126 85342
rect 74190 85278 75420 85342
rect 73984 85272 75420 85278
rect 76296 85272 76508 85408
rect 72760 84668 72972 84804
rect 74120 84798 74332 84804
rect 74120 84734 74262 84798
rect 74326 84734 74332 84798
rect 74120 84668 74332 84734
rect 72760 84662 74430 84668
rect 72760 84598 74398 84662
rect 74462 84598 74468 84662
rect 72760 84592 74430 84598
rect 1632 84452 1844 84532
rect 1632 84396 1718 84452
rect 1774 84396 1844 84452
rect 1224 84390 1844 84396
rect 1224 84326 1230 84390
rect 1294 84326 1844 84390
rect 1224 84320 1844 84326
rect 89080 84452 89428 84532
rect 89080 84396 89216 84452
rect 89272 84396 89428 84452
rect 89080 84390 89836 84396
rect 89080 84326 89766 84390
rect 89830 84326 89836 84390
rect 89080 84320 89836 84326
rect 72760 83172 72972 83308
rect 74120 83302 74332 83308
rect 74120 83238 74126 83302
rect 74190 83238 74332 83302
rect 74120 83172 74332 83238
rect 72760 83166 74332 83172
rect 72760 83102 74262 83166
rect 74326 83102 74332 83166
rect 72760 83096 74332 83102
rect 1632 82772 1844 82900
rect 1632 82764 1718 82772
rect 1224 82758 1718 82764
rect 1224 82694 1230 82758
rect 1294 82716 1718 82758
rect 1774 82716 1844 82772
rect 1294 82694 1844 82716
rect 1224 82688 1844 82694
rect 89080 82772 89428 82900
rect 89080 82716 89216 82772
rect 89272 82764 89428 82772
rect 89272 82758 89836 82764
rect 89272 82716 89766 82758
rect 89080 82694 89766 82716
rect 89830 82694 89836 82758
rect 89080 82688 89836 82694
rect 72760 81812 72972 81948
rect 74120 81942 74468 81948
rect 74120 81878 74398 81942
rect 74462 81878 74468 81942
rect 74120 81872 74468 81878
rect 74120 81812 74332 81872
rect 72760 81806 74332 81812
rect 72760 81742 74126 81806
rect 74190 81742 74332 81806
rect 72760 81736 74332 81742
rect 1632 81092 1844 81132
rect 1632 81036 1718 81092
rect 1774 81036 1844 81092
rect 1632 80996 1844 81036
rect 1224 80990 1844 80996
rect 1224 80926 1230 80990
rect 1294 80926 1844 80990
rect 1224 80920 1844 80926
rect 89080 81092 89428 81132
rect 89080 81036 89216 81092
rect 89272 81036 89428 81092
rect 89080 80996 89428 81036
rect 89080 80990 89836 80996
rect 89080 80926 89766 80990
rect 89830 80926 89836 80990
rect 89080 80920 89836 80926
rect 72760 80316 72972 80452
rect 74120 80446 74332 80452
rect 74120 80382 74262 80446
rect 74326 80382 74332 80446
rect 74120 80316 74332 80382
rect 72760 80310 74332 80316
rect 72760 80246 74262 80310
rect 74326 80246 74332 80310
rect 72760 80240 74332 80246
rect 79288 80174 79636 80316
rect 79288 80110 79294 80174
rect 79358 80110 79636 80174
rect 79288 80104 79636 80110
rect 88400 80180 88612 80316
rect 88400 80174 90516 80180
rect 88400 80110 90446 80174
rect 90510 80110 90516 80174
rect 88400 80104 90516 80110
rect 88128 79696 91060 79772
rect 85000 79530 85212 79636
rect 1632 79412 1844 79500
rect 85000 79474 85119 79530
rect 85175 79500 85212 79530
rect 88128 79635 88340 79696
rect 88128 79579 88256 79635
rect 88312 79579 88340 79635
rect 85175 79494 88068 79500
rect 85175 79474 87998 79494
rect 85000 79430 87998 79474
rect 88062 79430 88068 79494
rect 85000 79424 88068 79430
rect 88128 79424 88340 79579
rect 1632 79364 1718 79412
rect 1224 79358 1718 79364
rect 1224 79294 1230 79358
rect 1294 79356 1718 79358
rect 1774 79356 1844 79412
rect 1294 79294 1844 79356
rect 1224 79288 1844 79294
rect 89080 79412 89428 79500
rect 89080 79358 89216 79412
rect 89080 79294 89086 79358
rect 89150 79356 89216 79358
rect 89272 79364 89428 79412
rect 89272 79358 89836 79364
rect 89272 79356 89766 79358
rect 89150 79294 89766 79356
rect 89830 79294 89836 79358
rect 89080 79288 89836 79294
rect 88030 79222 91060 79228
rect 87992 79158 87998 79222
rect 88062 79158 91060 79222
rect 88030 79152 91060 79158
rect 72760 78956 72972 79092
rect 74120 79086 74332 79092
rect 74120 79022 74126 79086
rect 74190 79022 74332 79086
rect 74120 78956 74332 79022
rect 72760 78950 74332 78956
rect 72760 78886 74126 78950
rect 74190 78886 74332 78950
rect 72760 78880 74332 78886
rect 79288 78678 79636 78820
rect 79288 78614 79566 78678
rect 79630 78614 79636 78678
rect 79288 78608 79636 78614
rect 88400 78814 89156 78820
rect 88400 78750 89086 78814
rect 89150 78750 89156 78814
rect 88400 78744 89156 78750
rect 88400 78608 88612 78744
rect 25568 77998 25780 78004
rect 25568 77934 25574 77998
rect 25638 77934 25780 77998
rect 25976 77950 26052 78004
rect 25568 77910 25780 77934
rect 1632 77732 1844 77868
rect 25568 77854 25626 77910
rect 25682 77854 25780 77910
rect 25568 77792 25780 77854
rect 25859 77862 26052 77950
rect 25859 77852 25982 77862
rect 25976 77798 25982 77852
rect 26046 77798 26052 77862
rect 25976 77792 26052 77798
rect 30464 77998 30676 78004
rect 30464 77934 30606 77998
rect 30670 77934 30676 77998
rect 30872 77950 31084 78004
rect 30464 77931 30676 77934
rect 30464 77910 30695 77931
rect 30464 77854 30618 77910
rect 30674 77854 30695 77910
rect 30464 77833 30695 77854
rect 30851 77862 31084 77950
rect 30851 77852 30878 77862
rect 30464 77792 30676 77833
rect 30872 77798 30878 77852
rect 30942 77798 31084 77862
rect 30872 77792 31084 77798
rect 35496 77998 35708 78004
rect 35496 77934 35638 77998
rect 35702 77934 35708 77998
rect 35904 77950 35980 78004
rect 35496 77910 35708 77934
rect 35496 77854 35610 77910
rect 35666 77854 35708 77910
rect 35496 77792 35708 77854
rect 35843 77862 35980 77950
rect 35843 77852 35910 77862
rect 35904 77798 35910 77852
rect 35974 77798 35980 77862
rect 35904 77792 35980 77798
rect 40528 77998 40740 78004
rect 40528 77934 40670 77998
rect 40734 77934 40740 77998
rect 40936 77950 41012 78004
rect 40528 77910 40740 77934
rect 40528 77854 40602 77910
rect 40658 77854 40740 77910
rect 40528 77792 40740 77854
rect 40835 77868 41012 77950
rect 45560 77998 45636 78004
rect 45560 77934 45566 77998
rect 45630 77934 45636 77998
rect 45832 77950 46044 78004
rect 45560 77931 45636 77934
rect 45560 77910 45671 77931
rect 40835 77862 41148 77868
rect 40835 77852 41078 77862
rect 40936 77798 41078 77852
rect 41142 77798 41148 77862
rect 40936 77792 41148 77798
rect 45560 77854 45594 77910
rect 45650 77854 45671 77910
rect 45560 77833 45671 77854
rect 45827 77862 46044 77950
rect 45827 77852 45974 77862
rect 45560 77792 45636 77833
rect 45832 77798 45974 77852
rect 46038 77798 46044 77862
rect 45832 77792 46044 77798
rect 50456 77998 50668 78004
rect 50456 77934 50462 77998
rect 50526 77934 50668 77998
rect 50864 77950 50940 78004
rect 50456 77910 50668 77934
rect 50456 77854 50586 77910
rect 50642 77854 50668 77910
rect 50456 77792 50668 77854
rect 50819 77862 50940 77950
rect 50819 77852 50870 77862
rect 50864 77798 50870 77852
rect 50934 77798 50940 77862
rect 50864 77792 50940 77798
rect 55488 77998 55700 78004
rect 55488 77934 55630 77998
rect 55694 77934 55700 77998
rect 55896 77950 55972 78004
rect 55488 77910 55700 77934
rect 55488 77854 55578 77910
rect 55634 77854 55700 77910
rect 55488 77792 55700 77854
rect 55811 77868 55972 77950
rect 60520 77998 60732 78004
rect 60520 77934 60662 77998
rect 60726 77934 60732 77998
rect 60928 77950 61004 78004
rect 60520 77910 60732 77934
rect 55811 77862 56108 77868
rect 55811 77852 56038 77862
rect 55896 77798 56038 77852
rect 56102 77798 56108 77862
rect 55896 77792 56108 77798
rect 60520 77854 60570 77910
rect 60626 77854 60732 77910
rect 60520 77792 60732 77854
rect 60803 77862 61004 77950
rect 60803 77852 60934 77862
rect 60928 77798 60934 77852
rect 60998 77798 61004 77862
rect 60928 77792 61004 77798
rect 89080 77732 89428 77868
rect 1224 77726 1718 77732
rect 1224 77662 1230 77726
rect 1294 77676 1718 77726
rect 1774 77676 1844 77732
rect 1294 77662 1844 77676
rect 1224 77656 1844 77662
rect 1632 77520 1844 77656
rect 25840 77590 26052 77732
rect 25840 77526 25846 77590
rect 25910 77526 26052 77590
rect 25840 77520 26052 77526
rect 30736 77590 31084 77732
rect 30736 77526 30742 77590
rect 30806 77526 31084 77590
rect 30736 77520 31084 77526
rect 35768 77590 35980 77732
rect 35768 77526 35774 77590
rect 35838 77526 35980 77590
rect 35768 77520 35980 77526
rect 40800 77590 41012 77732
rect 40800 77526 40942 77590
rect 41006 77526 41012 77590
rect 40800 77520 41012 77526
rect 45696 77590 46044 77732
rect 45696 77526 45838 77590
rect 45902 77526 46044 77590
rect 45696 77520 46044 77526
rect 50728 77590 50940 77732
rect 50728 77526 50734 77590
rect 50798 77526 50940 77590
rect 50728 77520 50940 77526
rect 55760 77590 55972 77732
rect 55760 77526 55902 77590
rect 55966 77526 55972 77590
rect 55760 77520 55972 77526
rect 60792 77590 61004 77732
rect 60792 77526 60934 77590
rect 60998 77526 61004 77590
rect 60792 77520 61004 77526
rect 72760 77596 72972 77732
rect 74120 77726 74332 77732
rect 74120 77662 74262 77726
rect 74326 77662 74332 77726
rect 74120 77596 74332 77662
rect 72760 77590 74332 77596
rect 72760 77526 72902 77590
rect 72966 77526 74332 77590
rect 72760 77520 74332 77526
rect 89080 77676 89216 77732
rect 89272 77676 89428 77732
rect 89080 77596 89428 77676
rect 89080 77590 89836 77596
rect 89080 77526 89766 77590
rect 89830 77526 89836 77590
rect 89080 77520 89836 77526
rect 79288 77454 79636 77460
rect 79288 77390 79294 77454
rect 79358 77390 79636 77454
rect 79288 77318 79636 77390
rect 79288 77254 79294 77318
rect 79358 77254 79430 77318
rect 79494 77254 79636 77318
rect 79288 77248 79636 77254
rect 25840 76910 26052 76916
rect 25840 76846 25846 76910
rect 25910 76846 26052 76910
rect 25840 76638 26052 76846
rect 30736 76910 30948 76916
rect 30736 76846 30742 76910
rect 30806 76846 30948 76910
rect 30736 76644 30948 76846
rect 30366 76638 30948 76644
rect 25840 76574 25846 76638
rect 25910 76574 26052 76638
rect 30328 76574 30334 76638
rect 30398 76574 30948 76638
rect 25840 76568 26052 76574
rect 30366 76568 30948 76574
rect 35768 76910 35980 76916
rect 35768 76846 35774 76910
rect 35838 76846 35980 76910
rect 35768 76644 35980 76846
rect 40800 76910 41012 76916
rect 40800 76846 40942 76910
rect 41006 76846 41012 76910
rect 35768 76638 36932 76644
rect 35768 76574 36862 76638
rect 36926 76574 36932 76638
rect 35768 76568 36932 76574
rect 40800 76638 41012 76846
rect 40800 76574 40806 76638
rect 40870 76574 41012 76638
rect 40800 76568 41012 76574
rect 45696 76910 46044 76916
rect 45696 76846 45838 76910
rect 45902 76846 46044 76910
rect 45696 76638 46044 76846
rect 45696 76574 45702 76638
rect 45766 76574 46044 76638
rect 45696 76568 46044 76574
rect 50728 76910 50940 76916
rect 50728 76846 50734 76910
rect 50798 76846 50940 76910
rect 50728 76638 50940 76846
rect 55760 76910 55972 76916
rect 55760 76846 55902 76910
rect 55966 76846 55972 76910
rect 55760 76644 55972 76846
rect 55390 76638 55972 76644
rect 50728 76574 50734 76638
rect 50798 76574 50940 76638
rect 55352 76574 55358 76638
rect 55422 76574 55972 76638
rect 50728 76568 50940 76574
rect 55390 76568 55972 76574
rect 60656 76910 61004 76916
rect 60656 76846 60934 76910
rect 60998 76846 61004 76910
rect 60656 76644 61004 76846
rect 60656 76638 61548 76644
rect 60656 76574 61478 76638
rect 61542 76574 61548 76638
rect 60656 76568 61548 76574
rect 72760 76230 79364 76236
rect 72760 76166 74126 76230
rect 74190 76166 79294 76230
rect 79358 76166 79364 76230
rect 72760 76160 79364 76166
rect 72760 76100 72972 76160
rect 1632 76052 1844 76100
rect 1632 75996 1718 76052
rect 1774 75996 1844 76052
rect 25840 76094 26188 76100
rect 25840 76030 25982 76094
rect 26046 76030 26118 76094
rect 26182 76030 26188 76094
rect 25840 76024 26188 76030
rect 30872 76094 31084 76100
rect 30872 76030 30878 76094
rect 30942 76030 31014 76094
rect 31078 76030 31084 76094
rect 30872 76024 31084 76030
rect 35904 76094 36116 76100
rect 35904 76030 35910 76094
rect 35974 76030 36046 76094
rect 36110 76030 36116 76094
rect 35904 76024 36116 76030
rect 40800 76094 41110 76100
rect 45832 76094 46180 76100
rect 40800 76030 40942 76094
rect 41006 76030 41078 76094
rect 41142 76030 41148 76094
rect 45832 76030 45974 76094
rect 46038 76030 46110 76094
rect 46174 76030 46180 76094
rect 40800 76024 41110 76030
rect 45832 76024 46180 76030
rect 50864 76094 51076 76100
rect 50864 76030 50870 76094
rect 50934 76030 51006 76094
rect 51070 76030 51076 76094
rect 50864 76024 51076 76030
rect 55760 76094 56244 76100
rect 55760 76030 56038 76094
rect 56102 76030 56174 76094
rect 56238 76030 56244 76094
rect 55760 76024 56244 76030
rect 60792 76094 61004 76100
rect 60792 76030 60798 76094
rect 60862 76030 60934 76094
rect 60998 76030 61004 76094
rect 60792 76024 61004 76030
rect 72624 76094 72972 76100
rect 72624 76030 72630 76094
rect 72694 76030 72972 76094
rect 72624 76024 72972 76030
rect 74120 76024 74332 76160
rect 79288 76094 79636 76100
rect 79288 76030 79566 76094
rect 79630 76030 79636 76094
rect 1632 75964 1844 75996
rect 1224 75958 1844 75964
rect 1224 75894 1230 75958
rect 1294 75894 1844 75958
rect 25929 75918 26027 76024
rect 30921 75918 31019 76024
rect 35913 75918 36011 76024
rect 40905 75918 41003 76024
rect 45897 75918 45995 76024
rect 50889 75918 50987 76024
rect 55881 75918 55979 76024
rect 60873 75918 60971 76024
rect 1224 75888 1844 75894
rect 79288 75822 79636 76030
rect 89080 76052 89428 76100
rect 89080 75996 89216 76052
rect 89272 75996 89428 76052
rect 89080 75964 89428 75996
rect 89080 75958 89836 75964
rect 89080 75894 89766 75958
rect 89830 75894 89836 75958
rect 89080 75888 89836 75894
rect 79288 75758 79294 75822
rect 79358 75758 79566 75822
rect 79630 75758 79636 75822
rect 79288 75752 79636 75758
rect 67128 75254 67194 75259
rect 67128 75198 67133 75254
rect 67189 75253 67194 75254
rect 67189 75234 79405 75253
rect 67189 75198 79344 75234
rect 67128 75193 79344 75198
rect 79339 75178 79344 75193
rect 79400 75178 79405 75234
rect 79339 75173 79405 75178
rect 72760 74870 79364 74876
rect 72760 74806 72902 74870
rect 72966 74806 79294 74870
rect 79358 74806 79364 74870
rect 72760 74800 79364 74806
rect 72760 74734 72972 74800
rect 72760 74670 72766 74734
rect 72830 74670 72972 74734
rect 72760 74664 72972 74670
rect 74120 74664 74332 74800
rect 79288 74598 79636 74604
rect 79288 74534 79430 74598
rect 79494 74534 79636 74598
rect 1632 74372 1844 74468
rect 79288 74462 79636 74534
rect 79288 74398 79294 74462
rect 79358 74398 79636 74462
rect 79288 74392 79636 74398
rect 86904 74528 87932 74604
rect 86904 74392 87116 74528
rect 87720 74468 87932 74528
rect 87720 74462 89836 74468
rect 87720 74398 89766 74462
rect 89830 74398 89836 74462
rect 87720 74392 89836 74398
rect 1632 74332 1718 74372
rect 1224 74326 1718 74332
rect 1224 74262 1230 74326
rect 1294 74316 1718 74326
rect 1774 74316 1844 74372
rect 1294 74262 1844 74316
rect 1224 74256 1844 74262
rect 89080 74372 89428 74392
rect 89080 74316 89216 74372
rect 89272 74316 89428 74372
rect 89080 74256 89428 74316
rect 67252 73838 67318 73841
rect 79339 73838 79405 73841
rect 67252 73836 79405 73838
rect 67252 73780 67257 73836
rect 67313 73780 79344 73836
rect 79400 73780 79405 73836
rect 67252 73778 79405 73780
rect 67252 73775 67318 73778
rect 79339 73775 79405 73778
rect 25976 73646 26324 73652
rect 25976 73582 26118 73646
rect 26182 73582 26324 73646
rect 25976 73516 26324 73582
rect 27336 73516 27548 73652
rect 28560 73516 28772 73652
rect 25976 73440 28772 73516
rect 25976 73374 26324 73440
rect 25976 73310 25982 73374
rect 26046 73310 26324 73374
rect 25976 73304 26324 73310
rect 27336 73304 27548 73440
rect 28560 73380 28772 73440
rect 29784 73646 31220 73652
rect 29784 73582 31014 73646
rect 31078 73582 31220 73646
rect 29784 73576 31220 73582
rect 29784 73380 29996 73576
rect 28560 73304 29996 73380
rect 31008 73380 31220 73576
rect 32232 73576 33804 73652
rect 32232 73380 32444 73576
rect 31008 73304 32444 73380
rect 33456 73380 33804 73576
rect 34816 73516 35028 73652
rect 36040 73646 36252 73652
rect 36040 73582 36046 73646
rect 36110 73582 36252 73646
rect 36040 73516 36252 73582
rect 37264 73516 37476 73652
rect 34816 73440 37476 73516
rect 34816 73380 35028 73440
rect 33456 73304 35028 73380
rect 36040 73304 36252 73440
rect 37264 73380 37476 73440
rect 38488 73646 42508 73652
rect 38488 73582 41078 73646
rect 41142 73582 42508 73646
rect 38488 73576 42508 73582
rect 38488 73380 38700 73576
rect 37264 73304 38700 73380
rect 39712 73304 40060 73576
rect 41072 73304 41284 73576
rect 42296 73380 42508 73576
rect 43520 73516 43732 73652
rect 44744 73516 44956 73652
rect 45968 73646 46180 73652
rect 45968 73582 46110 73646
rect 46174 73582 46180 73646
rect 45968 73516 46180 73582
rect 43520 73440 46180 73516
rect 43520 73380 43732 73440
rect 42296 73304 43732 73380
rect 44744 73304 44956 73440
rect 45968 73380 46180 73440
rect 47192 73516 47540 73652
rect 48552 73646 51212 73652
rect 48552 73582 51006 73646
rect 51070 73582 51212 73646
rect 48552 73576 51212 73582
rect 48552 73516 48764 73576
rect 47192 73440 48764 73516
rect 47192 73380 47540 73440
rect 45968 73304 47540 73380
rect 48552 73304 48764 73440
rect 49776 73304 49988 73576
rect 51000 73516 51212 73576
rect 52224 73516 52436 73652
rect 53448 73516 53660 73652
rect 54672 73516 55020 73652
rect 56032 73646 56244 73652
rect 56032 73582 56174 73646
rect 56238 73582 56244 73646
rect 56032 73516 56244 73582
rect 57256 73576 59916 73652
rect 57256 73516 57468 73576
rect 51000 73440 57468 73516
rect 51000 73304 51212 73440
rect 52224 73304 52436 73440
rect 53448 73304 53660 73440
rect 54672 73304 55020 73440
rect 56032 73304 56244 73440
rect 57256 73304 57468 73440
rect 58480 73304 58692 73576
rect 59704 73380 59916 73576
rect 60928 73646 61276 73652
rect 60928 73582 60934 73646
rect 60998 73582 61276 73646
rect 60928 73380 61276 73582
rect 62288 73516 62500 73652
rect 63512 73516 63724 73652
rect 64736 73516 64948 73652
rect 62288 73440 64948 73516
rect 72662 73510 72972 73516
rect 72624 73446 72630 73510
rect 72694 73446 72972 73510
rect 72662 73440 72972 73446
rect 62288 73380 62500 73440
rect 59704 73304 62500 73380
rect 63512 73304 63724 73440
rect 64736 73380 64948 73440
rect 72760 73380 72972 73440
rect 74120 73380 74332 73516
rect 64736 73374 66852 73380
rect 64736 73310 66782 73374
rect 66846 73310 66852 73374
rect 64736 73304 66852 73310
rect 72760 73304 74332 73380
rect 72760 73168 72972 73304
rect 74120 73238 74332 73304
rect 74120 73174 74126 73238
rect 74190 73174 74332 73238
rect 74120 73168 74332 73174
rect 79288 73238 79636 73244
rect 79288 73174 79566 73238
rect 79630 73174 79636 73238
rect 79288 73032 79636 73174
rect 86904 73108 87116 73244
rect 87720 73238 90516 73244
rect 87720 73174 90446 73238
rect 90510 73174 90516 73238
rect 87720 73168 90516 73174
rect 87720 73108 87932 73168
rect 86904 73032 87932 73108
rect 1632 72700 1844 72836
rect 88459 72723 88465 72725
rect 1224 72694 1844 72700
rect 1224 72630 1230 72694
rect 1294 72692 1844 72694
rect 1294 72636 1718 72692
rect 1774 72636 1844 72692
rect 72344 72663 72404 72723
rect 79204 72663 88465 72723
rect 88459 72661 88465 72663
rect 88529 72661 88535 72725
rect 89080 72692 89428 72836
rect 1294 72630 1844 72636
rect 1224 72624 1844 72630
rect 1632 72488 1844 72624
rect 89080 72636 89216 72692
rect 89272 72636 89428 72692
rect 89080 72564 89428 72636
rect 89080 72558 89836 72564
rect 89080 72494 89086 72558
rect 89150 72494 89766 72558
rect 89830 72494 89836 72558
rect 89080 72488 89836 72494
rect 71113 72424 71179 72427
rect 79339 72424 79405 72427
rect 71113 72422 79405 72424
rect 71113 72366 71118 72422
rect 71174 72366 79344 72422
rect 79400 72366 79405 72422
rect 71113 72364 79405 72366
rect 71113 72361 71179 72364
rect 79339 72361 79405 72364
rect 25568 72014 25916 72020
rect 25568 71950 25846 72014
rect 25910 71950 25916 72014
rect 25568 71944 25916 71950
rect 25568 71878 25780 71944
rect 25568 71814 25574 71878
rect 25638 71814 25780 71878
rect 25568 71808 25780 71814
rect 26520 71884 26732 72020
rect 26792 71884 27140 72020
rect 27744 71944 28364 72020
rect 26520 71878 27684 71884
rect 26520 71814 26798 71878
rect 26862 71814 27614 71878
rect 27678 71814 27684 71878
rect 26520 71808 27684 71814
rect 27744 71878 27956 71944
rect 27744 71814 27750 71878
rect 27814 71814 27956 71878
rect 27744 71808 27956 71814
rect 28152 71808 28364 71944
rect 28968 71884 29180 72020
rect 29376 71884 29588 72020
rect 28968 71878 29588 71884
rect 28968 71814 28974 71878
rect 29038 71814 29518 71878
rect 29582 71814 29588 71878
rect 28968 71808 29588 71814
rect 30192 72014 30812 72020
rect 30192 71950 30334 72014
rect 30398 71950 30812 72014
rect 30192 71944 30812 71950
rect 30192 71808 30404 71944
rect 30600 71878 30812 71944
rect 30600 71814 30742 71878
rect 30806 71814 30812 71878
rect 30600 71808 30812 71814
rect 31416 71884 31628 72020
rect 31824 71884 32036 72020
rect 32640 71944 33260 72020
rect 32640 71884 32988 71944
rect 31416 71878 32036 71884
rect 32542 71878 32988 71884
rect 31416 71814 31422 71878
rect 31486 71814 31966 71878
rect 32030 71814 32036 71878
rect 32504 71814 32510 71878
rect 32574 71814 32988 71878
rect 31416 71808 32036 71814
rect 32542 71808 32988 71814
rect 33048 71878 33260 71944
rect 33048 71814 33054 71878
rect 33118 71814 33260 71878
rect 33048 71808 33260 71814
rect 34000 71944 34620 72020
rect 34000 71878 34212 71944
rect 34000 71814 34006 71878
rect 34070 71814 34212 71878
rect 34000 71808 34212 71814
rect 34272 71878 34620 71944
rect 34272 71814 34414 71878
rect 34478 71814 34620 71878
rect 34272 71808 34620 71814
rect 35224 71884 35436 72020
rect 35632 71884 35844 72020
rect 35224 71878 35844 71884
rect 35224 71814 35230 71878
rect 35294 71814 35774 71878
rect 35838 71814 35844 71878
rect 35224 71808 35844 71814
rect 36448 72014 37068 72020
rect 36448 71950 36862 72014
rect 36926 71950 37068 72014
rect 36448 71944 37068 71950
rect 36448 71878 36660 71944
rect 36448 71814 36454 71878
rect 36518 71814 36660 71878
rect 36448 71808 36660 71814
rect 36856 71878 37068 71944
rect 36856 71814 36998 71878
rect 37062 71814 37068 71878
rect 36856 71808 37068 71814
rect 37672 71884 37884 72020
rect 38080 71884 38292 72020
rect 37672 71878 38292 71884
rect 37672 71814 37678 71878
rect 37742 71814 38222 71878
rect 38286 71814 38292 71878
rect 37672 71808 38292 71814
rect 38896 71944 39516 72020
rect 38896 71808 39244 71944
rect 39304 71878 39516 71944
rect 39304 71814 39446 71878
rect 39510 71814 39516 71878
rect 39304 71808 39516 71814
rect 40256 72014 40876 72020
rect 40256 71950 40806 72014
rect 40870 71950 40876 72014
rect 40256 71944 40876 71950
rect 40256 71878 40468 71944
rect 40256 71814 40262 71878
rect 40326 71814 40468 71878
rect 40256 71808 40468 71814
rect 40528 71878 40876 71944
rect 40528 71814 40670 71878
rect 40734 71814 40876 71878
rect 40528 71808 40876 71814
rect 41480 71884 41692 72020
rect 41888 71884 42100 72020
rect 41480 71878 42100 71884
rect 41480 71814 41622 71878
rect 41686 71814 42100 71878
rect 41480 71808 42100 71814
rect 42704 71944 43324 72020
rect 42704 71878 42916 71944
rect 42704 71814 42710 71878
rect 42774 71814 42916 71878
rect 42704 71808 42916 71814
rect 43112 71878 43324 71944
rect 43112 71814 43254 71878
rect 43318 71814 43324 71878
rect 43112 71808 43324 71814
rect 43928 71884 44140 72020
rect 44336 71884 44548 72020
rect 43928 71878 44548 71884
rect 43928 71814 43934 71878
rect 43998 71814 44548 71878
rect 43928 71808 44548 71814
rect 45152 72014 45772 72020
rect 45152 71950 45702 72014
rect 45766 71950 45772 72014
rect 45152 71944 45772 71950
rect 45152 71878 45364 71944
rect 45152 71814 45158 71878
rect 45222 71814 45364 71878
rect 45152 71808 45364 71814
rect 45560 71878 45772 71944
rect 45560 71814 45702 71878
rect 45766 71814 45772 71878
rect 45560 71808 45772 71814
rect 46376 71884 46724 72020
rect 46784 71884 46996 72020
rect 46376 71878 46996 71884
rect 46376 71814 46926 71878
rect 46990 71814 46996 71878
rect 46376 71808 46996 71814
rect 47736 71884 47948 72020
rect 48008 71884 48356 72020
rect 47736 71878 48356 71884
rect 47736 71814 47742 71878
rect 47806 71814 48356 71878
rect 47736 71808 48356 71814
rect 48960 71944 49580 72020
rect 48960 71878 49172 71944
rect 48960 71814 48966 71878
rect 49030 71814 49172 71878
rect 48960 71808 49172 71814
rect 49368 71878 49580 71944
rect 49368 71814 49374 71878
rect 49438 71814 49580 71878
rect 49368 71808 49580 71814
rect 50184 71884 50396 72020
rect 50592 72014 50804 72020
rect 50592 71950 50734 72014
rect 50798 71950 50804 72014
rect 50592 71884 50804 71950
rect 50184 71878 50804 71884
rect 50184 71814 50190 71878
rect 50254 71814 50804 71878
rect 50184 71808 50804 71814
rect 51408 71944 52028 72020
rect 51408 71878 51620 71944
rect 51408 71814 51414 71878
rect 51478 71814 51620 71878
rect 51408 71808 51620 71814
rect 51816 71878 52028 71944
rect 51816 71814 51958 71878
rect 52022 71814 52028 71878
rect 51816 71808 52028 71814
rect 52632 71884 52844 72020
rect 53040 71944 54204 72020
rect 53040 71884 53252 71944
rect 52632 71878 53252 71884
rect 52632 71814 52638 71878
rect 52702 71814 53252 71878
rect 52632 71808 53252 71814
rect 53856 71884 54204 71944
rect 54264 71884 54476 72020
rect 53856 71878 54476 71884
rect 53856 71814 54134 71878
rect 54198 71814 54476 71878
rect 53856 71808 54476 71814
rect 55216 72014 55836 72020
rect 55216 71950 55358 72014
rect 55422 71950 55836 72014
rect 55216 71944 55836 71950
rect 55216 71808 55428 71944
rect 55488 71878 55836 71944
rect 55488 71814 55766 71878
rect 55830 71814 55836 71878
rect 55488 71808 55836 71814
rect 56440 71884 56652 72020
rect 56848 71884 57060 72020
rect 56440 71878 57060 71884
rect 56440 71814 56446 71878
rect 56510 71814 56990 71878
rect 57054 71814 57060 71878
rect 56440 71808 57060 71814
rect 57664 71944 58284 72020
rect 57664 71878 57876 71944
rect 57664 71814 57670 71878
rect 57734 71814 57876 71878
rect 57664 71808 57876 71814
rect 58072 71878 58284 71944
rect 58072 71814 58214 71878
rect 58278 71814 58284 71878
rect 58072 71808 58284 71814
rect 58888 71884 59100 72020
rect 59296 71884 59508 72020
rect 58888 71878 59508 71884
rect 58888 71814 58894 71878
rect 58958 71814 59508 71878
rect 58888 71808 59508 71814
rect 60112 71944 60732 72020
rect 60112 71808 60460 71944
rect 60520 71878 60732 71944
rect 60520 71814 60662 71878
rect 60726 71814 60732 71878
rect 60520 71808 60732 71814
rect 61472 72014 62092 72020
rect 61472 71950 61478 72014
rect 61542 71950 62092 72014
rect 61472 71944 62092 71950
rect 61472 71878 61684 71944
rect 61472 71814 61478 71878
rect 61542 71814 61684 71878
rect 61472 71808 61684 71814
rect 61744 71878 62092 71944
rect 61744 71814 62022 71878
rect 62086 71814 62092 71878
rect 61744 71808 62092 71814
rect 62696 71884 62908 72020
rect 63104 71884 63316 72020
rect 62696 71878 63316 71884
rect 62696 71814 62702 71878
rect 62766 71814 63110 71878
rect 63174 71814 63316 71878
rect 62696 71808 63316 71814
rect 63920 71944 64540 72020
rect 63920 71878 64132 71944
rect 63920 71814 63926 71878
rect 63990 71814 64132 71878
rect 63920 71808 64132 71814
rect 64328 71878 64540 71944
rect 64328 71814 64470 71878
rect 64534 71814 64540 71878
rect 64328 71808 64540 71814
rect 65144 71884 65356 72020
rect 65552 71884 65764 72020
rect 65144 71878 65764 71884
rect 65144 71814 65150 71878
rect 65214 71814 65694 71878
rect 65758 71814 65764 71878
rect 65144 71808 65764 71814
rect 79288 71742 79636 71748
rect 79288 71678 79294 71742
rect 79358 71678 79636 71742
rect 79288 71536 79636 71678
rect 86904 71612 87116 71748
rect 87720 71742 89156 71748
rect 87720 71678 89086 71742
rect 89150 71678 89156 71742
rect 87720 71672 89156 71678
rect 87720 71612 87932 71672
rect 86904 71536 87932 71612
rect 25160 71470 25644 71476
rect 25160 71406 25574 71470
rect 25638 71406 25644 71470
rect 25160 71400 25644 71406
rect 25160 71340 25372 71400
rect 25704 71340 25916 71476
rect 26384 71470 26868 71476
rect 26384 71406 26798 71470
rect 26862 71406 26868 71470
rect 26384 71400 26868 71406
rect 26384 71340 26596 71400
rect 26928 71340 27140 71476
rect 25160 71264 27140 71340
rect 27608 71470 27820 71476
rect 27608 71406 27614 71470
rect 27678 71406 27750 71470
rect 27814 71406 27820 71470
rect 27608 71340 27820 71406
rect 28152 71340 28500 71476
rect 28832 71470 29044 71476
rect 28832 71406 28974 71470
rect 29038 71406 29044 71470
rect 28832 71340 29044 71406
rect 27608 71264 29044 71340
rect 29512 71470 29724 71476
rect 29512 71406 29518 71470
rect 29582 71406 29724 71470
rect 29512 71340 29724 71406
rect 30056 71340 30268 71476
rect 30736 71470 31628 71476
rect 30736 71406 30742 71470
rect 30806 71406 31422 71470
rect 31486 71406 31628 71470
rect 30736 71400 31628 71406
rect 30736 71340 30948 71400
rect 29512 71264 30948 71340
rect 31280 71264 31628 71400
rect 31960 71470 32580 71476
rect 31960 71406 31966 71470
rect 32030 71406 32510 71470
rect 32574 71406 32580 71470
rect 31960 71400 32580 71406
rect 32640 71470 33124 71476
rect 32640 71406 33054 71470
rect 33118 71406 33124 71470
rect 32640 71400 33124 71406
rect 33184 71470 34076 71476
rect 33184 71406 34006 71470
rect 34070 71406 34076 71470
rect 33184 71400 34076 71406
rect 31960 71264 32172 71400
rect 32640 71340 32852 71400
rect 33184 71340 33396 71400
rect 32640 71264 33396 71340
rect 33864 71264 34076 71400
rect 34408 71470 35300 71476
rect 34408 71406 34414 71470
rect 34478 71406 35230 71470
rect 35294 71406 35300 71470
rect 34408 71400 35300 71406
rect 34408 71264 34756 71400
rect 35088 71264 35300 71400
rect 35768 71470 35980 71476
rect 35768 71406 35774 71470
rect 35838 71406 35980 71470
rect 35768 71340 35980 71406
rect 36312 71470 36524 71476
rect 36312 71406 36454 71470
rect 36518 71406 36524 71470
rect 36312 71340 36524 71406
rect 35768 71264 36524 71340
rect 36992 71470 37748 71476
rect 36992 71406 36998 71470
rect 37062 71406 37678 71470
rect 37742 71406 37748 71470
rect 36992 71400 37748 71406
rect 36992 71264 37204 71400
rect 37536 71264 37748 71400
rect 38216 71470 38428 71476
rect 38216 71406 38222 71470
rect 38286 71406 38428 71470
rect 38216 71340 38428 71406
rect 38760 71470 40332 71476
rect 38760 71406 39446 71470
rect 39510 71406 40262 71470
rect 40326 71406 40332 71470
rect 38760 71400 40332 71406
rect 38760 71340 39108 71400
rect 38216 71264 39108 71340
rect 39440 71264 39652 71400
rect 40120 71264 40332 71400
rect 40664 71470 40876 71476
rect 40664 71406 40670 71470
rect 40734 71406 40876 71470
rect 40664 71340 40876 71406
rect 41344 71470 42780 71476
rect 41344 71406 42710 71470
rect 42774 71406 42780 71470
rect 41344 71400 42780 71406
rect 41344 71340 41556 71400
rect 41888 71340 42236 71400
rect 40664 71264 41556 71340
rect 41654 71334 42236 71340
rect 41616 71270 41622 71334
rect 41686 71270 42236 71334
rect 41654 71264 42236 71270
rect 42568 71264 42780 71400
rect 43248 71470 44684 71476
rect 43248 71406 43254 71470
rect 43318 71406 43934 71470
rect 43998 71406 44684 71470
rect 43248 71400 44684 71406
rect 43248 71264 43460 71400
rect 43792 71264 44004 71400
rect 44472 71340 44684 71400
rect 45016 71470 45364 71476
rect 45016 71406 45158 71470
rect 45222 71406 45364 71470
rect 45016 71340 45364 71406
rect 44472 71264 45364 71340
rect 45696 71470 46588 71476
rect 45696 71406 45702 71470
rect 45766 71406 46588 71470
rect 45696 71400 46588 71406
rect 45696 71264 45908 71400
rect 46376 71340 46588 71400
rect 46920 71470 47132 71476
rect 46920 71406 46926 71470
rect 46990 71406 47132 71470
rect 46920 71340 47132 71406
rect 47600 71470 49036 71476
rect 47600 71406 47742 71470
rect 47806 71406 48966 71470
rect 49030 71406 49036 71470
rect 47600 71400 49036 71406
rect 47600 71340 47812 71400
rect 46376 71264 47812 71340
rect 48144 71264 48356 71400
rect 48824 71264 49036 71400
rect 49368 71470 49716 71476
rect 49368 71406 49374 71470
rect 49438 71406 49716 71470
rect 49368 71340 49716 71406
rect 50048 71470 50940 71476
rect 50048 71406 50190 71470
rect 50254 71406 50940 71470
rect 50048 71400 50940 71406
rect 50048 71340 50260 71400
rect 49368 71264 50260 71340
rect 50728 71340 50940 71400
rect 51272 71470 51484 71476
rect 51272 71406 51414 71470
rect 51478 71406 51484 71470
rect 51272 71340 51484 71406
rect 50728 71264 51484 71340
rect 51952 71470 52844 71476
rect 51952 71406 51958 71470
rect 52022 71406 52638 71470
rect 52702 71406 52844 71470
rect 51952 71400 52844 71406
rect 51952 71264 52164 71400
rect 52496 71340 52844 71400
rect 53176 71340 53388 71476
rect 52496 71264 53388 71340
rect 53856 71400 55292 71476
rect 53856 71264 54068 71400
rect 54400 71340 54612 71400
rect 54166 71334 54612 71340
rect 54128 71270 54134 71334
rect 54198 71270 54612 71334
rect 54166 71264 54612 71270
rect 55080 71340 55292 71400
rect 55624 71470 55972 71476
rect 55624 71406 55766 71470
rect 55830 71406 55972 71470
rect 55624 71340 55972 71406
rect 56304 71470 56516 71476
rect 56304 71406 56446 71470
rect 56510 71406 56516 71470
rect 56304 71340 56516 71406
rect 55080 71264 56516 71340
rect 56984 71470 57196 71476
rect 56984 71406 56990 71470
rect 57054 71406 57196 71470
rect 56984 71340 57196 71406
rect 57528 71470 57740 71476
rect 57528 71406 57670 71470
rect 57734 71406 57740 71470
rect 57528 71340 57740 71406
rect 56984 71264 57740 71340
rect 58208 71470 59644 71476
rect 58208 71406 58214 71470
rect 58278 71406 58894 71470
rect 58958 71406 59644 71470
rect 58208 71400 59644 71406
rect 58208 71264 58420 71400
rect 58752 71264 58964 71400
rect 59432 71340 59644 71400
rect 59976 71340 60324 71476
rect 60656 71470 61548 71476
rect 60656 71406 60662 71470
rect 60726 71406 61478 71470
rect 61542 71406 61548 71470
rect 60656 71400 61548 71406
rect 60656 71340 60868 71400
rect 59432 71264 60868 71340
rect 61336 71264 61548 71400
rect 61880 71470 62092 71476
rect 61880 71406 62022 71470
rect 62086 71406 62092 71470
rect 61880 71340 62092 71406
rect 62560 71470 62772 71476
rect 62560 71406 62702 71470
rect 62766 71406 62772 71470
rect 62560 71340 62772 71406
rect 61880 71264 62772 71340
rect 63104 71470 63996 71476
rect 63104 71406 63110 71470
rect 63174 71406 63926 71470
rect 63990 71406 63996 71470
rect 63104 71400 63996 71406
rect 63104 71264 63452 71400
rect 63784 71264 63996 71400
rect 64464 71470 65220 71476
rect 64464 71406 64470 71470
rect 64534 71406 65150 71470
rect 65214 71406 65220 71470
rect 64464 71400 65220 71406
rect 64464 71264 64676 71400
rect 65008 71264 65220 71400
rect 65688 71470 65900 71476
rect 65688 71406 65694 71470
rect 65758 71406 65900 71470
rect 65688 71340 65900 71406
rect 65688 71334 67804 71340
rect 65688 71270 67734 71334
rect 67798 71270 67804 71334
rect 65688 71264 67804 71270
rect 24072 71068 24284 71204
rect 66776 71198 66988 71204
rect 66776 71134 66782 71198
rect 66846 71134 66988 71198
rect 1224 71062 1844 71068
rect 1224 70998 1230 71062
rect 1294 71012 1844 71062
rect 1294 70998 1718 71012
rect 1224 70992 1718 70998
rect 1632 70956 1718 70992
rect 1774 70956 1844 71012
rect 24072 70992 24420 71068
rect 1632 70856 1844 70956
rect 24344 70932 24420 70992
rect 66776 70992 66988 71134
rect 67728 71062 70660 71068
rect 67728 70998 67734 71062
rect 67798 70998 70660 71062
rect 67728 70992 70660 70998
rect 66776 70932 66852 70992
rect 24344 70926 26052 70932
rect 24344 70862 25982 70926
rect 26046 70862 26052 70926
rect 24344 70856 26052 70862
rect 66368 70856 66852 70932
rect 67728 70856 67940 70992
rect 70448 70932 70660 70992
rect 71264 71062 72836 71068
rect 71264 70998 72766 71062
rect 72830 70998 72836 71062
rect 71264 70992 72836 70998
rect 89080 71012 89428 71068
rect 70448 70926 71204 70932
rect 70448 70862 71134 70926
rect 71198 70862 71204 70926
rect 70448 70856 71204 70862
rect 71264 70926 71476 70992
rect 71264 70862 71406 70926
rect 71470 70862 71476 70926
rect 71264 70856 71476 70862
rect 89080 70956 89216 71012
rect 89272 70956 89428 71012
rect 89080 70932 89428 70956
rect 89080 70926 89836 70932
rect 89080 70862 89766 70926
rect 89830 70862 89836 70926
rect 89080 70856 89836 70862
rect 24344 70720 24692 70856
rect 66368 70720 66580 70856
rect 24480 70660 24556 70720
rect 66368 70660 66444 70720
rect 17816 70382 18028 70524
rect 17816 70318 17958 70382
rect 18022 70318 18028 70382
rect 17816 70312 18028 70318
rect 18224 70382 18436 70524
rect 18224 70318 18230 70382
rect 18294 70318 18436 70382
rect 18224 70312 18436 70318
rect 18632 70382 18980 70524
rect 18632 70318 18910 70382
rect 18974 70318 18980 70382
rect 18632 70312 18980 70318
rect 19040 70382 19252 70524
rect 19040 70318 19046 70382
rect 19110 70318 19252 70382
rect 19040 70312 19252 70318
rect 19448 70382 19660 70524
rect 24344 70448 24692 70660
rect 66368 70518 66580 70660
rect 71166 70518 71476 70524
rect 66368 70454 66510 70518
rect 66574 70454 66580 70518
rect 71128 70454 71134 70518
rect 71198 70454 71406 70518
rect 71470 70454 71476 70518
rect 66368 70448 66580 70454
rect 71166 70448 71476 70454
rect 24480 70388 24556 70448
rect 66368 70388 66444 70448
rect 19448 70318 19590 70382
rect 19654 70318 19660 70382
rect 19448 70312 19660 70318
rect 17816 70110 18028 70116
rect 17816 70046 17958 70110
rect 18022 70046 18028 70110
rect 17816 69974 18028 70046
rect 17816 69910 17958 69974
rect 18022 69910 18028 69974
rect 17816 69904 18028 69910
rect 18224 70110 18436 70116
rect 18224 70046 18230 70110
rect 18294 70046 18436 70110
rect 18224 69974 18436 70046
rect 18224 69910 18230 69974
rect 18294 69910 18436 69974
rect 18224 69904 18436 69910
rect 18632 70110 18980 70116
rect 18632 70046 18910 70110
rect 18974 70046 18980 70110
rect 18632 69904 18980 70046
rect 19040 70110 19252 70116
rect 19040 70046 19046 70110
rect 19110 70046 19252 70110
rect 19040 69974 19252 70046
rect 19040 69910 19182 69974
rect 19246 69910 19252 69974
rect 19040 69904 19252 69910
rect 19448 70110 19660 70116
rect 19448 70046 19590 70110
rect 19654 70046 19660 70110
rect 19448 69974 19660 70046
rect 19448 69910 19590 69974
rect 19654 69910 19660 69974
rect 19448 69904 19660 69910
rect 24344 69904 24692 70388
rect 66368 70110 66580 70388
rect 71264 70382 71476 70448
rect 71264 70318 71270 70382
rect 71334 70318 71476 70382
rect 71264 70312 71476 70318
rect 71672 70382 71884 70524
rect 71672 70318 71678 70382
rect 71742 70318 71884 70382
rect 71672 70312 71884 70318
rect 72080 70382 72292 70524
rect 72488 70388 72700 70524
rect 72390 70382 72700 70388
rect 72080 70318 72222 70382
rect 72286 70318 72292 70382
rect 72352 70318 72358 70382
rect 72422 70318 72700 70382
rect 72080 70312 72292 70318
rect 72390 70312 72700 70318
rect 72896 70518 74196 70524
rect 72896 70454 74126 70518
rect 74190 70454 74196 70518
rect 72896 70448 74196 70454
rect 72896 70382 73108 70448
rect 72896 70318 73038 70382
rect 73102 70318 73108 70382
rect 72896 70312 73108 70318
rect 86904 70252 87116 70388
rect 87720 70252 87932 70388
rect 86904 70246 90516 70252
rect 86904 70182 90446 70246
rect 90510 70182 90516 70246
rect 86904 70176 90516 70182
rect 66368 70046 66510 70110
rect 66574 70046 66580 70110
rect 66368 69904 66580 70046
rect 71264 70110 71476 70116
rect 71264 70046 71270 70110
rect 71334 70046 71476 70110
rect 71264 69974 71476 70046
rect 71264 69910 71406 69974
rect 71470 69910 71476 69974
rect 71264 69904 71476 69910
rect 71672 70110 71884 70116
rect 71672 70046 71678 70110
rect 71742 70046 71884 70110
rect 71672 69974 71884 70046
rect 71672 69910 71814 69974
rect 71878 69910 71884 69974
rect 71672 69904 71884 69910
rect 72080 70110 72428 70116
rect 72080 70046 72222 70110
rect 72286 70046 72358 70110
rect 72422 70046 72428 70110
rect 72080 70040 72428 70046
rect 72080 69980 72292 70040
rect 72488 69980 72700 70116
rect 72080 69974 72700 69980
rect 72080 69910 72630 69974
rect 72694 69910 72700 69974
rect 72080 69904 72700 69910
rect 72896 70110 73108 70116
rect 72896 70046 73038 70110
rect 73102 70046 73108 70110
rect 72896 69974 73108 70046
rect 72896 69910 72902 69974
rect 72966 69910 73108 69974
rect 72896 69904 73108 69910
rect 18632 69844 18708 69904
rect 18360 69768 18708 69844
rect 24344 69844 24420 69904
rect 66368 69844 66444 69904
rect 18360 69708 18436 69768
rect 17816 69702 18028 69708
rect 17816 69638 17958 69702
rect 18022 69638 18028 69702
rect 17816 69566 18028 69638
rect 17816 69502 17822 69566
rect 17886 69502 18028 69566
rect 17816 69496 18028 69502
rect 18224 69702 18980 69708
rect 18224 69638 18230 69702
rect 18294 69638 18980 69702
rect 18224 69632 18980 69638
rect 18224 69566 18436 69632
rect 18224 69502 18230 69566
rect 18294 69502 18436 69566
rect 18224 69496 18436 69502
rect 18632 69496 18980 69632
rect 19040 69702 19252 69708
rect 19040 69638 19182 69702
rect 19246 69638 19252 69702
rect 19040 69566 19252 69638
rect 19040 69502 19182 69566
rect 19246 69502 19252 69566
rect 19040 69496 19252 69502
rect 19448 69702 19660 69708
rect 19448 69638 19590 69702
rect 19654 69638 19660 69702
rect 19448 69566 19660 69638
rect 19448 69502 19454 69566
rect 19518 69502 19660 69566
rect 19448 69496 19660 69502
rect 24344 69632 24692 69844
rect 66368 69632 66580 69844
rect 71264 69702 71476 69708
rect 71264 69638 71406 69702
rect 71470 69638 71476 69702
rect 24344 69572 24420 69632
rect 66368 69572 66444 69632
rect 1632 69332 1844 69436
rect 24344 69360 24692 69572
rect 1632 69300 1718 69332
rect 1224 69294 1718 69300
rect 1224 69230 1230 69294
rect 1294 69276 1718 69294
rect 1774 69276 1844 69332
rect 24616 69300 24692 69360
rect 1294 69230 1844 69276
rect 1224 69224 1844 69230
rect 17816 69294 18028 69300
rect 17816 69230 17822 69294
rect 17886 69230 18028 69294
rect 17816 69158 18028 69230
rect 17816 69094 17822 69158
rect 17886 69094 18028 69158
rect 17816 69088 18028 69094
rect 18224 69294 18436 69300
rect 18224 69230 18230 69294
rect 18294 69230 18436 69294
rect 18224 69158 18436 69230
rect 18632 69164 18980 69300
rect 18534 69158 18980 69164
rect 18224 69094 18230 69158
rect 18294 69094 18436 69158
rect 18496 69094 18502 69158
rect 18566 69094 18980 69158
rect 18224 69088 18436 69094
rect 18534 69088 18980 69094
rect 19040 69294 19252 69300
rect 19040 69230 19182 69294
rect 19246 69230 19252 69294
rect 19040 69158 19252 69230
rect 19040 69094 19046 69158
rect 19110 69094 19252 69158
rect 19040 69088 19252 69094
rect 19448 69294 19660 69300
rect 19448 69230 19454 69294
rect 19518 69230 19660 69294
rect 19448 69158 19660 69230
rect 19448 69094 19590 69158
rect 19654 69094 19660 69158
rect 19448 69088 19660 69094
rect 24344 69088 24692 69300
rect 66368 69360 66580 69572
rect 71264 69566 71476 69638
rect 71264 69502 71406 69566
rect 71470 69502 71476 69566
rect 71264 69496 71476 69502
rect 71672 69702 71884 69708
rect 71672 69638 71814 69702
rect 71878 69638 71884 69702
rect 71672 69566 71884 69638
rect 71672 69502 71678 69566
rect 71742 69502 71884 69566
rect 71672 69496 71884 69502
rect 72080 69566 72292 69708
rect 72080 69502 72222 69566
rect 72286 69502 72292 69566
rect 72080 69496 72292 69502
rect 72488 69702 72700 69708
rect 72488 69638 72630 69702
rect 72694 69638 72700 69702
rect 72488 69496 72700 69638
rect 72896 69702 73108 69708
rect 72896 69638 72902 69702
rect 72966 69638 73108 69702
rect 72896 69566 73108 69638
rect 72896 69502 72902 69566
rect 72966 69502 73108 69566
rect 72896 69496 73108 69502
rect 72488 69436 72564 69496
rect 72216 69360 72564 69436
rect 89080 69430 89836 69436
rect 89080 69366 89766 69430
rect 89830 69366 89836 69430
rect 89080 69360 89836 69366
rect 66368 69300 66444 69360
rect 72216 69300 72292 69360
rect 89080 69332 89428 69360
rect 66368 69088 66580 69300
rect 71264 69294 71476 69300
rect 71264 69230 71406 69294
rect 71470 69230 71476 69294
rect 71264 69158 71476 69230
rect 71264 69094 71270 69158
rect 71334 69094 71476 69158
rect 71264 69088 71476 69094
rect 71672 69294 71884 69300
rect 71672 69230 71678 69294
rect 71742 69230 71884 69294
rect 71672 69158 71884 69230
rect 71672 69094 71678 69158
rect 71742 69094 71884 69158
rect 71672 69088 71884 69094
rect 72080 69294 72700 69300
rect 72080 69230 72222 69294
rect 72286 69230 72700 69294
rect 72080 69224 72700 69230
rect 72080 69164 72292 69224
rect 72080 69158 72428 69164
rect 72080 69094 72358 69158
rect 72422 69094 72428 69158
rect 72080 69088 72428 69094
rect 72488 69088 72700 69224
rect 72896 69294 73108 69300
rect 72896 69230 72902 69294
rect 72966 69230 73108 69294
rect 72896 69158 73108 69230
rect 89080 69294 89216 69332
rect 89080 69230 89086 69294
rect 89150 69276 89216 69294
rect 89272 69276 89428 69332
rect 89150 69230 89428 69276
rect 89080 69224 89428 69230
rect 72896 69094 73038 69158
rect 73102 69094 73108 69158
rect 72896 69088 73108 69094
rect 24344 69028 24420 69088
rect 66504 69028 66580 69088
rect 17816 68886 18028 68892
rect 17816 68822 17822 68886
rect 17886 68822 18028 68886
rect 17816 68680 18028 68822
rect 18224 68886 18572 68892
rect 18224 68822 18230 68886
rect 18294 68822 18502 68886
rect 18566 68822 18572 68886
rect 18224 68816 18572 68822
rect 18224 68750 18436 68816
rect 18632 68756 18980 68892
rect 18534 68750 18980 68756
rect 18224 68686 18366 68750
rect 18430 68686 18436 68750
rect 18496 68686 18502 68750
rect 18566 68686 18980 68750
rect 18224 68680 18436 68686
rect 18534 68680 18980 68686
rect 19040 68886 19252 68892
rect 19040 68822 19046 68886
rect 19110 68822 19252 68886
rect 19040 68750 19252 68822
rect 19040 68686 19182 68750
rect 19246 68686 19252 68750
rect 19040 68680 19252 68686
rect 19448 68886 19660 68892
rect 19448 68822 19590 68886
rect 19654 68822 19660 68886
rect 19448 68750 19660 68822
rect 24344 68816 24692 69028
rect 24616 68756 24692 68816
rect 19448 68686 19454 68750
rect 19518 68686 19660 68750
rect 19448 68680 19660 68686
rect 17816 68620 17892 68680
rect 17816 68272 18028 68620
rect 18360 68544 18708 68620
rect 24344 68544 24692 68756
rect 66368 68816 66580 69028
rect 71264 68886 71476 68892
rect 71264 68822 71270 68886
rect 71334 68822 71476 68886
rect 66368 68756 66444 68816
rect 66368 68614 66580 68756
rect 71264 68750 71476 68822
rect 71264 68686 71406 68750
rect 71470 68686 71476 68750
rect 71264 68680 71476 68686
rect 71672 68886 71884 68892
rect 71672 68822 71678 68886
rect 71742 68822 71884 68886
rect 71672 68750 71884 68822
rect 71672 68686 71814 68750
rect 71878 68686 71884 68750
rect 71672 68680 71884 68686
rect 72080 68750 72292 68892
rect 72390 68886 72700 68892
rect 72352 68822 72358 68886
rect 72422 68822 72700 68886
rect 72390 68816 72700 68822
rect 72080 68686 72086 68750
rect 72150 68686 72292 68750
rect 72080 68680 72292 68686
rect 72488 68750 72700 68816
rect 72488 68686 72494 68750
rect 72558 68686 72700 68750
rect 72488 68680 72700 68686
rect 72896 68886 73108 68892
rect 72896 68822 73038 68886
rect 73102 68822 73108 68886
rect 72896 68680 73108 68822
rect 86904 68756 87116 69028
rect 87720 69022 89156 69028
rect 87720 68958 89086 69022
rect 89150 68958 89156 69022
rect 87720 68952 89156 68958
rect 87720 68756 87932 68952
rect 86904 68680 87932 68756
rect 66368 68550 66374 68614
rect 66438 68550 66580 68614
rect 66368 68544 66580 68550
rect 72896 68620 72972 68680
rect 18360 68484 18436 68544
rect 18632 68484 18708 68544
rect 24480 68484 24556 68544
rect 66368 68484 66444 68544
rect 18224 68478 18572 68484
rect 18224 68414 18366 68478
rect 18430 68414 18502 68478
rect 18566 68414 18572 68478
rect 18224 68408 18572 68414
rect 18224 68348 18436 68408
rect 18224 68272 18572 68348
rect 18632 68272 18980 68484
rect 19040 68478 19252 68484
rect 19040 68414 19182 68478
rect 19246 68414 19252 68478
rect 19040 68342 19252 68414
rect 19040 68278 19046 68342
rect 19110 68278 19252 68342
rect 19040 68272 19252 68278
rect 19448 68478 19660 68484
rect 19448 68414 19454 68478
rect 19518 68414 19660 68478
rect 19448 68342 19660 68414
rect 19448 68278 19590 68342
rect 19654 68278 19660 68342
rect 19448 68272 19660 68278
rect 17952 68212 18028 68272
rect 18360 68212 18436 68272
rect 17816 67864 18028 68212
rect 18224 67864 18436 68212
rect 18496 68212 18572 68272
rect 18496 68136 18980 68212
rect 18632 67940 18980 68136
rect 18534 67934 18980 67940
rect 18496 67870 18502 67934
rect 18566 67870 18980 67934
rect 18534 67864 18980 67870
rect 19040 68070 19252 68076
rect 19040 68006 19046 68070
rect 19110 68006 19252 68070
rect 19040 67934 19252 68006
rect 19040 67870 19046 67934
rect 19110 67870 19252 67934
rect 19040 67864 19252 67870
rect 19448 68070 19660 68076
rect 19448 68006 19590 68070
rect 19654 68006 19660 68070
rect 19448 67934 19660 68006
rect 19448 67870 19454 67934
rect 19518 67870 19660 67934
rect 19448 67864 19660 67870
rect 24344 68000 24692 68484
rect 66368 68342 66580 68484
rect 66368 68278 66374 68342
rect 66438 68278 66510 68342
rect 66574 68278 66580 68342
rect 66368 68000 66580 68278
rect 71264 68478 71476 68484
rect 71264 68414 71406 68478
rect 71470 68414 71476 68478
rect 71264 68342 71476 68414
rect 71264 68278 71270 68342
rect 71334 68278 71476 68342
rect 71264 68272 71476 68278
rect 71672 68478 71884 68484
rect 71672 68414 71814 68478
rect 71878 68414 71884 68478
rect 71672 68342 71884 68414
rect 71672 68278 71814 68342
rect 71878 68278 71884 68342
rect 71672 68272 71884 68278
rect 72080 68478 72292 68484
rect 72080 68414 72086 68478
rect 72150 68414 72292 68478
rect 72080 68272 72292 68414
rect 72216 68212 72292 68272
rect 72080 68076 72292 68212
rect 72488 68478 72700 68484
rect 72488 68414 72494 68478
rect 72558 68414 72700 68478
rect 72488 68272 72700 68414
rect 72896 68272 73108 68620
rect 72488 68212 72564 68272
rect 72896 68212 72972 68272
rect 72488 68076 72700 68212
rect 71264 68070 71476 68076
rect 71264 68006 71270 68070
rect 71334 68006 71476 68070
rect 24344 67940 24420 68000
rect 17816 67804 17892 67864
rect 1224 67798 1844 67804
rect 1224 67734 1230 67798
rect 1294 67734 1844 67798
rect 1224 67728 1844 67734
rect 1632 67652 1844 67728
rect 1632 67596 1718 67652
rect 1774 67596 1844 67652
rect 1632 67456 1844 67596
rect 17816 67662 18028 67804
rect 24344 67728 24692 67940
rect 66368 67934 66580 67940
rect 66368 67870 66510 67934
rect 66574 67870 66580 67934
rect 66368 67728 66580 67870
rect 71264 67934 71476 68006
rect 71264 67870 71270 67934
rect 71334 67870 71476 67934
rect 71264 67864 71476 67870
rect 71672 68070 71884 68076
rect 71672 68006 71814 68070
rect 71878 68006 71884 68070
rect 71672 67934 71884 68006
rect 71672 67870 71678 67934
rect 71742 67870 71884 67934
rect 71672 67864 71884 67870
rect 72080 68000 72700 68076
rect 72080 67940 72292 68000
rect 72080 67934 72428 67940
rect 72080 67870 72358 67934
rect 72422 67870 72428 67934
rect 72080 67864 72428 67870
rect 72488 67864 72700 68000
rect 72896 67864 73108 68212
rect 73032 67804 73108 67864
rect 24344 67668 24420 67728
rect 66504 67668 66580 67728
rect 17816 67598 17822 67662
rect 17886 67598 18028 67662
rect 17816 67592 18028 67598
rect 18224 67662 18572 67668
rect 18224 67598 18502 67662
rect 18566 67598 18572 67662
rect 18224 67592 18572 67598
rect 18224 67456 18436 67592
rect 18632 67456 18980 67668
rect 18360 67396 18436 67456
rect 18904 67396 18980 67456
rect 17816 67390 18028 67396
rect 17816 67326 17822 67390
rect 17886 67326 18028 67390
rect 17816 67254 18028 67326
rect 17816 67190 17822 67254
rect 17886 67190 18028 67254
rect 17816 67184 18028 67190
rect 18224 67320 18980 67396
rect 18224 67260 18436 67320
rect 18224 67254 18572 67260
rect 18224 67190 18502 67254
rect 18566 67190 18572 67254
rect 18224 67184 18572 67190
rect 18632 67184 18980 67320
rect 19040 67662 19252 67668
rect 19040 67598 19046 67662
rect 19110 67598 19252 67662
rect 19040 67456 19252 67598
rect 19448 67662 19660 67668
rect 19448 67598 19454 67662
rect 19518 67598 19660 67662
rect 19448 67456 19660 67598
rect 19040 67396 19116 67456
rect 19448 67396 19524 67456
rect 19040 67048 19252 67396
rect 19448 67048 19660 67396
rect 24344 67390 24692 67668
rect 24344 67326 24350 67390
rect 24414 67326 24692 67390
rect 24344 67320 24692 67326
rect 66368 67390 66580 67668
rect 71264 67662 71476 67668
rect 71264 67598 71270 67662
rect 71334 67598 71476 67662
rect 71264 67456 71476 67598
rect 71400 67396 71476 67456
rect 66368 67326 66510 67390
rect 66574 67326 66580 67390
rect 66368 67320 66580 67326
rect 24344 67118 24692 67124
rect 24344 67054 24350 67118
rect 24414 67054 24692 67118
rect 19040 66988 19116 67048
rect 19448 66988 19524 67048
rect 17816 66982 18028 66988
rect 17816 66918 17822 66982
rect 17886 66918 18028 66982
rect 17816 66846 18028 66918
rect 17816 66782 17822 66846
rect 17886 66782 18028 66846
rect 17816 66776 18028 66782
rect 18224 66640 18436 66988
rect 18534 66982 18980 66988
rect 18496 66918 18502 66982
rect 18566 66918 18980 66982
rect 18534 66912 18980 66918
rect 18632 66640 18980 66912
rect 19040 66640 19252 66988
rect 19448 66640 19660 66988
rect 18360 66580 18436 66640
rect 18768 66580 18844 66640
rect 19176 66580 19252 66640
rect 19584 66580 19660 66640
rect 17816 66574 18028 66580
rect 17816 66510 17822 66574
rect 17886 66510 18028 66574
rect 17816 66438 18028 66510
rect 17816 66374 17958 66438
rect 18022 66374 18028 66438
rect 17816 66368 18028 66374
rect 18224 66504 18980 66580
rect 18224 66368 18436 66504
rect 18632 66438 18980 66504
rect 18632 66374 18910 66438
rect 18974 66374 18980 66438
rect 18632 66368 18980 66374
rect 19040 66438 19252 66580
rect 19040 66374 19182 66438
rect 19246 66374 19252 66438
rect 19040 66368 19252 66374
rect 19448 66438 19660 66580
rect 24344 66982 24692 67054
rect 24344 66918 24622 66982
rect 24686 66918 24692 66982
rect 24344 66710 24692 66918
rect 24344 66646 24622 66710
rect 24686 66646 24692 66710
rect 24344 66504 24692 66646
rect 66368 67118 66580 67124
rect 66368 67054 66510 67118
rect 66574 67054 66580 67118
rect 66368 66982 66580 67054
rect 66368 66918 66510 66982
rect 66574 66918 66580 66982
rect 66368 66710 66580 66918
rect 66368 66646 66510 66710
rect 66574 66646 66580 66710
rect 66368 66504 66580 66646
rect 71264 67048 71476 67396
rect 71672 67662 71884 67668
rect 71672 67598 71678 67662
rect 71742 67598 71884 67662
rect 71672 67456 71884 67598
rect 72080 67456 72292 67668
rect 72390 67662 72700 67668
rect 72352 67598 72358 67662
rect 72422 67598 72700 67662
rect 72390 67592 72700 67598
rect 72896 67662 73108 67804
rect 72896 67598 72902 67662
rect 72966 67598 73108 67662
rect 72896 67592 73108 67598
rect 89080 67798 89836 67804
rect 89080 67734 89766 67798
rect 89830 67734 89836 67798
rect 89080 67728 89836 67734
rect 89080 67652 89428 67728
rect 89080 67596 89216 67652
rect 89272 67596 89428 67652
rect 72488 67456 72700 67592
rect 71672 67396 71748 67456
rect 72080 67396 72156 67456
rect 72488 67396 72564 67456
rect 86904 67396 87116 67532
rect 87720 67396 87932 67532
rect 89080 67456 89428 67596
rect 71672 67048 71884 67396
rect 72080 67254 72292 67396
rect 72080 67190 72086 67254
rect 72150 67190 72292 67254
rect 72080 67184 72292 67190
rect 72488 67254 72700 67396
rect 72488 67190 72630 67254
rect 72694 67190 72700 67254
rect 72488 67184 72700 67190
rect 72896 67390 73108 67396
rect 72896 67326 72902 67390
rect 72966 67326 73108 67390
rect 72896 67254 73108 67326
rect 86904 67390 87932 67396
rect 86904 67326 87726 67390
rect 87790 67326 87932 67390
rect 86904 67320 87932 67326
rect 72896 67190 72902 67254
rect 72966 67190 73108 67254
rect 72896 67184 73108 67190
rect 71264 66988 71340 67048
rect 71808 66988 71884 67048
rect 71264 66640 71476 66988
rect 71672 66640 71884 66988
rect 72080 66982 72292 66988
rect 72080 66918 72086 66982
rect 72150 66918 72292 66982
rect 72080 66716 72292 66918
rect 72488 66982 72700 66988
rect 72488 66918 72630 66982
rect 72694 66918 72700 66982
rect 72080 66710 72428 66716
rect 72080 66646 72086 66710
rect 72150 66646 72428 66710
rect 72080 66640 72428 66646
rect 71400 66580 71476 66640
rect 71808 66580 71884 66640
rect 72216 66580 72292 66640
rect 24480 66444 24556 66504
rect 66368 66444 66444 66504
rect 71264 66444 71476 66580
rect 19448 66374 19454 66438
rect 19518 66374 19660 66438
rect 19448 66368 19660 66374
rect 17816 66166 18028 66172
rect 17816 66102 17958 66166
rect 18022 66102 18028 66166
rect 1632 65972 1844 66036
rect 1632 65916 1718 65972
rect 1774 65916 1844 65972
rect 17816 66030 18028 66102
rect 17816 65966 17822 66030
rect 17886 65966 18028 66030
rect 17816 65960 18028 65966
rect 18224 66030 18436 66172
rect 18224 65966 18230 66030
rect 18294 65966 18436 66030
rect 18224 65960 18436 65966
rect 18632 66166 18980 66172
rect 18632 66102 18910 66166
rect 18974 66102 18980 66166
rect 18632 66030 18980 66102
rect 18632 65966 18774 66030
rect 18838 65966 18980 66030
rect 18632 65960 18980 65966
rect 19040 66166 19252 66172
rect 19040 66102 19182 66166
rect 19246 66102 19252 66166
rect 19040 66030 19252 66102
rect 19040 65966 19046 66030
rect 19110 65966 19252 66030
rect 19040 65960 19252 65966
rect 19448 66166 19660 66172
rect 19448 66102 19454 66166
rect 19518 66102 19660 66166
rect 19448 66030 19660 66102
rect 19448 65966 19454 66030
rect 19518 65966 19660 66030
rect 19448 65960 19660 65966
rect 24344 66166 24692 66444
rect 24344 66102 24622 66166
rect 24686 66102 24692 66166
rect 24344 65960 24692 66102
rect 66368 66166 66580 66444
rect 71264 66438 71612 66444
rect 71264 66374 71406 66438
rect 71470 66374 71612 66438
rect 71264 66368 71612 66374
rect 71672 66438 71884 66580
rect 71672 66374 71814 66438
rect 71878 66374 71884 66438
rect 71672 66368 71884 66374
rect 72080 66444 72292 66580
rect 72352 66580 72428 66640
rect 72488 66640 72700 66918
rect 72896 66982 73108 66988
rect 72896 66918 72902 66982
rect 72966 66918 73108 66982
rect 72896 66846 73108 66918
rect 72896 66782 72902 66846
rect 72966 66782 73108 66846
rect 72896 66776 73108 66782
rect 72488 66580 72564 66640
rect 72352 66504 72700 66580
rect 72080 66368 72428 66444
rect 72488 66368 72700 66504
rect 72896 66574 73108 66580
rect 72896 66510 72902 66574
rect 72966 66510 73108 66574
rect 72896 66438 73108 66510
rect 72896 66374 72902 66438
rect 72966 66374 73108 66438
rect 72896 66368 73108 66374
rect 71536 66308 71612 66368
rect 72352 66308 72428 66368
rect 71536 66302 72156 66308
rect 71536 66238 72086 66302
rect 72150 66238 72156 66302
rect 71536 66232 72156 66238
rect 72352 66232 72564 66308
rect 72488 66172 72564 66232
rect 66368 66102 66510 66166
rect 66574 66102 66580 66166
rect 66368 65960 66580 66102
rect 71264 66166 71476 66172
rect 71264 66102 71406 66166
rect 71470 66102 71476 66166
rect 71264 66030 71476 66102
rect 71264 65966 71270 66030
rect 71334 65966 71476 66030
rect 71264 65960 71476 65966
rect 71672 66166 71884 66172
rect 71672 66102 71814 66166
rect 71878 66102 71884 66166
rect 71672 66030 71884 66102
rect 71672 65966 71678 66030
rect 71742 65966 71884 66030
rect 71672 65960 71884 65966
rect 72080 66096 72700 66172
rect 72080 66036 72292 66096
rect 72080 66030 72428 66036
rect 72080 65966 72222 66030
rect 72286 65966 72358 66030
rect 72422 65966 72428 66030
rect 72080 65960 72428 65966
rect 72488 65960 72700 66096
rect 72896 66166 73108 66172
rect 72896 66102 72902 66166
rect 72966 66102 73108 66166
rect 72896 66030 73108 66102
rect 72896 65966 73038 66030
rect 73102 65966 73108 66030
rect 72896 65960 73108 65966
rect 86904 66096 87932 66172
rect 86904 65960 87116 66096
rect 87720 66036 87932 66096
rect 87720 65972 89428 66036
rect 87720 65960 89216 65972
rect 1632 65900 1844 65916
rect 24480 65900 24556 65960
rect 66504 65900 66580 65960
rect 1224 65894 1844 65900
rect 1224 65830 1230 65894
rect 1294 65830 1844 65894
rect 1224 65824 1844 65830
rect 24344 65894 24692 65900
rect 24344 65830 24622 65894
rect 24686 65830 24692 65894
rect 17816 65758 18028 65764
rect 17816 65694 17822 65758
rect 17886 65694 18028 65758
rect 17816 65622 18028 65694
rect 17816 65558 17822 65622
rect 17886 65558 18028 65622
rect 17816 65552 18028 65558
rect 18224 65758 18436 65764
rect 18224 65694 18230 65758
rect 18294 65694 18436 65758
rect 18224 65622 18436 65694
rect 18632 65758 18980 65764
rect 18632 65694 18774 65758
rect 18838 65694 18980 65758
rect 18632 65628 18980 65694
rect 18534 65622 18980 65628
rect 18224 65558 18230 65622
rect 18294 65558 18436 65622
rect 18496 65558 18502 65622
rect 18566 65558 18980 65622
rect 18224 65552 18436 65558
rect 18534 65552 18980 65558
rect 19040 65758 19252 65764
rect 19040 65694 19046 65758
rect 19110 65694 19252 65758
rect 19040 65622 19252 65694
rect 19040 65558 19046 65622
rect 19110 65558 19252 65622
rect 19040 65552 19252 65558
rect 19448 65758 19660 65764
rect 19448 65694 19454 65758
rect 19518 65694 19660 65758
rect 19448 65622 19660 65694
rect 19448 65558 19454 65622
rect 19518 65558 19660 65622
rect 19448 65552 19660 65558
rect 24344 65688 24692 65830
rect 66368 65894 66580 65900
rect 66368 65830 66510 65894
rect 66574 65830 66580 65894
rect 66368 65688 66580 65830
rect 89080 65916 89216 65960
rect 89272 65916 89428 65972
rect 89080 65900 89428 65916
rect 89080 65894 89836 65900
rect 89080 65830 89766 65894
rect 89830 65830 89836 65894
rect 89080 65824 89836 65830
rect 24344 65628 24420 65688
rect 66504 65628 66580 65688
rect 24344 65416 24692 65628
rect 24616 65356 24692 65416
rect 17816 65350 18028 65356
rect 17816 65286 17822 65350
rect 17886 65286 18028 65350
rect 17816 65214 18028 65286
rect 17816 65150 17822 65214
rect 17886 65150 18028 65214
rect 17816 65144 18028 65150
rect 18224 65350 18572 65356
rect 18224 65286 18230 65350
rect 18294 65286 18502 65350
rect 18566 65286 18572 65350
rect 18224 65280 18572 65286
rect 18224 65220 18436 65280
rect 18632 65220 18980 65356
rect 18224 65214 18980 65220
rect 18224 65150 18638 65214
rect 18702 65150 18980 65214
rect 18224 65144 18980 65150
rect 19040 65350 19252 65356
rect 19040 65286 19046 65350
rect 19110 65286 19252 65350
rect 19040 65214 19252 65286
rect 19040 65150 19182 65214
rect 19246 65150 19252 65214
rect 19040 65144 19252 65150
rect 19448 65350 19660 65356
rect 19448 65286 19454 65350
rect 19518 65286 19660 65350
rect 19448 65214 19660 65286
rect 19448 65150 19454 65214
rect 19518 65150 19660 65214
rect 19448 65144 19660 65150
rect 24344 65144 24692 65356
rect 24616 65084 24692 65144
rect 17816 64942 18028 64948
rect 17816 64878 17822 64942
rect 17886 64878 18028 64942
rect 17816 64736 18028 64878
rect 18224 64806 18436 64948
rect 18224 64742 18230 64806
rect 18294 64742 18436 64806
rect 18224 64736 18436 64742
rect 18632 64942 18980 64948
rect 18632 64878 18638 64942
rect 18702 64878 18980 64942
rect 18632 64806 18980 64878
rect 18632 64742 18910 64806
rect 18974 64742 18980 64806
rect 18632 64736 18980 64742
rect 19040 64942 19252 64948
rect 19040 64878 19182 64942
rect 19246 64878 19252 64942
rect 19040 64806 19252 64878
rect 19040 64742 19046 64806
rect 19110 64742 19252 64806
rect 19040 64736 19252 64742
rect 19448 64942 19660 64948
rect 19448 64878 19454 64942
rect 19518 64878 19660 64942
rect 19448 64806 19660 64878
rect 24344 64872 24692 65084
rect 66368 65416 66580 65628
rect 71264 65758 71476 65764
rect 71264 65694 71270 65758
rect 71334 65694 71476 65758
rect 71264 65622 71476 65694
rect 71264 65558 71406 65622
rect 71470 65558 71476 65622
rect 71264 65552 71476 65558
rect 71672 65758 71884 65764
rect 71672 65694 71678 65758
rect 71742 65694 71884 65758
rect 71672 65622 71884 65694
rect 71672 65558 71678 65622
rect 71742 65558 71884 65622
rect 71672 65552 71884 65558
rect 72080 65758 72292 65764
rect 72390 65758 72700 65764
rect 72080 65694 72222 65758
rect 72286 65694 72292 65758
rect 72352 65694 72358 65758
rect 72422 65694 72700 65758
rect 72080 65622 72292 65694
rect 72390 65688 72700 65694
rect 72080 65558 72086 65622
rect 72150 65558 72292 65622
rect 72080 65552 72292 65558
rect 72488 65622 72700 65688
rect 72488 65558 72494 65622
rect 72558 65558 72700 65622
rect 72488 65552 72700 65558
rect 72896 65758 73108 65764
rect 72896 65694 73038 65758
rect 73102 65694 73108 65758
rect 72896 65622 73108 65694
rect 72896 65558 72902 65622
rect 72966 65558 73108 65622
rect 72896 65552 73108 65558
rect 66368 65356 66444 65416
rect 66368 65144 66580 65356
rect 71264 65350 71476 65356
rect 71264 65286 71406 65350
rect 71470 65286 71476 65350
rect 71264 65214 71476 65286
rect 71264 65150 71406 65214
rect 71470 65150 71476 65214
rect 71264 65144 71476 65150
rect 71672 65350 71884 65356
rect 71672 65286 71678 65350
rect 71742 65286 71884 65350
rect 71672 65214 71884 65286
rect 71672 65150 71814 65214
rect 71878 65150 71884 65214
rect 71672 65144 71884 65150
rect 72080 65350 72292 65356
rect 72080 65286 72086 65350
rect 72150 65286 72292 65350
rect 72080 65144 72292 65286
rect 72488 65350 72700 65356
rect 72488 65286 72494 65350
rect 72558 65286 72700 65350
rect 72488 65220 72700 65286
rect 72390 65214 72700 65220
rect 72352 65150 72358 65214
rect 72422 65150 72700 65214
rect 72390 65144 72700 65150
rect 72896 65350 73108 65356
rect 72896 65286 72902 65350
rect 72966 65286 73108 65350
rect 72896 65214 73108 65286
rect 72896 65150 73038 65214
rect 73102 65150 73108 65214
rect 72896 65144 73108 65150
rect 66368 65084 66444 65144
rect 66368 64872 66580 65084
rect 24616 64812 24692 64872
rect 66504 64812 66580 64872
rect 19448 64742 19590 64806
rect 19654 64742 19660 64806
rect 19448 64736 19660 64742
rect 17816 64676 17892 64736
rect 1632 64292 1844 64404
rect 17816 64398 18028 64676
rect 24344 64600 24692 64812
rect 66368 64600 66580 64812
rect 71264 64942 71476 64948
rect 71264 64878 71406 64942
rect 71470 64878 71476 64942
rect 71264 64806 71476 64878
rect 71264 64742 71270 64806
rect 71334 64742 71476 64806
rect 71264 64736 71476 64742
rect 71672 64942 71884 64948
rect 71672 64878 71814 64942
rect 71878 64878 71884 64942
rect 71672 64806 71884 64878
rect 71672 64742 71678 64806
rect 71742 64742 71884 64806
rect 71672 64736 71884 64742
rect 72080 64942 72428 64948
rect 72080 64878 72358 64942
rect 72422 64878 72428 64942
rect 72080 64872 72428 64878
rect 72080 64812 72292 64872
rect 72488 64812 72700 64948
rect 72080 64806 72700 64812
rect 72080 64742 72222 64806
rect 72286 64742 72630 64806
rect 72694 64742 72700 64806
rect 72080 64736 72700 64742
rect 72896 64942 73108 64948
rect 72896 64878 73038 64942
rect 73102 64878 73108 64942
rect 72896 64736 73108 64878
rect 73032 64676 73108 64736
rect 24616 64540 24692 64600
rect 66504 64540 66580 64600
rect 17816 64334 17958 64398
rect 18022 64334 18028 64398
rect 17816 64328 18028 64334
rect 18224 64534 18436 64540
rect 18224 64470 18230 64534
rect 18294 64470 18436 64534
rect 18224 64398 18436 64470
rect 18224 64334 18366 64398
rect 18430 64334 18436 64398
rect 18224 64328 18436 64334
rect 18632 64534 18980 64540
rect 18632 64470 18910 64534
rect 18974 64470 18980 64534
rect 18632 64328 18980 64470
rect 19040 64534 19252 64540
rect 19040 64470 19046 64534
rect 19110 64470 19252 64534
rect 19040 64398 19252 64470
rect 19040 64334 19182 64398
rect 19246 64334 19252 64398
rect 19040 64328 19252 64334
rect 19448 64534 19660 64540
rect 19448 64470 19590 64534
rect 19654 64470 19660 64534
rect 19448 64398 19660 64470
rect 19448 64334 19590 64398
rect 19654 64334 19660 64398
rect 19448 64328 19660 64334
rect 24344 64328 24692 64540
rect 1632 64268 1718 64292
rect 1224 64262 1718 64268
rect 1224 64198 1230 64262
rect 1294 64236 1718 64262
rect 1774 64236 1844 64292
rect 18632 64268 18708 64328
rect 24616 64268 24692 64328
rect 1294 64198 1844 64236
rect 1224 64192 1844 64198
rect 18360 64192 18708 64268
rect 18360 64132 18436 64192
rect 17816 64126 18028 64132
rect 17816 64062 17958 64126
rect 18022 64062 18028 64126
rect 17816 63920 18028 64062
rect 18224 64126 18980 64132
rect 18224 64062 18366 64126
rect 18430 64062 18980 64126
rect 18224 64056 18980 64062
rect 18224 63920 18436 64056
rect 18632 63990 18980 64056
rect 18632 63926 18910 63990
rect 18974 63926 18980 63990
rect 18632 63920 18980 63926
rect 19040 64126 19252 64132
rect 19040 64062 19182 64126
rect 19246 64062 19252 64126
rect 19040 63990 19252 64062
rect 19040 63926 19182 63990
rect 19246 63926 19252 63990
rect 19040 63920 19252 63926
rect 19448 64126 19660 64132
rect 19448 64062 19590 64126
rect 19654 64062 19660 64126
rect 19448 63990 19660 64062
rect 24344 64056 24692 64268
rect 66368 64328 66580 64540
rect 71264 64534 71476 64540
rect 71264 64470 71270 64534
rect 71334 64470 71476 64534
rect 71264 64398 71476 64470
rect 71264 64334 71406 64398
rect 71470 64334 71476 64398
rect 71264 64328 71476 64334
rect 71672 64534 71884 64540
rect 71672 64470 71678 64534
rect 71742 64470 71884 64534
rect 71672 64398 71884 64470
rect 71672 64334 71678 64398
rect 71742 64334 71884 64398
rect 71672 64328 71884 64334
rect 72080 64534 72292 64540
rect 72080 64470 72222 64534
rect 72286 64470 72292 64534
rect 72080 64328 72292 64470
rect 72488 64534 72700 64540
rect 72488 64470 72630 64534
rect 72694 64470 72700 64534
rect 72488 64398 72700 64470
rect 72488 64334 72494 64398
rect 72558 64334 72700 64398
rect 72488 64328 72700 64334
rect 72896 64398 73108 64676
rect 86904 64670 87932 64676
rect 86904 64606 87726 64670
rect 87790 64606 87932 64670
rect 86904 64600 87932 64606
rect 86904 64540 87116 64600
rect 87720 64540 87932 64600
rect 86904 64534 87660 64540
rect 86904 64470 87590 64534
rect 87654 64470 87660 64534
rect 86904 64464 87660 64470
rect 87720 64534 90516 64540
rect 87720 64470 90446 64534
rect 90510 64470 90516 64534
rect 87720 64464 90516 64470
rect 72896 64334 72902 64398
rect 72966 64334 73108 64398
rect 72896 64328 73108 64334
rect 66368 64268 66444 64328
rect 89080 64292 89428 64404
rect 66368 64056 66580 64268
rect 89080 64236 89216 64292
rect 89272 64268 89428 64292
rect 89272 64262 89836 64268
rect 89272 64236 89766 64262
rect 89080 64198 89766 64236
rect 89830 64198 89836 64262
rect 89080 64192 89836 64198
rect 71264 64126 71476 64132
rect 71264 64062 71406 64126
rect 71470 64062 71476 64126
rect 24480 63996 24556 64056
rect 66368 63996 66444 64056
rect 19448 63926 19590 63990
rect 19654 63926 19660 63990
rect 19448 63920 19660 63926
rect 17952 63860 18028 63920
rect 17816 63718 18028 63860
rect 24344 63854 24692 63996
rect 24344 63790 24486 63854
rect 24550 63790 24692 63854
rect 24344 63784 24692 63790
rect 66368 63854 66580 63996
rect 71264 63990 71476 64062
rect 71264 63926 71270 63990
rect 71334 63926 71476 63990
rect 71264 63920 71476 63926
rect 71672 64126 71884 64132
rect 71672 64062 71678 64126
rect 71742 64062 71884 64126
rect 71672 63990 71884 64062
rect 71672 63926 71678 63990
rect 71742 63926 71884 63990
rect 71672 63920 71884 63926
rect 72080 63990 72292 64132
rect 72488 64126 72700 64132
rect 72488 64062 72494 64126
rect 72558 64062 72700 64126
rect 72488 63996 72700 64062
rect 72390 63990 72700 63996
rect 72080 63926 72086 63990
rect 72150 63926 72292 63990
rect 72352 63926 72358 63990
rect 72422 63926 72700 63990
rect 72080 63920 72292 63926
rect 72390 63920 72700 63926
rect 72896 64126 73108 64132
rect 72896 64062 72902 64126
rect 72966 64062 73108 64126
rect 72896 63920 73108 64062
rect 66368 63790 66510 63854
rect 66574 63790 66580 63854
rect 66368 63784 66580 63790
rect 24344 63724 24420 63784
rect 66504 63724 66580 63784
rect 72896 63860 72972 63920
rect 17816 63654 17822 63718
rect 17886 63654 18028 63718
rect 17816 63648 18028 63654
rect 18224 63512 18436 63724
rect 18632 63718 18980 63724
rect 18632 63654 18910 63718
rect 18974 63654 18980 63718
rect 18632 63588 18980 63654
rect 18496 63512 18980 63588
rect 19040 63718 19252 63724
rect 19040 63654 19182 63718
rect 19246 63654 19252 63718
rect 19040 63512 19252 63654
rect 19448 63718 19660 63724
rect 19448 63654 19590 63718
rect 19654 63654 19660 63718
rect 19448 63512 19660 63654
rect 18224 63452 18300 63512
rect 18496 63452 18572 63512
rect 17816 63446 18028 63452
rect 17816 63382 17822 63446
rect 17886 63382 18028 63446
rect 17816 63310 18028 63382
rect 17816 63246 17958 63310
rect 18022 63246 18028 63310
rect 17816 63240 18028 63246
rect 18224 63376 18572 63452
rect 18632 63452 18708 63512
rect 19040 63452 19116 63512
rect 19584 63452 19660 63512
rect 18224 63316 18436 63376
rect 18224 63310 18572 63316
rect 18224 63246 18502 63310
rect 18566 63246 18572 63310
rect 18224 63240 18572 63246
rect 18632 63240 18980 63452
rect 19040 63104 19252 63452
rect 19176 63044 19252 63104
rect 17816 63038 18028 63044
rect 17816 62974 17958 63038
rect 18022 62974 18028 63038
rect 17816 62902 18028 62974
rect 17816 62838 17958 62902
rect 18022 62838 18028 62902
rect 17816 62832 18028 62838
rect 18224 62696 18436 63044
rect 18534 63038 18980 63044
rect 18496 62974 18502 63038
rect 18566 62974 18980 63038
rect 18534 62968 18980 62974
rect 18752 62772 18850 62968
rect 18360 62636 18436 62696
rect 1632 62612 1844 62636
rect 1632 62556 1718 62612
rect 1774 62556 1844 62612
rect 1632 62500 1844 62556
rect 1224 62494 1844 62500
rect 1224 62430 1230 62494
rect 1294 62430 1844 62494
rect 1224 62424 1844 62430
rect 17816 62630 18028 62636
rect 17816 62566 17958 62630
rect 18022 62566 18028 62630
rect 17816 62494 18028 62566
rect 17816 62430 17822 62494
rect 17886 62430 18028 62494
rect 17816 62424 18028 62430
rect 18224 62494 18436 62636
rect 18224 62430 18366 62494
rect 18430 62430 18436 62494
rect 18224 62424 18436 62430
rect 18632 62696 18980 62772
rect 19040 62696 19252 63044
rect 19448 63104 19660 63452
rect 24344 63582 24692 63724
rect 24344 63518 24486 63582
rect 24550 63518 24692 63582
rect 24344 63446 24692 63518
rect 24344 63382 24622 63446
rect 24686 63382 24692 63446
rect 24344 63376 24692 63382
rect 66368 63582 66580 63724
rect 66368 63518 66510 63582
rect 66574 63518 66580 63582
rect 66368 63446 66580 63518
rect 66368 63382 66374 63446
rect 66438 63382 66580 63446
rect 66368 63376 66580 63382
rect 71264 63718 71476 63724
rect 71264 63654 71270 63718
rect 71334 63654 71476 63718
rect 71264 63512 71476 63654
rect 71672 63718 71884 63724
rect 71672 63654 71678 63718
rect 71742 63654 71884 63718
rect 71672 63512 71884 63654
rect 72080 63718 72428 63724
rect 72080 63654 72086 63718
rect 72150 63654 72358 63718
rect 72422 63654 72428 63718
rect 72080 63648 72428 63654
rect 72080 63588 72292 63648
rect 72488 63588 72700 63724
rect 72896 63718 73108 63860
rect 72896 63654 73038 63718
rect 73102 63654 73108 63718
rect 72896 63648 73108 63654
rect 72080 63512 72700 63588
rect 71264 63452 71340 63512
rect 71808 63452 71884 63512
rect 72216 63452 72292 63512
rect 24344 63174 24692 63180
rect 24344 63110 24622 63174
rect 24686 63110 24692 63174
rect 19448 63044 19524 63104
rect 19448 62696 19660 63044
rect 24344 63038 24692 63110
rect 24344 62974 24350 63038
rect 24414 62974 24692 63038
rect 24344 62766 24692 62974
rect 24344 62702 24350 62766
rect 24414 62702 24692 62766
rect 18632 62636 18708 62696
rect 19040 62636 19116 62696
rect 19448 62636 19524 62696
rect 18632 62424 18980 62636
rect 19040 62494 19252 62636
rect 19040 62430 19046 62494
rect 19110 62430 19252 62494
rect 19040 62424 19252 62430
rect 19448 62494 19660 62636
rect 24344 62560 24692 62702
rect 24616 62500 24692 62560
rect 19448 62430 19590 62494
rect 19654 62430 19660 62494
rect 19448 62424 19660 62430
rect 18632 62364 18708 62424
rect 18360 62288 18708 62364
rect 18360 62228 18436 62288
rect 17816 62222 18028 62228
rect 17816 62158 17822 62222
rect 17886 62158 18028 62222
rect 17816 62086 18028 62158
rect 17816 62022 17822 62086
rect 17886 62022 18028 62086
rect 17816 62016 18028 62022
rect 18224 62222 18980 62228
rect 18224 62158 18366 62222
rect 18430 62158 18980 62222
rect 18224 62152 18980 62158
rect 18224 62016 18436 62152
rect 18632 62086 18980 62152
rect 18632 62022 18910 62086
rect 18974 62022 18980 62086
rect 18632 62016 18980 62022
rect 19040 62222 19252 62228
rect 19040 62158 19046 62222
rect 19110 62158 19252 62222
rect 19040 62086 19252 62158
rect 19040 62022 19182 62086
rect 19246 62022 19252 62086
rect 19040 62016 19252 62022
rect 19448 62222 19660 62228
rect 19448 62158 19590 62222
rect 19654 62158 19660 62222
rect 19448 62086 19660 62158
rect 19448 62022 19454 62086
rect 19518 62022 19660 62086
rect 19448 62016 19660 62022
rect 24344 62016 24692 62500
rect 66368 63174 66580 63180
rect 66368 63110 66374 63174
rect 66438 63110 66580 63174
rect 66368 63038 66580 63110
rect 71264 63104 71476 63452
rect 71400 63044 71476 63104
rect 66368 62974 66374 63038
rect 66438 62974 66580 63038
rect 66368 62766 66580 62974
rect 66368 62702 66374 62766
rect 66438 62702 66510 62766
rect 66574 62702 66580 62766
rect 66368 62560 66580 62702
rect 71264 62696 71476 63044
rect 71672 63104 71884 63452
rect 72080 63310 72292 63452
rect 72080 63246 72086 63310
rect 72150 63246 72292 63310
rect 72080 63240 72292 63246
rect 72488 63452 72564 63512
rect 72488 63240 72700 63452
rect 72896 63446 73108 63452
rect 72896 63382 73038 63446
rect 73102 63382 73108 63446
rect 72896 63310 73108 63382
rect 72896 63246 72902 63310
rect 72966 63246 73108 63310
rect 72896 63240 73108 63246
rect 86904 63180 87116 63316
rect 87720 63180 87932 63316
rect 86904 63174 89156 63180
rect 86904 63110 89086 63174
rect 89150 63110 89156 63174
rect 86904 63104 89156 63110
rect 71672 63044 71748 63104
rect 71672 62696 71884 63044
rect 72080 63038 72292 63044
rect 72080 62974 72086 63038
rect 72150 62974 72292 63038
rect 72080 62696 72292 62974
rect 72488 62696 72700 63044
rect 72896 63038 73108 63044
rect 72896 62974 72902 63038
rect 72966 62974 73108 63038
rect 72896 62902 73108 62974
rect 72896 62838 72902 62902
rect 72966 62838 73108 62902
rect 72896 62832 73108 62838
rect 71264 62636 71340 62696
rect 71672 62636 71748 62696
rect 72216 62636 72292 62696
rect 72624 62636 72700 62696
rect 66368 62500 66444 62560
rect 66368 62494 66580 62500
rect 66368 62430 66510 62494
rect 66574 62430 66580 62494
rect 66368 62016 66580 62430
rect 71264 62494 71476 62636
rect 71264 62430 71406 62494
rect 71470 62430 71476 62494
rect 71264 62424 71476 62430
rect 71672 62494 71884 62636
rect 71672 62430 71678 62494
rect 71742 62430 71884 62494
rect 71672 62424 71884 62430
rect 72080 62560 72700 62636
rect 72080 62424 72292 62560
rect 72488 62494 72700 62560
rect 72488 62430 72494 62494
rect 72558 62430 72700 62494
rect 72488 62424 72700 62430
rect 72896 62630 73108 62636
rect 72896 62566 72902 62630
rect 72966 62566 73108 62630
rect 72896 62494 73108 62566
rect 72896 62430 72902 62494
rect 72966 62430 73108 62494
rect 89080 62630 89836 62636
rect 89080 62566 89086 62630
rect 89150 62612 89766 62630
rect 89150 62566 89216 62612
rect 89080 62556 89216 62566
rect 89272 62566 89766 62612
rect 89830 62566 89836 62630
rect 89272 62560 89836 62566
rect 89272 62556 89428 62560
rect 88464 62490 88530 62491
rect 72896 62424 73108 62430
rect 88422 62426 88465 62490
rect 88529 62426 88572 62490
rect 88464 62425 88530 62426
rect 89080 62424 89428 62556
rect 71264 62222 71476 62228
rect 71264 62158 71406 62222
rect 71470 62158 71476 62222
rect 71264 62086 71476 62158
rect 71264 62022 71406 62086
rect 71470 62022 71476 62086
rect 71264 62016 71476 62022
rect 71672 62222 71884 62228
rect 71672 62158 71678 62222
rect 71742 62158 71884 62222
rect 71672 62086 71884 62158
rect 71672 62022 71678 62086
rect 71742 62022 71884 62086
rect 71672 62016 71884 62022
rect 72080 62086 72292 62228
rect 72488 62222 72700 62228
rect 72488 62158 72494 62222
rect 72558 62158 72700 62222
rect 72488 62092 72700 62158
rect 72390 62086 72700 62092
rect 72080 62022 72086 62086
rect 72150 62022 72292 62086
rect 72352 62022 72358 62086
rect 72422 62022 72700 62086
rect 72080 62016 72292 62022
rect 72390 62016 72700 62022
rect 72896 62222 73108 62228
rect 72896 62158 72902 62222
rect 72966 62158 73108 62222
rect 72896 62086 73108 62158
rect 72896 62022 72902 62086
rect 72966 62022 73108 62086
rect 72896 62016 73108 62022
rect 24480 61956 24556 62016
rect 66368 61956 66444 62016
rect 17816 61814 18028 61820
rect 17816 61750 17822 61814
rect 17886 61750 18028 61814
rect 17816 61678 18028 61750
rect 17816 61614 17822 61678
rect 17886 61614 18028 61678
rect 17816 61608 18028 61614
rect 18224 61678 18436 61820
rect 18224 61614 18230 61678
rect 18294 61614 18436 61678
rect 18224 61608 18436 61614
rect 18632 61814 18980 61820
rect 18632 61750 18910 61814
rect 18974 61750 18980 61814
rect 18632 61678 18980 61750
rect 18632 61614 18774 61678
rect 18838 61614 18980 61678
rect 18632 61608 18980 61614
rect 19040 61814 19252 61820
rect 19040 61750 19182 61814
rect 19246 61750 19252 61814
rect 19040 61678 19252 61750
rect 19040 61614 19046 61678
rect 19110 61614 19252 61678
rect 19040 61608 19252 61614
rect 19448 61814 19660 61820
rect 19448 61750 19454 61814
rect 19518 61750 19660 61814
rect 19448 61678 19660 61750
rect 24344 61744 24692 61956
rect 66368 61744 66580 61956
rect 86904 61950 87932 61956
rect 86904 61886 87726 61950
rect 87790 61886 87932 61950
rect 86904 61880 87932 61886
rect 24616 61684 24692 61744
rect 66504 61684 66580 61744
rect 19448 61614 19454 61678
rect 19518 61614 19660 61678
rect 19448 61608 19660 61614
rect 24344 61472 24692 61684
rect 66368 61472 66580 61684
rect 71264 61814 71476 61820
rect 71264 61750 71406 61814
rect 71470 61750 71476 61814
rect 71264 61678 71476 61750
rect 71264 61614 71270 61678
rect 71334 61614 71476 61678
rect 71264 61608 71476 61614
rect 71672 61814 71884 61820
rect 71672 61750 71678 61814
rect 71742 61750 71884 61814
rect 71672 61678 71884 61750
rect 71672 61614 71814 61678
rect 71878 61614 71884 61678
rect 71672 61608 71884 61614
rect 72080 61814 72428 61820
rect 72080 61750 72086 61814
rect 72150 61750 72358 61814
rect 72422 61750 72428 61814
rect 72080 61744 72428 61750
rect 72080 61684 72292 61744
rect 72080 61678 72428 61684
rect 72080 61614 72222 61678
rect 72286 61614 72358 61678
rect 72422 61614 72428 61678
rect 72080 61608 72428 61614
rect 72488 61608 72700 61820
rect 72896 61814 73108 61820
rect 72896 61750 72902 61814
rect 72966 61750 73108 61814
rect 72896 61678 73108 61750
rect 72896 61614 73038 61678
rect 73102 61614 73108 61678
rect 72896 61608 73108 61614
rect 86904 61608 87116 61880
rect 87720 61608 87932 61880
rect 72216 61548 72292 61608
rect 72488 61548 72564 61608
rect 72216 61472 72564 61548
rect 24344 61412 24420 61472
rect 66504 61412 66580 61472
rect 17816 61406 18028 61412
rect 17816 61342 17822 61406
rect 17886 61342 18028 61406
rect 17816 61270 18028 61342
rect 17816 61206 17958 61270
rect 18022 61206 18028 61270
rect 17816 61200 18028 61206
rect 18224 61406 18436 61412
rect 18224 61342 18230 61406
rect 18294 61342 18436 61406
rect 18224 61270 18436 61342
rect 18224 61206 18366 61270
rect 18430 61206 18436 61270
rect 18224 61200 18436 61206
rect 18632 61406 18980 61412
rect 18632 61342 18774 61406
rect 18838 61342 18980 61406
rect 18632 61270 18980 61342
rect 18632 61206 18774 61270
rect 18838 61206 18980 61270
rect 18632 61200 18980 61206
rect 19040 61406 19252 61412
rect 19040 61342 19046 61406
rect 19110 61342 19252 61406
rect 19040 61270 19252 61342
rect 19040 61206 19046 61270
rect 19110 61206 19252 61270
rect 19040 61200 19252 61206
rect 19448 61406 19660 61412
rect 19448 61342 19454 61406
rect 19518 61342 19660 61406
rect 19448 61270 19660 61342
rect 19448 61206 19590 61270
rect 19654 61206 19660 61270
rect 19448 61200 19660 61206
rect 24344 61200 24692 61412
rect 66368 61200 66580 61412
rect 71264 61406 71476 61412
rect 71264 61342 71270 61406
rect 71334 61342 71476 61406
rect 71264 61270 71476 61342
rect 71264 61206 71406 61270
rect 71470 61206 71476 61270
rect 71264 61200 71476 61206
rect 71672 61406 71884 61412
rect 71672 61342 71814 61406
rect 71878 61342 71884 61406
rect 71672 61270 71884 61342
rect 71672 61206 71814 61270
rect 71878 61206 71884 61270
rect 71672 61200 71884 61206
rect 72080 61406 72292 61412
rect 72390 61406 72700 61412
rect 72080 61342 72222 61406
rect 72286 61342 72292 61406
rect 72352 61342 72358 61406
rect 72422 61342 72700 61406
rect 72080 61270 72292 61342
rect 72390 61336 72700 61342
rect 72080 61206 72086 61270
rect 72150 61206 72292 61270
rect 72080 61200 72292 61206
rect 72488 61270 72700 61336
rect 72488 61206 72630 61270
rect 72694 61206 72700 61270
rect 72488 61200 72700 61206
rect 72896 61406 73108 61412
rect 72896 61342 73038 61406
rect 73102 61342 73108 61406
rect 72896 61270 73108 61342
rect 72896 61206 73038 61270
rect 73102 61206 73108 61270
rect 72896 61200 73108 61206
rect 24344 61140 24420 61200
rect 66504 61140 66580 61200
rect 1632 60932 1844 61004
rect 1632 60876 1718 60932
rect 1774 60876 1844 60932
rect 1632 60868 1844 60876
rect 1224 60862 1844 60868
rect 1224 60798 1230 60862
rect 1294 60798 1844 60862
rect 1224 60792 1844 60798
rect 17816 60998 18028 61004
rect 17816 60934 17958 60998
rect 18022 60934 18028 60998
rect 17816 60792 18028 60934
rect 18224 60998 18980 61004
rect 18224 60934 18366 60998
rect 18430 60934 18774 60998
rect 18838 60934 18980 60998
rect 18224 60928 18980 60934
rect 18224 60792 18436 60928
rect 18632 60862 18980 60928
rect 18632 60798 18638 60862
rect 18702 60798 18980 60862
rect 18632 60792 18980 60798
rect 19040 60998 19252 61004
rect 19040 60934 19046 60998
rect 19110 60934 19252 60998
rect 19040 60862 19252 60934
rect 19040 60798 19046 60862
rect 19110 60798 19252 60862
rect 19040 60792 19252 60798
rect 19448 60998 19660 61004
rect 19448 60934 19590 60998
rect 19654 60934 19660 60998
rect 19448 60862 19660 60934
rect 19448 60798 19454 60862
rect 19518 60798 19660 60862
rect 19448 60792 19660 60798
rect 24344 60928 24692 61140
rect 66368 60928 66580 61140
rect 71264 60998 71476 61004
rect 71264 60934 71406 60998
rect 71470 60934 71476 60998
rect 24344 60868 24420 60928
rect 66368 60868 66444 60928
rect 17816 60732 17892 60792
rect 17816 60454 18028 60732
rect 24344 60656 24692 60868
rect 24616 60596 24692 60656
rect 17816 60390 17958 60454
rect 18022 60390 18028 60454
rect 17816 60384 18028 60390
rect 18224 60454 18436 60596
rect 18224 60390 18230 60454
rect 18294 60390 18436 60454
rect 18224 60384 18436 60390
rect 18632 60590 18980 60596
rect 18632 60526 18638 60590
rect 18702 60526 18980 60590
rect 18632 60454 18980 60526
rect 18632 60390 18910 60454
rect 18974 60390 18980 60454
rect 18632 60384 18980 60390
rect 19040 60590 19252 60596
rect 19040 60526 19046 60590
rect 19110 60526 19252 60590
rect 19040 60454 19252 60526
rect 19040 60390 19046 60454
rect 19110 60390 19252 60454
rect 19040 60384 19252 60390
rect 19448 60590 19660 60596
rect 19448 60526 19454 60590
rect 19518 60526 19660 60590
rect 19448 60454 19660 60526
rect 19448 60390 19454 60454
rect 19518 60390 19660 60454
rect 19448 60384 19660 60390
rect 24344 60384 24692 60596
rect 66368 60656 66580 60868
rect 71264 60862 71476 60934
rect 71264 60798 71270 60862
rect 71334 60798 71476 60862
rect 71264 60792 71476 60798
rect 71672 60998 71884 61004
rect 71672 60934 71814 60998
rect 71878 60934 71884 60998
rect 71672 60862 71884 60934
rect 71672 60798 71678 60862
rect 71742 60798 71884 60862
rect 71672 60792 71884 60798
rect 72080 60998 72292 61004
rect 72080 60934 72086 60998
rect 72150 60934 72292 60998
rect 72080 60792 72292 60934
rect 72488 60998 72700 61004
rect 72488 60934 72630 60998
rect 72694 60934 72700 60998
rect 72488 60792 72700 60934
rect 72896 60998 73108 61004
rect 72896 60934 73038 60998
rect 73102 60934 73108 60998
rect 72896 60792 73108 60934
rect 89080 60998 89836 61004
rect 89080 60934 89766 60998
rect 89830 60934 89836 60998
rect 89080 60932 89836 60934
rect 89080 60876 89216 60932
rect 89272 60928 89836 60932
rect 89272 60876 89428 60928
rect 89080 60792 89428 60876
rect 72488 60732 72564 60792
rect 72216 60656 72564 60732
rect 72896 60732 72972 60792
rect 66368 60596 66444 60656
rect 72216 60596 72292 60656
rect 66368 60384 66580 60596
rect 71264 60590 71476 60596
rect 71264 60526 71270 60590
rect 71334 60526 71476 60590
rect 71264 60454 71476 60526
rect 71264 60390 71270 60454
rect 71334 60390 71476 60454
rect 71264 60384 71476 60390
rect 71672 60590 71884 60596
rect 71672 60526 71678 60590
rect 71742 60526 71884 60590
rect 71672 60454 71884 60526
rect 71672 60390 71678 60454
rect 71742 60390 71884 60454
rect 71672 60384 71884 60390
rect 72080 60520 72700 60596
rect 72080 60454 72292 60520
rect 72080 60390 72222 60454
rect 72286 60390 72292 60454
rect 72080 60384 72292 60390
rect 72488 60454 72700 60520
rect 72488 60390 72630 60454
rect 72694 60390 72700 60454
rect 72488 60384 72700 60390
rect 72896 60454 73108 60732
rect 72896 60390 73038 60454
rect 73102 60390 73108 60454
rect 72896 60384 73108 60390
rect 24344 60324 24420 60384
rect 66504 60324 66580 60384
rect 17816 60182 18028 60188
rect 17816 60118 17958 60182
rect 18022 60118 18028 60182
rect 17816 59976 18028 60118
rect 18224 60182 18436 60188
rect 18224 60118 18230 60182
rect 18294 60118 18436 60182
rect 18224 60052 18436 60118
rect 18632 60182 18980 60188
rect 18632 60118 18910 60182
rect 18974 60118 18980 60182
rect 18224 60046 18572 60052
rect 18224 59982 18366 60046
rect 18430 59982 18502 60046
rect 18566 59982 18572 60046
rect 18224 59976 18572 59982
rect 18632 60046 18980 60118
rect 18632 59982 18774 60046
rect 18838 59982 18980 60046
rect 18632 59976 18980 59982
rect 19040 60182 19252 60188
rect 19040 60118 19046 60182
rect 19110 60118 19252 60182
rect 19040 60046 19252 60118
rect 19040 59982 19182 60046
rect 19246 59982 19252 60046
rect 19040 59976 19252 59982
rect 19448 60182 19660 60188
rect 19448 60118 19454 60182
rect 19518 60118 19660 60182
rect 19448 60046 19660 60118
rect 24344 60112 24692 60324
rect 24616 60052 24692 60112
rect 19448 59982 19454 60046
rect 19518 59982 19660 60046
rect 19448 59976 19660 59982
rect 17816 59916 17892 59976
rect 17816 59774 18028 59916
rect 24344 59910 24692 60052
rect 24344 59846 24622 59910
rect 24686 59846 24692 59910
rect 24344 59840 24692 59846
rect 24616 59780 24692 59840
rect 17816 59710 17822 59774
rect 17886 59710 18028 59774
rect 17816 59704 18028 59710
rect 18224 59774 18436 59780
rect 18534 59774 18980 59780
rect 18224 59710 18366 59774
rect 18430 59710 18436 59774
rect 18496 59710 18502 59774
rect 18566 59710 18774 59774
rect 18838 59710 18980 59774
rect 18224 59568 18436 59710
rect 18534 59704 18980 59710
rect 18632 59568 18980 59704
rect 19040 59774 19252 59780
rect 19040 59710 19182 59774
rect 19246 59710 19252 59774
rect 19040 59638 19252 59710
rect 19040 59574 19182 59638
rect 19246 59574 19252 59638
rect 19040 59568 19252 59574
rect 19448 59774 19660 59780
rect 19448 59710 19454 59774
rect 19518 59710 19660 59774
rect 19448 59638 19660 59710
rect 19448 59574 19590 59638
rect 19654 59574 19660 59638
rect 19448 59568 19660 59574
rect 24344 59638 24692 59780
rect 24344 59574 24622 59638
rect 24686 59574 24692 59638
rect 18224 59508 18300 59568
rect 18904 59508 18980 59568
rect 17816 59502 18028 59508
rect 17816 59438 17822 59502
rect 17886 59438 18028 59502
rect 1632 59252 1844 59372
rect 1632 59236 1718 59252
rect 1224 59230 1718 59236
rect 1224 59166 1230 59230
rect 1294 59196 1718 59230
rect 1774 59196 1844 59252
rect 1294 59166 1844 59196
rect 1224 59160 1844 59166
rect 17816 59160 18028 59438
rect 18224 59160 18436 59508
rect 18632 59230 18980 59508
rect 18632 59166 18910 59230
rect 18974 59166 18980 59230
rect 18632 59160 18980 59166
rect 19040 59366 19252 59372
rect 19040 59302 19182 59366
rect 19246 59302 19252 59366
rect 19040 59160 19252 59302
rect 19448 59366 19660 59372
rect 19448 59302 19590 59366
rect 19654 59302 19660 59366
rect 19448 59160 19660 59302
rect 24344 59296 24692 59574
rect 66368 60112 66580 60324
rect 71264 60182 71476 60188
rect 71264 60118 71270 60182
rect 71334 60118 71476 60182
rect 66368 60052 66444 60112
rect 66368 59910 66580 60052
rect 71264 60046 71476 60118
rect 71264 59982 71406 60046
rect 71470 59982 71476 60046
rect 71264 59976 71476 59982
rect 71672 60182 71884 60188
rect 71672 60118 71678 60182
rect 71742 60118 71884 60182
rect 71672 60046 71884 60118
rect 71672 59982 71678 60046
rect 71742 59982 71884 60046
rect 71672 59976 71884 59982
rect 72080 60182 72292 60188
rect 72080 60118 72222 60182
rect 72286 60118 72292 60182
rect 72080 60046 72292 60118
rect 72080 59982 72086 60046
rect 72150 59982 72292 60046
rect 72080 59976 72292 59982
rect 72488 60182 72700 60188
rect 72488 60118 72630 60182
rect 72694 60118 72700 60182
rect 72488 59976 72700 60118
rect 72896 60182 73108 60188
rect 72896 60118 73038 60182
rect 73102 60118 73108 60182
rect 72896 59976 73108 60118
rect 66368 59846 66374 59910
rect 66438 59846 66580 59910
rect 66368 59840 66580 59846
rect 72896 59916 72972 59976
rect 66368 59780 66444 59840
rect 66368 59638 66580 59780
rect 66368 59574 66374 59638
rect 66438 59574 66510 59638
rect 66574 59574 66580 59638
rect 66368 59296 66580 59574
rect 71264 59774 71476 59780
rect 71264 59710 71406 59774
rect 71470 59710 71476 59774
rect 71264 59638 71476 59710
rect 71264 59574 71270 59638
rect 71334 59574 71476 59638
rect 71264 59568 71476 59574
rect 71672 59774 71884 59780
rect 71672 59710 71678 59774
rect 71742 59710 71884 59774
rect 71672 59638 71884 59710
rect 71672 59574 71814 59638
rect 71878 59574 71884 59638
rect 71672 59568 71884 59574
rect 72080 59774 72292 59780
rect 72080 59710 72086 59774
rect 72150 59710 72292 59774
rect 72080 59568 72292 59710
rect 72488 59644 72700 59780
rect 72896 59774 73108 59916
rect 72896 59710 72902 59774
rect 72966 59710 73108 59774
rect 72896 59704 73108 59710
rect 72216 59508 72292 59568
rect 72352 59568 72700 59644
rect 72352 59508 72428 59568
rect 72080 59432 72428 59508
rect 72080 59372 72292 59432
rect 72488 59372 72700 59508
rect 71264 59366 71476 59372
rect 71264 59302 71270 59366
rect 71334 59302 71476 59366
rect 24480 59236 24556 59296
rect 17952 59100 18028 59160
rect 17816 58958 18028 59100
rect 19040 59100 19116 59160
rect 19448 59100 19524 59160
rect 17816 58894 17822 58958
rect 17886 58894 18028 58958
rect 17816 58888 18028 58894
rect 18224 58752 18436 58964
rect 18632 58958 18980 58964
rect 18632 58894 18910 58958
rect 18974 58894 18980 58958
rect 18632 58828 18980 58894
rect 18534 58822 18980 58828
rect 18496 58758 18502 58822
rect 18566 58758 18980 58822
rect 18534 58752 18980 58758
rect 19040 58752 19252 59100
rect 19448 58752 19660 59100
rect 18360 58692 18436 58752
rect 19176 58692 19252 58752
rect 19584 58692 19660 58752
rect 17816 58686 18028 58692
rect 17816 58622 17822 58686
rect 17886 58622 18028 58686
rect 17816 58550 18028 58622
rect 17816 58486 17822 58550
rect 17886 58486 18028 58550
rect 17816 58480 18028 58486
rect 18224 58616 18980 58692
rect 18224 58556 18436 58616
rect 18224 58550 18572 58556
rect 18224 58486 18502 58550
rect 18566 58486 18572 58550
rect 18224 58480 18572 58486
rect 18632 58550 18980 58616
rect 18632 58486 18774 58550
rect 18838 58486 18980 58550
rect 18632 58480 18980 58486
rect 19040 58344 19252 58692
rect 19448 58344 19660 58692
rect 24344 58686 24692 59236
rect 24344 58622 24350 58686
rect 24414 58622 24692 58686
rect 24344 58616 24692 58622
rect 66368 59230 66580 59236
rect 66368 59166 66510 59230
rect 66574 59166 66580 59230
rect 66368 59094 66580 59166
rect 66368 59030 66374 59094
rect 66438 59030 66580 59094
rect 66368 58822 66580 59030
rect 66368 58758 66374 58822
rect 66438 58758 66580 58822
rect 66368 58686 66580 58758
rect 66368 58622 66510 58686
rect 66574 58622 66580 58686
rect 66368 58616 66580 58622
rect 71264 59160 71476 59302
rect 71672 59366 71884 59372
rect 71672 59302 71814 59366
rect 71878 59302 71884 59366
rect 71672 59160 71884 59302
rect 72080 59296 72700 59372
rect 72080 59236 72292 59296
rect 72080 59230 72428 59236
rect 72080 59166 72358 59230
rect 72422 59166 72428 59230
rect 72080 59160 72428 59166
rect 72488 59160 72700 59296
rect 72896 59502 73108 59508
rect 72896 59438 72902 59502
rect 72966 59438 73108 59502
rect 72896 59160 73108 59438
rect 89080 59252 89428 59372
rect 89080 59196 89216 59252
rect 89272 59236 89428 59252
rect 89272 59230 89836 59236
rect 89272 59196 89766 59230
rect 89080 59166 89766 59196
rect 89830 59166 89836 59230
rect 89080 59160 89836 59166
rect 71264 59100 71340 59160
rect 71808 59100 71884 59160
rect 73032 59100 73108 59160
rect 71264 58752 71476 59100
rect 71672 58752 71884 59100
rect 72080 58752 72292 58964
rect 72390 58958 72700 58964
rect 72352 58894 72358 58958
rect 72422 58894 72700 58958
rect 72390 58888 72700 58894
rect 72896 58958 73108 59100
rect 72896 58894 72902 58958
rect 72966 58894 73108 58958
rect 72896 58888 73108 58894
rect 72488 58752 72700 58888
rect 71264 58692 71340 58752
rect 71672 58692 71748 58752
rect 72080 58692 72156 58752
rect 72488 58692 72564 58752
rect 24344 58414 24692 58420
rect 24344 58350 24350 58414
rect 24414 58350 24692 58414
rect 19040 58284 19116 58344
rect 19448 58284 19524 58344
rect 17816 58278 18028 58284
rect 17816 58214 17822 58278
rect 17886 58214 18028 58278
rect 17816 58142 18028 58214
rect 17816 58078 17822 58142
rect 17886 58078 18028 58142
rect 17816 58072 18028 58078
rect 18224 57936 18436 58284
rect 18632 58278 18980 58284
rect 18632 58214 18774 58278
rect 18838 58214 18980 58278
rect 18632 57936 18980 58214
rect 19040 58142 19252 58284
rect 19040 58078 19046 58142
rect 19110 58078 19252 58142
rect 19040 58072 19252 58078
rect 19448 58142 19660 58284
rect 19448 58078 19454 58142
rect 19518 58078 19660 58142
rect 19448 58072 19660 58078
rect 24344 58072 24692 58350
rect 66368 58414 66580 58420
rect 66368 58350 66510 58414
rect 66574 58350 66580 58414
rect 66368 58072 66580 58350
rect 71264 58344 71476 58692
rect 71672 58344 71884 58692
rect 72080 58550 72292 58692
rect 72488 58556 72700 58692
rect 72390 58550 72700 58556
rect 72080 58486 72086 58550
rect 72150 58486 72292 58550
rect 72352 58486 72358 58550
rect 72422 58486 72700 58550
rect 72080 58480 72292 58486
rect 72390 58480 72700 58486
rect 72896 58686 73108 58692
rect 72896 58622 72902 58686
rect 72966 58622 73108 58686
rect 72896 58550 73108 58622
rect 72896 58486 73038 58550
rect 73102 58486 73108 58550
rect 72896 58480 73108 58486
rect 71264 58284 71340 58344
rect 71672 58284 71748 58344
rect 71264 58142 71476 58284
rect 71264 58078 71270 58142
rect 71334 58078 71476 58142
rect 71264 58072 71476 58078
rect 71672 58142 71884 58284
rect 71672 58078 71814 58142
rect 71878 58078 71884 58142
rect 71672 58072 71884 58078
rect 72080 58278 72428 58284
rect 72080 58214 72086 58278
rect 72150 58214 72358 58278
rect 72422 58214 72428 58278
rect 72080 58208 72428 58214
rect 24480 58012 24556 58072
rect 66504 58012 66580 58072
rect 18360 57876 18436 57936
rect 18768 57876 18844 57936
rect 17816 57870 18028 57876
rect 17816 57806 17822 57870
rect 17886 57806 18028 57870
rect 17816 57734 18028 57806
rect 17816 57670 17822 57734
rect 17886 57670 18028 57734
rect 17816 57664 18028 57670
rect 18224 57800 18980 57876
rect 18224 57664 18436 57800
rect 18632 57734 18980 57800
rect 18632 57670 18638 57734
rect 18702 57670 18980 57734
rect 18632 57664 18980 57670
rect 19040 57870 19252 57876
rect 19040 57806 19046 57870
rect 19110 57806 19252 57870
rect 19040 57734 19252 57806
rect 19040 57670 19182 57734
rect 19246 57670 19252 57734
rect 19040 57664 19252 57670
rect 19448 57870 19660 57876
rect 19448 57806 19454 57870
rect 19518 57806 19660 57870
rect 19448 57734 19660 57806
rect 24344 57800 24692 58012
rect 66368 57800 66580 58012
rect 72080 58012 72292 58208
rect 72080 57936 72428 58012
rect 72216 57876 72292 57936
rect 71264 57870 71476 57876
rect 71264 57806 71270 57870
rect 71334 57806 71476 57870
rect 24480 57740 24556 57800
rect 66368 57740 66444 57800
rect 19448 57670 19454 57734
rect 19518 57670 19660 57734
rect 19448 57664 19660 57670
rect 1632 57572 1844 57604
rect 1632 57516 1718 57572
rect 1774 57516 1844 57572
rect 24344 57528 24692 57740
rect 1632 57468 1844 57516
rect 24616 57468 24692 57528
rect 1224 57462 1844 57468
rect 1224 57398 1230 57462
rect 1294 57398 1844 57462
rect 1224 57392 1844 57398
rect 17816 57462 18028 57468
rect 17816 57398 17822 57462
rect 17886 57398 18028 57462
rect 17816 57326 18028 57398
rect 17816 57262 17822 57326
rect 17886 57262 18028 57326
rect 17816 57256 18028 57262
rect 18224 57462 18980 57468
rect 18224 57398 18638 57462
rect 18702 57398 18980 57462
rect 18224 57392 18980 57398
rect 18224 57326 18436 57392
rect 18224 57262 18230 57326
rect 18294 57262 18436 57326
rect 18224 57256 18436 57262
rect 18632 57256 18980 57392
rect 19040 57462 19252 57468
rect 19040 57398 19182 57462
rect 19246 57398 19252 57462
rect 19040 57326 19252 57398
rect 19040 57262 19046 57326
rect 19110 57262 19252 57326
rect 19040 57256 19252 57262
rect 19448 57462 19660 57468
rect 19448 57398 19454 57462
rect 19518 57398 19660 57462
rect 19448 57326 19660 57398
rect 19448 57262 19590 57326
rect 19654 57262 19660 57326
rect 19448 57256 19660 57262
rect 24344 57256 24692 57468
rect 66368 57528 66580 57740
rect 71264 57734 71476 57806
rect 71264 57670 71406 57734
rect 71470 57670 71476 57734
rect 71264 57664 71476 57670
rect 71672 57870 71884 57876
rect 71672 57806 71814 57870
rect 71878 57806 71884 57870
rect 71672 57734 71884 57806
rect 71672 57670 71814 57734
rect 71878 57670 71884 57734
rect 71672 57664 71884 57670
rect 72080 57664 72292 57876
rect 72352 57876 72428 57936
rect 72488 57936 72700 58284
rect 72896 58278 73108 58284
rect 72896 58214 73038 58278
rect 73102 58214 73108 58278
rect 72896 58142 73108 58214
rect 72896 58078 72902 58142
rect 72966 58078 73108 58142
rect 72896 58072 73108 58078
rect 72488 57876 72564 57936
rect 72352 57800 72700 57876
rect 72488 57740 72700 57800
rect 72390 57734 72700 57740
rect 72352 57670 72358 57734
rect 72422 57670 72700 57734
rect 72390 57664 72700 57670
rect 72896 57870 73108 57876
rect 72896 57806 72902 57870
rect 72966 57806 73108 57870
rect 72896 57734 73108 57806
rect 72896 57670 72902 57734
rect 72966 57670 73108 57734
rect 72896 57664 73108 57670
rect 71944 57528 72972 57604
rect 66368 57468 66444 57528
rect 71944 57468 72020 57528
rect 72896 57468 72972 57528
rect 89080 57572 89428 57604
rect 89080 57516 89216 57572
rect 89272 57516 89428 57572
rect 89080 57468 89428 57516
rect 66368 57256 66580 57468
rect 71264 57462 71476 57468
rect 71264 57398 71406 57462
rect 71470 57398 71476 57462
rect 71264 57326 71476 57398
rect 71264 57262 71270 57326
rect 71334 57262 71476 57326
rect 71264 57256 71476 57262
rect 71672 57462 72020 57468
rect 71672 57398 71814 57462
rect 71878 57398 72020 57462
rect 71672 57392 72020 57398
rect 72080 57462 72428 57468
rect 72080 57398 72358 57462
rect 72422 57398 72428 57462
rect 72080 57392 72428 57398
rect 71672 57326 71884 57392
rect 71672 57262 71814 57326
rect 71878 57262 71884 57326
rect 71672 57256 71884 57262
rect 72080 57326 72292 57392
rect 72080 57262 72222 57326
rect 72286 57262 72292 57326
rect 72080 57256 72292 57262
rect 72488 57256 72700 57468
rect 72896 57462 73108 57468
rect 72896 57398 72902 57462
rect 72966 57398 73108 57462
rect 72896 57326 73108 57398
rect 89080 57462 89836 57468
rect 89080 57398 89766 57462
rect 89830 57398 89836 57462
rect 89080 57392 89836 57398
rect 72896 57262 73038 57326
rect 73102 57262 73108 57326
rect 72896 57256 73108 57262
rect 24480 57196 24556 57256
rect 66504 57196 66580 57256
rect 72488 57196 72564 57256
rect 17816 57054 18028 57060
rect 17816 56990 17822 57054
rect 17886 56990 18028 57054
rect 17816 56918 18028 56990
rect 17816 56854 17958 56918
rect 18022 56854 18028 56918
rect 17816 56848 18028 56854
rect 18224 57054 18436 57060
rect 18224 56990 18230 57054
rect 18294 56990 18436 57054
rect 18224 56918 18436 56990
rect 18632 56924 18980 57060
rect 18534 56918 18980 56924
rect 18224 56854 18366 56918
rect 18430 56854 18436 56918
rect 18496 56854 18502 56918
rect 18566 56854 18980 56918
rect 18224 56848 18436 56854
rect 18534 56848 18980 56854
rect 19040 57054 19252 57060
rect 19040 56990 19046 57054
rect 19110 56990 19252 57054
rect 19040 56918 19252 56990
rect 19040 56854 19182 56918
rect 19246 56854 19252 56918
rect 19040 56848 19252 56854
rect 19448 57054 19660 57060
rect 19448 56990 19590 57054
rect 19654 56990 19660 57054
rect 19448 56918 19660 56990
rect 19448 56854 19590 56918
rect 19654 56854 19660 56918
rect 19448 56848 19660 56854
rect 24344 56984 24692 57196
rect 66368 56984 66580 57196
rect 72216 57120 72564 57196
rect 72216 57060 72292 57120
rect 24344 56924 24420 56984
rect 66504 56924 66580 56984
rect 18360 56712 18708 56788
rect 24344 56712 24692 56924
rect 18360 56652 18436 56712
rect 18632 56652 18708 56712
rect 24616 56652 24692 56712
rect 17816 56646 18028 56652
rect 17816 56582 17958 56646
rect 18022 56582 18028 56646
rect 17816 56510 18028 56582
rect 17816 56446 17822 56510
rect 17886 56446 18028 56510
rect 17816 56440 18028 56446
rect 18224 56646 18572 56652
rect 18224 56582 18366 56646
rect 18430 56582 18502 56646
rect 18566 56582 18572 56646
rect 18224 56576 18572 56582
rect 18224 56516 18436 56576
rect 18224 56510 18572 56516
rect 18224 56446 18366 56510
rect 18430 56446 18502 56510
rect 18566 56446 18572 56510
rect 18224 56440 18572 56446
rect 18632 56440 18980 56652
rect 19040 56646 19252 56652
rect 19040 56582 19182 56646
rect 19246 56582 19252 56646
rect 19040 56510 19252 56582
rect 19040 56446 19182 56510
rect 19246 56446 19252 56510
rect 19040 56440 19252 56446
rect 19448 56646 19660 56652
rect 19448 56582 19590 56646
rect 19654 56582 19660 56646
rect 19448 56510 19660 56582
rect 19448 56446 19590 56510
rect 19654 56446 19660 56510
rect 19448 56440 19660 56446
rect 24344 56440 24692 56652
rect 66368 56712 66580 56924
rect 71264 57054 71476 57060
rect 71264 56990 71270 57054
rect 71334 56990 71476 57054
rect 71264 56918 71476 56990
rect 71264 56854 71270 56918
rect 71334 56854 71476 56918
rect 71264 56848 71476 56854
rect 71672 57054 71884 57060
rect 71672 56990 71814 57054
rect 71878 56990 71884 57054
rect 71672 56918 71884 56990
rect 71672 56854 71678 56918
rect 71742 56854 71884 56918
rect 71672 56848 71884 56854
rect 72080 57054 72700 57060
rect 72080 56990 72222 57054
rect 72286 56990 72700 57054
rect 72080 56984 72700 56990
rect 72080 56918 72292 56984
rect 72080 56854 72086 56918
rect 72150 56854 72292 56918
rect 72080 56848 72292 56854
rect 72488 56918 72700 56984
rect 72488 56854 72494 56918
rect 72558 56854 72700 56918
rect 72488 56848 72700 56854
rect 72896 57054 73108 57060
rect 72896 56990 73038 57054
rect 73102 56990 73108 57054
rect 72896 56918 73108 56990
rect 72896 56854 72902 56918
rect 72966 56854 73108 56918
rect 72896 56848 73108 56854
rect 66368 56652 66444 56712
rect 66368 56440 66580 56652
rect 71264 56646 71476 56652
rect 71264 56582 71270 56646
rect 71334 56582 71476 56646
rect 71264 56510 71476 56582
rect 71264 56446 71406 56510
rect 71470 56446 71476 56510
rect 71264 56440 71476 56446
rect 71672 56646 71884 56652
rect 71672 56582 71678 56646
rect 71742 56582 71884 56646
rect 71672 56510 71884 56582
rect 71672 56446 71678 56510
rect 71742 56446 71884 56510
rect 71672 56440 71884 56446
rect 72080 56646 72292 56652
rect 72080 56582 72086 56646
rect 72150 56582 72292 56646
rect 72080 56440 72292 56582
rect 72488 56646 72700 56652
rect 72488 56582 72494 56646
rect 72558 56582 72700 56646
rect 72488 56516 72700 56582
rect 72390 56510 72700 56516
rect 72352 56446 72358 56510
rect 72422 56446 72700 56510
rect 72390 56440 72700 56446
rect 72896 56646 73108 56652
rect 72896 56582 72902 56646
rect 72966 56582 73108 56646
rect 72896 56510 73108 56582
rect 72896 56446 72902 56510
rect 72966 56446 73108 56510
rect 72896 56440 73108 56446
rect 24344 56380 24420 56440
rect 66368 56380 66444 56440
rect 17816 56238 18028 56244
rect 17816 56174 17822 56238
rect 17886 56174 18028 56238
rect 17816 56032 18028 56174
rect 18224 56238 18436 56244
rect 18534 56238 18980 56244
rect 18224 56174 18366 56238
rect 18430 56174 18436 56238
rect 18496 56174 18502 56238
rect 18566 56174 18980 56238
rect 18224 56032 18436 56174
rect 18534 56168 18980 56174
rect 18632 56102 18980 56168
rect 18632 56038 18910 56102
rect 18974 56038 18980 56102
rect 18632 56032 18980 56038
rect 19040 56238 19252 56244
rect 19040 56174 19182 56238
rect 19246 56174 19252 56238
rect 19040 56102 19252 56174
rect 19040 56038 19046 56102
rect 19110 56038 19252 56102
rect 19040 56032 19252 56038
rect 19448 56238 19660 56244
rect 19448 56174 19590 56238
rect 19654 56174 19660 56238
rect 19448 56102 19660 56174
rect 24344 56168 24692 56380
rect 66368 56168 66580 56380
rect 24480 56108 24556 56168
rect 66504 56108 66580 56168
rect 19448 56038 19590 56102
rect 19654 56038 19660 56102
rect 19448 56032 19660 56038
rect 17816 55972 17892 56032
rect 1632 55892 1844 55972
rect 1632 55836 1718 55892
rect 1774 55836 1844 55892
rect 1224 55830 1844 55836
rect 1224 55766 1230 55830
rect 1294 55766 1844 55830
rect 1224 55760 1844 55766
rect 17816 55624 18028 55972
rect 24344 55896 24692 56108
rect 66368 55896 66580 56108
rect 71264 56238 71476 56244
rect 71264 56174 71406 56238
rect 71470 56174 71476 56238
rect 71264 56102 71476 56174
rect 71264 56038 71270 56102
rect 71334 56038 71476 56102
rect 71264 56032 71476 56038
rect 71672 56238 71884 56244
rect 71672 56174 71678 56238
rect 71742 56174 71884 56238
rect 71672 56102 71884 56174
rect 71672 56038 71678 56102
rect 71742 56038 71884 56102
rect 71672 56032 71884 56038
rect 72080 56238 72428 56244
rect 72080 56174 72358 56238
rect 72422 56174 72428 56238
rect 72080 56168 72428 56174
rect 72080 56108 72292 56168
rect 72488 56108 72700 56244
rect 72080 56102 72700 56108
rect 72080 56038 72630 56102
rect 72694 56038 72700 56102
rect 72080 56032 72700 56038
rect 72896 56238 73108 56244
rect 72896 56174 72902 56238
rect 72966 56174 73108 56238
rect 72896 56032 73108 56174
rect 73032 55972 73108 56032
rect 24344 55836 24420 55896
rect 66504 55836 66580 55896
rect 17952 55564 18028 55624
rect 17816 55216 18028 55564
rect 18224 55624 18436 55836
rect 18632 55830 18980 55836
rect 18632 55766 18910 55830
rect 18974 55766 18980 55830
rect 18632 55624 18980 55766
rect 19040 55830 19252 55836
rect 19040 55766 19046 55830
rect 19110 55766 19252 55830
rect 19040 55694 19252 55766
rect 19040 55630 19182 55694
rect 19246 55630 19252 55694
rect 19040 55624 19252 55630
rect 19448 55830 19660 55836
rect 19448 55766 19590 55830
rect 19654 55766 19660 55830
rect 19448 55694 19660 55766
rect 19448 55630 19590 55694
rect 19654 55630 19660 55694
rect 19448 55624 19660 55630
rect 18224 55564 18300 55624
rect 18632 55564 18708 55624
rect 18224 55292 18436 55564
rect 18632 55292 18980 55564
rect 18224 55286 18980 55292
rect 18224 55222 18638 55286
rect 18702 55222 18980 55286
rect 18224 55216 18980 55222
rect 19040 55422 19252 55428
rect 19040 55358 19182 55422
rect 19246 55358 19252 55422
rect 19040 55216 19252 55358
rect 19448 55422 19660 55428
rect 19448 55358 19590 55422
rect 19654 55358 19660 55422
rect 19448 55216 19660 55358
rect 24344 55352 24692 55836
rect 66368 55352 66580 55836
rect 71264 55830 71476 55836
rect 71264 55766 71270 55830
rect 71334 55766 71476 55830
rect 71264 55694 71476 55766
rect 71264 55630 71406 55694
rect 71470 55630 71476 55694
rect 71264 55624 71476 55630
rect 71672 55830 71884 55836
rect 71672 55766 71678 55830
rect 71742 55766 71884 55830
rect 71672 55694 71884 55766
rect 71672 55630 71814 55694
rect 71878 55630 71884 55694
rect 71672 55624 71884 55630
rect 72080 55830 72700 55836
rect 72080 55766 72630 55830
rect 72694 55766 72700 55830
rect 72080 55760 72700 55766
rect 72080 55624 72292 55760
rect 72488 55624 72700 55760
rect 72896 55624 73108 55972
rect 89080 55892 89428 55972
rect 89080 55836 89216 55892
rect 89272 55836 89428 55892
rect 89080 55830 89836 55836
rect 89080 55766 89766 55830
rect 89830 55766 89836 55830
rect 89080 55760 89836 55766
rect 72216 55564 72292 55624
rect 72896 55564 72972 55624
rect 71264 55422 71476 55428
rect 71264 55358 71406 55422
rect 71470 55358 71476 55422
rect 24480 55292 24556 55352
rect 66368 55292 66444 55352
rect 17816 55156 17892 55216
rect 19176 55156 19252 55216
rect 19584 55156 19660 55216
rect 17816 55014 18028 55156
rect 17816 54950 17958 55014
rect 18022 54950 18028 55014
rect 17816 54944 18028 54950
rect 18224 54808 18436 55020
rect 18632 55014 18980 55020
rect 18632 54950 18638 55014
rect 18702 54950 18980 55014
rect 18632 54884 18980 54950
rect 18496 54808 18980 54884
rect 18224 54748 18300 54808
rect 18496 54748 18572 54808
rect 18904 54748 18980 54808
rect 17816 54742 18028 54748
rect 17816 54678 17958 54742
rect 18022 54678 18028 54742
rect 17816 54606 18028 54678
rect 17816 54542 17822 54606
rect 17886 54542 18028 54606
rect 17816 54536 18028 54542
rect 18224 54672 18572 54748
rect 18224 54612 18436 54672
rect 18224 54606 18572 54612
rect 18224 54542 18366 54606
rect 18430 54542 18502 54606
rect 18566 54542 18572 54606
rect 18224 54536 18572 54542
rect 18632 54536 18980 54748
rect 19040 54808 19252 55156
rect 19448 54808 19660 55156
rect 19040 54748 19116 54808
rect 19584 54748 19660 54808
rect 19040 54400 19252 54748
rect 19448 54400 19660 54748
rect 24344 54742 24692 55292
rect 24344 54678 24622 54742
rect 24686 54678 24692 54742
rect 24344 54672 24692 54678
rect 66368 55150 66580 55292
rect 71264 55216 71476 55358
rect 71672 55422 71884 55428
rect 71672 55358 71814 55422
rect 71878 55358 71884 55422
rect 71672 55216 71884 55358
rect 72080 55286 72292 55564
rect 72488 55292 72700 55564
rect 72390 55286 72700 55292
rect 72080 55222 72222 55286
rect 72286 55222 72292 55286
rect 72352 55222 72358 55286
rect 72422 55222 72700 55286
rect 72080 55216 72292 55222
rect 72390 55216 72700 55222
rect 72896 55216 73108 55564
rect 71400 55156 71476 55216
rect 71808 55156 71884 55216
rect 73032 55156 73108 55216
rect 66368 55086 66510 55150
rect 66574 55086 66580 55150
rect 66368 54878 66580 55086
rect 66368 54814 66510 54878
rect 66574 54814 66580 54878
rect 66368 54742 66580 54814
rect 66368 54678 66510 54742
rect 66574 54678 66580 54742
rect 66368 54672 66580 54678
rect 71264 54808 71476 55156
rect 71672 54808 71884 55156
rect 72080 55014 72428 55020
rect 72080 54950 72222 55014
rect 72286 54950 72358 55014
rect 72422 54950 72428 55014
rect 72080 54944 72428 54950
rect 72080 54884 72292 54944
rect 72080 54808 72428 54884
rect 72488 54808 72700 55020
rect 72896 55014 73108 55156
rect 72896 54950 73038 55014
rect 73102 54950 73108 55014
rect 72896 54944 73108 54950
rect 71264 54748 71340 54808
rect 71808 54748 71884 54808
rect 72216 54748 72292 54808
rect 19176 54340 19252 54400
rect 19584 54340 19660 54400
rect 1632 54212 1844 54340
rect 1632 54204 1718 54212
rect 1224 54198 1718 54204
rect 1224 54134 1230 54198
rect 1294 54156 1718 54198
rect 1774 54156 1844 54212
rect 1294 54134 1844 54156
rect 1224 54128 1844 54134
rect 17816 54334 18028 54340
rect 17816 54270 17822 54334
rect 17886 54270 18028 54334
rect 17816 54198 18028 54270
rect 17816 54134 17958 54198
rect 18022 54134 18028 54198
rect 17816 54128 18028 54134
rect 18224 54334 18436 54340
rect 18534 54334 18980 54340
rect 18224 54270 18366 54334
rect 18430 54270 18436 54334
rect 18496 54270 18502 54334
rect 18566 54270 18980 54334
rect 18224 53992 18436 54270
rect 18534 54264 18980 54270
rect 18360 53932 18436 53992
rect 17816 53926 18028 53932
rect 17816 53862 17958 53926
rect 18022 53862 18028 53926
rect 17816 53790 18028 53862
rect 17816 53726 17822 53790
rect 17886 53726 18028 53790
rect 17816 53720 18028 53726
rect 18224 53720 18436 53932
rect 18632 53992 18980 54264
rect 19040 54198 19252 54340
rect 19040 54134 19182 54198
rect 19246 54134 19252 54198
rect 19040 54128 19252 54134
rect 19448 54198 19660 54340
rect 19448 54134 19454 54198
rect 19518 54134 19660 54198
rect 19448 54128 19660 54134
rect 24344 54470 24692 54476
rect 24344 54406 24622 54470
rect 24686 54406 24692 54470
rect 24344 54334 24692 54406
rect 24344 54270 24350 54334
rect 24414 54270 24692 54334
rect 24344 54128 24692 54270
rect 66368 54470 66580 54476
rect 66368 54406 66510 54470
rect 66574 54406 66580 54470
rect 66368 54128 66580 54406
rect 71264 54400 71476 54748
rect 71672 54400 71884 54748
rect 72080 54612 72292 54748
rect 72352 54748 72428 54808
rect 72624 54748 72700 54808
rect 72352 54672 72700 54748
rect 72080 54606 72428 54612
rect 72080 54542 72358 54606
rect 72422 54542 72428 54606
rect 72080 54536 72428 54542
rect 72488 54536 72700 54672
rect 72896 54742 73108 54748
rect 72896 54678 73038 54742
rect 73102 54678 73108 54742
rect 72896 54606 73108 54678
rect 72896 54542 72902 54606
rect 72966 54542 73108 54606
rect 72896 54536 73108 54542
rect 71400 54340 71476 54400
rect 71808 54340 71884 54400
rect 71264 54198 71476 54340
rect 71264 54134 71406 54198
rect 71470 54134 71476 54198
rect 71264 54128 71476 54134
rect 71672 54198 71884 54340
rect 71672 54134 71814 54198
rect 71878 54134 71884 54198
rect 71672 54128 71884 54134
rect 24480 54068 24556 54128
rect 66368 54068 66444 54128
rect 72080 54068 72292 54340
rect 72390 54334 72700 54340
rect 72352 54270 72358 54334
rect 72422 54270 72700 54334
rect 72390 54264 72700 54270
rect 24344 54062 24692 54068
rect 24344 53998 24350 54062
rect 24414 53998 24692 54062
rect 18632 53932 18708 53992
rect 18632 53720 18980 53932
rect 19040 53926 19252 53932
rect 19040 53862 19182 53926
rect 19246 53862 19252 53926
rect 19040 53790 19252 53862
rect 19040 53726 19182 53790
rect 19246 53726 19252 53790
rect 19040 53720 19252 53726
rect 19448 53926 19660 53932
rect 19448 53862 19454 53926
rect 19518 53862 19660 53926
rect 19448 53790 19660 53862
rect 24344 53856 24692 53998
rect 24616 53796 24692 53856
rect 19448 53726 19454 53790
rect 19518 53726 19660 53790
rect 19448 53720 19660 53726
rect 18632 53660 18708 53720
rect 18360 53584 18708 53660
rect 18360 53524 18436 53584
rect 17816 53518 18028 53524
rect 17816 53454 17822 53518
rect 17886 53454 18028 53518
rect 17816 53382 18028 53454
rect 17816 53318 17822 53382
rect 17886 53318 18028 53382
rect 17816 53312 18028 53318
rect 18224 53448 18980 53524
rect 18224 53388 18436 53448
rect 18224 53382 18572 53388
rect 18224 53318 18502 53382
rect 18566 53318 18572 53382
rect 18224 53312 18572 53318
rect 18632 53312 18980 53448
rect 19040 53518 19252 53524
rect 19040 53454 19182 53518
rect 19246 53454 19252 53518
rect 19040 53382 19252 53454
rect 19040 53318 19182 53382
rect 19246 53318 19252 53382
rect 19040 53312 19252 53318
rect 19448 53518 19660 53524
rect 19448 53454 19454 53518
rect 19518 53454 19660 53518
rect 19448 53382 19660 53454
rect 19448 53318 19454 53382
rect 19518 53318 19660 53382
rect 19448 53312 19660 53318
rect 24344 53312 24692 53796
rect 66368 53856 66580 54068
rect 72080 53992 72428 54068
rect 72488 53992 72700 54264
rect 72896 54334 73108 54340
rect 72896 54270 72902 54334
rect 72966 54270 73108 54334
rect 72896 54198 73108 54270
rect 72896 54134 73038 54198
rect 73102 54134 73108 54198
rect 72896 54128 73108 54134
rect 89080 54212 89428 54340
rect 89080 54156 89216 54212
rect 89272 54204 89428 54212
rect 89272 54198 89836 54204
rect 89272 54156 89766 54198
rect 89080 54134 89766 54156
rect 89830 54134 89836 54198
rect 89080 54128 89836 54134
rect 72216 53932 72292 53992
rect 71264 53926 71476 53932
rect 71264 53862 71406 53926
rect 71470 53862 71476 53926
rect 66368 53796 66444 53856
rect 66368 53312 66580 53796
rect 71264 53790 71476 53862
rect 71264 53726 71406 53790
rect 71470 53726 71476 53790
rect 71264 53720 71476 53726
rect 71672 53926 71884 53932
rect 71672 53862 71814 53926
rect 71878 53862 71884 53926
rect 71672 53790 71884 53862
rect 71672 53726 71678 53790
rect 71742 53726 71884 53790
rect 71672 53720 71884 53726
rect 72080 53790 72292 53932
rect 72352 53932 72428 53992
rect 72624 53932 72700 53992
rect 72352 53856 72700 53932
rect 72080 53726 72086 53790
rect 72150 53726 72292 53790
rect 72080 53720 72292 53726
rect 72488 53720 72700 53856
rect 72896 53926 73108 53932
rect 72896 53862 73038 53926
rect 73102 53862 73108 53926
rect 72896 53790 73108 53862
rect 72896 53726 73038 53790
rect 73102 53726 73108 53790
rect 72896 53720 73108 53726
rect 71264 53518 71476 53524
rect 71264 53454 71406 53518
rect 71470 53454 71476 53518
rect 71264 53382 71476 53454
rect 71264 53318 71406 53382
rect 71470 53318 71476 53382
rect 71264 53312 71476 53318
rect 71672 53518 71884 53524
rect 71672 53454 71678 53518
rect 71742 53454 71884 53518
rect 71672 53382 71884 53454
rect 71672 53318 71678 53382
rect 71742 53318 71884 53382
rect 71672 53312 71884 53318
rect 72080 53518 72292 53524
rect 72080 53454 72086 53518
rect 72150 53454 72292 53518
rect 72080 53382 72292 53454
rect 72488 53388 72700 53524
rect 72390 53382 72700 53388
rect 72080 53318 72086 53382
rect 72150 53318 72292 53382
rect 72352 53318 72358 53382
rect 72422 53318 72700 53382
rect 72080 53312 72292 53318
rect 72390 53312 72700 53318
rect 72896 53518 73108 53524
rect 72896 53454 73038 53518
rect 73102 53454 73108 53518
rect 72896 53382 73108 53454
rect 72896 53318 72902 53382
rect 72966 53318 73108 53382
rect 72896 53312 73108 53318
rect 24480 53252 24556 53312
rect 66368 53252 66444 53312
rect 17816 53110 18028 53116
rect 17816 53046 17822 53110
rect 17886 53046 18028 53110
rect 17816 52974 18028 53046
rect 17816 52910 17822 52974
rect 17886 52910 18028 52974
rect 17816 52904 18028 52910
rect 18224 52974 18436 53116
rect 18534 53110 18980 53116
rect 18496 53046 18502 53110
rect 18566 53046 18980 53110
rect 18534 53040 18980 53046
rect 18224 52910 18230 52974
rect 18294 52910 18436 52974
rect 18224 52904 18436 52910
rect 18632 52974 18980 53040
rect 18632 52910 18910 52974
rect 18974 52910 18980 52974
rect 18632 52904 18980 52910
rect 19040 53110 19252 53116
rect 19040 53046 19182 53110
rect 19246 53046 19252 53110
rect 19040 52974 19252 53046
rect 19040 52910 19046 52974
rect 19110 52910 19252 52974
rect 19040 52904 19252 52910
rect 19448 53110 19660 53116
rect 19448 53046 19454 53110
rect 19518 53046 19660 53110
rect 19448 52974 19660 53046
rect 24344 53040 24692 53252
rect 24616 52980 24692 53040
rect 19448 52910 19454 52974
rect 19518 52910 19660 52974
rect 19448 52904 19660 52910
rect 24344 52768 24692 52980
rect 66368 53040 66580 53252
rect 71264 53110 71476 53116
rect 71264 53046 71406 53110
rect 71470 53046 71476 53110
rect 66368 52980 66444 53040
rect 66368 52768 66580 52980
rect 71264 52974 71476 53046
rect 71264 52910 71270 52974
rect 71334 52910 71476 52974
rect 71264 52904 71476 52910
rect 71672 53110 71884 53116
rect 71672 53046 71678 53110
rect 71742 53046 71884 53110
rect 71672 52974 71884 53046
rect 71672 52910 71678 52974
rect 71742 52910 71884 52974
rect 71672 52904 71884 52910
rect 72080 53110 72428 53116
rect 72080 53046 72086 53110
rect 72150 53046 72358 53110
rect 72422 53046 72428 53110
rect 72080 53040 72428 53046
rect 72080 52974 72292 53040
rect 72080 52910 72222 52974
rect 72286 52910 72292 52974
rect 72080 52904 72292 52910
rect 72488 52904 72700 53116
rect 72896 53110 73108 53116
rect 72896 53046 72902 53110
rect 72966 53046 73108 53110
rect 72896 52974 73108 53046
rect 72896 52910 73038 52974
rect 73102 52910 73108 52974
rect 72896 52904 73108 52910
rect 72488 52844 72564 52904
rect 24344 52708 24420 52768
rect 66504 52708 66580 52768
rect 72216 52768 72564 52844
rect 72216 52708 72292 52768
rect 17816 52702 18028 52708
rect 17816 52638 17822 52702
rect 17886 52638 18028 52702
rect 1224 52566 1844 52572
rect 1224 52502 1230 52566
rect 1294 52532 1844 52566
rect 1294 52502 1718 52532
rect 1224 52496 1718 52502
rect 1632 52476 1718 52496
rect 1774 52476 1844 52532
rect 17816 52566 18028 52638
rect 17816 52502 17822 52566
rect 17886 52502 18028 52566
rect 17816 52496 18028 52502
rect 18224 52702 18436 52708
rect 18224 52638 18230 52702
rect 18294 52638 18436 52702
rect 18224 52566 18436 52638
rect 18632 52702 18980 52708
rect 18632 52638 18910 52702
rect 18974 52638 18980 52702
rect 18632 52572 18980 52638
rect 18534 52566 18980 52572
rect 18224 52502 18366 52566
rect 18430 52502 18436 52566
rect 18496 52502 18502 52566
rect 18566 52502 18980 52566
rect 18224 52496 18436 52502
rect 18534 52496 18980 52502
rect 19040 52702 19252 52708
rect 19040 52638 19046 52702
rect 19110 52638 19252 52702
rect 19040 52566 19252 52638
rect 19040 52502 19046 52566
rect 19110 52502 19252 52566
rect 19040 52496 19252 52502
rect 19448 52702 19660 52708
rect 19448 52638 19454 52702
rect 19518 52638 19660 52702
rect 19448 52566 19660 52638
rect 19448 52502 19590 52566
rect 19654 52502 19660 52566
rect 19448 52496 19660 52502
rect 24344 52496 24692 52708
rect 66368 52496 66580 52708
rect 71264 52702 71476 52708
rect 71264 52638 71270 52702
rect 71334 52638 71476 52702
rect 71264 52566 71476 52638
rect 71264 52502 71270 52566
rect 71334 52502 71476 52566
rect 71264 52496 71476 52502
rect 71672 52702 71884 52708
rect 71672 52638 71678 52702
rect 71742 52638 71884 52702
rect 71672 52566 71884 52638
rect 71672 52502 71678 52566
rect 71742 52502 71884 52566
rect 71672 52496 71884 52502
rect 72080 52702 72700 52708
rect 72080 52638 72222 52702
rect 72286 52638 72700 52702
rect 72080 52632 72700 52638
rect 72080 52566 72292 52632
rect 72080 52502 72086 52566
rect 72150 52502 72292 52566
rect 72080 52496 72292 52502
rect 72488 52566 72700 52632
rect 72488 52502 72630 52566
rect 72694 52502 72700 52566
rect 72488 52496 72700 52502
rect 72896 52702 73108 52708
rect 72896 52638 73038 52702
rect 73102 52638 73108 52702
rect 72896 52566 73108 52638
rect 72896 52502 72902 52566
rect 72966 52502 73108 52566
rect 72896 52496 73108 52502
rect 89080 52532 89428 52572
rect 1632 52360 1844 52476
rect 24344 52436 24420 52496
rect 66504 52436 66580 52496
rect 17816 52294 18028 52300
rect 17816 52230 17822 52294
rect 17886 52230 18028 52294
rect 17816 52088 18028 52230
rect 18224 52294 18572 52300
rect 18224 52230 18366 52294
rect 18430 52230 18502 52294
rect 18566 52230 18572 52294
rect 18224 52224 18572 52230
rect 18224 52164 18436 52224
rect 18632 52164 18980 52300
rect 18224 52158 18980 52164
rect 18224 52094 18910 52158
rect 18974 52094 18980 52158
rect 18224 52088 18980 52094
rect 19040 52294 19252 52300
rect 19040 52230 19046 52294
rect 19110 52230 19252 52294
rect 19040 52158 19252 52230
rect 19040 52094 19182 52158
rect 19246 52094 19252 52158
rect 19040 52088 19252 52094
rect 19448 52294 19660 52300
rect 19448 52230 19590 52294
rect 19654 52230 19660 52294
rect 19448 52158 19660 52230
rect 19448 52094 19454 52158
rect 19518 52094 19660 52158
rect 19448 52088 19660 52094
rect 24344 52224 24692 52436
rect 66368 52224 66580 52436
rect 89080 52476 89216 52532
rect 89272 52476 89428 52532
rect 89080 52436 89428 52476
rect 89080 52430 89836 52436
rect 89080 52366 89766 52430
rect 89830 52366 89836 52430
rect 89080 52360 89836 52366
rect 71264 52294 71476 52300
rect 71264 52230 71270 52294
rect 71334 52230 71476 52294
rect 24344 52164 24420 52224
rect 66368 52164 66444 52224
rect 17952 52028 18028 52088
rect 17816 51680 18028 52028
rect 24344 51952 24692 52164
rect 24616 51892 24692 51952
rect 18224 51886 18980 51892
rect 18224 51822 18910 51886
rect 18974 51822 18980 51886
rect 18224 51816 18980 51822
rect 18224 51680 18436 51816
rect 18632 51680 18980 51816
rect 19040 51886 19252 51892
rect 19040 51822 19182 51886
rect 19246 51822 19252 51886
rect 19040 51750 19252 51822
rect 19040 51686 19046 51750
rect 19110 51686 19252 51750
rect 19040 51680 19252 51686
rect 19448 51886 19660 51892
rect 19448 51822 19454 51886
rect 19518 51822 19660 51886
rect 19448 51750 19660 51822
rect 19448 51686 19590 51750
rect 19654 51686 19660 51750
rect 19448 51680 19660 51686
rect 17816 51620 17892 51680
rect 18632 51620 18708 51680
rect 17816 51272 18028 51620
rect 18224 51348 18436 51620
rect 18224 51342 18572 51348
rect 18224 51278 18502 51342
rect 18566 51278 18572 51342
rect 18224 51272 18572 51278
rect 18632 51272 18980 51620
rect 19040 51478 19252 51484
rect 19040 51414 19046 51478
rect 19110 51414 19252 51478
rect 19040 51342 19252 51414
rect 19040 51278 19182 51342
rect 19246 51278 19252 51342
rect 19040 51272 19252 51278
rect 19448 51478 19660 51484
rect 19448 51414 19590 51478
rect 19654 51414 19660 51478
rect 19448 51342 19660 51414
rect 24344 51408 24692 51892
rect 66368 51952 66580 52164
rect 71264 52158 71476 52230
rect 71264 52094 71270 52158
rect 71334 52094 71476 52158
rect 71264 52088 71476 52094
rect 71672 52294 71884 52300
rect 71672 52230 71678 52294
rect 71742 52230 71884 52294
rect 71672 52158 71884 52230
rect 71672 52094 71678 52158
rect 71742 52094 71884 52158
rect 71672 52088 71884 52094
rect 72080 52294 72292 52300
rect 72080 52230 72086 52294
rect 72150 52230 72292 52294
rect 72080 52088 72292 52230
rect 72488 52294 72700 52300
rect 72488 52230 72630 52294
rect 72694 52230 72700 52294
rect 72488 52164 72700 52230
rect 72390 52158 72700 52164
rect 72352 52094 72358 52158
rect 72422 52094 72700 52158
rect 72390 52088 72700 52094
rect 72896 52294 73108 52300
rect 72896 52230 72902 52294
rect 72966 52230 73108 52294
rect 72896 52088 73108 52230
rect 73032 52028 73108 52088
rect 66368 51892 66444 51952
rect 66368 51408 66580 51892
rect 71264 51886 71476 51892
rect 71264 51822 71270 51886
rect 71334 51822 71476 51886
rect 71264 51750 71476 51822
rect 71264 51686 71270 51750
rect 71334 51686 71476 51750
rect 71264 51680 71476 51686
rect 71672 51886 71884 51892
rect 71672 51822 71678 51886
rect 71742 51822 71884 51886
rect 71672 51750 71884 51822
rect 71672 51686 71678 51750
rect 71742 51686 71884 51750
rect 71672 51680 71884 51686
rect 72080 51886 72428 51892
rect 72080 51822 72358 51886
rect 72422 51822 72428 51886
rect 72080 51816 72428 51822
rect 72080 51756 72292 51816
rect 72080 51680 72428 51756
rect 72488 51750 72700 51892
rect 72488 51686 72494 51750
rect 72558 51686 72700 51750
rect 72488 51680 72700 51686
rect 72352 51620 72428 51680
rect 72624 51620 72700 51680
rect 72080 51484 72292 51620
rect 72352 51544 72700 51620
rect 24616 51348 24692 51408
rect 66504 51348 66580 51408
rect 19448 51278 19454 51342
rect 19518 51278 19660 51342
rect 19448 51272 19660 51278
rect 17952 51212 18028 51272
rect 18632 51212 18708 51272
rect 17816 51070 18028 51212
rect 18360 51136 18708 51212
rect 18942 51206 19524 51212
rect 18904 51142 18910 51206
rect 18974 51142 19524 51206
rect 18942 51136 19524 51142
rect 24344 51206 24692 51348
rect 24344 51142 24622 51206
rect 24686 51142 24692 51206
rect 24344 51136 24692 51142
rect 18360 51076 18436 51136
rect 19448 51076 19524 51136
rect 24616 51076 24692 51136
rect 17816 51006 17822 51070
rect 17886 51006 18028 51070
rect 17816 51000 18028 51006
rect 18224 50940 18436 51076
rect 18534 51070 18980 51076
rect 18496 51006 18502 51070
rect 18566 51006 18980 51070
rect 18534 51000 18980 51006
rect 1632 50852 1844 50940
rect 1632 50804 1718 50852
rect 1224 50798 1718 50804
rect 1224 50734 1230 50798
rect 1294 50796 1718 50798
rect 1774 50796 1844 50852
rect 18224 50864 18572 50940
rect 18632 50864 18980 51000
rect 19040 51070 19252 51076
rect 19040 51006 19182 51070
rect 19246 51006 19252 51070
rect 19040 50864 19252 51006
rect 18224 50804 18300 50864
rect 18496 50804 18572 50864
rect 18768 50804 18844 50864
rect 19176 50804 19252 50864
rect 1294 50734 1844 50796
rect 1224 50728 1844 50734
rect 17816 50798 18028 50804
rect 17816 50734 17822 50798
rect 17886 50734 18028 50798
rect 17816 50662 18028 50734
rect 17816 50598 17958 50662
rect 18022 50598 18028 50662
rect 17816 50592 18028 50598
rect 18224 50592 18436 50804
rect 18496 50798 18980 50804
rect 18496 50734 18910 50798
rect 18974 50734 18980 50798
rect 18496 50728 18980 50734
rect 18632 50662 18980 50728
rect 18632 50598 18638 50662
rect 18702 50598 18980 50662
rect 18632 50592 18980 50598
rect 19040 50456 19252 50804
rect 19448 51070 19660 51076
rect 19448 51006 19454 51070
rect 19518 51006 19660 51070
rect 19448 50864 19660 51006
rect 24344 50934 24692 51076
rect 24344 50870 24486 50934
rect 24550 50870 24622 50934
rect 24686 50870 24692 50934
rect 19448 50804 19524 50864
rect 19448 50456 19660 50804
rect 24344 50728 24692 50870
rect 66368 51206 66580 51348
rect 71264 51478 71476 51484
rect 71264 51414 71270 51478
rect 71334 51414 71476 51478
rect 71264 51342 71476 51414
rect 71264 51278 71406 51342
rect 71470 51278 71476 51342
rect 71264 51272 71476 51278
rect 71672 51478 71884 51484
rect 71672 51414 71678 51478
rect 71742 51414 71884 51478
rect 71672 51342 71884 51414
rect 71672 51278 71678 51342
rect 71742 51278 71884 51342
rect 71672 51272 71884 51278
rect 72080 51478 72428 51484
rect 72080 51414 72358 51478
rect 72422 51414 72428 51478
rect 72080 51408 72428 51414
rect 72080 51272 72292 51408
rect 72488 51342 72700 51544
rect 72488 51278 72494 51342
rect 72558 51278 72700 51342
rect 72488 51272 72700 51278
rect 72896 51680 73108 52028
rect 72896 51620 72972 51680
rect 72896 51272 73108 51620
rect 66368 51142 66374 51206
rect 66438 51142 66580 51206
rect 66368 51136 66580 51142
rect 72896 51212 72972 51272
rect 66368 51076 66444 51136
rect 66368 50934 66580 51076
rect 66368 50870 66374 50934
rect 66438 50870 66580 50934
rect 66368 50798 66580 50870
rect 71264 51070 71476 51076
rect 71264 51006 71406 51070
rect 71470 51006 71476 51070
rect 71264 50864 71476 51006
rect 71400 50804 71476 50864
rect 66368 50734 66374 50798
rect 66438 50734 66510 50798
rect 66574 50734 66580 50798
rect 66368 50728 66580 50734
rect 19040 50396 19116 50456
rect 19584 50396 19660 50456
rect 17816 50390 18028 50396
rect 17816 50326 17958 50390
rect 18022 50326 18028 50390
rect 17816 50254 18028 50326
rect 17816 50190 17958 50254
rect 18022 50190 18028 50254
rect 17816 50184 18028 50190
rect 18224 50260 18436 50396
rect 18632 50390 18980 50396
rect 18632 50326 18638 50390
rect 18702 50326 18980 50390
rect 18632 50260 18980 50326
rect 18224 50184 18980 50260
rect 18224 50124 18436 50184
rect 18224 50048 18572 50124
rect 18632 50048 18980 50184
rect 19040 50048 19252 50396
rect 19448 50048 19660 50396
rect 24344 50526 24692 50532
rect 24344 50462 24486 50526
rect 24550 50462 24692 50526
rect 24344 50320 24692 50462
rect 66368 50526 66580 50532
rect 66368 50462 66374 50526
rect 66438 50462 66580 50526
rect 66368 50390 66580 50462
rect 71264 50456 71476 50804
rect 71672 51070 71884 51076
rect 71672 51006 71678 51070
rect 71742 51006 71884 51070
rect 71672 50864 71884 51006
rect 72080 50864 72292 51076
rect 72488 51070 72700 51076
rect 72488 51006 72494 51070
rect 72558 51006 72700 51070
rect 72488 50940 72700 51006
rect 72896 51070 73108 51212
rect 72896 51006 72902 51070
rect 72966 51006 73108 51070
rect 72896 51000 73108 51006
rect 72352 50864 72700 50940
rect 71672 50804 71748 50864
rect 72080 50804 72156 50864
rect 72352 50804 72428 50864
rect 89080 50852 89428 50940
rect 71672 50456 71884 50804
rect 72080 50728 72428 50804
rect 72080 50668 72292 50728
rect 72080 50662 72428 50668
rect 72080 50598 72358 50662
rect 72422 50598 72428 50662
rect 72080 50592 72428 50598
rect 72488 50592 72700 50804
rect 72896 50798 73108 50804
rect 72896 50734 72902 50798
rect 72966 50734 73108 50798
rect 72896 50662 73108 50734
rect 89080 50796 89216 50852
rect 89272 50804 89428 50852
rect 89272 50798 89836 50804
rect 89272 50796 89766 50798
rect 89080 50734 89766 50796
rect 89830 50734 89836 50798
rect 89080 50728 89836 50734
rect 72896 50598 73038 50662
rect 73102 50598 73108 50662
rect 72896 50592 73108 50598
rect 72216 50532 72292 50592
rect 72488 50532 72564 50592
rect 72216 50456 72564 50532
rect 71400 50396 71476 50456
rect 71808 50396 71884 50456
rect 66368 50326 66510 50390
rect 66574 50326 66580 50390
rect 24470 50124 24568 50320
rect 18224 49988 18300 50048
rect 18496 49988 18572 50048
rect 19176 49988 19252 50048
rect 19584 49988 19660 50048
rect 17816 49982 18028 49988
rect 17816 49918 17958 49982
rect 18022 49918 18028 49982
rect 17816 49846 18028 49918
rect 17816 49782 17958 49846
rect 18022 49782 18028 49846
rect 17816 49776 18028 49782
rect 18224 49846 18436 49988
rect 18496 49912 18980 49988
rect 18224 49782 18230 49846
rect 18294 49782 18436 49846
rect 18224 49776 18436 49782
rect 18632 49846 18980 49912
rect 18632 49782 18774 49846
rect 18838 49782 18980 49846
rect 18632 49776 18980 49782
rect 19040 49846 19252 49988
rect 19040 49782 19182 49846
rect 19246 49782 19252 49846
rect 19040 49776 19252 49782
rect 19448 49846 19660 49988
rect 24344 49912 24692 50124
rect 66368 49912 66580 50326
rect 71264 50048 71476 50396
rect 71672 50048 71884 50396
rect 71400 49988 71476 50048
rect 71808 49988 71884 50048
rect 24480 49852 24556 49912
rect 66368 49852 66444 49912
rect 19448 49782 19590 49846
rect 19654 49782 19660 49846
rect 19448 49776 19660 49782
rect 17816 49574 18028 49580
rect 17816 49510 17958 49574
rect 18022 49510 18028 49574
rect 17816 49438 18028 49510
rect 17816 49374 17822 49438
rect 17886 49374 18028 49438
rect 17816 49368 18028 49374
rect 18224 49574 18436 49580
rect 18224 49510 18230 49574
rect 18294 49510 18436 49574
rect 18224 49368 18436 49510
rect 18632 49574 18980 49580
rect 18632 49510 18774 49574
rect 18838 49510 18980 49574
rect 18632 49438 18980 49510
rect 18632 49374 18774 49438
rect 18838 49374 18980 49438
rect 18632 49368 18980 49374
rect 19040 49574 19252 49580
rect 19040 49510 19182 49574
rect 19246 49510 19252 49574
rect 19040 49438 19252 49510
rect 19040 49374 19182 49438
rect 19246 49374 19252 49438
rect 19040 49368 19252 49374
rect 19448 49574 19660 49580
rect 19448 49510 19590 49574
rect 19654 49510 19660 49574
rect 19448 49438 19660 49510
rect 19448 49374 19454 49438
rect 19518 49374 19660 49438
rect 19448 49368 19660 49374
rect 24344 49368 24692 49852
rect 66368 49368 66580 49852
rect 71264 49846 71476 49988
rect 71264 49782 71270 49846
rect 71334 49782 71476 49846
rect 71264 49776 71476 49782
rect 71672 49846 71884 49988
rect 71672 49782 71678 49846
rect 71742 49782 71884 49846
rect 71672 49776 71884 49782
rect 72080 50048 72292 50396
rect 72390 50390 72700 50396
rect 72352 50326 72358 50390
rect 72422 50326 72700 50390
rect 72390 50320 72700 50326
rect 72488 50048 72700 50320
rect 72896 50390 73108 50396
rect 72896 50326 73038 50390
rect 73102 50326 73108 50390
rect 72896 50254 73108 50326
rect 72896 50190 72902 50254
rect 72966 50190 73108 50254
rect 72896 50184 73108 50190
rect 72080 49988 72156 50048
rect 72488 49988 72564 50048
rect 72080 49846 72292 49988
rect 72080 49782 72086 49846
rect 72150 49782 72292 49846
rect 72080 49776 72292 49782
rect 72488 49846 72700 49988
rect 72488 49782 72630 49846
rect 72694 49782 72700 49846
rect 72488 49776 72700 49782
rect 72896 49982 73108 49988
rect 72896 49918 72902 49982
rect 72966 49918 73108 49982
rect 72896 49846 73108 49918
rect 72896 49782 73038 49846
rect 73102 49782 73108 49846
rect 72896 49776 73108 49782
rect 71264 49574 71476 49580
rect 71264 49510 71270 49574
rect 71334 49510 71476 49574
rect 71264 49438 71476 49510
rect 71264 49374 71270 49438
rect 71334 49374 71476 49438
rect 71264 49368 71476 49374
rect 71672 49574 71884 49580
rect 71672 49510 71678 49574
rect 71742 49510 71884 49574
rect 71672 49438 71884 49510
rect 71672 49374 71678 49438
rect 71742 49374 71884 49438
rect 71672 49368 71884 49374
rect 72080 49574 72700 49580
rect 72080 49510 72086 49574
rect 72150 49510 72630 49574
rect 72694 49510 72700 49574
rect 72080 49504 72700 49510
rect 72080 49368 72292 49504
rect 72488 49438 72700 49504
rect 72488 49374 72630 49438
rect 72694 49374 72700 49438
rect 72488 49368 72700 49374
rect 72896 49574 73108 49580
rect 72896 49510 73038 49574
rect 73102 49510 73108 49574
rect 72896 49438 73108 49510
rect 72896 49374 73038 49438
rect 73102 49374 73108 49438
rect 72896 49368 73108 49374
rect 24480 49308 24556 49368
rect 66504 49308 66580 49368
rect 1632 49172 1844 49308
rect 1632 49116 1718 49172
rect 1774 49116 1844 49172
rect 1632 49036 1844 49116
rect 1224 49030 1844 49036
rect 1224 48966 1230 49030
rect 1294 48966 1844 49030
rect 1224 48960 1844 48966
rect 17816 49166 18028 49172
rect 17816 49102 17822 49166
rect 17886 49102 18028 49166
rect 17816 49030 18028 49102
rect 17816 48966 17958 49030
rect 18022 48966 18028 49030
rect 17816 48960 18028 48966
rect 18224 49166 18980 49172
rect 18224 49102 18774 49166
rect 18838 49102 18980 49166
rect 18224 49096 18980 49102
rect 18224 48960 18436 49096
rect 18632 49030 18980 49096
rect 18632 48966 18638 49030
rect 18702 48966 18980 49030
rect 18632 48960 18980 48966
rect 19040 49166 19252 49172
rect 19040 49102 19182 49166
rect 19246 49102 19252 49166
rect 19040 49030 19252 49102
rect 19040 48966 19182 49030
rect 19246 48966 19252 49030
rect 19040 48960 19252 48966
rect 19448 49166 19660 49172
rect 19448 49102 19454 49166
rect 19518 49102 19660 49166
rect 19448 49030 19660 49102
rect 24344 49096 24692 49308
rect 66368 49096 66580 49308
rect 89080 49172 89428 49308
rect 71264 49166 71476 49172
rect 71264 49102 71270 49166
rect 71334 49102 71476 49166
rect 24480 49036 24556 49096
rect 66368 49036 66444 49096
rect 19448 48966 19454 49030
rect 19518 48966 19660 49030
rect 19448 48960 19660 48966
rect 24344 48824 24692 49036
rect 24616 48764 24692 48824
rect 17816 48758 18028 48764
rect 17816 48694 17958 48758
rect 18022 48694 18028 48758
rect 17816 48622 18028 48694
rect 17816 48558 17822 48622
rect 17886 48558 18028 48622
rect 17816 48552 18028 48558
rect 18224 48622 18436 48764
rect 18224 48558 18230 48622
rect 18294 48558 18436 48622
rect 18224 48552 18436 48558
rect 18632 48758 18980 48764
rect 18632 48694 18638 48758
rect 18702 48694 18980 48758
rect 18632 48622 18980 48694
rect 18632 48558 18910 48622
rect 18974 48558 18980 48622
rect 18632 48552 18980 48558
rect 19040 48758 19252 48764
rect 19040 48694 19182 48758
rect 19246 48694 19252 48758
rect 19040 48622 19252 48694
rect 19040 48558 19046 48622
rect 19110 48558 19252 48622
rect 19040 48552 19252 48558
rect 19448 48758 19660 48764
rect 19448 48694 19454 48758
rect 19518 48694 19660 48758
rect 19448 48622 19660 48694
rect 19448 48558 19590 48622
rect 19654 48558 19660 48622
rect 19448 48552 19660 48558
rect 24344 48552 24692 48764
rect 66368 48824 66580 49036
rect 71264 49030 71476 49102
rect 71264 48966 71406 49030
rect 71470 48966 71476 49030
rect 71264 48960 71476 48966
rect 71672 49166 71884 49172
rect 71672 49102 71678 49166
rect 71742 49102 71884 49166
rect 71672 49030 71884 49102
rect 71672 48966 71814 49030
rect 71878 48966 71884 49030
rect 71672 48960 71884 48966
rect 72080 49030 72292 49172
rect 72080 48966 72086 49030
rect 72150 48966 72292 49030
rect 72080 48960 72292 48966
rect 72488 49166 72700 49172
rect 72488 49102 72630 49166
rect 72694 49102 72700 49166
rect 72488 49030 72700 49102
rect 72488 48966 72494 49030
rect 72558 48966 72700 49030
rect 72488 48960 72700 48966
rect 72896 49166 73108 49172
rect 72896 49102 73038 49166
rect 73102 49102 73108 49166
rect 72896 49030 73108 49102
rect 72896 48966 72902 49030
rect 72966 48966 73108 49030
rect 72896 48960 73108 48966
rect 89080 49116 89216 49172
rect 89272 49166 89836 49172
rect 89272 49116 89766 49166
rect 89080 49102 89766 49116
rect 89830 49102 89836 49166
rect 89080 49096 89836 49102
rect 89080 48960 89428 49096
rect 66368 48764 66444 48824
rect 66368 48552 66580 48764
rect 71264 48758 71476 48764
rect 71264 48694 71406 48758
rect 71470 48694 71476 48758
rect 71264 48622 71476 48694
rect 71264 48558 71270 48622
rect 71334 48558 71476 48622
rect 71264 48552 71476 48558
rect 71672 48758 71884 48764
rect 71672 48694 71814 48758
rect 71878 48694 71884 48758
rect 71672 48622 71884 48694
rect 71672 48558 71678 48622
rect 71742 48558 71884 48622
rect 71672 48552 71884 48558
rect 72080 48758 72292 48764
rect 72080 48694 72086 48758
rect 72150 48694 72292 48758
rect 72080 48628 72292 48694
rect 72488 48758 72700 48764
rect 72488 48694 72494 48758
rect 72558 48694 72700 48758
rect 72488 48628 72700 48694
rect 72080 48622 72700 48628
rect 72080 48558 72222 48622
rect 72286 48558 72700 48622
rect 72080 48552 72700 48558
rect 72896 48758 73108 48764
rect 72896 48694 72902 48758
rect 72966 48694 73108 48758
rect 72896 48622 73108 48694
rect 72896 48558 73038 48622
rect 73102 48558 73108 48622
rect 72896 48552 73108 48558
rect 24480 48492 24556 48552
rect 66504 48492 66580 48552
rect 17816 48350 18028 48356
rect 17816 48286 17822 48350
rect 17886 48286 18028 48350
rect 17816 48144 18028 48286
rect 18224 48350 18436 48356
rect 18224 48286 18230 48350
rect 18294 48286 18436 48350
rect 18224 48214 18436 48286
rect 18224 48150 18230 48214
rect 18294 48150 18436 48214
rect 18224 48144 18436 48150
rect 18632 48350 18980 48356
rect 18632 48286 18910 48350
rect 18974 48286 18980 48350
rect 18632 48144 18980 48286
rect 19040 48350 19252 48356
rect 19040 48286 19046 48350
rect 19110 48286 19252 48350
rect 19040 48214 19252 48286
rect 19040 48150 19046 48214
rect 19110 48150 19252 48214
rect 19040 48144 19252 48150
rect 19448 48350 19660 48356
rect 19448 48286 19590 48350
rect 19654 48286 19660 48350
rect 19448 48214 19660 48286
rect 19448 48150 19454 48214
rect 19518 48150 19660 48214
rect 19448 48144 19660 48150
rect 24344 48280 24692 48492
rect 66368 48280 66580 48492
rect 72216 48492 72292 48552
rect 72216 48416 72564 48492
rect 72488 48356 72564 48416
rect 24344 48220 24420 48280
rect 66504 48220 66580 48280
rect 17952 48084 18028 48144
rect 18632 48084 18708 48144
rect 17816 47736 18028 48084
rect 18360 48008 18708 48084
rect 24344 48008 24692 48220
rect 18360 47948 18436 48008
rect 24616 47948 24692 48008
rect 17952 47676 18028 47736
rect 1632 47492 1844 47540
rect 1632 47436 1718 47492
rect 1774 47436 1844 47492
rect 1632 47404 1844 47436
rect 1224 47398 1844 47404
rect 1224 47334 1230 47398
rect 1294 47334 1844 47398
rect 1224 47328 1844 47334
rect 17816 47328 18028 47676
rect 18224 47942 18980 47948
rect 18224 47878 18230 47942
rect 18294 47878 18980 47942
rect 18224 47872 18980 47878
rect 18224 47736 18436 47872
rect 18632 47736 18980 47872
rect 19040 47942 19252 47948
rect 19040 47878 19046 47942
rect 19110 47878 19252 47942
rect 19040 47806 19252 47878
rect 19040 47742 19182 47806
rect 19246 47742 19252 47806
rect 19040 47736 19252 47742
rect 19448 47942 19660 47948
rect 19448 47878 19454 47942
rect 19518 47878 19660 47942
rect 19448 47806 19660 47878
rect 19448 47742 19454 47806
rect 19518 47742 19660 47806
rect 19448 47736 19660 47742
rect 24344 47736 24692 47948
rect 66368 48008 66580 48220
rect 71264 48350 71476 48356
rect 71264 48286 71270 48350
rect 71334 48286 71476 48350
rect 71264 48214 71476 48286
rect 71264 48150 71270 48214
rect 71334 48150 71476 48214
rect 71264 48144 71476 48150
rect 71672 48350 71884 48356
rect 71672 48286 71678 48350
rect 71742 48286 71884 48350
rect 71672 48214 71884 48286
rect 71672 48150 71814 48214
rect 71878 48150 71884 48214
rect 71672 48144 71884 48150
rect 72080 48350 72292 48356
rect 72080 48286 72222 48350
rect 72286 48286 72292 48350
rect 72080 48214 72292 48286
rect 72080 48150 72086 48214
rect 72150 48150 72292 48214
rect 72080 48144 72292 48150
rect 72488 48144 72700 48356
rect 72896 48350 73108 48356
rect 72896 48286 73038 48350
rect 73102 48286 73108 48350
rect 72896 48144 73108 48286
rect 72896 48084 72972 48144
rect 66368 47948 66444 48008
rect 66368 47736 66580 47948
rect 71264 47942 71476 47948
rect 71264 47878 71270 47942
rect 71334 47878 71476 47942
rect 71264 47806 71476 47878
rect 71264 47742 71270 47806
rect 71334 47742 71476 47806
rect 71264 47736 71476 47742
rect 71672 47942 71884 47948
rect 71672 47878 71814 47942
rect 71878 47878 71884 47942
rect 71672 47806 71884 47878
rect 71672 47742 71814 47806
rect 71878 47742 71884 47806
rect 71672 47736 71884 47742
rect 72080 47942 72292 47948
rect 72080 47878 72086 47942
rect 72150 47878 72292 47942
rect 72080 47736 72292 47878
rect 72488 47736 72700 47948
rect 72896 47736 73108 48084
rect 18224 47676 18300 47736
rect 18632 47676 18708 47736
rect 24344 47676 24420 47736
rect 66368 47676 66444 47736
rect 72080 47676 72156 47736
rect 72488 47676 72564 47736
rect 72896 47676 72972 47736
rect 18224 47328 18436 47676
rect 18632 47600 18980 47676
rect 18752 47404 18850 47600
rect 19040 47534 19252 47540
rect 19040 47470 19182 47534
rect 19246 47470 19252 47534
rect 18632 47398 18980 47404
rect 18632 47334 18910 47398
rect 18974 47334 18980 47398
rect 18632 47328 18980 47334
rect 19040 47398 19252 47470
rect 19040 47334 19046 47398
rect 19110 47334 19252 47398
rect 19040 47328 19252 47334
rect 19448 47534 19660 47540
rect 19448 47470 19454 47534
rect 19518 47470 19660 47534
rect 19448 47398 19660 47470
rect 24344 47464 24692 47676
rect 66368 47464 66580 47676
rect 24480 47404 24556 47464
rect 66504 47404 66580 47464
rect 19448 47334 19590 47398
rect 19654 47334 19660 47398
rect 19448 47328 19660 47334
rect 17952 47268 18028 47328
rect 17816 47126 18028 47268
rect 24344 47192 24692 47404
rect 66368 47192 66580 47404
rect 71264 47534 71476 47540
rect 71264 47470 71270 47534
rect 71334 47470 71476 47534
rect 71264 47398 71476 47470
rect 71264 47334 71270 47398
rect 71334 47334 71476 47398
rect 71264 47328 71476 47334
rect 71672 47534 71884 47540
rect 71672 47470 71814 47534
rect 71878 47470 71884 47534
rect 71672 47398 71884 47470
rect 71672 47334 71814 47398
rect 71878 47334 71884 47398
rect 71672 47328 71884 47334
rect 72080 47404 72292 47676
rect 72488 47404 72700 47676
rect 72080 47398 72700 47404
rect 72080 47334 72222 47398
rect 72286 47334 72700 47398
rect 72080 47328 72700 47334
rect 72896 47328 73108 47676
rect 89080 47492 89428 47540
rect 89080 47436 89216 47492
rect 89272 47436 89428 47492
rect 89080 47404 89428 47436
rect 89080 47398 89836 47404
rect 89080 47334 89766 47398
rect 89830 47334 89836 47398
rect 89080 47328 89836 47334
rect 73032 47268 73108 47328
rect 24344 47132 24420 47192
rect 66504 47132 66580 47192
rect 17816 47062 17958 47126
rect 18022 47062 18028 47126
rect 17816 47056 18028 47062
rect 18224 46920 18436 47132
rect 18632 47126 18980 47132
rect 18632 47062 18910 47126
rect 18974 47062 18980 47126
rect 18632 46996 18980 47062
rect 18534 46990 18980 46996
rect 18496 46926 18502 46990
rect 18566 46926 18980 46990
rect 18534 46920 18980 46926
rect 19040 47126 19252 47132
rect 19040 47062 19046 47126
rect 19110 47062 19252 47126
rect 19040 46920 19252 47062
rect 19448 47126 19660 47132
rect 19448 47062 19590 47126
rect 19654 47062 19660 47126
rect 19448 46920 19660 47062
rect 18360 46860 18436 46920
rect 19040 46860 19116 46920
rect 19448 46860 19524 46920
rect 17816 46854 18028 46860
rect 17816 46790 17958 46854
rect 18022 46790 18028 46854
rect 17816 46718 18028 46790
rect 17816 46654 17822 46718
rect 17886 46654 18028 46718
rect 17816 46648 18028 46654
rect 18224 46784 18980 46860
rect 18224 46724 18436 46784
rect 18224 46718 18572 46724
rect 18224 46654 18502 46718
rect 18566 46654 18572 46718
rect 18224 46648 18572 46654
rect 18632 46718 18980 46784
rect 18632 46654 18774 46718
rect 18838 46654 18980 46718
rect 18632 46648 18980 46654
rect 19040 46512 19252 46860
rect 19448 46512 19660 46860
rect 24344 46854 24692 47132
rect 24344 46790 24486 46854
rect 24550 46790 24692 46854
rect 24344 46784 24692 46790
rect 66368 46854 66580 47132
rect 71264 47126 71476 47132
rect 71264 47062 71270 47126
rect 71334 47062 71476 47126
rect 71264 46920 71476 47062
rect 71400 46860 71476 46920
rect 66368 46790 66374 46854
rect 66438 46790 66580 46854
rect 66368 46784 66580 46790
rect 24344 46582 24692 46588
rect 24344 46518 24486 46582
rect 24550 46518 24692 46582
rect 19040 46452 19116 46512
rect 19448 46452 19524 46512
rect 17816 46446 18028 46452
rect 17816 46382 17822 46446
rect 17886 46382 18028 46446
rect 17816 46310 18028 46382
rect 17816 46246 17958 46310
rect 18022 46246 18028 46310
rect 17816 46240 18028 46246
rect 18224 46104 18436 46452
rect 18632 46446 18980 46452
rect 18632 46382 18774 46446
rect 18838 46382 18980 46446
rect 18632 46104 18980 46382
rect 18360 46044 18436 46104
rect 18904 46044 18980 46104
rect 17816 46038 18028 46044
rect 17816 45974 17958 46038
rect 18022 45974 18028 46038
rect 1632 45812 1844 45908
rect 17816 45902 18028 45974
rect 17816 45838 17958 45902
rect 18022 45838 18028 45902
rect 17816 45832 18028 45838
rect 18224 45902 18436 46044
rect 18632 45908 18980 46044
rect 18534 45902 18980 45908
rect 18224 45838 18366 45902
rect 18430 45838 18436 45902
rect 18496 45838 18502 45902
rect 18566 45838 18980 45902
rect 18224 45832 18436 45838
rect 18534 45832 18980 45838
rect 19040 46104 19252 46452
rect 19448 46104 19660 46452
rect 24344 46180 24692 46518
rect 22886 46174 24692 46180
rect 22848 46110 22854 46174
rect 22918 46110 24486 46174
rect 24550 46110 24692 46174
rect 22886 46104 24692 46110
rect 19040 46044 19116 46104
rect 19584 46044 19660 46104
rect 19040 45902 19252 46044
rect 19040 45838 19182 45902
rect 19246 45838 19252 45902
rect 19040 45832 19252 45838
rect 19448 45902 19660 46044
rect 24344 45968 24692 46104
rect 66368 46582 66580 46588
rect 66368 46518 66374 46582
rect 66438 46518 66580 46582
rect 66368 46446 66580 46518
rect 66368 46382 66510 46446
rect 66574 46382 66580 46446
rect 66368 46174 66580 46382
rect 66368 46110 66510 46174
rect 66574 46110 66580 46174
rect 66368 46044 66580 46110
rect 71264 46512 71476 46860
rect 71672 47126 71884 47132
rect 71672 47062 71814 47126
rect 71878 47062 71884 47126
rect 71672 46920 71884 47062
rect 72080 47126 72700 47132
rect 72080 47062 72222 47126
rect 72286 47062 72700 47126
rect 72080 47056 72700 47062
rect 72896 47126 73108 47268
rect 72896 47062 72902 47126
rect 72966 47062 73108 47126
rect 72896 47056 73108 47062
rect 72080 46920 72292 47056
rect 72488 46920 72700 47056
rect 71672 46860 71748 46920
rect 72080 46860 72156 46920
rect 72488 46860 72564 46920
rect 71672 46512 71884 46860
rect 72080 46648 72292 46860
rect 72488 46718 72700 46860
rect 72488 46654 72494 46718
rect 72558 46654 72700 46718
rect 72488 46648 72700 46654
rect 72896 46854 73108 46860
rect 72896 46790 72902 46854
rect 72966 46790 73108 46854
rect 72896 46718 73108 46790
rect 72896 46654 72902 46718
rect 72966 46654 73108 46718
rect 72896 46648 73108 46654
rect 71264 46452 71340 46512
rect 71672 46452 71748 46512
rect 71264 46104 71476 46452
rect 71672 46104 71884 46452
rect 72080 46104 72292 46452
rect 71400 46044 71476 46104
rect 71808 46044 71884 46104
rect 72216 46044 72292 46104
rect 66368 46038 69436 46044
rect 66368 45974 69366 46038
rect 69430 45974 69436 46038
rect 66368 45968 69436 45974
rect 66504 45908 66580 45968
rect 19448 45838 19454 45902
rect 19518 45838 19660 45902
rect 19448 45832 19660 45838
rect 24344 45902 24692 45908
rect 24344 45838 24486 45902
rect 24550 45838 24692 45902
rect 1632 45772 1718 45812
rect 1224 45766 1718 45772
rect 1224 45702 1230 45766
rect 1294 45756 1718 45766
rect 1774 45756 1844 45812
rect 1294 45702 1844 45756
rect 1224 45696 1844 45702
rect 19312 45696 19932 45772
rect 19312 45636 19388 45696
rect 19856 45636 19932 45696
rect 20128 45696 21428 45772
rect 20128 45636 20204 45696
rect 21352 45636 21428 45696
rect 17816 45630 18028 45636
rect 17816 45566 17958 45630
rect 18022 45566 18028 45630
rect 17816 45494 18028 45566
rect 17816 45430 17958 45494
rect 18022 45430 18028 45494
rect 17816 45424 18028 45430
rect 18224 45630 18572 45636
rect 18224 45566 18366 45630
rect 18430 45566 18502 45630
rect 18566 45566 18572 45630
rect 18224 45560 18572 45566
rect 18224 45500 18436 45560
rect 18632 45500 18980 45636
rect 18224 45424 18980 45500
rect 19040 45630 19388 45636
rect 19040 45566 19182 45630
rect 19246 45566 19388 45630
rect 19040 45560 19388 45566
rect 19448 45630 19660 45636
rect 19448 45566 19454 45630
rect 19518 45566 19660 45630
rect 19040 45494 19252 45560
rect 19040 45430 19046 45494
rect 19110 45430 19252 45494
rect 19040 45424 19252 45430
rect 19448 45500 19660 45566
rect 19856 45560 20204 45636
rect 19448 45494 19796 45500
rect 19448 45430 19454 45494
rect 19518 45430 19796 45494
rect 19448 45424 19796 45430
rect 19856 45424 20068 45560
rect 20264 45500 20612 45636
rect 21352 45630 22924 45636
rect 21352 45566 22854 45630
rect 22918 45566 22924 45630
rect 21352 45560 22924 45566
rect 20264 45424 21292 45500
rect 21352 45424 21564 45560
rect 22984 45424 23196 45636
rect 24344 45630 24692 45838
rect 24344 45566 24350 45630
rect 24414 45566 24692 45630
rect 24344 45424 24692 45566
rect 66368 45424 66580 45908
rect 71264 45902 71476 46044
rect 71264 45838 71406 45902
rect 71470 45838 71476 45902
rect 71264 45832 71476 45838
rect 71672 45902 71884 46044
rect 71672 45838 71678 45902
rect 71742 45838 71884 45902
rect 71672 45832 71884 45838
rect 72080 45902 72292 46044
rect 72080 45838 72086 45902
rect 72150 45838 72292 45902
rect 72080 45832 72292 45838
rect 72488 46446 72700 46452
rect 72488 46382 72494 46446
rect 72558 46382 72700 46446
rect 72488 46104 72700 46382
rect 72896 46446 73108 46452
rect 72896 46382 72902 46446
rect 72966 46382 73108 46446
rect 72896 46310 73108 46382
rect 72896 46246 73038 46310
rect 73102 46246 73108 46310
rect 72896 46240 73108 46246
rect 72488 46044 72564 46104
rect 72488 45902 72700 46044
rect 72488 45838 72494 45902
rect 72558 45838 72700 45902
rect 72488 45832 72700 45838
rect 72896 46038 73108 46044
rect 72896 45974 73038 46038
rect 73102 45974 73108 46038
rect 72896 45902 73108 45974
rect 72896 45838 72902 45902
rect 72966 45838 73108 45902
rect 72896 45832 73108 45838
rect 89080 45812 89428 45908
rect 69224 45696 70524 45772
rect 89080 45756 89216 45812
rect 89272 45772 89428 45812
rect 89272 45766 89836 45772
rect 89272 45756 89766 45766
rect 89080 45702 89766 45756
rect 89830 45702 89836 45766
rect 89080 45696 89836 45702
rect 69224 45636 69300 45696
rect 70448 45636 70524 45696
rect 67728 45560 69300 45636
rect 69360 45630 69572 45636
rect 69360 45566 69366 45630
rect 69430 45566 69572 45630
rect 67728 45424 67940 45560
rect 69360 45500 69572 45566
rect 70448 45500 70660 45636
rect 70856 45500 71068 45636
rect 71264 45630 71476 45636
rect 71264 45566 71406 45630
rect 71470 45566 71476 45630
rect 69360 45424 70388 45500
rect 70448 45494 70796 45500
rect 70448 45430 70726 45494
rect 70790 45430 70796 45494
rect 70448 45424 70796 45430
rect 70856 45424 71204 45500
rect 71264 45494 71476 45566
rect 71264 45430 71270 45494
rect 71334 45430 71476 45494
rect 71264 45424 71476 45430
rect 71672 45630 71884 45636
rect 71672 45566 71678 45630
rect 71742 45566 71884 45630
rect 71672 45494 71884 45566
rect 71672 45430 71678 45494
rect 71742 45430 71884 45494
rect 71672 45424 71884 45430
rect 72080 45630 72292 45636
rect 72080 45566 72086 45630
rect 72150 45566 72292 45630
rect 72080 45494 72292 45566
rect 72488 45630 72700 45636
rect 72488 45566 72494 45630
rect 72558 45566 72700 45630
rect 72488 45500 72700 45566
rect 72390 45494 72700 45500
rect 72080 45430 72222 45494
rect 72286 45430 72292 45494
rect 72352 45430 72358 45494
rect 72422 45430 72700 45494
rect 72080 45424 72292 45430
rect 72390 45424 72700 45430
rect 72896 45630 73108 45636
rect 72896 45566 72902 45630
rect 72966 45566 73108 45630
rect 72896 45494 73108 45566
rect 72896 45430 73038 45494
rect 73102 45430 73108 45494
rect 72896 45424 73108 45430
rect 18632 45364 18708 45424
rect 18496 45288 18708 45364
rect 19720 45364 19796 45424
rect 20264 45364 20340 45424
rect 19720 45288 20340 45364
rect 21216 45364 21292 45424
rect 22984 45364 23060 45424
rect 24480 45364 24556 45424
rect 66368 45364 66444 45424
rect 70312 45364 70388 45424
rect 70856 45364 70932 45424
rect 21216 45288 23060 45364
rect 24344 45358 24692 45364
rect 24344 45294 24350 45358
rect 24414 45294 24692 45358
rect 18496 45228 18572 45288
rect 17816 45222 18028 45228
rect 17816 45158 17958 45222
rect 18022 45158 18028 45222
rect 17816 45086 18028 45158
rect 17816 45022 17822 45086
rect 17886 45022 18028 45086
rect 17816 45016 18028 45022
rect 18224 45152 18572 45228
rect 18224 45086 18436 45152
rect 18224 45022 18366 45086
rect 18430 45022 18436 45086
rect 18224 45016 18436 45022
rect 18632 45016 18980 45228
rect 19040 45222 19252 45228
rect 19040 45158 19046 45222
rect 19110 45158 19252 45222
rect 19040 45086 19252 45158
rect 19040 45022 19046 45086
rect 19110 45022 19252 45086
rect 19040 45016 19252 45022
rect 19448 45222 19660 45228
rect 19448 45158 19454 45222
rect 19518 45158 19660 45222
rect 19448 45086 19660 45158
rect 24344 45152 24692 45294
rect 66368 45152 66580 45364
rect 70312 45288 70932 45364
rect 71128 45364 71204 45424
rect 71672 45364 71748 45424
rect 71128 45288 71748 45364
rect 70758 45222 71476 45228
rect 70720 45158 70726 45222
rect 70790 45158 71270 45222
rect 71334 45158 71476 45222
rect 70758 45152 71476 45158
rect 24616 45092 24692 45152
rect 66504 45092 66580 45152
rect 19448 45022 19454 45086
rect 19518 45022 19660 45086
rect 19448 45016 19660 45022
rect 18632 44956 18708 45016
rect 18360 44880 18708 44956
rect 24344 44880 24692 45092
rect 66368 44880 66580 45092
rect 71264 45086 71476 45152
rect 71264 45022 71270 45086
rect 71334 45022 71476 45086
rect 71264 45016 71476 45022
rect 71672 45222 71884 45228
rect 71672 45158 71678 45222
rect 71742 45158 71884 45222
rect 71672 45086 71884 45158
rect 71672 45022 71678 45086
rect 71742 45022 71884 45086
rect 71672 45016 71884 45022
rect 72080 45222 72428 45228
rect 72080 45158 72222 45222
rect 72286 45158 72358 45222
rect 72422 45158 72428 45222
rect 72080 45152 72428 45158
rect 72080 45092 72292 45152
rect 72488 45092 72700 45228
rect 72080 45086 72700 45092
rect 72080 45022 72494 45086
rect 72558 45022 72700 45086
rect 72080 45016 72700 45022
rect 72896 45222 73108 45228
rect 72896 45158 73038 45222
rect 73102 45158 73108 45222
rect 72896 45086 73108 45158
rect 72896 45022 73038 45086
rect 73102 45022 73108 45086
rect 72896 45016 73108 45022
rect 18360 44820 18436 44880
rect 24480 44820 24556 44880
rect 66368 44820 66444 44880
rect 17816 44814 18028 44820
rect 17816 44750 17822 44814
rect 17886 44750 18028 44814
rect 17816 44678 18028 44750
rect 17816 44614 17822 44678
rect 17886 44614 18028 44678
rect 17816 44608 18028 44614
rect 18224 44814 18980 44820
rect 18224 44750 18366 44814
rect 18430 44750 18980 44814
rect 18224 44744 18980 44750
rect 18224 44608 18436 44744
rect 18632 44678 18980 44744
rect 18632 44614 18638 44678
rect 18702 44614 18980 44678
rect 18632 44608 18980 44614
rect 19040 44814 19252 44820
rect 19040 44750 19046 44814
rect 19110 44750 19252 44814
rect 19040 44678 19252 44750
rect 19040 44614 19182 44678
rect 19246 44614 19252 44678
rect 19040 44608 19252 44614
rect 19448 44814 19660 44820
rect 19448 44750 19454 44814
rect 19518 44750 19660 44814
rect 19448 44678 19660 44750
rect 19448 44614 19590 44678
rect 19654 44614 19660 44678
rect 19448 44608 19660 44614
rect 24344 44608 24692 44820
rect 66368 44608 66580 44820
rect 71264 44814 71476 44820
rect 71264 44750 71270 44814
rect 71334 44750 71476 44814
rect 71264 44678 71476 44750
rect 71264 44614 71406 44678
rect 71470 44614 71476 44678
rect 71264 44608 71476 44614
rect 71672 44814 71884 44820
rect 71672 44750 71678 44814
rect 71742 44750 71884 44814
rect 71672 44678 71884 44750
rect 71672 44614 71814 44678
rect 71878 44614 71884 44678
rect 71672 44608 71884 44614
rect 72080 44678 72292 44820
rect 72488 44814 72700 44820
rect 72488 44750 72494 44814
rect 72558 44750 72700 44814
rect 72488 44684 72700 44750
rect 72390 44678 72700 44684
rect 72080 44614 72086 44678
rect 72150 44614 72292 44678
rect 72352 44614 72358 44678
rect 72422 44614 72700 44678
rect 72080 44608 72292 44614
rect 72390 44608 72700 44614
rect 72896 44814 73108 44820
rect 72896 44750 73038 44814
rect 73102 44750 73108 44814
rect 72896 44678 73108 44750
rect 72896 44614 72902 44678
rect 72966 44614 73108 44678
rect 72896 44608 73108 44614
rect 24480 44548 24556 44608
rect 66368 44548 66444 44608
rect 17816 44406 18028 44412
rect 17816 44342 17822 44406
rect 17886 44342 18028 44406
rect 1224 44270 1844 44276
rect 1224 44206 1230 44270
rect 1294 44206 1844 44270
rect 1224 44200 1844 44206
rect 1632 44132 1844 44200
rect 1632 44076 1718 44132
rect 1774 44076 1844 44132
rect 1632 43928 1844 44076
rect 17816 44200 18028 44342
rect 18224 44270 18436 44412
rect 18224 44206 18230 44270
rect 18294 44206 18436 44270
rect 18224 44200 18436 44206
rect 18632 44406 18980 44412
rect 18632 44342 18638 44406
rect 18702 44342 18980 44406
rect 18632 44270 18980 44342
rect 18632 44206 18910 44270
rect 18974 44206 18980 44270
rect 18632 44200 18980 44206
rect 19040 44406 19252 44412
rect 19040 44342 19182 44406
rect 19246 44342 19252 44406
rect 19040 44270 19252 44342
rect 19040 44206 19046 44270
rect 19110 44206 19252 44270
rect 19040 44200 19252 44206
rect 19448 44406 19660 44412
rect 19448 44342 19590 44406
rect 19654 44342 19660 44406
rect 19448 44270 19660 44342
rect 24344 44336 24692 44548
rect 24616 44276 24692 44336
rect 19448 44206 19590 44270
rect 19654 44206 19660 44270
rect 19448 44200 19660 44206
rect 17816 44140 17892 44200
rect 17816 43862 18028 44140
rect 24344 44064 24692 44276
rect 66368 44336 66580 44548
rect 71264 44406 71476 44412
rect 71264 44342 71406 44406
rect 71470 44342 71476 44406
rect 66368 44276 66444 44336
rect 66368 44064 66580 44276
rect 71264 44270 71476 44342
rect 71264 44206 71270 44270
rect 71334 44206 71476 44270
rect 71264 44200 71476 44206
rect 71672 44406 71884 44412
rect 71672 44342 71814 44406
rect 71878 44342 71884 44406
rect 71672 44270 71884 44342
rect 71672 44206 71678 44270
rect 71742 44206 71884 44270
rect 71672 44200 71884 44206
rect 72080 44406 72428 44412
rect 72080 44342 72086 44406
rect 72150 44342 72358 44406
rect 72422 44342 72428 44406
rect 72080 44336 72428 44342
rect 72080 44270 72292 44336
rect 72080 44206 72222 44270
rect 72286 44206 72292 44270
rect 72080 44200 72292 44206
rect 72488 44200 72700 44412
rect 72896 44406 73108 44412
rect 72896 44342 72902 44406
rect 72966 44342 73108 44406
rect 72896 44200 73108 44342
rect 72488 44140 72564 44200
rect 73032 44140 73108 44200
rect 24344 44004 24420 44064
rect 66504 44004 66580 44064
rect 72216 44064 72564 44140
rect 72216 44004 72292 44064
rect 17816 43798 17958 43862
rect 18022 43798 18028 43862
rect 17816 43792 18028 43798
rect 18224 43998 18436 44004
rect 18224 43934 18230 43998
rect 18294 43934 18436 43998
rect 18224 43862 18436 43934
rect 18224 43798 18366 43862
rect 18430 43798 18436 43862
rect 18224 43792 18436 43798
rect 18632 43998 18980 44004
rect 18632 43934 18910 43998
rect 18974 43934 18980 43998
rect 18632 43792 18980 43934
rect 19040 43998 19252 44004
rect 19040 43934 19046 43998
rect 19110 43934 19252 43998
rect 19040 43862 19252 43934
rect 19040 43798 19046 43862
rect 19110 43798 19252 43862
rect 19040 43792 19252 43798
rect 19448 43998 19660 44004
rect 19448 43934 19590 43998
rect 19654 43934 19660 43998
rect 19448 43862 19660 43934
rect 19448 43798 19590 43862
rect 19654 43798 19660 43862
rect 19448 43792 19660 43798
rect 24344 43792 24692 44004
rect 66368 43792 66580 44004
rect 71264 43998 71476 44004
rect 71264 43934 71270 43998
rect 71334 43934 71476 43998
rect 71264 43862 71476 43934
rect 71264 43798 71270 43862
rect 71334 43798 71476 43862
rect 71264 43792 71476 43798
rect 71672 43998 71884 44004
rect 71672 43934 71678 43998
rect 71742 43934 71884 43998
rect 71672 43862 71884 43934
rect 71672 43798 71678 43862
rect 71742 43798 71884 43862
rect 71672 43792 71884 43798
rect 72080 43998 72700 44004
rect 72080 43934 72222 43998
rect 72286 43934 72700 43998
rect 72080 43928 72700 43934
rect 72080 43792 72292 43928
rect 72488 43862 72700 43928
rect 72488 43798 72630 43862
rect 72694 43798 72700 43862
rect 72488 43792 72700 43798
rect 72896 43862 73108 44140
rect 89080 44132 89428 44276
rect 89080 44076 89216 44132
rect 89272 44076 89428 44132
rect 89080 44004 89428 44076
rect 89080 43998 89836 44004
rect 89080 43934 89766 43998
rect 89830 43934 89836 43998
rect 89080 43928 89836 43934
rect 72896 43798 73038 43862
rect 73102 43798 73108 43862
rect 72896 43792 73108 43798
rect 18632 43732 18708 43792
rect 18360 43656 18708 43732
rect 24344 43732 24420 43792
rect 66368 43732 66444 43792
rect 18360 43596 18436 43656
rect 17816 43590 18028 43596
rect 17816 43526 17958 43590
rect 18022 43526 18028 43590
rect 17816 43384 18028 43526
rect 18224 43590 18980 43596
rect 18224 43526 18366 43590
rect 18430 43526 18980 43590
rect 18224 43520 18980 43526
rect 18224 43384 18436 43520
rect 18632 43454 18980 43520
rect 18632 43390 18910 43454
rect 18974 43390 18980 43454
rect 18632 43384 18980 43390
rect 19040 43590 19252 43596
rect 19040 43526 19046 43590
rect 19110 43526 19252 43590
rect 19040 43454 19252 43526
rect 19040 43390 19046 43454
rect 19110 43390 19252 43454
rect 19040 43384 19252 43390
rect 19448 43590 19660 43596
rect 19448 43526 19590 43590
rect 19654 43526 19660 43590
rect 19448 43454 19660 43526
rect 19448 43390 19454 43454
rect 19518 43390 19660 43454
rect 19448 43384 19660 43390
rect 24344 43520 24692 43732
rect 66368 43520 66580 43732
rect 71264 43590 71476 43596
rect 71264 43526 71270 43590
rect 71334 43526 71476 43590
rect 24344 43460 24420 43520
rect 66368 43460 66444 43520
rect 17952 43324 18028 43384
rect 17816 43182 18028 43324
rect 24344 43248 24692 43460
rect 66368 43248 66580 43460
rect 71264 43454 71476 43526
rect 71264 43390 71406 43454
rect 71470 43390 71476 43454
rect 71264 43384 71476 43390
rect 71672 43590 71884 43596
rect 71672 43526 71678 43590
rect 71742 43526 71884 43590
rect 71672 43454 71884 43526
rect 71672 43390 71814 43454
rect 71878 43390 71884 43454
rect 71672 43384 71884 43390
rect 72080 43454 72292 43596
rect 72488 43590 72700 43596
rect 72488 43526 72630 43590
rect 72694 43526 72700 43590
rect 72488 43460 72700 43526
rect 72390 43454 72700 43460
rect 72080 43390 72222 43454
rect 72286 43390 72292 43454
rect 72352 43390 72358 43454
rect 72422 43390 72700 43454
rect 72080 43384 72292 43390
rect 72390 43384 72700 43390
rect 72896 43590 73108 43596
rect 72896 43526 73038 43590
rect 73102 43526 73108 43590
rect 72896 43384 73108 43526
rect 24616 43188 24692 43248
rect 66504 43188 66580 43248
rect 72896 43324 72972 43384
rect 17816 43118 17822 43182
rect 17886 43118 18028 43182
rect 17816 43112 18028 43118
rect 18224 42976 18436 43188
rect 18632 43182 18980 43188
rect 18632 43118 18910 43182
rect 18974 43118 18980 43182
rect 18632 42976 18980 43118
rect 19040 43182 19252 43188
rect 19040 43118 19046 43182
rect 19110 43118 19252 43182
rect 19040 43046 19252 43118
rect 19040 42982 19046 43046
rect 19110 42982 19252 43046
rect 19040 42976 19252 42982
rect 19448 43182 19660 43188
rect 19448 43118 19454 43182
rect 19518 43118 19660 43182
rect 19448 43046 19660 43118
rect 19448 42982 19454 43046
rect 19518 42982 19660 43046
rect 19448 42976 19660 42982
rect 18224 42916 18300 42976
rect 18904 42916 18980 42976
rect 17816 42910 18028 42916
rect 17816 42846 17822 42910
rect 17886 42846 18028 42910
rect 17816 42568 18028 42846
rect 18224 42638 18436 42916
rect 18224 42574 18366 42638
rect 18430 42574 18436 42638
rect 18224 42568 18436 42574
rect 18632 42568 18980 42916
rect 19040 42774 19252 42780
rect 19040 42710 19046 42774
rect 19110 42710 19252 42774
rect 19040 42568 19252 42710
rect 17952 42508 18028 42568
rect 18632 42508 18708 42568
rect 19176 42508 19252 42568
rect 1632 42452 1844 42508
rect 1632 42396 1718 42452
rect 1774 42396 1844 42452
rect 1632 42372 1844 42396
rect 1224 42366 1844 42372
rect 1224 42302 1230 42366
rect 1294 42302 1844 42366
rect 1224 42296 1844 42302
rect 17816 42366 18028 42508
rect 18360 42432 18708 42508
rect 18360 42372 18436 42432
rect 17816 42302 17822 42366
rect 17886 42302 18028 42366
rect 17816 42296 18028 42302
rect 18224 42366 18980 42372
rect 18224 42302 18366 42366
rect 18430 42302 18980 42366
rect 18224 42296 18980 42302
rect 18224 42236 18436 42296
rect 18224 42160 18572 42236
rect 18632 42160 18980 42296
rect 19040 42160 19252 42508
rect 19448 42774 19660 42780
rect 19448 42710 19454 42774
rect 19518 42710 19660 42774
rect 19448 42568 19660 42710
rect 24344 42774 24692 43188
rect 24344 42710 24350 42774
rect 24414 42710 24692 42774
rect 24344 42704 24692 42710
rect 24616 42644 24692 42704
rect 19448 42508 19524 42568
rect 19448 42160 19660 42508
rect 24344 42502 24692 42644
rect 24344 42438 24350 42502
rect 24414 42438 24622 42502
rect 24686 42438 24692 42502
rect 24344 42230 24692 42438
rect 24344 42166 24622 42230
rect 24686 42166 24692 42230
rect 18224 42100 18300 42160
rect 18496 42100 18572 42160
rect 19040 42100 19116 42160
rect 19448 42100 19524 42160
rect 17816 42094 18028 42100
rect 17816 42030 17822 42094
rect 17886 42030 18028 42094
rect 17816 41958 18028 42030
rect 17816 41894 17822 41958
rect 17886 41894 18028 41958
rect 17816 41888 18028 41894
rect 18224 41958 18436 42100
rect 18496 42024 18980 42100
rect 18224 41894 18230 41958
rect 18294 41894 18436 41958
rect 18224 41888 18436 41894
rect 18632 41888 18980 42024
rect 19040 41958 19252 42100
rect 19040 41894 19182 41958
rect 19246 41894 19252 41958
rect 19040 41888 19252 41894
rect 19448 41958 19660 42100
rect 19448 41894 19454 41958
rect 19518 41894 19660 41958
rect 19448 41888 19660 41894
rect 24344 42024 24692 42166
rect 66368 42704 66580 43188
rect 71264 43182 71476 43188
rect 71264 43118 71406 43182
rect 71470 43118 71476 43182
rect 71264 43046 71476 43118
rect 71264 42982 71270 43046
rect 71334 42982 71476 43046
rect 71264 42976 71476 42982
rect 71672 43182 71884 43188
rect 71672 43118 71814 43182
rect 71878 43118 71884 43182
rect 71672 43046 71884 43118
rect 71672 42982 71814 43046
rect 71878 42982 71884 43046
rect 71672 42976 71884 42982
rect 72080 43182 72428 43188
rect 72080 43118 72222 43182
rect 72286 43118 72358 43182
rect 72422 43118 72428 43182
rect 72080 43112 72428 43118
rect 72080 42976 72292 43112
rect 72488 43052 72700 43188
rect 72896 43182 73108 43324
rect 72896 43118 73038 43182
rect 73102 43118 73108 43182
rect 72896 43112 73108 43118
rect 72216 42916 72292 42976
rect 72352 42976 72700 43052
rect 72352 42916 72428 42976
rect 72624 42916 72700 42976
rect 72080 42840 72428 42916
rect 71264 42774 71476 42780
rect 71264 42710 71270 42774
rect 71334 42710 71476 42774
rect 66368 42644 66444 42704
rect 66368 42502 66580 42644
rect 71264 42568 71476 42710
rect 71400 42508 71476 42568
rect 66368 42438 66510 42502
rect 66574 42438 66580 42502
rect 66368 42230 66580 42438
rect 66368 42166 66374 42230
rect 66438 42166 66510 42230
rect 66574 42166 66580 42230
rect 66368 42024 66580 42166
rect 71264 42160 71476 42508
rect 71672 42774 71884 42780
rect 71672 42710 71814 42774
rect 71878 42710 71884 42774
rect 71672 42568 71884 42710
rect 72080 42638 72292 42840
rect 72080 42574 72086 42638
rect 72150 42574 72292 42638
rect 72080 42568 72292 42574
rect 72488 42568 72700 42916
rect 72896 42910 73108 42916
rect 72896 42846 73038 42910
rect 73102 42846 73108 42910
rect 72896 42568 73108 42846
rect 71672 42508 71748 42568
rect 72896 42508 72972 42568
rect 71672 42160 71884 42508
rect 72080 42366 72292 42372
rect 72080 42302 72086 42366
rect 72150 42302 72292 42366
rect 72080 42160 72292 42302
rect 72488 42236 72700 42372
rect 72896 42366 73108 42508
rect 72896 42302 72902 42366
rect 72966 42302 73108 42366
rect 72896 42296 73108 42302
rect 89080 42452 89428 42508
rect 89080 42396 89216 42452
rect 89272 42396 89428 42452
rect 89080 42372 89428 42396
rect 89080 42366 89836 42372
rect 89080 42302 89766 42366
rect 89830 42302 89836 42366
rect 89080 42296 89836 42302
rect 72352 42160 72700 42236
rect 71264 42100 71340 42160
rect 71672 42100 71748 42160
rect 72080 42100 72156 42160
rect 72352 42100 72428 42160
rect 24344 41964 24420 42024
rect 18088 41822 19116 41828
rect 18088 41758 19046 41822
rect 19110 41758 19116 41822
rect 18088 41752 19116 41758
rect 18088 41692 18164 41752
rect 17816 41686 18164 41692
rect 17816 41622 17822 41686
rect 17886 41622 18164 41686
rect 17816 41616 18164 41622
rect 18224 41686 18436 41692
rect 18224 41622 18230 41686
rect 18294 41622 18436 41686
rect 17816 41550 18028 41616
rect 17816 41486 17958 41550
rect 18022 41486 18028 41550
rect 17816 41480 18028 41486
rect 18224 41344 18436 41622
rect 18632 41616 18980 41692
rect 19040 41686 19252 41692
rect 19040 41622 19182 41686
rect 19246 41622 19252 41686
rect 18752 41420 18850 41616
rect 19040 41550 19252 41622
rect 19040 41486 19182 41550
rect 19246 41486 19252 41550
rect 19040 41480 19252 41486
rect 19448 41686 19660 41692
rect 19448 41622 19454 41686
rect 19518 41622 19660 41686
rect 19448 41550 19660 41622
rect 19448 41486 19590 41550
rect 19654 41486 19660 41550
rect 19448 41480 19660 41486
rect 24344 41480 24692 41964
rect 24616 41420 24692 41480
rect 18534 41414 18980 41420
rect 18496 41350 18502 41414
rect 18566 41350 18980 41414
rect 18534 41344 18980 41350
rect 18224 41284 18300 41344
rect 17816 41278 18028 41284
rect 17816 41214 17958 41278
rect 18022 41214 18028 41278
rect 17816 41142 18028 41214
rect 17816 41078 17958 41142
rect 18022 41078 18028 41142
rect 17816 41072 18028 41078
rect 18224 41208 18980 41284
rect 18224 41148 18436 41208
rect 18224 41142 18572 41148
rect 18224 41078 18502 41142
rect 18566 41078 18572 41142
rect 18224 41072 18572 41078
rect 18632 41072 18980 41208
rect 19040 41278 19252 41284
rect 19040 41214 19046 41278
rect 19110 41214 19182 41278
rect 19246 41214 19252 41278
rect 19040 41142 19252 41214
rect 19040 41078 19182 41142
rect 19246 41078 19252 41142
rect 19040 41072 19252 41078
rect 19448 41278 19660 41284
rect 19448 41214 19590 41278
rect 19654 41214 19660 41278
rect 19448 41142 19660 41214
rect 24344 41208 24692 41420
rect 24616 41148 24692 41208
rect 19448 41078 19454 41142
rect 19518 41078 19660 41142
rect 19448 41072 19660 41078
rect 18632 41012 18708 41072
rect 18496 40936 18708 41012
rect 24344 40936 24692 41148
rect 66368 41958 66580 41964
rect 66368 41894 66374 41958
rect 66438 41894 66580 41958
rect 66368 41686 66580 41894
rect 71264 41958 71476 42100
rect 71264 41894 71270 41958
rect 71334 41894 71476 41958
rect 71264 41888 71476 41894
rect 71672 41958 71884 42100
rect 71672 41894 71678 41958
rect 71742 41894 71884 41958
rect 71672 41888 71884 41894
rect 72080 42024 72428 42100
rect 72488 42100 72564 42160
rect 72080 41888 72292 42024
rect 72488 41958 72700 42100
rect 72488 41894 72630 41958
rect 72694 41894 72700 41958
rect 72488 41888 72700 41894
rect 72896 42094 73108 42100
rect 72896 42030 72902 42094
rect 72966 42030 73108 42094
rect 72896 41958 73108 42030
rect 72896 41894 73038 41958
rect 73102 41894 73108 41958
rect 72896 41888 73108 41894
rect 66368 41622 66374 41686
rect 66438 41622 66580 41686
rect 66368 41480 66580 41622
rect 71264 41686 71476 41692
rect 71264 41622 71270 41686
rect 71334 41622 71476 41686
rect 71264 41550 71476 41622
rect 71264 41486 71406 41550
rect 71470 41486 71476 41550
rect 71264 41480 71476 41486
rect 71672 41686 71884 41692
rect 71672 41622 71678 41686
rect 71742 41622 71884 41686
rect 71672 41550 71884 41622
rect 71672 41486 71814 41550
rect 71878 41486 71884 41550
rect 71672 41480 71884 41486
rect 66368 41420 66444 41480
rect 66368 41414 66580 41420
rect 66368 41350 66374 41414
rect 66438 41350 66580 41414
rect 66368 41208 66580 41350
rect 72080 41344 72292 41692
rect 72488 41686 72700 41692
rect 72488 41622 72630 41686
rect 72694 41622 72700 41686
rect 72488 41344 72700 41622
rect 72896 41686 73108 41692
rect 72896 41622 73038 41686
rect 73102 41622 73108 41686
rect 72896 41550 73108 41622
rect 72896 41486 72902 41550
rect 72966 41486 73108 41550
rect 72896 41480 73108 41486
rect 72080 41284 72156 41344
rect 72488 41284 72564 41344
rect 71264 41278 71476 41284
rect 71264 41214 71406 41278
rect 71470 41214 71476 41278
rect 66368 41148 66444 41208
rect 66368 40936 66580 41148
rect 71264 41142 71476 41214
rect 71264 41078 71406 41142
rect 71470 41078 71476 41142
rect 71264 41072 71476 41078
rect 71672 41278 71884 41284
rect 71672 41214 71814 41278
rect 71878 41214 71884 41278
rect 71672 41142 71884 41214
rect 71672 41078 71814 41142
rect 71878 41078 71884 41142
rect 71672 41072 71884 41078
rect 72080 41142 72292 41284
rect 72080 41078 72086 41142
rect 72150 41078 72292 41142
rect 72080 41072 72292 41078
rect 72488 41072 72700 41284
rect 72896 41278 73108 41284
rect 72896 41214 72902 41278
rect 72966 41214 73108 41278
rect 72896 41142 73108 41214
rect 72896 41078 72902 41142
rect 72966 41078 73108 41142
rect 72896 41072 73108 41078
rect 72488 41012 72564 41072
rect 18496 40876 18572 40936
rect 24616 40876 24692 40936
rect 66504 40876 66580 40936
rect 72216 40936 72564 41012
rect 72216 40876 72292 40936
rect 1632 40772 1844 40876
rect 1632 40740 1718 40772
rect 1224 40734 1718 40740
rect 1224 40670 1230 40734
rect 1294 40716 1718 40734
rect 1774 40716 1844 40772
rect 1294 40670 1844 40716
rect 1224 40664 1844 40670
rect 17816 40870 18028 40876
rect 17816 40806 17958 40870
rect 18022 40806 18028 40870
rect 17816 40734 18028 40806
rect 17816 40670 17822 40734
rect 17886 40670 18028 40734
rect 17816 40664 18028 40670
rect 18224 40800 18572 40876
rect 18224 40734 18436 40800
rect 18632 40740 18980 40876
rect 18534 40734 18980 40740
rect 18224 40670 18366 40734
rect 18430 40670 18436 40734
rect 18496 40670 18502 40734
rect 18566 40670 18980 40734
rect 18224 40664 18436 40670
rect 18534 40664 18980 40670
rect 19040 40870 19252 40876
rect 19040 40806 19182 40870
rect 19246 40806 19252 40870
rect 19040 40734 19252 40806
rect 19040 40670 19182 40734
rect 19246 40670 19252 40734
rect 19040 40664 19252 40670
rect 19448 40870 19660 40876
rect 19448 40806 19454 40870
rect 19518 40806 19660 40870
rect 19448 40734 19660 40806
rect 19448 40670 19454 40734
rect 19518 40670 19660 40734
rect 19448 40664 19660 40670
rect 24344 40664 24692 40876
rect 66368 40664 66580 40876
rect 71264 40870 71476 40876
rect 71264 40806 71406 40870
rect 71470 40806 71476 40870
rect 71264 40734 71476 40806
rect 71264 40670 71406 40734
rect 71470 40670 71476 40734
rect 71264 40664 71476 40670
rect 71672 40870 71884 40876
rect 71672 40806 71814 40870
rect 71878 40806 71884 40870
rect 71672 40734 71884 40806
rect 71672 40670 71678 40734
rect 71742 40670 71884 40734
rect 71672 40664 71884 40670
rect 72080 40870 72700 40876
rect 72080 40806 72086 40870
rect 72150 40806 72700 40870
rect 72080 40800 72700 40806
rect 72080 40664 72292 40800
rect 72488 40734 72700 40800
rect 72488 40670 72494 40734
rect 72558 40670 72700 40734
rect 72488 40664 72700 40670
rect 72896 40870 73108 40876
rect 72896 40806 72902 40870
rect 72966 40806 73108 40870
rect 72896 40734 73108 40806
rect 72896 40670 72902 40734
rect 72966 40670 73108 40734
rect 72896 40664 73108 40670
rect 89080 40870 89836 40876
rect 89080 40806 89766 40870
rect 89830 40806 89836 40870
rect 89080 40800 89836 40806
rect 89080 40772 89428 40800
rect 89080 40716 89216 40772
rect 89272 40716 89428 40772
rect 89080 40664 89428 40716
rect 24616 40604 24692 40664
rect 66504 40604 66580 40664
rect 17816 40462 18028 40468
rect 17816 40398 17822 40462
rect 17886 40398 18028 40462
rect 17816 40326 18028 40398
rect 17816 40262 17958 40326
rect 18022 40262 18028 40326
rect 17816 40256 18028 40262
rect 18224 40462 18572 40468
rect 18224 40398 18366 40462
rect 18430 40398 18502 40462
rect 18566 40398 18572 40462
rect 18224 40392 18572 40398
rect 18224 40332 18436 40392
rect 18632 40332 18980 40468
rect 18224 40326 18980 40332
rect 18224 40262 18638 40326
rect 18702 40262 18980 40326
rect 18224 40256 18980 40262
rect 19040 40462 19252 40468
rect 19040 40398 19182 40462
rect 19246 40398 19252 40462
rect 19040 40326 19252 40398
rect 19040 40262 19182 40326
rect 19246 40262 19252 40326
rect 19040 40256 19252 40262
rect 19448 40462 19660 40468
rect 19448 40398 19454 40462
rect 19518 40398 19660 40462
rect 19448 40326 19660 40398
rect 24344 40392 24692 40604
rect 66368 40392 66580 40604
rect 71264 40462 71476 40468
rect 71264 40398 71406 40462
rect 71470 40398 71476 40462
rect 24480 40332 24556 40392
rect 66368 40332 66444 40392
rect 19448 40262 19590 40326
rect 19654 40262 19660 40326
rect 19448 40256 19660 40262
rect 24344 40120 24692 40332
rect 24616 40060 24692 40120
rect 17816 40054 18028 40060
rect 17816 39990 17958 40054
rect 18022 39990 18028 40054
rect 17816 39918 18028 39990
rect 17816 39854 17822 39918
rect 17886 39854 18028 39918
rect 17816 39848 18028 39854
rect 18224 39918 18436 40060
rect 18224 39854 18230 39918
rect 18294 39854 18436 39918
rect 18224 39848 18436 39854
rect 18632 40054 18980 40060
rect 18632 39990 18638 40054
rect 18702 39990 18980 40054
rect 18632 39918 18980 39990
rect 18632 39854 18910 39918
rect 18974 39854 18980 39918
rect 18632 39848 18980 39854
rect 19040 40054 19252 40060
rect 19040 39990 19182 40054
rect 19246 39990 19252 40054
rect 19040 39918 19252 39990
rect 19040 39854 19046 39918
rect 19110 39854 19252 39918
rect 19040 39848 19252 39854
rect 19448 40054 19660 40060
rect 19448 39990 19590 40054
rect 19654 39990 19660 40054
rect 19448 39918 19660 39990
rect 19448 39854 19590 39918
rect 19654 39854 19660 39918
rect 19448 39848 19660 39854
rect 24344 39848 24692 40060
rect 66368 40120 66580 40332
rect 71264 40326 71476 40398
rect 71264 40262 71406 40326
rect 71470 40262 71476 40326
rect 71264 40256 71476 40262
rect 71672 40462 71884 40468
rect 71672 40398 71678 40462
rect 71742 40398 71884 40462
rect 71672 40326 71884 40398
rect 71672 40262 71678 40326
rect 71742 40262 71884 40326
rect 71672 40256 71884 40262
rect 72080 40326 72292 40468
rect 72488 40462 72700 40468
rect 72488 40398 72494 40462
rect 72558 40398 72700 40462
rect 72488 40332 72700 40398
rect 72390 40326 72700 40332
rect 72080 40262 72086 40326
rect 72150 40262 72292 40326
rect 72352 40262 72358 40326
rect 72422 40262 72700 40326
rect 72080 40256 72292 40262
rect 72390 40256 72700 40262
rect 72896 40462 73108 40468
rect 72896 40398 72902 40462
rect 72966 40398 73108 40462
rect 72896 40326 73108 40398
rect 72896 40262 72902 40326
rect 72966 40262 73108 40326
rect 72896 40256 73108 40262
rect 66368 40060 66444 40120
rect 66368 39848 66580 40060
rect 71264 40054 71476 40060
rect 71264 39990 71406 40054
rect 71470 39990 71476 40054
rect 71264 39918 71476 39990
rect 71264 39854 71270 39918
rect 71334 39854 71476 39918
rect 71264 39848 71476 39854
rect 71672 40054 71884 40060
rect 71672 39990 71678 40054
rect 71742 39990 71884 40054
rect 71672 39918 71884 39990
rect 71672 39854 71814 39918
rect 71878 39854 71884 39918
rect 71672 39848 71884 39854
rect 72080 40054 72428 40060
rect 72080 39990 72086 40054
rect 72150 39990 72358 40054
rect 72422 39990 72428 40054
rect 72080 39984 72428 39990
rect 72080 39924 72292 39984
rect 72080 39918 72428 39924
rect 72080 39854 72222 39918
rect 72286 39854 72358 39918
rect 72422 39854 72428 39918
rect 72080 39848 72428 39854
rect 72488 39848 72700 40060
rect 72896 40054 73108 40060
rect 72896 39990 72902 40054
rect 72966 39990 73108 40054
rect 72896 39918 73108 39990
rect 72896 39854 73038 39918
rect 73102 39854 73108 39918
rect 72896 39848 73108 39854
rect 24480 39788 24556 39848
rect 66504 39788 66580 39848
rect 17816 39646 18028 39652
rect 17816 39582 17822 39646
rect 17886 39582 18028 39646
rect 17816 39440 18028 39582
rect 18224 39646 18436 39652
rect 18224 39582 18230 39646
rect 18294 39582 18436 39646
rect 18224 39510 18436 39582
rect 18632 39646 18980 39652
rect 18632 39582 18910 39646
rect 18974 39582 18980 39646
rect 18632 39516 18980 39582
rect 18534 39510 18980 39516
rect 18224 39446 18366 39510
rect 18430 39446 18436 39510
rect 18496 39446 18502 39510
rect 18566 39446 18774 39510
rect 18838 39446 18980 39510
rect 18224 39440 18436 39446
rect 18534 39440 18980 39446
rect 19040 39646 19252 39652
rect 19040 39582 19046 39646
rect 19110 39582 19252 39646
rect 19040 39510 19252 39582
rect 19040 39446 19182 39510
rect 19246 39446 19252 39510
rect 19040 39440 19252 39446
rect 19448 39646 19660 39652
rect 19448 39582 19590 39646
rect 19654 39582 19660 39646
rect 19448 39510 19660 39582
rect 19448 39446 19454 39510
rect 19518 39446 19660 39510
rect 19448 39440 19660 39446
rect 24344 39576 24692 39788
rect 66368 39576 66580 39788
rect 72216 39788 72292 39848
rect 72488 39788 72564 39848
rect 72216 39712 72564 39788
rect 24344 39516 24420 39576
rect 66504 39516 66580 39576
rect 17816 39380 17892 39440
rect 1224 39238 1844 39244
rect 1224 39174 1230 39238
rect 1294 39174 1844 39238
rect 1224 39168 1844 39174
rect 1632 39092 1844 39168
rect 1632 39036 1718 39092
rect 1774 39036 1844 39092
rect 1632 38896 1844 39036
rect 17816 39032 18028 39380
rect 24344 39374 24692 39516
rect 24344 39310 24350 39374
rect 24414 39310 24692 39374
rect 24344 39304 24692 39310
rect 66368 39374 66580 39516
rect 71264 39646 71476 39652
rect 71264 39582 71270 39646
rect 71334 39582 71476 39646
rect 71264 39510 71476 39582
rect 71264 39446 71270 39510
rect 71334 39446 71476 39510
rect 71264 39440 71476 39446
rect 71672 39646 71884 39652
rect 71672 39582 71814 39646
rect 71878 39582 71884 39646
rect 71672 39510 71884 39582
rect 71672 39446 71814 39510
rect 71878 39446 71884 39510
rect 71672 39440 71884 39446
rect 72080 39646 72292 39652
rect 72390 39646 72700 39652
rect 72080 39582 72222 39646
rect 72286 39582 72292 39646
rect 72352 39582 72358 39646
rect 72422 39582 72700 39646
rect 72080 39510 72292 39582
rect 72390 39576 72700 39582
rect 72080 39446 72086 39510
rect 72150 39446 72292 39510
rect 72080 39440 72292 39446
rect 72488 39440 72700 39576
rect 72896 39646 73108 39652
rect 72896 39582 73038 39646
rect 73102 39582 73108 39646
rect 72896 39440 73108 39582
rect 73032 39380 73108 39440
rect 66368 39310 66374 39374
rect 66438 39310 66580 39374
rect 66368 39304 66580 39310
rect 24480 39244 24556 39304
rect 66368 39244 66444 39304
rect 18224 39238 18572 39244
rect 18224 39174 18366 39238
rect 18430 39174 18502 39238
rect 18566 39174 18572 39238
rect 18224 39168 18572 39174
rect 18632 39238 18980 39244
rect 18632 39174 18774 39238
rect 18838 39174 18980 39238
rect 18224 39032 18436 39168
rect 17952 38972 18028 39032
rect 18360 38972 18436 39032
rect 17816 38624 18028 38972
rect 18224 38624 18436 38972
rect 18632 39032 18980 39174
rect 19040 39238 19252 39244
rect 19040 39174 19182 39238
rect 19246 39174 19252 39238
rect 19040 39102 19252 39174
rect 19040 39038 19046 39102
rect 19110 39038 19252 39102
rect 19040 39032 19252 39038
rect 19448 39238 19660 39244
rect 19448 39174 19454 39238
rect 19518 39174 19660 39238
rect 19448 39102 19660 39174
rect 19448 39038 19454 39102
rect 19518 39038 19660 39102
rect 19448 39032 19660 39038
rect 24344 39102 24692 39244
rect 24344 39038 24350 39102
rect 24414 39038 24692 39102
rect 18632 38972 18708 39032
rect 18632 38694 18980 38972
rect 18632 38630 18910 38694
rect 18974 38630 18980 38694
rect 18632 38624 18980 38630
rect 19040 38830 19252 38836
rect 19040 38766 19046 38830
rect 19110 38766 19252 38830
rect 19040 38624 19252 38766
rect 19448 38830 19660 38836
rect 19448 38766 19454 38830
rect 19518 38766 19660 38830
rect 19448 38624 19660 38766
rect 24344 38760 24692 39038
rect 66368 39102 66580 39244
rect 66368 39038 66374 39102
rect 66438 39038 66580 39102
rect 66368 38830 66580 39038
rect 71264 39238 71476 39244
rect 71264 39174 71270 39238
rect 71334 39174 71476 39238
rect 71264 39102 71476 39174
rect 71264 39038 71270 39102
rect 71334 39038 71476 39102
rect 71264 39032 71476 39038
rect 71672 39238 71884 39244
rect 71672 39174 71814 39238
rect 71878 39174 71884 39238
rect 71672 39102 71884 39174
rect 71672 39038 71814 39102
rect 71878 39038 71884 39102
rect 71672 39032 71884 39038
rect 72080 39238 72292 39244
rect 72080 39174 72086 39238
rect 72150 39174 72292 39238
rect 72080 39032 72292 39174
rect 72488 39032 72700 39244
rect 72896 39032 73108 39380
rect 89080 39238 89836 39244
rect 89080 39174 89766 39238
rect 89830 39174 89836 39238
rect 89080 39168 89836 39174
rect 89080 39092 89428 39168
rect 89080 39036 89216 39092
rect 89272 39036 89428 39092
rect 72080 38972 72156 39032
rect 72488 38972 72564 39032
rect 72896 38972 72972 39032
rect 66368 38766 66510 38830
rect 66574 38766 66580 38830
rect 66368 38760 66580 38766
rect 71264 38830 71476 38836
rect 71264 38766 71270 38830
rect 71334 38766 71476 38830
rect 24480 38700 24556 38760
rect 66368 38700 66444 38760
rect 17952 38564 18028 38624
rect 17816 38422 18028 38564
rect 19040 38564 19116 38624
rect 19448 38564 19524 38624
rect 17816 38358 17822 38422
rect 17886 38358 18028 38422
rect 17816 38352 18028 38358
rect 18224 38216 18436 38428
rect 18632 38422 18980 38428
rect 18632 38358 18910 38422
rect 18974 38358 18980 38422
rect 18632 38216 18980 38358
rect 19040 38216 19252 38564
rect 18360 38156 18436 38216
rect 18768 38156 18844 38216
rect 19176 38156 19252 38216
rect 11016 38014 11228 38156
rect 11016 37950 11158 38014
rect 11222 37950 11228 38014
rect 11016 37944 11228 37950
rect 17816 38150 18028 38156
rect 17816 38086 17822 38150
rect 17886 38086 18028 38150
rect 17816 38014 18028 38086
rect 17816 37950 17822 38014
rect 17886 37950 18028 38014
rect 17816 37944 18028 37950
rect 18224 38080 18980 38156
rect 18224 38020 18436 38080
rect 18224 38014 18572 38020
rect 18224 37950 18502 38014
rect 18566 37950 18572 38014
rect 18224 37944 18572 37950
rect 18632 37944 18980 38080
rect 19040 37808 19252 38156
rect 19448 38216 19660 38564
rect 19448 38156 19524 38216
rect 19448 37808 19660 38156
rect 24344 38150 24692 38700
rect 24344 38086 24622 38150
rect 24686 38086 24692 38150
rect 24344 38080 24692 38086
rect 66368 38558 66580 38700
rect 66368 38494 66510 38558
rect 66574 38494 66580 38558
rect 66368 38150 66580 38494
rect 71264 38624 71476 38766
rect 71672 38830 71884 38836
rect 71672 38766 71814 38830
rect 71878 38766 71884 38830
rect 71672 38624 71884 38766
rect 72080 38700 72292 38972
rect 72488 38700 72700 38972
rect 72080 38694 72700 38700
rect 72080 38630 72222 38694
rect 72286 38630 72700 38694
rect 72080 38624 72700 38630
rect 72896 38624 73108 38972
rect 89080 38896 89428 39036
rect 71264 38564 71340 38624
rect 71672 38564 71748 38624
rect 73032 38564 73108 38624
rect 71264 38216 71476 38564
rect 71400 38156 71476 38216
rect 66368 38086 66374 38150
rect 66438 38086 66510 38150
rect 66574 38086 66580 38150
rect 66368 38080 66580 38086
rect 19040 37748 19116 37808
rect 19584 37748 19660 37808
rect 17816 37742 18028 37748
rect 17816 37678 17822 37742
rect 17886 37678 18028 37742
rect 17816 37606 18028 37678
rect 17816 37542 17958 37606
rect 18022 37542 18028 37606
rect 17816 37536 18028 37542
rect 1632 37412 1844 37476
rect 1632 37356 1718 37412
rect 1774 37356 1844 37412
rect 1632 37340 1844 37356
rect 18224 37400 18436 37748
rect 18534 37742 18980 37748
rect 18496 37678 18502 37742
rect 18566 37678 18980 37742
rect 18534 37672 18980 37678
rect 18632 37400 18980 37672
rect 19040 37606 19252 37748
rect 19040 37542 19046 37606
rect 19110 37542 19252 37606
rect 19040 37536 19252 37542
rect 19448 37606 19660 37748
rect 19448 37542 19590 37606
rect 19654 37542 19660 37606
rect 19448 37536 19660 37542
rect 24344 37878 24692 37884
rect 24344 37814 24622 37878
rect 24686 37814 24692 37878
rect 24344 37536 24692 37814
rect 66368 37878 66580 37884
rect 66368 37814 66374 37878
rect 66438 37814 66580 37878
rect 66368 37742 66580 37814
rect 66368 37678 66510 37742
rect 66574 37678 66580 37742
rect 66368 37536 66580 37678
rect 71264 37808 71476 38156
rect 71672 38216 71884 38564
rect 72080 38422 72292 38428
rect 72080 38358 72222 38422
rect 72286 38358 72292 38422
rect 72080 38292 72292 38358
rect 72080 38216 72428 38292
rect 71672 38156 71748 38216
rect 72080 38156 72156 38216
rect 72352 38156 72428 38216
rect 72488 38216 72700 38428
rect 72896 38422 73108 38564
rect 72896 38358 72902 38422
rect 72966 38358 73108 38422
rect 72896 38352 73108 38358
rect 72488 38156 72564 38216
rect 71672 37808 71884 38156
rect 72080 38014 72292 38156
rect 72352 38080 72700 38156
rect 72080 37950 72086 38014
rect 72150 37950 72292 38014
rect 72080 37944 72292 37950
rect 72488 37944 72700 38080
rect 72896 38150 73108 38156
rect 72896 38086 72902 38150
rect 72966 38086 73108 38150
rect 72896 38014 73108 38086
rect 72896 37950 72902 38014
rect 72966 37950 73108 38014
rect 72896 37944 73108 37950
rect 71264 37748 71340 37808
rect 71808 37748 71884 37808
rect 71264 37606 71476 37748
rect 71264 37542 71270 37606
rect 71334 37542 71476 37606
rect 71264 37536 71476 37542
rect 71672 37606 71884 37748
rect 71672 37542 71678 37606
rect 71742 37542 71884 37606
rect 71672 37536 71884 37542
rect 72080 37742 72292 37748
rect 72080 37678 72086 37742
rect 72150 37678 72292 37742
rect 72080 37612 72292 37678
rect 72488 37612 72700 37748
rect 72080 37536 72700 37612
rect 72896 37742 73108 37748
rect 72896 37678 72902 37742
rect 72966 37678 73108 37742
rect 72896 37606 73108 37678
rect 72896 37542 73038 37606
rect 73102 37542 73108 37606
rect 72896 37536 73108 37542
rect 24480 37476 24556 37536
rect 66504 37476 66580 37536
rect 18224 37340 18300 37400
rect 18904 37340 18980 37400
rect 1224 37334 1844 37340
rect 1224 37270 1230 37334
rect 1294 37270 1844 37334
rect 1224 37264 1844 37270
rect 10608 37189 10820 37340
rect 17816 37334 18028 37340
rect 17816 37270 17958 37334
rect 18022 37270 18028 37334
rect 11616 37262 11682 37265
rect 12350 37262 12416 37265
rect 11616 37260 12416 37262
rect 11616 37204 11621 37260
rect 11677 37204 12355 37260
rect 12411 37204 12416 37260
rect 11616 37202 12416 37204
rect 11616 37199 11682 37202
rect 12350 37199 12416 37202
rect 10608 37133 10676 37189
rect 10732 37133 10820 37189
rect 10608 37068 10820 37133
rect 17816 37198 18028 37270
rect 17816 37134 17822 37198
rect 17886 37134 18028 37198
rect 17816 37128 18028 37134
rect 18224 37204 18436 37340
rect 18632 37204 18980 37340
rect 18224 37198 18980 37204
rect 18224 37134 18366 37198
rect 18430 37134 18980 37198
rect 18224 37128 18980 37134
rect 19040 37334 19252 37340
rect 19040 37270 19046 37334
rect 19110 37270 19252 37334
rect 19040 37198 19252 37270
rect 19040 37134 19182 37198
rect 19246 37134 19252 37198
rect 19040 37128 19252 37134
rect 19448 37334 19660 37340
rect 19448 37270 19590 37334
rect 19654 37270 19660 37334
rect 19448 37198 19660 37270
rect 24344 37264 24692 37476
rect 66368 37264 66580 37476
rect 72080 37476 72292 37536
rect 72080 37400 72428 37476
rect 72488 37400 72700 37536
rect 89080 37412 89428 37476
rect 72080 37340 72156 37400
rect 72352 37340 72428 37400
rect 89080 37356 89216 37412
rect 89272 37356 89428 37412
rect 89080 37340 89428 37356
rect 71264 37334 71476 37340
rect 71264 37270 71270 37334
rect 71334 37270 71476 37334
rect 24480 37204 24556 37264
rect 66368 37204 66444 37264
rect 19448 37134 19454 37198
rect 19518 37134 19660 37198
rect 19448 37128 19660 37134
rect 0 36992 10820 37068
rect 18360 37068 18436 37128
rect 18360 36992 18708 37068
rect 18632 36932 18708 36992
rect 17816 36926 18028 36932
rect 17816 36862 17822 36926
rect 17886 36862 18028 36926
rect 17816 36790 18028 36862
rect 17816 36726 17958 36790
rect 18022 36726 18028 36790
rect 17816 36720 18028 36726
rect 18224 36926 18436 36932
rect 18224 36862 18366 36926
rect 18430 36862 18436 36926
rect 18224 36790 18436 36862
rect 18224 36726 18230 36790
rect 18294 36726 18436 36790
rect 18224 36720 18436 36726
rect 18632 36790 18980 36932
rect 18632 36726 18910 36790
rect 18974 36726 18980 36790
rect 18632 36720 18980 36726
rect 19040 36926 19252 36932
rect 19040 36862 19182 36926
rect 19246 36862 19252 36926
rect 19040 36790 19252 36862
rect 19040 36726 19182 36790
rect 19246 36726 19252 36790
rect 19040 36720 19252 36726
rect 19448 36926 19660 36932
rect 19448 36862 19454 36926
rect 19518 36862 19660 36926
rect 19448 36790 19660 36862
rect 19448 36726 19590 36790
rect 19654 36726 19660 36790
rect 19448 36720 19660 36726
rect 24344 36926 24692 37204
rect 24344 36862 24622 36926
rect 24686 36862 24692 36926
rect 24344 36720 24692 36862
rect 66368 36926 66580 37204
rect 71264 37198 71476 37270
rect 71264 37134 71406 37198
rect 71470 37134 71476 37198
rect 71264 37128 71476 37134
rect 71672 37334 71884 37340
rect 71672 37270 71678 37334
rect 71742 37270 71884 37334
rect 71672 37198 71884 37270
rect 71672 37134 71678 37198
rect 71742 37134 71884 37198
rect 71672 37128 71884 37134
rect 72080 37128 72292 37340
rect 72352 37264 72700 37340
rect 72488 37198 72700 37264
rect 72488 37134 72494 37198
rect 72558 37134 72700 37198
rect 72488 37128 72700 37134
rect 72896 37334 73108 37340
rect 72896 37270 73038 37334
rect 73102 37270 73108 37334
rect 72896 37198 73108 37270
rect 89080 37334 89836 37340
rect 89080 37270 89766 37334
rect 89830 37270 89836 37334
rect 89080 37264 89836 37270
rect 72896 37134 72902 37198
rect 72966 37134 73108 37198
rect 72896 37128 73108 37134
rect 66368 36862 66374 36926
rect 66438 36862 66580 36926
rect 66368 36720 66580 36862
rect 71264 36926 71476 36932
rect 71264 36862 71406 36926
rect 71470 36862 71476 36926
rect 71264 36790 71476 36862
rect 71264 36726 71270 36790
rect 71334 36726 71476 36790
rect 71264 36720 71476 36726
rect 71672 36926 71884 36932
rect 71672 36862 71678 36926
rect 71742 36862 71884 36926
rect 71672 36790 71884 36862
rect 71672 36726 71678 36790
rect 71742 36726 71884 36790
rect 71672 36720 71884 36726
rect 72080 36790 72292 36932
rect 72488 36926 72700 36932
rect 72488 36862 72494 36926
rect 72558 36862 72700 36926
rect 72488 36796 72700 36862
rect 72390 36790 72700 36796
rect 72080 36726 72086 36790
rect 72150 36726 72292 36790
rect 72352 36726 72358 36790
rect 72422 36726 72700 36790
rect 72080 36720 72292 36726
rect 72390 36720 72700 36726
rect 72896 36926 73108 36932
rect 72896 36862 72902 36926
rect 72966 36862 73108 36926
rect 72896 36790 73108 36862
rect 72896 36726 73038 36790
rect 73102 36726 73108 36790
rect 72896 36720 73108 36726
rect 24344 36660 24420 36720
rect 66504 36660 66580 36720
rect 11016 36524 11228 36660
rect 24344 36654 24692 36660
rect 24344 36590 24622 36654
rect 24686 36590 24692 36654
rect 11016 36518 11326 36524
rect 17816 36518 18028 36524
rect 11016 36454 11294 36518
rect 11358 36454 11364 36518
rect 17816 36454 17958 36518
rect 18022 36454 18028 36518
rect 11016 36448 11326 36454
rect 17816 36382 18028 36454
rect 17816 36318 17822 36382
rect 17886 36318 18028 36382
rect 17816 36312 18028 36318
rect 18224 36518 18436 36524
rect 18224 36454 18230 36518
rect 18294 36454 18436 36518
rect 18224 36312 18436 36454
rect 18632 36518 18980 36524
rect 18632 36454 18910 36518
rect 18974 36454 18980 36518
rect 18632 36312 18980 36454
rect 19040 36518 19252 36524
rect 19040 36454 19182 36518
rect 19246 36454 19252 36518
rect 19040 36382 19252 36454
rect 19040 36318 19046 36382
rect 19110 36318 19252 36382
rect 19040 36312 19252 36318
rect 19448 36518 19660 36524
rect 19448 36454 19590 36518
rect 19654 36454 19660 36518
rect 19448 36382 19660 36454
rect 24344 36448 24692 36590
rect 66368 36654 66580 36660
rect 66368 36590 66374 36654
rect 66438 36590 66580 36654
rect 66368 36448 66580 36590
rect 24616 36388 24692 36448
rect 66504 36388 66580 36448
rect 19448 36318 19454 36382
rect 19518 36318 19660 36382
rect 19448 36312 19660 36318
rect 18632 36252 18708 36312
rect 18360 36176 18708 36252
rect 24344 36176 24692 36388
rect 66368 36176 66580 36388
rect 71264 36518 71476 36524
rect 71264 36454 71270 36518
rect 71334 36454 71476 36518
rect 71264 36382 71476 36454
rect 71264 36318 71270 36382
rect 71334 36318 71476 36382
rect 71264 36312 71476 36318
rect 71672 36518 71884 36524
rect 71672 36454 71678 36518
rect 71742 36454 71884 36518
rect 71672 36382 71884 36454
rect 71672 36318 71678 36382
rect 71742 36318 71884 36382
rect 71672 36312 71884 36318
rect 72080 36518 72428 36524
rect 72080 36454 72086 36518
rect 72150 36454 72358 36518
rect 72422 36454 72428 36518
rect 72080 36448 72428 36454
rect 72080 36388 72292 36448
rect 72488 36388 72700 36524
rect 72080 36382 72700 36388
rect 72080 36318 72494 36382
rect 72558 36318 72700 36382
rect 72080 36312 72700 36318
rect 72896 36518 73108 36524
rect 72896 36454 73038 36518
rect 73102 36454 73108 36518
rect 72896 36382 73108 36454
rect 72896 36318 72902 36382
rect 72966 36318 73108 36382
rect 72896 36312 73108 36318
rect 18360 36116 18436 36176
rect 24480 36116 24556 36176
rect 66368 36116 66444 36176
rect 10608 36061 10820 36116
rect 10608 36005 10676 36061
rect 10732 36005 10820 36061
rect 10608 35980 10820 36005
rect 17816 36110 18028 36116
rect 17816 36046 17822 36110
rect 17886 36046 18028 36110
rect 0 35904 10820 35980
rect 11616 35992 11682 35995
rect 12270 35992 12336 35995
rect 11616 35990 12336 35992
rect 11616 35934 11621 35990
rect 11677 35934 12275 35990
rect 12331 35934 12336 35990
rect 11616 35932 12336 35934
rect 11616 35929 11682 35932
rect 12270 35929 12336 35932
rect 17816 35974 18028 36046
rect 17816 35910 17822 35974
rect 17886 35910 18028 35974
rect 17816 35904 18028 35910
rect 18224 36040 18980 36116
rect 18224 35904 18436 36040
rect 18632 35974 18980 36040
rect 18632 35910 18910 35974
rect 18974 35910 18980 35974
rect 18632 35904 18980 35910
rect 19040 36110 19252 36116
rect 19040 36046 19046 36110
rect 19110 36046 19252 36110
rect 19040 35974 19252 36046
rect 19040 35910 19182 35974
rect 19246 35910 19252 35974
rect 19040 35904 19252 35910
rect 19448 36110 19660 36116
rect 19448 36046 19454 36110
rect 19518 36046 19660 36110
rect 19448 35974 19660 36046
rect 19448 35910 19454 35974
rect 19518 35910 19660 35974
rect 19448 35904 19660 35910
rect 24344 35904 24692 36116
rect 66368 35904 66580 36116
rect 71264 36110 71476 36116
rect 71264 36046 71270 36110
rect 71334 36046 71476 36110
rect 71264 35974 71476 36046
rect 71264 35910 71406 35974
rect 71470 35910 71476 35974
rect 71264 35904 71476 35910
rect 71672 36110 71884 36116
rect 71672 36046 71678 36110
rect 71742 36046 71884 36110
rect 71672 35974 71884 36046
rect 71672 35910 71678 35974
rect 71742 35910 71884 35974
rect 71672 35904 71884 35910
rect 72080 35974 72292 36116
rect 72488 36110 72700 36116
rect 72488 36046 72494 36110
rect 72558 36046 72700 36110
rect 72488 35980 72700 36046
rect 72390 35974 72700 35980
rect 72080 35910 72086 35974
rect 72150 35910 72292 35974
rect 72352 35910 72358 35974
rect 72422 35910 72700 35974
rect 72080 35904 72292 35910
rect 72390 35904 72700 35910
rect 72896 36110 73108 36116
rect 72896 36046 72902 36110
rect 72966 36046 73108 36110
rect 72896 35974 73108 36046
rect 72896 35910 72902 35974
rect 72966 35910 73108 35974
rect 72896 35904 73108 35910
rect 24480 35844 24556 35904
rect 66368 35844 66444 35904
rect 1632 35732 1844 35844
rect 1632 35708 1718 35732
rect 1224 35702 1718 35708
rect 1224 35638 1230 35702
rect 1294 35676 1718 35702
rect 1774 35676 1844 35732
rect 1294 35638 1844 35676
rect 1224 35632 1844 35638
rect 17816 35702 18028 35708
rect 17816 35638 17822 35702
rect 17886 35638 18028 35702
rect 17816 35496 18028 35638
rect 18224 35572 18436 35708
rect 18632 35702 18980 35708
rect 18632 35638 18910 35702
rect 18974 35638 18980 35702
rect 18224 35566 18572 35572
rect 18224 35502 18502 35566
rect 18566 35502 18572 35566
rect 18224 35496 18572 35502
rect 18632 35566 18980 35638
rect 18632 35502 18910 35566
rect 18974 35502 18980 35566
rect 18632 35496 18980 35502
rect 19040 35702 19252 35708
rect 19040 35638 19182 35702
rect 19246 35638 19252 35702
rect 19040 35566 19252 35638
rect 19040 35502 19046 35566
rect 19110 35502 19252 35566
rect 19040 35496 19252 35502
rect 19448 35702 19660 35708
rect 19448 35638 19454 35702
rect 19518 35638 19660 35702
rect 19448 35566 19660 35638
rect 24344 35632 24692 35844
rect 24616 35572 24692 35632
rect 19448 35502 19590 35566
rect 19654 35502 19660 35566
rect 19448 35496 19660 35502
rect 17816 35436 17892 35496
rect 11016 35294 11228 35300
rect 11016 35230 11158 35294
rect 11222 35230 11228 35294
rect 11016 35158 11228 35230
rect 11016 35094 11022 35158
rect 11086 35094 11228 35158
rect 11016 35088 11228 35094
rect 17816 35088 18028 35436
rect 24344 35360 24692 35572
rect 66368 35632 66580 35844
rect 89080 35732 89428 35844
rect 71264 35702 71476 35708
rect 71264 35638 71406 35702
rect 71470 35638 71476 35702
rect 66368 35572 66444 35632
rect 66368 35360 66580 35572
rect 71264 35566 71476 35638
rect 71264 35502 71270 35566
rect 71334 35502 71476 35566
rect 71264 35496 71476 35502
rect 71672 35702 71884 35708
rect 71672 35638 71678 35702
rect 71742 35638 71884 35702
rect 71672 35566 71884 35638
rect 71672 35502 71814 35566
rect 71878 35502 71884 35566
rect 71672 35496 71884 35502
rect 72080 35702 72428 35708
rect 72080 35638 72086 35702
rect 72150 35638 72358 35702
rect 72422 35638 72428 35702
rect 72080 35632 72428 35638
rect 72080 35566 72292 35632
rect 72488 35572 72700 35708
rect 72390 35566 72700 35572
rect 72080 35502 72222 35566
rect 72286 35502 72292 35566
rect 72352 35502 72358 35566
rect 72422 35502 72700 35566
rect 72080 35496 72292 35502
rect 72390 35496 72700 35502
rect 72896 35702 73108 35708
rect 72896 35638 72902 35702
rect 72966 35638 73108 35702
rect 72896 35496 73108 35638
rect 89080 35676 89216 35732
rect 89272 35708 89428 35732
rect 89272 35702 89836 35708
rect 89272 35676 89766 35702
rect 89080 35638 89766 35676
rect 89830 35638 89836 35702
rect 89080 35632 89836 35638
rect 73032 35436 73108 35496
rect 24480 35300 24556 35360
rect 66504 35300 66580 35360
rect 18224 35088 18436 35300
rect 18534 35294 18980 35300
rect 18496 35230 18502 35294
rect 18566 35230 18910 35294
rect 18974 35230 18980 35294
rect 18534 35224 18980 35230
rect 18632 35164 18980 35224
rect 17952 35028 18028 35088
rect 18360 35028 18436 35088
rect 18496 35088 18980 35164
rect 19040 35294 19252 35300
rect 19040 35230 19046 35294
rect 19110 35230 19252 35294
rect 19040 35158 19252 35230
rect 19040 35094 19046 35158
rect 19110 35094 19252 35158
rect 19040 35088 19252 35094
rect 19448 35294 19660 35300
rect 19448 35230 19590 35294
rect 19654 35230 19660 35294
rect 19448 35158 19660 35230
rect 19448 35094 19454 35158
rect 19518 35094 19660 35158
rect 19448 35088 19660 35094
rect 18496 35028 18572 35088
rect 17816 34680 18028 35028
rect 18224 34952 18572 35028
rect 18632 35028 18708 35088
rect 18224 34680 18436 34952
rect 18632 34750 18980 35028
rect 18632 34686 18638 34750
rect 18702 34686 18980 34750
rect 18632 34680 18980 34686
rect 19040 34886 19252 34892
rect 19040 34822 19046 34886
rect 19110 34822 19252 34886
rect 19040 34750 19252 34822
rect 19040 34686 19046 34750
rect 19110 34686 19252 34750
rect 19040 34680 19252 34686
rect 19448 34886 19660 34892
rect 19448 34822 19454 34886
rect 19518 34822 19660 34886
rect 19448 34750 19660 34822
rect 19448 34686 19454 34750
rect 19518 34686 19660 34750
rect 19448 34680 19660 34686
rect 24344 34816 24692 35300
rect 66368 34816 66580 35300
rect 71264 35294 71476 35300
rect 71264 35230 71270 35294
rect 71334 35230 71476 35294
rect 71264 35158 71476 35230
rect 71264 35094 71270 35158
rect 71334 35094 71476 35158
rect 71264 35088 71476 35094
rect 71672 35294 71884 35300
rect 71672 35230 71814 35294
rect 71878 35230 71884 35294
rect 71672 35158 71884 35230
rect 71672 35094 71814 35158
rect 71878 35094 71884 35158
rect 71672 35088 71884 35094
rect 72080 35294 72428 35300
rect 72080 35230 72222 35294
rect 72286 35230 72358 35294
rect 72422 35230 72428 35294
rect 72080 35224 72428 35230
rect 72080 35088 72292 35224
rect 72488 35088 72700 35300
rect 72216 35028 72292 35088
rect 72624 35028 72700 35088
rect 24344 34756 24420 34816
rect 66504 34756 66580 34816
rect 17952 34620 18028 34680
rect 10608 34361 10820 34484
rect 17816 34478 18028 34620
rect 24344 34614 24692 34756
rect 24344 34550 24622 34614
rect 24686 34550 24692 34614
rect 24344 34544 24692 34550
rect 66368 34544 66580 34756
rect 71264 34886 71476 34892
rect 71264 34822 71270 34886
rect 71334 34822 71476 34886
rect 71264 34750 71476 34822
rect 71264 34686 71270 34750
rect 71334 34686 71476 34750
rect 71264 34680 71476 34686
rect 71672 34886 71884 34892
rect 71672 34822 71814 34886
rect 71878 34822 71884 34886
rect 71672 34750 71884 34822
rect 71672 34686 71678 34750
rect 71742 34686 71884 34750
rect 71672 34680 71884 34686
rect 72080 34750 72292 35028
rect 72080 34686 72222 34750
rect 72286 34686 72292 34750
rect 72080 34680 72292 34686
rect 72488 34680 72700 35028
rect 72896 35088 73108 35436
rect 72896 35028 72972 35088
rect 72896 34680 73108 35028
rect 72488 34620 72564 34680
rect 24616 34484 24692 34544
rect 66504 34484 66580 34544
rect 72216 34544 72564 34620
rect 72896 34620 72972 34680
rect 72216 34484 72292 34544
rect 11616 34434 11682 34437
rect 12190 34434 12256 34437
rect 11616 34432 12256 34434
rect 11616 34376 11621 34432
rect 11677 34376 12195 34432
rect 12251 34376 12256 34432
rect 17816 34414 17958 34478
rect 18022 34414 18028 34478
rect 17816 34408 18028 34414
rect 11616 34374 12256 34376
rect 11616 34371 11682 34374
rect 12190 34371 12256 34374
rect 10608 34348 10676 34361
rect 0 34305 10676 34348
rect 10732 34305 10820 34361
rect 0 34272 10820 34305
rect 18224 34272 18436 34484
rect 18632 34478 18980 34484
rect 18632 34414 18638 34478
rect 18702 34414 18980 34478
rect 18632 34272 18980 34414
rect 19040 34478 19252 34484
rect 19040 34414 19046 34478
rect 19110 34414 19252 34478
rect 19040 34272 19252 34414
rect 19448 34478 19660 34484
rect 19448 34414 19454 34478
rect 19518 34414 19660 34478
rect 19448 34272 19660 34414
rect 24344 34342 24692 34484
rect 24344 34278 24622 34342
rect 24686 34278 24692 34342
rect 18224 34212 18300 34272
rect 18632 34212 18708 34272
rect 19040 34212 19116 34272
rect 19448 34212 19524 34272
rect 17816 34206 18028 34212
rect 17816 34142 17958 34206
rect 18022 34142 18028 34206
rect 1224 34070 1844 34076
rect 1224 34006 1230 34070
rect 1294 34052 1844 34070
rect 1294 34006 1718 34052
rect 1224 34000 1718 34006
rect 1632 33996 1718 34000
rect 1774 33996 1844 34052
rect 17816 34070 18028 34142
rect 17816 34006 17822 34070
rect 17886 34006 18028 34070
rect 17816 34000 18028 34006
rect 18224 34070 18436 34212
rect 18224 34006 18230 34070
rect 18294 34006 18436 34070
rect 18224 34000 18436 34006
rect 18632 34070 18980 34212
rect 18632 34006 18638 34070
rect 18702 34006 18980 34070
rect 18632 34000 18980 34006
rect 1632 33864 1844 33996
rect 11016 33934 11364 33940
rect 11016 33870 11294 33934
rect 11358 33870 11364 33934
rect 11016 33864 11364 33870
rect 19040 33864 19252 34212
rect 19448 33864 19660 34212
rect 24344 34206 24692 34278
rect 24344 34142 24622 34206
rect 24686 34142 24692 34206
rect 24344 34136 24692 34142
rect 66368 34206 66580 34484
rect 66368 34142 66510 34206
rect 66574 34142 66580 34206
rect 66368 34136 66580 34142
rect 71264 34478 71476 34484
rect 71264 34414 71270 34478
rect 71334 34414 71476 34478
rect 71264 34272 71476 34414
rect 71672 34478 71884 34484
rect 71672 34414 71678 34478
rect 71742 34414 71884 34478
rect 71672 34272 71884 34414
rect 72080 34478 72700 34484
rect 72080 34414 72222 34478
rect 72286 34414 72700 34478
rect 72080 34408 72700 34414
rect 72896 34478 73108 34620
rect 72896 34414 73038 34478
rect 73102 34414 73108 34478
rect 72896 34408 73108 34414
rect 72080 34348 72292 34408
rect 72080 34272 72428 34348
rect 72488 34272 72700 34408
rect 71264 34212 71340 34272
rect 71672 34212 71748 34272
rect 72216 34212 72292 34272
rect 11016 33662 11228 33864
rect 19176 33804 19252 33864
rect 19584 33804 19660 33864
rect 11016 33598 11158 33662
rect 11222 33598 11228 33662
rect 11016 33592 11228 33598
rect 17816 33798 18028 33804
rect 17816 33734 17822 33798
rect 17886 33734 18028 33798
rect 17816 33662 18028 33734
rect 17816 33598 17822 33662
rect 17886 33598 18028 33662
rect 17816 33592 18028 33598
rect 18224 33798 18436 33804
rect 18224 33734 18230 33798
rect 18294 33734 18436 33798
rect 18224 33668 18436 33734
rect 18632 33798 18980 33804
rect 18632 33734 18638 33798
rect 18702 33734 18980 33798
rect 18224 33662 18572 33668
rect 18224 33598 18502 33662
rect 18566 33598 18572 33662
rect 18224 33592 18572 33598
rect 18224 33532 18436 33592
rect 18632 33532 18980 33734
rect 19040 33662 19252 33804
rect 19040 33598 19182 33662
rect 19246 33598 19252 33662
rect 19040 33592 19252 33598
rect 19448 33662 19660 33804
rect 19448 33598 19590 33662
rect 19654 33598 19660 33662
rect 19448 33592 19660 33598
rect 24344 33798 24692 33940
rect 24344 33734 24486 33798
rect 24550 33734 24622 33798
rect 24686 33734 24692 33798
rect 24344 33592 24692 33734
rect 66368 33934 66580 33940
rect 66368 33870 66510 33934
rect 66574 33870 66580 33934
rect 66368 33798 66580 33870
rect 71264 33864 71476 34212
rect 71400 33804 71476 33864
rect 66368 33734 66374 33798
rect 66438 33734 66580 33798
rect 66368 33592 66580 33734
rect 71264 33662 71476 33804
rect 71264 33598 71406 33662
rect 71470 33598 71476 33662
rect 71264 33592 71476 33598
rect 71672 33864 71884 34212
rect 72080 34000 72292 34212
rect 72352 34212 72428 34272
rect 72352 34136 72700 34212
rect 72488 34070 72700 34136
rect 72488 34006 72630 34070
rect 72694 34006 72700 34070
rect 72488 34000 72700 34006
rect 72896 34206 73108 34212
rect 72896 34142 73038 34206
rect 73102 34142 73108 34206
rect 72896 34070 73108 34142
rect 72896 34006 72902 34070
rect 72966 34006 73108 34070
rect 72896 34000 73108 34006
rect 89080 34070 89836 34076
rect 89080 34052 89766 34070
rect 89080 33996 89216 34052
rect 89272 34006 89766 34052
rect 89830 34006 89836 34070
rect 89272 34000 89836 34006
rect 89272 33996 89428 34000
rect 89080 33864 89428 33996
rect 71672 33804 71748 33864
rect 71672 33662 71884 33804
rect 71672 33598 71814 33662
rect 71878 33598 71884 33662
rect 71672 33592 71884 33598
rect 24480 33532 24556 33592
rect 66368 33532 66444 33592
rect 18224 33456 18980 33532
rect 24344 33526 24692 33532
rect 24344 33462 24486 33526
rect 24550 33462 24692 33526
rect 18224 33396 18300 33456
rect 17816 33390 18028 33396
rect 17816 33326 17822 33390
rect 17886 33326 18028 33390
rect 0 33233 10820 33260
rect 0 33184 10676 33233
rect 10608 33177 10676 33184
rect 10732 33177 10820 33233
rect 17816 33254 18028 33326
rect 17816 33190 17958 33254
rect 18022 33190 18028 33254
rect 17816 33184 18028 33190
rect 18224 33184 18436 33396
rect 18534 33390 18980 33396
rect 18496 33326 18502 33390
rect 18566 33326 18980 33390
rect 18534 33320 18980 33326
rect 18632 33254 18980 33320
rect 18632 33190 18638 33254
rect 18702 33190 18980 33254
rect 18632 33184 18980 33190
rect 19040 33390 19252 33396
rect 19040 33326 19182 33390
rect 19246 33326 19252 33390
rect 19040 33254 19252 33326
rect 19040 33190 19046 33254
rect 19110 33190 19252 33254
rect 19040 33184 19252 33190
rect 19448 33390 19660 33396
rect 19448 33326 19590 33390
rect 19654 33326 19660 33390
rect 19448 33254 19660 33326
rect 19448 33190 19590 33254
rect 19654 33190 19660 33254
rect 19448 33184 19660 33190
rect 24344 33320 24692 33462
rect 66368 33526 66580 33532
rect 66368 33462 66374 33526
rect 66438 33462 66580 33526
rect 66368 33320 66580 33462
rect 72080 33456 72292 33804
rect 72488 33798 72700 33804
rect 72488 33734 72630 33798
rect 72694 33734 72700 33798
rect 72488 33532 72700 33734
rect 72896 33798 73108 33804
rect 72896 33734 72902 33798
rect 72966 33734 73108 33798
rect 72896 33662 73108 33734
rect 72896 33598 72902 33662
rect 72966 33598 73108 33662
rect 72896 33592 73108 33598
rect 72390 33526 72700 33532
rect 72352 33462 72358 33526
rect 72422 33462 72700 33526
rect 72390 33456 72700 33462
rect 72216 33396 72292 33456
rect 24344 33260 24420 33320
rect 66504 33260 66580 33320
rect 10608 33048 10820 33177
rect 11616 33164 11682 33167
rect 12110 33164 12176 33167
rect 11616 33162 12176 33164
rect 11616 33106 11621 33162
rect 11677 33106 12115 33162
rect 12171 33106 12176 33162
rect 11616 33104 12176 33106
rect 11616 33101 11682 33104
rect 12110 33101 12176 33104
rect 17816 32982 18028 32988
rect 17816 32918 17958 32982
rect 18022 32918 18028 32982
rect 17816 32846 18028 32918
rect 17816 32782 17822 32846
rect 17886 32782 18028 32846
rect 17816 32776 18028 32782
rect 18224 32846 18436 32988
rect 18224 32782 18366 32846
rect 18430 32782 18436 32846
rect 18224 32776 18436 32782
rect 18632 32982 18980 32988
rect 18632 32918 18638 32982
rect 18702 32918 18980 32982
rect 18632 32776 18980 32918
rect 19040 32982 19252 32988
rect 19040 32918 19046 32982
rect 19110 32918 19252 32982
rect 19040 32846 19252 32918
rect 19040 32782 19182 32846
rect 19246 32782 19252 32846
rect 19040 32776 19252 32782
rect 19448 32982 19660 32988
rect 19448 32918 19590 32982
rect 19654 32918 19660 32982
rect 19448 32846 19660 32918
rect 19448 32782 19454 32846
rect 19518 32782 19660 32846
rect 19448 32776 19660 32782
rect 24344 32776 24692 33260
rect 18632 32716 18708 32776
rect 24616 32716 24692 32776
rect 18360 32640 18708 32716
rect 18360 32580 18436 32640
rect 17816 32574 18028 32580
rect 17816 32510 17822 32574
rect 17886 32510 18028 32574
rect 1632 32372 1844 32444
rect 1632 32316 1718 32372
rect 1774 32316 1844 32372
rect 1632 32308 1844 32316
rect 1224 32302 1844 32308
rect 1224 32238 1230 32302
rect 1294 32238 1844 32302
rect 1224 32232 1844 32238
rect 11016 32438 11228 32444
rect 11016 32374 11022 32438
rect 11086 32374 11228 32438
rect 11016 32302 11228 32374
rect 17816 32438 18028 32510
rect 17816 32374 17958 32438
rect 18022 32374 18028 32438
rect 17816 32368 18028 32374
rect 18224 32574 18980 32580
rect 18224 32510 18366 32574
rect 18430 32510 18980 32574
rect 18224 32504 18980 32510
rect 18224 32438 18436 32504
rect 18224 32374 18366 32438
rect 18430 32374 18436 32438
rect 18224 32368 18436 32374
rect 18632 32438 18980 32504
rect 18632 32374 18774 32438
rect 18838 32374 18980 32438
rect 18632 32368 18980 32374
rect 19040 32574 19252 32580
rect 19040 32510 19182 32574
rect 19246 32510 19252 32574
rect 19040 32438 19252 32510
rect 19040 32374 19182 32438
rect 19246 32374 19252 32438
rect 19040 32368 19252 32374
rect 19448 32574 19660 32580
rect 19448 32510 19454 32574
rect 19518 32510 19660 32574
rect 19448 32438 19660 32510
rect 24344 32504 24692 32716
rect 24616 32444 24692 32504
rect 19448 32374 19590 32438
rect 19654 32374 19660 32438
rect 19448 32368 19660 32374
rect 11016 32238 11022 32302
rect 11086 32238 11228 32302
rect 11016 32232 11228 32238
rect 24344 32232 24692 32444
rect 66368 32982 66580 33260
rect 71264 33390 71476 33396
rect 71264 33326 71406 33390
rect 71470 33326 71476 33390
rect 71264 33254 71476 33326
rect 71264 33190 71270 33254
rect 71334 33190 71476 33254
rect 71264 33184 71476 33190
rect 71672 33390 71884 33396
rect 71672 33326 71814 33390
rect 71878 33326 71884 33390
rect 71672 33254 71884 33326
rect 71672 33190 71814 33254
rect 71878 33190 71884 33254
rect 71672 33184 71884 33190
rect 72080 33320 72700 33396
rect 72080 33260 72292 33320
rect 72080 33254 72428 33260
rect 72080 33190 72358 33254
rect 72422 33190 72428 33254
rect 72080 33184 72428 33190
rect 72488 33254 72700 33320
rect 72488 33190 72630 33254
rect 72694 33190 72700 33254
rect 72488 33184 72700 33190
rect 72896 33390 73108 33396
rect 72896 33326 72902 33390
rect 72966 33326 73108 33390
rect 72896 33254 73108 33326
rect 72896 33190 73038 33254
rect 73102 33190 73108 33254
rect 72896 33184 73108 33190
rect 66368 32918 66374 32982
rect 66438 32918 66580 32982
rect 66368 32776 66580 32918
rect 71264 32982 71476 32988
rect 71264 32918 71270 32982
rect 71334 32918 71476 32982
rect 71264 32846 71476 32918
rect 71264 32782 71406 32846
rect 71470 32782 71476 32846
rect 71264 32776 71476 32782
rect 71672 32982 71884 32988
rect 71672 32918 71814 32982
rect 71878 32918 71884 32982
rect 71672 32846 71884 32918
rect 71672 32782 71678 32846
rect 71742 32782 71884 32846
rect 71672 32776 71884 32782
rect 72080 32982 72700 32988
rect 72080 32918 72630 32982
rect 72694 32918 72700 32982
rect 72080 32912 72700 32918
rect 72080 32852 72292 32912
rect 72080 32846 72428 32852
rect 72080 32782 72358 32846
rect 72422 32782 72428 32846
rect 72080 32776 72428 32782
rect 72488 32776 72700 32912
rect 72896 32982 73108 32988
rect 72896 32918 73038 32982
rect 73102 32918 73108 32982
rect 72896 32846 73108 32918
rect 72896 32782 72902 32846
rect 72966 32782 73108 32846
rect 72896 32776 73108 32782
rect 66368 32716 66444 32776
rect 66368 32710 66580 32716
rect 66368 32646 66374 32710
rect 66438 32646 66580 32710
rect 66368 32504 66580 32646
rect 71264 32574 71476 32580
rect 71264 32510 71406 32574
rect 71470 32510 71476 32574
rect 66368 32444 66444 32504
rect 66368 32232 66580 32444
rect 71264 32438 71476 32510
rect 71264 32374 71406 32438
rect 71470 32374 71476 32438
rect 71264 32368 71476 32374
rect 71672 32574 71884 32580
rect 71672 32510 71678 32574
rect 71742 32510 71884 32574
rect 71672 32438 71884 32510
rect 71672 32374 71814 32438
rect 71878 32374 71884 32438
rect 71672 32368 71884 32374
rect 72080 32438 72292 32580
rect 72390 32574 72700 32580
rect 72352 32510 72358 32574
rect 72422 32510 72700 32574
rect 72390 32504 72700 32510
rect 72080 32374 72086 32438
rect 72150 32374 72292 32438
rect 72080 32368 72292 32374
rect 72488 32438 72700 32504
rect 72488 32374 72630 32438
rect 72694 32374 72700 32438
rect 72488 32368 72700 32374
rect 72896 32574 73108 32580
rect 72896 32510 72902 32574
rect 72966 32510 73108 32574
rect 72896 32438 73108 32510
rect 72896 32374 73038 32438
rect 73102 32374 73108 32438
rect 72896 32368 73108 32374
rect 89080 32438 89836 32444
rect 89080 32374 89766 32438
rect 89830 32374 89836 32438
rect 89080 32372 89836 32374
rect 89080 32316 89216 32372
rect 89272 32368 89836 32372
rect 89272 32316 89428 32368
rect 89080 32232 89428 32316
rect 24616 32172 24692 32232
rect 66504 32172 66580 32232
rect 17816 32166 18028 32172
rect 17816 32102 17958 32166
rect 18022 32102 18028 32166
rect 17816 32030 18028 32102
rect 17816 31966 17958 32030
rect 18022 31966 18028 32030
rect 17816 31960 18028 31966
rect 18224 32166 18436 32172
rect 18224 32102 18366 32166
rect 18430 32102 18436 32166
rect 18224 31960 18436 32102
rect 18632 32166 18980 32172
rect 18632 32102 18774 32166
rect 18838 32102 18980 32166
rect 18632 32036 18980 32102
rect 18534 32030 18980 32036
rect 18496 31966 18502 32030
rect 18566 31966 18980 32030
rect 18534 31960 18980 31966
rect 19040 32166 19252 32172
rect 19040 32102 19182 32166
rect 19246 32102 19252 32166
rect 19040 32030 19252 32102
rect 19040 31966 19046 32030
rect 19110 31966 19252 32030
rect 19040 31960 19252 31966
rect 19448 32166 19660 32172
rect 19448 32102 19590 32166
rect 19654 32102 19660 32166
rect 19448 32030 19660 32102
rect 19448 31966 19454 32030
rect 19518 31966 19660 32030
rect 19448 31960 19660 31966
rect 24344 31960 24692 32172
rect 66368 31960 66580 32172
rect 71264 32166 71476 32172
rect 71264 32102 71406 32166
rect 71470 32102 71476 32166
rect 71264 32030 71476 32102
rect 71264 31966 71406 32030
rect 71470 31966 71476 32030
rect 71264 31960 71476 31966
rect 71672 32166 71884 32172
rect 71672 32102 71814 32166
rect 71878 32102 71884 32166
rect 71672 32030 71884 32102
rect 71672 31966 71678 32030
rect 71742 31966 71884 32030
rect 71672 31960 71884 31966
rect 72080 32166 72700 32172
rect 72080 32102 72086 32166
rect 72150 32102 72630 32166
rect 72694 32102 72700 32166
rect 72080 32096 72700 32102
rect 72080 31960 72292 32096
rect 72488 32030 72700 32096
rect 72488 31966 72494 32030
rect 72558 31966 72700 32030
rect 72488 31960 72700 31966
rect 72896 32166 73108 32172
rect 72896 32102 73038 32166
rect 73102 32102 73108 32166
rect 72896 32030 73108 32102
rect 72896 31966 73038 32030
rect 73102 31966 73108 32030
rect 72896 31960 73108 31966
rect 24480 31900 24556 31960
rect 66504 31900 66580 31960
rect 17816 31758 18028 31764
rect 17816 31694 17958 31758
rect 18022 31694 18028 31758
rect 0 31552 10820 31628
rect 10608 31533 10820 31552
rect 11616 31606 11682 31609
rect 12030 31606 12096 31609
rect 11616 31604 12096 31606
rect 11616 31548 11621 31604
rect 11677 31548 12035 31604
rect 12091 31548 12096 31604
rect 17816 31552 18028 31694
rect 18224 31758 18572 31764
rect 18224 31694 18502 31758
rect 18566 31694 18572 31758
rect 18224 31688 18572 31694
rect 18224 31628 18436 31688
rect 18632 31628 18980 31764
rect 18224 31622 18980 31628
rect 18224 31558 18366 31622
rect 18430 31558 18980 31622
rect 18224 31552 18980 31558
rect 19040 31758 19252 31764
rect 19040 31694 19046 31758
rect 19110 31694 19252 31758
rect 19040 31622 19252 31694
rect 19040 31558 19182 31622
rect 19246 31558 19252 31622
rect 19040 31552 19252 31558
rect 19448 31758 19660 31764
rect 19448 31694 19454 31758
rect 19518 31694 19660 31758
rect 19448 31622 19660 31694
rect 24344 31688 24692 31900
rect 66368 31688 66580 31900
rect 71264 31758 71476 31764
rect 71264 31694 71406 31758
rect 71470 31694 71476 31758
rect 24480 31628 24556 31688
rect 66368 31628 66444 31688
rect 19448 31558 19454 31622
rect 19518 31558 19660 31622
rect 19448 31552 19660 31558
rect 11616 31546 12096 31548
rect 11616 31543 11682 31546
rect 12030 31543 12096 31546
rect 10608 31477 10676 31533
rect 10732 31477 10820 31533
rect 17952 31492 18028 31552
rect 10608 31416 10820 31477
rect 17816 31144 18028 31492
rect 18360 31492 18436 31552
rect 18360 31416 18708 31492
rect 24344 31486 24692 31628
rect 24344 31422 24486 31486
rect 24550 31422 24692 31486
rect 24344 31416 24692 31422
rect 18632 31356 18708 31416
rect 24616 31356 24692 31416
rect 18224 31350 18436 31356
rect 18224 31286 18366 31350
rect 18430 31286 18436 31350
rect 18224 31220 18436 31286
rect 18224 31144 18572 31220
rect 18632 31144 18980 31356
rect 19040 31350 19252 31356
rect 19040 31286 19182 31350
rect 19246 31286 19252 31350
rect 19040 31214 19252 31286
rect 19040 31150 19046 31214
rect 19110 31150 19252 31214
rect 19040 31144 19252 31150
rect 19448 31350 19660 31356
rect 19448 31286 19454 31350
rect 19518 31286 19660 31350
rect 19448 31214 19660 31286
rect 19448 31150 19454 31214
rect 19518 31150 19660 31214
rect 19448 31144 19660 31150
rect 24344 31214 24692 31356
rect 24344 31150 24486 31214
rect 24550 31150 24692 31214
rect 17816 31084 17892 31144
rect 18224 31084 18300 31144
rect 18496 31084 18572 31144
rect 11016 31078 11228 31084
rect 11016 31014 11158 31078
rect 11222 31014 11228 31078
rect 11016 30942 11228 31014
rect 11016 30878 11158 30942
rect 11222 30878 11228 30942
rect 11016 30872 11228 30878
rect 1224 30806 1844 30812
rect 1224 30742 1230 30806
rect 1294 30742 1844 30806
rect 1224 30736 1844 30742
rect 1632 30692 1844 30736
rect 1632 30636 1718 30692
rect 1774 30636 1844 30692
rect 1632 30600 1844 30636
rect 17816 30736 18028 31084
rect 18224 30736 18436 31084
rect 18496 31008 18980 31084
rect 18632 30812 18980 31008
rect 18534 30806 18980 30812
rect 18496 30742 18502 30806
rect 18566 30742 18980 30806
rect 18534 30736 18980 30742
rect 19040 30942 19252 30948
rect 19040 30878 19046 30942
rect 19110 30878 19252 30942
rect 19040 30806 19252 30878
rect 19040 30742 19182 30806
rect 19246 30742 19252 30806
rect 19040 30736 19252 30742
rect 19448 30942 19660 30948
rect 19448 30878 19454 30942
rect 19518 30878 19660 30942
rect 19448 30806 19660 30878
rect 19448 30742 19590 30806
rect 19654 30742 19660 30806
rect 19448 30736 19660 30742
rect 24344 30872 24692 31150
rect 66368 31416 66580 31628
rect 71264 31622 71476 31694
rect 71264 31558 71406 31622
rect 71470 31558 71476 31622
rect 71264 31552 71476 31558
rect 71672 31758 71884 31764
rect 71672 31694 71678 31758
rect 71742 31694 71884 31758
rect 71672 31622 71884 31694
rect 71672 31558 71678 31622
rect 71742 31558 71884 31622
rect 71672 31552 71884 31558
rect 72080 31758 72700 31764
rect 72080 31694 72494 31758
rect 72558 31694 72700 31758
rect 72080 31688 72700 31694
rect 72080 31622 72292 31688
rect 72080 31558 72086 31622
rect 72150 31558 72292 31622
rect 72080 31552 72292 31558
rect 72488 31552 72700 31688
rect 72896 31758 73108 31764
rect 72896 31694 73038 31758
rect 73102 31694 73108 31758
rect 72896 31552 73108 31694
rect 72896 31492 72972 31552
rect 66368 31356 66444 31416
rect 66368 30872 66580 31356
rect 71264 31350 71476 31356
rect 71264 31286 71406 31350
rect 71470 31286 71476 31350
rect 71264 31214 71476 31286
rect 71264 31150 71270 31214
rect 71334 31150 71476 31214
rect 71264 31144 71476 31150
rect 71672 31350 71884 31356
rect 71672 31286 71678 31350
rect 71742 31286 71884 31350
rect 71672 31214 71884 31286
rect 71672 31150 71814 31214
rect 71878 31150 71884 31214
rect 71672 31144 71884 31150
rect 72080 31350 72292 31356
rect 72080 31286 72086 31350
rect 72150 31286 72292 31350
rect 72080 31220 72292 31286
rect 72488 31220 72700 31356
rect 72080 31144 72700 31220
rect 72896 31144 73108 31492
rect 72216 31084 72292 31144
rect 72624 31084 72700 31144
rect 73032 31084 73108 31144
rect 24344 30812 24420 30872
rect 66504 30812 66580 30872
rect 17816 30676 17892 30736
rect 10608 30405 10820 30540
rect 17816 30534 18028 30676
rect 18360 30600 18708 30676
rect 24344 30670 24692 30812
rect 24344 30606 24622 30670
rect 24686 30606 24692 30670
rect 24344 30600 24692 30606
rect 66368 30600 66580 30812
rect 71264 30942 71476 30948
rect 71264 30878 71270 30942
rect 71334 30878 71476 30942
rect 71264 30806 71476 30878
rect 71264 30742 71406 30806
rect 71470 30742 71476 30806
rect 71264 30736 71476 30742
rect 71672 30942 71884 30948
rect 71672 30878 71814 30942
rect 71878 30878 71884 30942
rect 71672 30806 71884 30878
rect 71672 30742 71814 30806
rect 71878 30742 71884 30806
rect 71672 30736 71884 30742
rect 72080 30806 72292 31084
rect 72080 30742 72086 30806
rect 72150 30742 72292 30806
rect 72080 30736 72292 30742
rect 72488 30736 72700 31084
rect 72896 30736 73108 31084
rect 73032 30676 73108 30736
rect 18360 30540 18436 30600
rect 18632 30540 18708 30600
rect 24480 30540 24556 30600
rect 66368 30540 66444 30600
rect 17816 30470 17822 30534
rect 17886 30470 18028 30534
rect 17816 30464 18028 30470
rect 18224 30534 18572 30540
rect 18224 30470 18502 30534
rect 18566 30470 18572 30534
rect 18224 30464 18572 30470
rect 10608 30349 10676 30405
rect 10732 30349 10820 30405
rect 10608 30268 10820 30349
rect 18224 30404 18436 30464
rect 11616 30336 11682 30339
rect 11950 30336 12016 30339
rect 11616 30334 12016 30336
rect 11616 30278 11621 30334
rect 11677 30278 11955 30334
rect 12011 30278 12016 30334
rect 18224 30328 18572 30404
rect 18632 30328 18980 30540
rect 19040 30534 19252 30540
rect 19040 30470 19182 30534
rect 19246 30470 19252 30534
rect 19040 30328 19252 30470
rect 11616 30276 12016 30278
rect 11616 30273 11682 30276
rect 11950 30273 12016 30276
rect 18360 30268 18436 30328
rect 0 30192 10820 30268
rect 17816 30262 18028 30268
rect 17816 30198 17822 30262
rect 17886 30198 18028 30262
rect 17816 30126 18028 30198
rect 17816 30062 17822 30126
rect 17886 30062 18028 30126
rect 17816 30056 18028 30062
rect 18224 30056 18436 30268
rect 18496 30268 18572 30328
rect 19176 30268 19252 30328
rect 18496 30192 18980 30268
rect 18632 30126 18980 30192
rect 18632 30062 18638 30126
rect 18702 30062 18980 30126
rect 18632 30056 18980 30062
rect 19040 29920 19252 30268
rect 19448 30534 19660 30540
rect 19448 30470 19590 30534
rect 19654 30470 19660 30534
rect 19448 30328 19660 30470
rect 24344 30398 24692 30540
rect 24344 30334 24622 30398
rect 24686 30334 24692 30398
rect 19448 30268 19524 30328
rect 19448 29920 19660 30268
rect 24344 30262 24692 30334
rect 24344 30198 24486 30262
rect 24550 30198 24692 30262
rect 24344 30192 24692 30198
rect 66368 30262 66580 30540
rect 71264 30534 71476 30540
rect 71264 30470 71406 30534
rect 71470 30470 71476 30534
rect 71264 30328 71476 30470
rect 71672 30534 71884 30540
rect 71672 30470 71814 30534
rect 71878 30470 71884 30534
rect 71672 30328 71884 30470
rect 71400 30268 71476 30328
rect 71808 30268 71884 30328
rect 66368 30198 66374 30262
rect 66438 30198 66580 30262
rect 66368 30192 66580 30198
rect 24344 29990 24692 29996
rect 24344 29926 24486 29990
rect 24550 29926 24692 29990
rect 19040 29860 19116 29920
rect 19448 29860 19524 29920
rect 17816 29854 18028 29860
rect 17816 29790 17822 29854
rect 17886 29790 18028 29854
rect 17816 29718 18028 29790
rect 17816 29654 17822 29718
rect 17886 29654 18028 29718
rect 17816 29648 18028 29654
rect 11016 29582 11228 29588
rect 11016 29518 11022 29582
rect 11086 29518 11228 29582
rect 11016 29452 11228 29518
rect 18224 29512 18436 29860
rect 18632 29854 18980 29860
rect 18632 29790 18638 29854
rect 18702 29790 18980 29854
rect 18632 29588 18980 29790
rect 18360 29452 18436 29512
rect 18496 29512 18980 29588
rect 19040 29512 19252 29860
rect 18496 29452 18572 29512
rect 11016 29446 14900 29452
rect 11016 29382 14830 29446
rect 14894 29382 14900 29446
rect 11016 29376 14900 29382
rect 17816 29446 18028 29452
rect 17816 29382 17822 29446
rect 17886 29382 18028 29446
rect 17816 29310 18028 29382
rect 17816 29246 17822 29310
rect 17886 29246 18028 29310
rect 17816 29240 18028 29246
rect 18224 29376 18572 29452
rect 18632 29452 18708 29512
rect 19176 29452 19252 29512
rect 18224 29240 18436 29376
rect 18632 29310 18980 29452
rect 18632 29246 18774 29310
rect 18838 29246 18980 29310
rect 18632 29240 18980 29246
rect 19040 29310 19252 29452
rect 19040 29246 19046 29310
rect 19110 29246 19252 29310
rect 19040 29240 19252 29246
rect 19448 29512 19660 29860
rect 19448 29452 19524 29512
rect 19448 29310 19660 29452
rect 24344 29376 24692 29926
rect 24616 29316 24692 29376
rect 19448 29246 19454 29310
rect 19518 29246 19660 29310
rect 19448 29240 19660 29246
rect 1632 29012 1844 29044
rect 1632 28956 1718 29012
rect 1774 28956 1844 29012
rect 1632 28908 1844 28956
rect 1224 28902 1844 28908
rect 1224 28838 1230 28902
rect 1294 28838 1844 28902
rect 1224 28832 1844 28838
rect 17816 29038 18028 29044
rect 17816 28974 17822 29038
rect 17886 28974 18028 29038
rect 17816 28902 18028 28974
rect 17816 28838 17822 28902
rect 17886 28838 18028 28902
rect 17816 28832 18028 28838
rect 18224 28902 18436 29044
rect 18632 29038 18980 29044
rect 18632 28974 18774 29038
rect 18838 28974 18980 29038
rect 18632 28908 18980 28974
rect 18534 28902 18980 28908
rect 18224 28838 18230 28902
rect 18294 28838 18436 28902
rect 18496 28838 18502 28902
rect 18566 28838 18980 28902
rect 18224 28832 18436 28838
rect 18534 28832 18980 28838
rect 19040 29038 19252 29044
rect 19040 28974 19046 29038
rect 19110 28974 19252 29038
rect 19040 28902 19252 28974
rect 19040 28838 19046 28902
rect 19110 28838 19252 28902
rect 19040 28832 19252 28838
rect 19448 29038 19660 29044
rect 19448 28974 19454 29038
rect 19518 28974 19660 29038
rect 19448 28902 19660 28974
rect 19448 28838 19590 28902
rect 19654 28838 19660 28902
rect 19448 28832 19660 28838
rect 24344 28832 24692 29316
rect 66368 29990 66580 29996
rect 66368 29926 66374 29990
rect 66438 29926 66580 29990
rect 66368 29854 66580 29926
rect 71264 29920 71476 30268
rect 71672 29920 71884 30268
rect 72080 30534 72292 30540
rect 72080 30470 72086 30534
rect 72150 30470 72292 30534
rect 72080 30328 72292 30470
rect 72488 30404 72700 30540
rect 72896 30534 73108 30676
rect 89080 30692 89428 30812
rect 89080 30636 89216 30692
rect 89272 30676 89428 30692
rect 89272 30670 89836 30676
rect 89272 30636 89766 30670
rect 89080 30606 89766 30636
rect 89830 30606 89836 30670
rect 89080 30600 89836 30606
rect 72896 30470 72902 30534
rect 72966 30470 73108 30534
rect 72896 30464 73108 30470
rect 72352 30328 72700 30404
rect 72080 30268 72156 30328
rect 72352 30268 72428 30328
rect 72080 30192 72428 30268
rect 72488 30268 72564 30328
rect 72080 30126 72292 30192
rect 72080 30062 72222 30126
rect 72286 30062 72292 30126
rect 72080 30056 72292 30062
rect 72488 30126 72700 30268
rect 72488 30062 72630 30126
rect 72694 30062 72700 30126
rect 72488 30056 72700 30062
rect 72896 30262 73108 30268
rect 72896 30198 72902 30262
rect 72966 30198 73108 30262
rect 72896 30126 73108 30198
rect 72896 30062 73038 30126
rect 73102 30062 73108 30126
rect 72896 30056 73108 30062
rect 71400 29860 71476 29920
rect 71808 29860 71884 29920
rect 66368 29790 66510 29854
rect 66574 29790 66580 29854
rect 66368 29582 66580 29790
rect 66368 29518 66510 29582
rect 66574 29518 66580 29582
rect 66368 29376 66580 29518
rect 71264 29512 71476 29860
rect 71400 29452 71476 29512
rect 66368 29316 66444 29376
rect 66368 29038 66580 29316
rect 71264 29310 71476 29452
rect 71264 29246 71406 29310
rect 71470 29246 71476 29310
rect 71264 29240 71476 29246
rect 71672 29512 71884 29860
rect 72080 29854 72292 29860
rect 72080 29790 72222 29854
rect 72286 29790 72292 29854
rect 72080 29512 72292 29790
rect 72488 29854 72700 29860
rect 72488 29790 72630 29854
rect 72694 29790 72700 29854
rect 72488 29512 72700 29790
rect 72896 29854 73108 29860
rect 72896 29790 73038 29854
rect 73102 29790 73108 29854
rect 72896 29718 73108 29790
rect 72896 29654 73038 29718
rect 73102 29654 73108 29718
rect 72896 29648 73108 29654
rect 71672 29452 71748 29512
rect 72080 29452 72156 29512
rect 72488 29452 72564 29512
rect 71672 29310 71884 29452
rect 71672 29246 71814 29310
rect 71878 29246 71884 29310
rect 71672 29240 71884 29246
rect 72080 29240 72292 29452
rect 72488 29240 72700 29452
rect 72896 29446 73108 29452
rect 72896 29382 73038 29446
rect 73102 29382 73108 29446
rect 72896 29310 73108 29382
rect 72896 29246 73038 29310
rect 73102 29246 73108 29310
rect 72896 29240 73108 29246
rect 72488 29180 72564 29240
rect 72216 29104 72564 29180
rect 72216 29044 72292 29104
rect 66368 28974 66510 29038
rect 66574 28974 66580 29038
rect 66368 28832 66580 28974
rect 71264 29038 71476 29044
rect 71264 28974 71406 29038
rect 71470 28974 71476 29038
rect 71264 28902 71476 28974
rect 71264 28838 71270 28902
rect 71334 28838 71476 28902
rect 71264 28832 71476 28838
rect 71672 29038 71884 29044
rect 71672 28974 71814 29038
rect 71878 28974 71884 29038
rect 71672 28902 71884 28974
rect 71672 28838 71814 28902
rect 71878 28838 71884 28902
rect 71672 28832 71884 28838
rect 72080 28968 72700 29044
rect 72080 28832 72292 28968
rect 72488 28902 72700 28968
rect 72488 28838 72494 28902
rect 72558 28838 72700 28902
rect 72488 28832 72700 28838
rect 72896 29038 73108 29044
rect 72896 28974 73038 29038
rect 73102 28974 73108 29038
rect 72896 28902 73108 28974
rect 72896 28838 73038 28902
rect 73102 28838 73108 28902
rect 72896 28832 73108 28838
rect 89080 29038 89836 29044
rect 89080 29012 89766 29038
rect 89080 28956 89216 29012
rect 89272 28974 89766 29012
rect 89830 28974 89836 29038
rect 89272 28968 89836 28974
rect 89272 28956 89428 28968
rect 89080 28832 89428 28956
rect 11616 28778 11682 28781
rect 11870 28778 11936 28781
rect 11616 28776 11936 28778
rect 10608 28705 10820 28772
rect 11616 28720 11621 28776
rect 11677 28720 11875 28776
rect 11931 28720 11936 28776
rect 11616 28718 11936 28720
rect 11616 28715 11682 28718
rect 11870 28715 11936 28718
rect 24344 28772 24420 28832
rect 66504 28772 66580 28832
rect 10608 28649 10676 28705
rect 10732 28649 10820 28705
rect 10608 28636 10820 28649
rect 0 28560 10820 28636
rect 17816 28630 18028 28636
rect 17816 28566 17822 28630
rect 17886 28566 18028 28630
rect 17816 28494 18028 28566
rect 11702 28454 11786 28458
rect 11702 28449 11819 28454
rect 11702 28393 11758 28449
rect 11814 28393 11819 28449
rect 17816 28430 17822 28494
rect 17886 28430 18028 28494
rect 17816 28424 18028 28430
rect 18224 28630 18572 28636
rect 18224 28566 18230 28630
rect 18294 28566 18502 28630
rect 18566 28566 18572 28630
rect 18224 28560 18572 28566
rect 18224 28500 18436 28560
rect 18632 28500 18980 28636
rect 18224 28494 18980 28500
rect 18224 28430 18366 28494
rect 18430 28430 18980 28494
rect 18224 28424 18980 28430
rect 19040 28630 19252 28636
rect 19040 28566 19046 28630
rect 19110 28566 19252 28630
rect 19040 28494 19252 28566
rect 19040 28430 19182 28494
rect 19246 28430 19252 28494
rect 19040 28424 19252 28430
rect 19448 28630 19660 28636
rect 19448 28566 19590 28630
rect 19654 28566 19660 28630
rect 19448 28494 19660 28566
rect 24344 28560 24692 28772
rect 66368 28766 66580 28772
rect 66368 28702 66510 28766
rect 66574 28702 66580 28766
rect 66368 28560 66580 28702
rect 71264 28630 71476 28636
rect 71264 28566 71270 28630
rect 71334 28566 71476 28630
rect 24480 28500 24556 28560
rect 66368 28500 66444 28560
rect 19448 28430 19590 28494
rect 19654 28430 19660 28494
rect 19448 28424 19660 28430
rect 11702 28388 11819 28393
rect 11702 28384 11786 28388
rect 18360 28364 18436 28424
rect 18360 28288 18708 28364
rect 24344 28288 24692 28500
rect 18632 28228 18708 28288
rect 24616 28228 24692 28288
rect 11016 28222 11228 28228
rect 11016 28158 11158 28222
rect 11222 28158 11228 28222
rect 11016 28092 11228 28158
rect 17816 28222 18028 28228
rect 17816 28158 17822 28222
rect 17886 28158 18028 28222
rect 11016 28086 12996 28092
rect 11016 28022 12926 28086
rect 12990 28022 12996 28086
rect 11016 28016 12996 28022
rect 17816 28086 18028 28158
rect 17816 28022 17822 28086
rect 17886 28022 18028 28086
rect 17816 28016 18028 28022
rect 18224 28222 18436 28228
rect 18224 28158 18366 28222
rect 18430 28158 18436 28222
rect 18224 28086 18436 28158
rect 18224 28022 18230 28086
rect 18294 28022 18436 28086
rect 18224 28016 18436 28022
rect 18632 28086 18980 28228
rect 18632 28022 18774 28086
rect 18838 28022 18980 28086
rect 18632 28016 18980 28022
rect 19040 28222 19252 28228
rect 19040 28158 19182 28222
rect 19246 28158 19252 28222
rect 19040 28086 19252 28158
rect 19040 28022 19046 28086
rect 19110 28022 19252 28086
rect 19040 28016 19252 28022
rect 19448 28222 19660 28228
rect 19448 28158 19590 28222
rect 19654 28158 19660 28222
rect 19448 28086 19660 28158
rect 19448 28022 19590 28086
rect 19654 28022 19660 28086
rect 19448 28016 19660 28022
rect 24344 28016 24692 28228
rect 66368 28288 66580 28500
rect 71264 28494 71476 28566
rect 71264 28430 71406 28494
rect 71470 28430 71476 28494
rect 71264 28424 71476 28430
rect 71672 28630 71884 28636
rect 71672 28566 71814 28630
rect 71878 28566 71884 28630
rect 71672 28494 71884 28566
rect 71672 28430 71678 28494
rect 71742 28430 71884 28494
rect 71672 28424 71884 28430
rect 72080 28494 72292 28636
rect 72080 28430 72086 28494
rect 72150 28430 72292 28494
rect 72080 28424 72292 28430
rect 72488 28630 72700 28636
rect 72488 28566 72494 28630
rect 72558 28566 72700 28630
rect 72488 28494 72700 28566
rect 72488 28430 72494 28494
rect 72558 28430 72700 28494
rect 72488 28424 72700 28430
rect 72896 28630 73108 28636
rect 72896 28566 73038 28630
rect 73102 28566 73108 28630
rect 72896 28494 73108 28566
rect 72896 28430 72902 28494
rect 72966 28430 73108 28494
rect 72896 28424 73108 28430
rect 66368 28228 66444 28288
rect 66368 28016 66580 28228
rect 71264 28222 71476 28228
rect 71264 28158 71406 28222
rect 71470 28158 71476 28222
rect 71264 28086 71476 28158
rect 71264 28022 71270 28086
rect 71334 28022 71476 28086
rect 71264 28016 71476 28022
rect 71672 28222 71884 28228
rect 71672 28158 71678 28222
rect 71742 28158 71884 28222
rect 71672 28086 71884 28158
rect 71672 28022 71678 28086
rect 71742 28022 71884 28086
rect 71672 28016 71884 28022
rect 72080 28222 72292 28228
rect 72080 28158 72086 28222
rect 72150 28158 72292 28222
rect 72080 28086 72292 28158
rect 72080 28022 72222 28086
rect 72286 28022 72292 28086
rect 72080 28016 72292 28022
rect 72488 28222 72700 28228
rect 72488 28158 72494 28222
rect 72558 28158 72700 28222
rect 72488 28016 72700 28158
rect 72896 28222 73108 28228
rect 72896 28158 72902 28222
rect 72966 28158 73108 28222
rect 72896 28086 73108 28158
rect 72896 28022 72902 28086
rect 72966 28022 73108 28086
rect 72896 28016 73108 28022
rect 24344 27956 24420 28016
rect 66504 27956 66580 28016
rect 72488 27956 72564 28016
rect 14416 27678 14628 27820
rect 14416 27614 14558 27678
rect 14622 27614 14628 27678
rect 14416 27608 14628 27614
rect 14824 27814 15444 27820
rect 14824 27750 14830 27814
rect 14894 27750 15444 27814
rect 14824 27744 15444 27750
rect 14824 27608 15036 27744
rect 15232 27684 15444 27744
rect 15232 27678 15580 27684
rect 15232 27614 15374 27678
rect 15438 27614 15580 27678
rect 15232 27608 15580 27614
rect 15640 27678 15852 27820
rect 15640 27614 15782 27678
rect 15846 27614 15852 27678
rect 15640 27608 15852 27614
rect 16048 27608 16260 27820
rect 17816 27814 18028 27820
rect 17816 27750 17822 27814
rect 17886 27750 18028 27814
rect 17816 27608 18028 27750
rect 18224 27814 18436 27820
rect 18224 27750 18230 27814
rect 18294 27750 18436 27814
rect 18224 27608 18436 27750
rect 18632 27814 18980 27820
rect 18632 27750 18774 27814
rect 18838 27750 18980 27814
rect 18632 27684 18980 27750
rect 18534 27678 18980 27684
rect 18496 27614 18502 27678
rect 18566 27614 18774 27678
rect 18838 27614 18980 27678
rect 18534 27608 18980 27614
rect 19040 27814 19252 27820
rect 19040 27750 19046 27814
rect 19110 27750 19252 27814
rect 19040 27678 19252 27750
rect 19040 27614 19046 27678
rect 19110 27614 19252 27678
rect 19040 27608 19252 27614
rect 19448 27814 19660 27820
rect 19448 27750 19590 27814
rect 19654 27750 19660 27814
rect 19448 27678 19660 27750
rect 24344 27744 24692 27956
rect 66368 27744 66580 27956
rect 72216 27880 72564 27956
rect 74936 27880 75556 27956
rect 72216 27820 72292 27880
rect 74936 27820 75012 27880
rect 75480 27820 75556 27880
rect 24616 27684 24692 27744
rect 66504 27684 66580 27744
rect 19448 27614 19454 27678
rect 19518 27614 19660 27678
rect 19448 27608 19660 27614
rect 15504 27548 15580 27608
rect 16048 27548 16124 27608
rect 17952 27548 18028 27608
rect 15504 27472 16124 27548
rect 1632 27332 1844 27412
rect 1632 27276 1718 27332
rect 1774 27276 1844 27332
rect 1224 27270 1844 27276
rect 1224 27206 1230 27270
rect 1294 27206 1844 27270
rect 1224 27200 1844 27206
rect 17816 27270 18028 27548
rect 24344 27472 24692 27684
rect 66368 27472 66580 27684
rect 71264 27814 71476 27820
rect 71264 27750 71270 27814
rect 71334 27750 71476 27814
rect 71264 27678 71476 27750
rect 71264 27614 71270 27678
rect 71334 27614 71476 27678
rect 71264 27608 71476 27614
rect 71672 27814 71884 27820
rect 71672 27750 71678 27814
rect 71742 27750 71884 27814
rect 71672 27678 71884 27750
rect 71672 27614 71678 27678
rect 71742 27614 71884 27678
rect 71672 27608 71884 27614
rect 72080 27814 72700 27820
rect 72080 27750 72222 27814
rect 72286 27750 72700 27814
rect 72080 27744 72700 27750
rect 72080 27608 72292 27744
rect 72488 27678 72700 27744
rect 72488 27614 72630 27678
rect 72694 27614 72700 27678
rect 72488 27608 72700 27614
rect 72896 27814 73108 27820
rect 72896 27750 72902 27814
rect 72966 27750 73108 27814
rect 72896 27608 73108 27750
rect 74664 27744 75012 27820
rect 74664 27678 74876 27744
rect 74664 27614 74806 27678
rect 74870 27614 74876 27678
rect 74664 27608 74876 27614
rect 75072 27678 75284 27820
rect 75072 27614 75214 27678
rect 75278 27614 75284 27678
rect 75072 27608 75284 27614
rect 75480 27744 76100 27820
rect 75480 27608 75692 27744
rect 75888 27608 76100 27744
rect 76296 27678 76644 27820
rect 76296 27614 76438 27678
rect 76502 27614 76644 27678
rect 76296 27608 76644 27614
rect 73032 27548 73108 27608
rect 24480 27412 24556 27472
rect 66368 27412 66444 27472
rect 17816 27206 17822 27270
rect 17886 27206 18028 27270
rect 17816 27200 18028 27206
rect 18224 27406 18572 27412
rect 18224 27342 18502 27406
rect 18566 27342 18572 27406
rect 18224 27336 18572 27342
rect 18632 27406 18980 27412
rect 18632 27342 18774 27406
rect 18838 27342 18980 27406
rect 18224 27200 18436 27336
rect 18632 27270 18980 27342
rect 18632 27206 18638 27270
rect 18702 27206 18980 27270
rect 18632 27200 18980 27206
rect 19040 27406 19252 27412
rect 19040 27342 19046 27406
rect 19110 27342 19252 27406
rect 19040 27270 19252 27342
rect 19040 27206 19182 27270
rect 19246 27206 19252 27270
rect 19040 27200 19252 27206
rect 19448 27406 19660 27412
rect 19448 27342 19454 27406
rect 19518 27342 19660 27406
rect 19448 27270 19660 27342
rect 19448 27206 19590 27270
rect 19654 27206 19660 27270
rect 19448 27200 19660 27206
rect 24344 27200 24692 27412
rect 24616 27140 24692 27200
rect 14416 26998 14628 27004
rect 14416 26934 14558 26998
rect 14622 26934 14628 26998
rect 14416 26868 14628 26934
rect 14824 26998 15444 27004
rect 14824 26934 15374 26998
rect 15438 26934 15444 26998
rect 14824 26928 15444 26934
rect 14416 26862 14764 26868
rect 14416 26798 14422 26862
rect 14486 26798 14764 26862
rect 14416 26792 14764 26798
rect 14824 26792 15036 26928
rect 15232 26868 15444 26928
rect 15134 26862 15444 26868
rect 15096 26798 15102 26862
rect 15166 26798 15444 26862
rect 15134 26792 15444 26798
rect 15640 26998 15852 27004
rect 15640 26934 15782 26998
rect 15846 26934 15852 26998
rect 15640 26862 15852 26934
rect 15640 26798 15646 26862
rect 15710 26798 15852 26862
rect 15640 26792 15852 26798
rect 16048 26862 16260 27004
rect 16048 26798 16190 26862
rect 16254 26798 16260 26862
rect 16048 26792 16260 26798
rect 17816 26998 18028 27004
rect 17816 26934 17822 26998
rect 17886 26934 18028 26998
rect 17816 26792 18028 26934
rect 18224 26868 18436 27004
rect 18632 26998 18980 27004
rect 18632 26934 18638 26998
rect 18702 26934 18980 26998
rect 18224 26862 18572 26868
rect 18224 26798 18502 26862
rect 18566 26798 18572 26862
rect 18224 26792 18572 26798
rect 18632 26862 18980 26934
rect 18632 26798 18910 26862
rect 18974 26798 18980 26862
rect 18632 26792 18980 26798
rect 19040 26998 19252 27004
rect 19040 26934 19182 26998
rect 19246 26934 19252 26998
rect 19040 26862 19252 26934
rect 19040 26798 19046 26862
rect 19110 26798 19252 26862
rect 19040 26792 19252 26798
rect 19448 26998 19660 27004
rect 19448 26934 19590 26998
rect 19654 26934 19660 26998
rect 19448 26862 19660 26934
rect 24344 26928 24692 27140
rect 24616 26868 24692 26928
rect 19448 26798 19454 26862
rect 19518 26798 19660 26862
rect 19448 26792 19660 26798
rect 14688 26732 14764 26792
rect 15640 26732 15716 26792
rect 14688 26656 15716 26732
rect 17816 26732 17892 26792
rect 17816 26590 18028 26732
rect 24344 26656 24692 26868
rect 66368 27200 66580 27412
rect 71264 27406 71476 27412
rect 71264 27342 71270 27406
rect 71334 27342 71476 27406
rect 71264 27270 71476 27342
rect 71264 27206 71406 27270
rect 71470 27206 71476 27270
rect 71264 27200 71476 27206
rect 71672 27406 71884 27412
rect 71672 27342 71678 27406
rect 71742 27342 71884 27406
rect 71672 27270 71884 27342
rect 71672 27206 71678 27270
rect 71742 27206 71884 27270
rect 71672 27200 71884 27206
rect 72080 27406 72700 27412
rect 72080 27342 72630 27406
rect 72694 27342 72700 27406
rect 72080 27336 72700 27342
rect 72080 27200 72292 27336
rect 72488 27270 72700 27336
rect 72488 27206 72494 27270
rect 72558 27206 72700 27270
rect 72488 27200 72700 27206
rect 72896 27270 73108 27548
rect 72896 27206 72902 27270
rect 72966 27206 73108 27270
rect 72896 27200 73108 27206
rect 89080 27406 89836 27412
rect 89080 27342 89766 27406
rect 89830 27342 89836 27406
rect 89080 27336 89836 27342
rect 89080 27332 89428 27336
rect 89080 27276 89216 27332
rect 89272 27276 89428 27332
rect 89080 27200 89428 27276
rect 66368 27140 66444 27200
rect 66368 26928 66580 27140
rect 71264 26998 71476 27004
rect 71264 26934 71406 26998
rect 71470 26934 71476 26998
rect 66368 26868 66444 26928
rect 66368 26656 66580 26868
rect 71264 26862 71476 26934
rect 71264 26798 71270 26862
rect 71334 26798 71476 26862
rect 71264 26792 71476 26798
rect 71672 26998 71884 27004
rect 71672 26934 71678 26998
rect 71742 26934 71884 26998
rect 71672 26862 71884 26934
rect 71672 26798 71814 26862
rect 71878 26798 71884 26862
rect 71672 26792 71884 26798
rect 72080 26868 72292 27004
rect 72488 26998 72700 27004
rect 72488 26934 72494 26998
rect 72558 26934 72700 26998
rect 72080 26862 72428 26868
rect 72080 26798 72358 26862
rect 72422 26798 72428 26862
rect 72080 26792 72428 26798
rect 72488 26792 72700 26934
rect 72896 26998 73108 27004
rect 72896 26934 72902 26998
rect 72966 26934 73108 26998
rect 72896 26792 73108 26934
rect 74664 26998 74876 27004
rect 74664 26934 74806 26998
rect 74870 26934 74876 26998
rect 74664 26868 74876 26934
rect 75072 26998 75284 27004
rect 75072 26934 75214 26998
rect 75278 26934 75284 26998
rect 74664 26792 75012 26868
rect 75072 26862 75284 26934
rect 75072 26798 75214 26862
rect 75278 26798 75284 26862
rect 75072 26792 75284 26798
rect 75480 26868 75692 27004
rect 75888 26868 76100 27004
rect 75480 26862 76100 26868
rect 75480 26798 76030 26862
rect 76094 26798 76100 26862
rect 75480 26792 76100 26798
rect 76296 26998 76644 27004
rect 76296 26934 76438 26998
rect 76502 26934 76644 26998
rect 76296 26862 76644 26934
rect 76296 26798 76302 26862
rect 76366 26798 76644 26862
rect 76296 26792 76644 26798
rect 72488 26732 72564 26792
rect 73032 26732 73108 26792
rect 24344 26596 24420 26656
rect 66504 26596 66580 26656
rect 72216 26656 72564 26732
rect 72216 26596 72292 26656
rect 17816 26526 17958 26590
rect 18022 26526 18028 26590
rect 17816 26520 18028 26526
rect 3128 26324 3340 26460
rect 3808 26324 4020 26460
rect 18224 26384 18436 26596
rect 18534 26590 18980 26596
rect 18496 26526 18502 26590
rect 18566 26526 18910 26590
rect 18974 26526 18980 26590
rect 18534 26520 18980 26526
rect 18632 26460 18980 26520
rect 18360 26324 18436 26384
rect 18496 26384 18980 26460
rect 19040 26590 19252 26596
rect 19040 26526 19046 26590
rect 19110 26526 19252 26590
rect 19040 26454 19252 26526
rect 19040 26390 19182 26454
rect 19246 26390 19252 26454
rect 19040 26384 19252 26390
rect 19448 26590 19660 26596
rect 19448 26526 19454 26590
rect 19518 26526 19660 26590
rect 19448 26454 19660 26526
rect 19448 26390 19454 26454
rect 19518 26390 19660 26454
rect 19448 26384 19660 26390
rect 18496 26324 18572 26384
rect 544 26318 4020 26324
rect 544 26254 550 26318
rect 614 26254 4020 26318
rect 544 26248 4020 26254
rect 14416 26318 14628 26324
rect 14416 26254 14422 26318
rect 14486 26254 14628 26318
rect 14416 26046 14628 26254
rect 14416 25982 14422 26046
rect 14486 25982 14628 26046
rect 14416 25976 14628 25982
rect 14824 26318 15172 26324
rect 14824 26254 15102 26318
rect 15166 26254 15172 26318
rect 14824 26248 15172 26254
rect 14824 26188 15036 26248
rect 15232 26188 15444 26324
rect 15950 26318 18028 26324
rect 15912 26254 15918 26318
rect 15982 26254 17958 26318
rect 18022 26254 18028 26318
rect 15950 26248 18028 26254
rect 14824 26112 15444 26188
rect 14824 26052 15036 26112
rect 14824 26046 15172 26052
rect 14824 25982 14830 26046
rect 14894 25982 15102 26046
rect 15166 25982 15172 26046
rect 14824 25976 15172 25982
rect 15232 25976 15444 26112
rect 15640 26182 15852 26188
rect 15640 26118 15646 26182
rect 15710 26118 15852 26182
rect 15640 26046 15852 26118
rect 15640 25982 15782 26046
rect 15846 25982 15852 26046
rect 15640 25976 15852 25982
rect 16048 26182 16260 26188
rect 16048 26118 16190 26182
rect 16254 26118 16260 26182
rect 16048 26052 16260 26118
rect 16048 26046 17756 26052
rect 16048 25982 16054 26046
rect 16118 25982 17686 26046
rect 17750 25982 17756 26046
rect 16048 25976 17756 25982
rect 17816 25976 18028 26248
rect 18224 26248 18572 26324
rect 18632 26324 18708 26384
rect 18632 26248 18980 26324
rect 18224 25976 18436 26248
rect 18752 26052 18850 26248
rect 19040 26182 19252 26188
rect 19040 26118 19182 26182
rect 19246 26118 19252 26182
rect 18632 26046 18980 26052
rect 18632 25982 18638 26046
rect 18702 25982 18980 26046
rect 18632 25976 18980 25982
rect 19040 25976 19252 26118
rect 19448 26182 19660 26188
rect 19448 26118 19454 26182
rect 19518 26118 19660 26182
rect 19448 25976 19660 26118
rect 17952 25916 18028 25976
rect 19176 25916 19252 25976
rect 19584 25916 19660 25976
rect 1632 25652 1844 25780
rect 17816 25774 18028 25916
rect 2460 25732 2526 25733
rect 2418 25668 2461 25732
rect 2525 25668 2568 25732
rect 17816 25710 17958 25774
rect 18022 25710 18028 25774
rect 17816 25704 18028 25710
rect 2460 25667 2526 25668
rect 1632 25644 1718 25652
rect 1224 25638 1718 25644
rect 1224 25574 1230 25638
rect 1294 25596 1718 25638
rect 1774 25644 1844 25652
rect 18224 25644 18436 25780
rect 1774 25638 2252 25644
rect 1774 25596 2182 25638
rect 1294 25574 2182 25596
rect 2246 25574 2252 25638
rect 1224 25568 2252 25574
rect 14280 25638 14900 25644
rect 14280 25574 14830 25638
rect 14894 25574 14900 25638
rect 14280 25568 14900 25574
rect 15504 25568 16124 25644
rect 17718 25638 18436 25644
rect 17680 25574 17686 25638
rect 17750 25574 18436 25638
rect 17718 25568 18436 25574
rect 18632 25774 18980 25780
rect 18632 25710 18638 25774
rect 18702 25710 18980 25774
rect 18632 25568 18980 25710
rect 19040 25568 19252 25916
rect 19448 25568 19660 25916
rect 14280 25508 14356 25568
rect 15504 25508 15580 25568
rect 16048 25508 16124 25568
rect 18224 25508 18300 25568
rect 18632 25508 18708 25568
rect 19040 25508 19116 25568
rect 19584 25508 19660 25568
rect 12920 25502 13132 25508
rect 12920 25438 12926 25502
rect 12990 25438 13132 25502
rect 12920 25372 13132 25438
rect 13328 25432 14356 25508
rect 14416 25502 14628 25508
rect 14416 25438 14422 25502
rect 14486 25438 14628 25502
rect 12920 25296 13268 25372
rect 13328 25296 13540 25432
rect 14416 25372 14628 25438
rect 14824 25372 15036 25508
rect 15134 25502 15580 25508
rect 15096 25438 15102 25502
rect 15166 25438 15580 25502
rect 15134 25432 15580 25438
rect 15640 25502 15988 25508
rect 15640 25438 15782 25502
rect 15846 25438 15918 25502
rect 15982 25438 15988 25502
rect 15640 25432 15988 25438
rect 16048 25502 16260 25508
rect 16048 25438 16054 25502
rect 16118 25438 16260 25502
rect 15232 25372 15444 25432
rect 14416 25366 14764 25372
rect 14416 25302 14694 25366
rect 14758 25302 14764 25366
rect 14416 25296 14764 25302
rect 14824 25296 15444 25372
rect 15640 25296 15852 25432
rect 16048 25296 16260 25438
rect 17816 25502 18028 25508
rect 17816 25438 17958 25502
rect 18022 25438 18028 25502
rect 17816 25366 18028 25438
rect 17816 25302 17822 25366
rect 17886 25302 18028 25366
rect 17816 25296 18028 25302
rect 18224 25366 18436 25508
rect 18632 25372 18980 25508
rect 18534 25366 18980 25372
rect 18224 25302 18230 25366
rect 18294 25302 18436 25366
rect 18496 25302 18502 25366
rect 18566 25302 18980 25366
rect 18224 25296 18436 25302
rect 18534 25296 18980 25302
rect 19040 25366 19252 25508
rect 19040 25302 19046 25366
rect 19110 25302 19252 25366
rect 19040 25296 19252 25302
rect 19448 25366 19660 25508
rect 24344 26112 24692 26596
rect 66368 26112 66580 26596
rect 71264 26590 71476 26596
rect 71264 26526 71270 26590
rect 71334 26526 71476 26590
rect 71264 26454 71476 26526
rect 71264 26390 71270 26454
rect 71334 26390 71476 26454
rect 71264 26384 71476 26390
rect 71672 26590 71884 26596
rect 71672 26526 71814 26590
rect 71878 26526 71884 26590
rect 71672 26454 71884 26526
rect 71672 26390 71678 26454
rect 71742 26390 71884 26454
rect 71672 26384 71884 26390
rect 72080 26460 72292 26596
rect 72390 26590 72700 26596
rect 72352 26526 72358 26590
rect 72422 26526 72700 26590
rect 72390 26520 72700 26526
rect 72896 26590 73108 26732
rect 74936 26732 75012 26792
rect 75480 26732 75556 26792
rect 74936 26656 75556 26732
rect 72896 26526 73038 26590
rect 73102 26526 73108 26590
rect 72896 26520 73108 26526
rect 72488 26460 72700 26520
rect 72080 26454 74740 26460
rect 72080 26390 74670 26454
rect 74734 26390 74740 26454
rect 72080 26384 74740 26390
rect 72216 26324 72292 26384
rect 72624 26324 72700 26384
rect 71264 26182 71476 26188
rect 71264 26118 71270 26182
rect 71334 26118 71476 26182
rect 24344 26052 24420 26112
rect 66368 26052 66444 26112
rect 24344 25910 24692 26052
rect 24344 25846 24622 25910
rect 24686 25846 24692 25910
rect 24344 25638 24692 25846
rect 24344 25574 24622 25638
rect 24686 25574 24692 25638
rect 24344 25432 24692 25574
rect 66368 25910 66580 26052
rect 71264 25976 71476 26118
rect 71672 26182 71884 26188
rect 71672 26118 71678 26182
rect 71742 26118 71884 26182
rect 71672 25976 71884 26118
rect 72080 26046 72292 26324
rect 72080 25982 72222 26046
rect 72286 25982 72292 26046
rect 72080 25976 72292 25982
rect 72488 25976 72700 26324
rect 72896 26318 73108 26324
rect 72896 26254 73038 26318
rect 73102 26254 73108 26318
rect 72896 25976 73108 26254
rect 75480 26318 76100 26324
rect 75480 26254 76030 26318
rect 76094 26254 76100 26318
rect 75480 26248 76100 26254
rect 76296 26318 76644 26324
rect 76296 26254 76302 26318
rect 76366 26254 76644 26318
rect 76296 26248 76644 26254
rect 74664 26182 74876 26188
rect 74664 26118 74670 26182
rect 74734 26118 74876 26182
rect 74664 26046 74876 26118
rect 74664 25982 74670 26046
rect 74734 25982 74876 26046
rect 74664 25976 74876 25982
rect 75072 26182 75284 26188
rect 75072 26118 75214 26182
rect 75278 26118 75284 26182
rect 75072 26046 75284 26118
rect 75072 25982 75078 26046
rect 75142 25982 75284 26046
rect 75072 25976 75284 25982
rect 75480 26052 75692 26248
rect 75888 26052 76100 26248
rect 76411 26052 76509 26248
rect 75480 26046 75828 26052
rect 75480 25982 75758 26046
rect 75822 25982 75828 26046
rect 75480 25976 75828 25982
rect 75888 25976 76236 26052
rect 76296 26046 76644 26052
rect 76296 25982 76302 26046
rect 76366 25982 76438 26046
rect 76502 25982 76644 26046
rect 76296 25976 76644 25982
rect 71400 25916 71476 25976
rect 71808 25916 71884 25976
rect 66368 25846 66374 25910
rect 66438 25846 66580 25910
rect 66368 25638 66580 25846
rect 66368 25574 66374 25638
rect 66438 25574 66580 25638
rect 66368 25432 66580 25574
rect 24616 25372 24692 25432
rect 66504 25372 66580 25432
rect 19448 25302 19590 25366
rect 19654 25302 19660 25366
rect 19448 25296 19660 25302
rect 13192 25236 13268 25296
rect 14416 25236 14492 25296
rect 13192 25160 14492 25236
rect 14960 25236 15036 25296
rect 14960 25230 15308 25236
rect 14960 25166 15238 25230
rect 15302 25166 15308 25230
rect 14960 25160 15308 25166
rect 2214 25094 4020 25100
rect 2176 25030 2182 25094
rect 2246 25030 4020 25094
rect 2214 25024 4020 25030
rect 3128 24888 3340 25024
rect 3808 24888 4020 25024
rect 17816 25094 18028 25100
rect 17816 25030 17822 25094
rect 17886 25030 18028 25094
rect 17816 24958 18028 25030
rect 17816 24894 17822 24958
rect 17886 24894 18028 24958
rect 17816 24888 18028 24894
rect 18224 25094 18572 25100
rect 18224 25030 18230 25094
rect 18294 25030 18502 25094
rect 18566 25030 18572 25094
rect 18224 25024 18572 25030
rect 18224 24964 18436 25024
rect 18632 24964 18980 25100
rect 18224 24958 18980 24964
rect 18224 24894 18774 24958
rect 18838 24894 18980 24958
rect 18224 24888 18980 24894
rect 19040 25094 19252 25100
rect 19040 25030 19046 25094
rect 19110 25030 19252 25094
rect 19040 24958 19252 25030
rect 19040 24894 19182 24958
rect 19246 24894 19252 24958
rect 19040 24888 19252 24894
rect 19448 25094 19660 25100
rect 19448 25030 19590 25094
rect 19654 25030 19660 25094
rect 19448 24958 19660 25030
rect 19448 24894 19454 24958
rect 19518 24894 19660 24958
rect 19448 24888 19660 24894
rect 24344 25094 24692 25372
rect 24344 25030 24622 25094
rect 24686 25030 24692 25094
rect 24344 24888 24692 25030
rect 66368 25094 66580 25372
rect 71264 25568 71476 25916
rect 71672 25568 71884 25916
rect 72896 25916 72972 25976
rect 76160 25916 76236 25976
rect 72080 25774 72292 25780
rect 72080 25710 72222 25774
rect 72286 25710 72292 25774
rect 72080 25568 72292 25710
rect 72488 25644 72700 25780
rect 72896 25774 73108 25916
rect 76160 25910 77460 25916
rect 76160 25846 77390 25910
rect 77454 25846 77460 25910
rect 76160 25840 77460 25846
rect 72896 25710 73038 25774
rect 73102 25710 73108 25774
rect 72896 25704 73108 25710
rect 89080 25652 89428 25780
rect 71264 25508 71340 25568
rect 71808 25508 71884 25568
rect 72216 25508 72292 25568
rect 72352 25568 72700 25644
rect 72352 25508 72428 25568
rect 72624 25508 72700 25568
rect 75344 25638 76372 25644
rect 75344 25574 76302 25638
rect 76366 25574 76372 25638
rect 75344 25568 76372 25574
rect 77248 25568 77868 25644
rect 89080 25596 89216 25652
rect 89272 25644 89428 25652
rect 89272 25638 89836 25644
rect 89272 25596 89766 25638
rect 89080 25574 89766 25596
rect 89830 25574 89836 25638
rect 89080 25568 89836 25574
rect 75344 25508 75420 25568
rect 77248 25508 77324 25568
rect 77792 25508 77868 25568
rect 71264 25366 71476 25508
rect 71264 25302 71406 25366
rect 71470 25302 71476 25366
rect 71264 25296 71476 25302
rect 71672 25366 71884 25508
rect 71672 25302 71678 25366
rect 71742 25302 71884 25366
rect 71672 25296 71884 25302
rect 72080 25432 72428 25508
rect 72080 25366 72292 25432
rect 72080 25302 72222 25366
rect 72286 25302 72292 25366
rect 72080 25296 72292 25302
rect 72488 25296 72700 25508
rect 72896 25502 73108 25508
rect 72896 25438 73038 25502
rect 73102 25438 73108 25502
rect 72896 25366 73108 25438
rect 72896 25302 72902 25366
rect 72966 25302 73108 25366
rect 72896 25296 73108 25302
rect 74664 25502 74876 25508
rect 74664 25438 74670 25502
rect 74734 25438 74876 25502
rect 74664 25372 74876 25438
rect 75072 25502 75420 25508
rect 75072 25438 75078 25502
rect 75142 25438 75420 25502
rect 75072 25432 75420 25438
rect 74664 25366 75012 25372
rect 74664 25302 74670 25366
rect 74734 25302 75012 25366
rect 74664 25296 75012 25302
rect 75072 25296 75284 25432
rect 75480 25372 75692 25508
rect 75790 25502 76100 25508
rect 75752 25438 75758 25502
rect 75822 25438 76100 25502
rect 75790 25432 76100 25438
rect 75888 25372 76100 25432
rect 75480 25296 76100 25372
rect 76296 25502 77324 25508
rect 76296 25438 76438 25502
rect 76502 25438 77324 25502
rect 76296 25432 77324 25438
rect 77384 25502 77596 25508
rect 77384 25438 77390 25502
rect 77454 25438 77596 25502
rect 76296 25366 76644 25432
rect 76296 25302 76302 25366
rect 76366 25302 76644 25366
rect 76296 25296 76644 25302
rect 77384 25296 77596 25438
rect 77792 25296 78004 25508
rect 74936 25236 75012 25296
rect 75480 25236 75556 25296
rect 74936 25160 75556 25236
rect 66368 25030 66374 25094
rect 66438 25030 66580 25094
rect 66368 24888 66580 25030
rect 71264 25094 71476 25100
rect 71264 25030 71406 25094
rect 71470 25030 71476 25094
rect 71264 24958 71476 25030
rect 71264 24894 71406 24958
rect 71470 24894 71476 24958
rect 71264 24888 71476 24894
rect 71672 25094 71884 25100
rect 71672 25030 71678 25094
rect 71742 25030 71884 25094
rect 71672 24958 71884 25030
rect 71672 24894 71678 24958
rect 71742 24894 71884 24958
rect 71672 24888 71884 24894
rect 72080 25094 72292 25100
rect 72080 25030 72222 25094
rect 72286 25030 72292 25094
rect 72080 24958 72292 25030
rect 72080 24894 72222 24958
rect 72286 24894 72292 24958
rect 72080 24888 72292 24894
rect 72488 24888 72700 25100
rect 72896 25094 73108 25100
rect 72896 25030 72902 25094
rect 72966 25030 73108 25094
rect 72896 24958 73108 25030
rect 72896 24894 73038 24958
rect 73102 24894 73108 24958
rect 72896 24888 73108 24894
rect 24480 24828 24556 24888
rect 66368 24828 66444 24888
rect 72488 24828 72564 24888
rect 24344 24822 24692 24828
rect 24344 24758 24622 24822
rect 24686 24758 24692 24822
rect 17816 24686 18028 24692
rect 17816 24622 17822 24686
rect 17886 24622 18028 24686
rect 17816 24550 18028 24622
rect 17816 24486 17958 24550
rect 18022 24486 18028 24550
rect 17816 24480 18028 24486
rect 18224 24550 18436 24692
rect 18224 24486 18230 24550
rect 18294 24486 18436 24550
rect 18224 24480 18436 24486
rect 18632 24686 18980 24692
rect 18632 24622 18774 24686
rect 18838 24622 18980 24686
rect 18632 24550 18980 24622
rect 18632 24486 18638 24550
rect 18702 24486 18980 24550
rect 18632 24480 18980 24486
rect 19040 24686 19252 24692
rect 19040 24622 19182 24686
rect 19246 24622 19252 24686
rect 19040 24550 19252 24622
rect 19040 24486 19046 24550
rect 19110 24486 19252 24550
rect 19040 24480 19252 24486
rect 19448 24686 19660 24692
rect 19448 24622 19454 24686
rect 19518 24622 19660 24686
rect 19448 24550 19660 24622
rect 19448 24486 19590 24550
rect 19654 24486 19660 24550
rect 19448 24480 19660 24486
rect 24344 24616 24692 24758
rect 66368 24822 66580 24828
rect 66368 24758 66374 24822
rect 66438 24758 66580 24822
rect 66368 24616 66580 24758
rect 72216 24752 72564 24828
rect 72216 24692 72292 24752
rect 24344 24556 24420 24616
rect 66504 24556 66580 24616
rect 24344 24344 24692 24556
rect 66368 24344 66580 24556
rect 71264 24686 71476 24692
rect 71264 24622 71406 24686
rect 71470 24622 71476 24686
rect 71264 24550 71476 24622
rect 71264 24486 71270 24550
rect 71334 24486 71476 24550
rect 71264 24480 71476 24486
rect 71672 24686 71884 24692
rect 71672 24622 71678 24686
rect 71742 24622 71884 24686
rect 71672 24550 71884 24622
rect 71672 24486 71678 24550
rect 71742 24486 71884 24550
rect 71672 24480 71884 24486
rect 72080 24686 72700 24692
rect 72080 24622 72222 24686
rect 72286 24622 72700 24686
rect 72080 24616 72700 24622
rect 72080 24480 72292 24616
rect 72488 24550 72700 24616
rect 72488 24486 72630 24550
rect 72694 24486 72700 24550
rect 72488 24480 72700 24486
rect 72896 24686 73108 24692
rect 72896 24622 73038 24686
rect 73102 24622 73108 24686
rect 72896 24550 73108 24622
rect 72896 24486 73038 24550
rect 73102 24486 73108 24550
rect 72896 24480 73108 24486
rect 24480 24284 24556 24344
rect 66504 24284 66580 24344
rect 17816 24278 18028 24284
rect 17816 24214 17958 24278
rect 18022 24214 18028 24278
rect 17816 24142 18028 24214
rect 17816 24078 17822 24142
rect 17886 24078 18028 24142
rect 17816 24072 18028 24078
rect 18224 24278 18980 24284
rect 18224 24214 18230 24278
rect 18294 24214 18638 24278
rect 18702 24214 18980 24278
rect 18224 24208 18980 24214
rect 18224 24148 18436 24208
rect 18224 24142 18572 24148
rect 18224 24078 18366 24142
rect 18430 24078 18502 24142
rect 18566 24078 18572 24142
rect 18224 24072 18572 24078
rect 18632 24072 18980 24208
rect 19040 24278 19252 24284
rect 19040 24214 19046 24278
rect 19110 24214 19252 24278
rect 19040 24142 19252 24214
rect 19040 24078 19182 24142
rect 19246 24078 19252 24142
rect 19040 24072 19252 24078
rect 19448 24278 19660 24284
rect 19448 24214 19590 24278
rect 19654 24214 19660 24278
rect 19448 24142 19660 24214
rect 19448 24078 19454 24142
rect 19518 24078 19660 24142
rect 19448 24072 19660 24078
rect 24344 24072 24692 24284
rect 66368 24072 66580 24284
rect 71264 24278 71476 24284
rect 71264 24214 71270 24278
rect 71334 24214 71476 24278
rect 71264 24142 71476 24214
rect 71264 24078 71406 24142
rect 71470 24078 71476 24142
rect 71264 24072 71476 24078
rect 71672 24278 71884 24284
rect 71672 24214 71678 24278
rect 71742 24214 71884 24278
rect 71672 24142 71884 24214
rect 71672 24078 71678 24142
rect 71742 24078 71884 24142
rect 71672 24072 71884 24078
rect 72080 24142 72292 24284
rect 72080 24078 72086 24142
rect 72150 24078 72292 24142
rect 72080 24072 72292 24078
rect 72488 24278 72700 24284
rect 72488 24214 72630 24278
rect 72694 24214 72700 24278
rect 72488 24142 72700 24214
rect 72488 24078 72494 24142
rect 72558 24078 72700 24142
rect 72488 24072 72700 24078
rect 72896 24278 73108 24284
rect 72896 24214 73038 24278
rect 73102 24214 73108 24278
rect 72896 24148 73108 24214
rect 72896 24142 75148 24148
rect 72896 24078 72902 24142
rect 72966 24078 75078 24142
rect 75142 24078 75148 24142
rect 72896 24072 75148 24078
rect 24344 24012 24420 24072
rect 66368 24012 66444 24072
rect 1632 23972 1844 24012
rect 1632 23916 1718 23972
rect 1774 23916 1844 23972
rect 1632 23876 1844 23916
rect 15504 23936 16124 24012
rect 15504 23876 15580 23936
rect 16048 23876 16124 23936
rect 1224 23870 1844 23876
rect 14726 23870 15036 23876
rect 1224 23806 1230 23870
rect 1294 23806 1844 23870
rect 14688 23806 14694 23870
rect 14758 23806 15036 23870
rect 1224 23800 1844 23806
rect 14726 23800 15036 23806
rect 14824 23740 15036 23800
rect 15232 23870 15580 23876
rect 15232 23806 15238 23870
rect 15302 23806 15580 23870
rect 15232 23800 15580 23806
rect 14824 23664 15172 23740
rect 15232 23734 15444 23800
rect 15232 23670 15238 23734
rect 15302 23670 15444 23734
rect 15232 23664 15444 23670
rect 15640 23734 15852 23876
rect 15640 23670 15782 23734
rect 15846 23670 15852 23734
rect 15640 23664 15852 23670
rect 16048 23734 16260 23876
rect 16048 23670 16190 23734
rect 16254 23670 16260 23734
rect 16048 23664 16260 23670
rect 17816 23870 18028 23876
rect 17816 23806 17822 23870
rect 17886 23806 18028 23870
rect 17816 23734 18028 23806
rect 17816 23670 17822 23734
rect 17886 23670 18028 23734
rect 17816 23664 18028 23670
rect 18224 23870 18436 23876
rect 18534 23870 18980 23876
rect 18224 23806 18366 23870
rect 18430 23806 18436 23870
rect 18496 23806 18502 23870
rect 18566 23806 18980 23870
rect 18224 23734 18436 23806
rect 18534 23800 18980 23806
rect 18224 23670 18230 23734
rect 18294 23670 18436 23734
rect 18224 23664 18436 23670
rect 18632 23664 18980 23800
rect 19040 23870 19252 23876
rect 19040 23806 19182 23870
rect 19246 23806 19252 23870
rect 19040 23734 19252 23806
rect 19040 23670 19182 23734
rect 19246 23670 19252 23734
rect 19040 23664 19252 23670
rect 19448 23870 19660 23876
rect 19448 23806 19454 23870
rect 19518 23806 19660 23870
rect 19448 23734 19660 23806
rect 24344 23800 24692 24012
rect 66368 23800 66580 24012
rect 75344 23936 75964 24012
rect 75344 23876 75420 23936
rect 75888 23876 75964 23936
rect 89080 23972 89428 24012
rect 89080 23916 89216 23972
rect 89272 23916 89428 23972
rect 89080 23876 89428 23916
rect 71264 23870 71476 23876
rect 71264 23806 71406 23870
rect 71470 23806 71476 23870
rect 24480 23740 24556 23800
rect 66368 23740 66444 23800
rect 19448 23670 19454 23734
rect 19518 23670 19660 23734
rect 19448 23664 19660 23670
rect 15096 23604 15172 23664
rect 15640 23604 15716 23664
rect 3128 23528 4020 23604
rect 15096 23528 15716 23604
rect 24344 23528 24692 23740
rect 66368 23528 66580 23740
rect 71264 23734 71476 23806
rect 71264 23670 71270 23734
rect 71334 23670 71476 23734
rect 71264 23664 71476 23670
rect 71672 23870 71884 23876
rect 71672 23806 71678 23870
rect 71742 23806 71884 23870
rect 71672 23734 71884 23806
rect 71672 23670 71678 23734
rect 71742 23670 71884 23734
rect 71672 23664 71884 23670
rect 72080 23870 72292 23876
rect 72080 23806 72086 23870
rect 72150 23806 72292 23870
rect 72080 23734 72292 23806
rect 72080 23670 72086 23734
rect 72150 23670 72292 23734
rect 72080 23664 72292 23670
rect 72488 23870 72700 23876
rect 72488 23806 72494 23870
rect 72558 23806 72700 23870
rect 72488 23664 72700 23806
rect 72896 23870 73108 23876
rect 72896 23806 72902 23870
rect 72966 23806 73108 23870
rect 72896 23734 73108 23806
rect 72896 23670 73038 23734
rect 73102 23670 73108 23734
rect 72896 23664 73108 23670
rect 74664 23870 74876 23876
rect 74664 23806 74670 23870
rect 74734 23806 74876 23870
rect 74664 23740 74876 23806
rect 75072 23870 75420 23876
rect 75072 23806 75078 23870
rect 75142 23806 75420 23870
rect 75072 23800 75420 23806
rect 74664 23734 75012 23740
rect 74664 23670 74670 23734
rect 74734 23670 75012 23734
rect 74664 23664 75012 23670
rect 75072 23664 75284 23800
rect 75480 23734 75692 23876
rect 75480 23670 75486 23734
rect 75550 23670 75692 23734
rect 75480 23664 75692 23670
rect 75888 23870 76372 23876
rect 75888 23806 76302 23870
rect 76366 23806 76372 23870
rect 75888 23800 76372 23806
rect 89080 23870 89836 23876
rect 89080 23806 89766 23870
rect 89830 23806 89836 23870
rect 89080 23800 89836 23806
rect 75888 23734 76100 23800
rect 75888 23670 76030 23734
rect 76094 23670 76100 23734
rect 75888 23664 76100 23670
rect 72488 23604 72564 23664
rect 3128 23392 3340 23528
rect 3808 23468 4020 23528
rect 24344 23468 24420 23528
rect 66504 23468 66580 23528
rect 72216 23528 72564 23604
rect 74936 23604 75012 23664
rect 75480 23604 75556 23664
rect 74936 23528 75556 23604
rect 72216 23468 72292 23528
rect 3710 23462 4020 23468
rect 3672 23398 3678 23462
rect 3742 23398 4020 23462
rect 3710 23392 4020 23398
rect 17816 23462 18028 23468
rect 17816 23398 17822 23462
rect 17886 23398 18028 23462
rect 17816 23326 18028 23398
rect 17816 23262 17822 23326
rect 17886 23262 18028 23326
rect 17816 23256 18028 23262
rect 18224 23462 18980 23468
rect 18224 23398 18230 23462
rect 18294 23398 18980 23462
rect 18224 23392 18980 23398
rect 18224 23256 18436 23392
rect 18632 23332 18980 23392
rect 18534 23326 18980 23332
rect 18496 23262 18502 23326
rect 18566 23262 18980 23326
rect 18534 23256 18980 23262
rect 19040 23462 19252 23468
rect 19040 23398 19182 23462
rect 19246 23398 19252 23462
rect 19040 23326 19252 23398
rect 19040 23262 19182 23326
rect 19246 23262 19252 23326
rect 19040 23256 19252 23262
rect 19448 23462 19660 23468
rect 19448 23398 19454 23462
rect 19518 23398 19660 23462
rect 19448 23326 19660 23398
rect 19448 23262 19590 23326
rect 19654 23262 19660 23326
rect 19448 23256 19660 23262
rect 24344 23256 24692 23468
rect 66368 23256 66580 23468
rect 71264 23462 71476 23468
rect 71264 23398 71270 23462
rect 71334 23398 71476 23462
rect 71264 23326 71476 23398
rect 71264 23262 71270 23326
rect 71334 23262 71476 23326
rect 71264 23256 71476 23262
rect 71672 23462 71884 23468
rect 71672 23398 71678 23462
rect 71742 23398 71884 23462
rect 71672 23326 71884 23398
rect 71672 23262 71678 23326
rect 71742 23262 71884 23326
rect 71672 23256 71884 23262
rect 72080 23462 72700 23468
rect 72080 23398 72086 23462
rect 72150 23398 72700 23462
rect 72080 23392 72700 23398
rect 72080 23326 72292 23392
rect 72080 23262 72086 23326
rect 72150 23262 72292 23326
rect 72080 23256 72292 23262
rect 72488 23256 72700 23392
rect 72896 23462 73108 23468
rect 72896 23398 73038 23462
rect 73102 23398 73108 23462
rect 72896 23326 73108 23398
rect 72896 23262 72902 23326
rect 72966 23262 73108 23326
rect 72896 23256 73108 23262
rect 24480 23196 24556 23256
rect 66504 23196 66580 23256
rect 13872 23120 14900 23196
rect 13872 23060 13948 23120
rect 14824 23060 14900 23120
rect 15096 23120 15716 23196
rect 15096 23060 15172 23120
rect 15640 23060 15716 23120
rect 13600 22984 13948 23060
rect 13600 22848 13812 22984
rect 14008 22924 14220 23060
rect 14824 22984 15172 23060
rect 15232 23054 15444 23060
rect 15232 22990 15238 23054
rect 15302 22990 15444 23054
rect 14008 22848 14764 22924
rect 14824 22848 15036 22984
rect 15232 22918 15444 22990
rect 15232 22854 15238 22918
rect 15302 22854 15444 22918
rect 15232 22848 15444 22854
rect 15640 23054 15852 23060
rect 15640 22990 15782 23054
rect 15846 22990 15852 23054
rect 15640 22918 15852 22990
rect 15640 22854 15646 22918
rect 15710 22854 15852 22918
rect 15640 22848 15852 22854
rect 16048 23054 16260 23060
rect 16048 22990 16190 23054
rect 16254 22990 16260 23054
rect 16048 22848 16260 22990
rect 17816 23054 18028 23060
rect 17816 22990 17822 23054
rect 17886 22990 18028 23054
rect 17816 22848 18028 22990
rect 18224 23054 18572 23060
rect 18224 22990 18502 23054
rect 18566 22990 18572 23054
rect 18224 22984 18572 22990
rect 18224 22924 18436 22984
rect 18632 22924 18980 23060
rect 18224 22848 18980 22924
rect 19040 23054 19252 23060
rect 19040 22990 19182 23054
rect 19246 22990 19252 23054
rect 19040 22918 19252 22990
rect 19040 22854 19182 22918
rect 19246 22854 19252 22918
rect 19040 22848 19252 22854
rect 19448 23054 19660 23060
rect 19448 22990 19590 23054
rect 19654 22990 19660 23054
rect 19448 22918 19660 22990
rect 24344 22984 24692 23196
rect 66368 22984 66580 23196
rect 75344 23120 75964 23196
rect 75344 23060 75420 23120
rect 75888 23060 75964 23120
rect 76704 23120 77324 23196
rect 76704 23060 76780 23120
rect 77248 23060 77324 23120
rect 71264 23054 71476 23060
rect 71264 22990 71270 23054
rect 71334 22990 71476 23054
rect 24480 22924 24556 22984
rect 66368 22924 66444 22984
rect 19448 22854 19590 22918
rect 19654 22854 19660 22918
rect 19448 22848 19660 22854
rect 14688 22788 14764 22848
rect 15232 22788 15308 22848
rect 14688 22712 15308 22788
rect 17816 22788 17892 22848
rect 18360 22788 18436 22848
rect 15134 22646 15716 22652
rect 15096 22582 15102 22646
rect 15166 22582 15646 22646
rect 15710 22582 15716 22646
rect 15134 22576 15716 22582
rect 17816 22646 18028 22788
rect 18360 22712 18708 22788
rect 24344 22712 24692 22924
rect 18632 22652 18708 22712
rect 24616 22652 24692 22712
rect 17816 22582 17958 22646
rect 18022 22582 18028 22646
rect 17816 22576 18028 22582
rect 18224 22440 18436 22652
rect 18632 22440 18980 22652
rect 19040 22646 19252 22652
rect 19040 22582 19182 22646
rect 19246 22582 19252 22646
rect 19040 22510 19252 22582
rect 19040 22446 19046 22510
rect 19110 22446 19252 22510
rect 19040 22440 19252 22446
rect 19448 22646 19660 22652
rect 19448 22582 19590 22646
rect 19654 22582 19660 22646
rect 19448 22510 19660 22582
rect 19448 22446 19454 22510
rect 19518 22446 19660 22510
rect 19448 22440 19660 22446
rect 18224 22380 18300 22440
rect 18904 22380 18980 22440
rect 1632 22292 1844 22380
rect 1632 22244 1718 22292
rect 1224 22238 1718 22244
rect 1224 22174 1230 22238
rect 1294 22236 1718 22238
rect 1774 22244 1844 22292
rect 17816 22374 18028 22380
rect 17816 22310 17958 22374
rect 18022 22310 18028 22374
rect 1774 22236 3340 22244
rect 1294 22174 3340 22236
rect 1224 22168 3340 22174
rect 3128 22108 3340 22168
rect 3808 22108 4020 22244
rect 3128 22032 4020 22108
rect 17816 22032 18028 22310
rect 18224 22102 18436 22380
rect 18224 22038 18366 22102
rect 18430 22038 18436 22102
rect 18224 22032 18436 22038
rect 18632 22102 18980 22380
rect 18632 22038 18774 22102
rect 18838 22038 18980 22102
rect 18632 22032 18980 22038
rect 19040 22238 19252 22244
rect 19040 22174 19046 22238
rect 19110 22174 19252 22238
rect 19040 22032 19252 22174
rect 19448 22238 19660 22244
rect 19448 22174 19454 22238
rect 19518 22174 19660 22238
rect 19448 22032 19660 22174
rect 17952 21972 18028 22032
rect 17816 21830 18028 21972
rect 19040 21972 19116 22032
rect 19584 21972 19660 22032
rect 17816 21766 17822 21830
rect 17886 21766 18028 21830
rect 17816 21760 18028 21766
rect 18224 21830 18436 21836
rect 18224 21766 18366 21830
rect 18430 21766 18436 21830
rect 18224 21700 18436 21766
rect 18632 21830 18980 21836
rect 18632 21766 18774 21830
rect 18838 21766 18980 21830
rect 15504 21624 16124 21700
rect 18224 21624 18572 21700
rect 18632 21624 18980 21766
rect 15504 21564 15580 21624
rect 16048 21564 16124 21624
rect 18360 21564 18436 21624
rect 14824 21558 15172 21564
rect 14824 21494 15102 21558
rect 15166 21494 15172 21558
rect 14824 21488 15172 21494
rect 15232 21558 15580 21564
rect 15232 21494 15238 21558
rect 15302 21494 15580 21558
rect 15232 21488 15580 21494
rect 14824 21428 15036 21488
rect 14824 21352 15172 21428
rect 15232 21352 15444 21488
rect 15096 21292 15172 21352
rect 15640 21292 15852 21564
rect 15096 21286 15852 21292
rect 15096 21222 15782 21286
rect 15846 21222 15852 21286
rect 15096 21216 15852 21222
rect 16048 21286 16260 21564
rect 17816 21558 18028 21564
rect 17816 21494 17822 21558
rect 17886 21494 18028 21558
rect 17816 21422 18028 21494
rect 17816 21358 17958 21422
rect 18022 21358 18028 21422
rect 17816 21352 18028 21358
rect 18224 21352 18436 21564
rect 18496 21564 18572 21624
rect 18904 21564 18980 21624
rect 18496 21488 18980 21564
rect 18632 21422 18980 21488
rect 18632 21358 18910 21422
rect 18974 21358 18980 21422
rect 18632 21352 18980 21358
rect 19040 21624 19252 21972
rect 19448 21624 19660 21972
rect 19040 21564 19116 21624
rect 19584 21564 19660 21624
rect 16048 21222 16190 21286
rect 16254 21222 16260 21286
rect 16048 21216 16260 21222
rect 19040 21216 19252 21564
rect 19448 21216 19660 21564
rect 24344 22168 24692 22652
rect 66368 22712 66580 22924
rect 71264 22918 71476 22990
rect 71264 22854 71406 22918
rect 71470 22854 71476 22918
rect 71264 22848 71476 22854
rect 71672 23054 71884 23060
rect 71672 22990 71678 23054
rect 71742 22990 71884 23054
rect 71672 22918 71884 22990
rect 71672 22854 71814 22918
rect 71878 22854 71884 22918
rect 71672 22848 71884 22854
rect 72080 23054 72292 23060
rect 72080 22990 72086 23054
rect 72150 22990 72292 23054
rect 72080 22918 72292 22990
rect 72080 22854 72086 22918
rect 72150 22854 72292 22918
rect 72080 22848 72292 22854
rect 72488 22918 72700 23060
rect 72488 22854 72494 22918
rect 72558 22854 72700 22918
rect 72488 22848 72700 22854
rect 72896 23054 73108 23060
rect 72896 22990 72902 23054
rect 72966 22990 73108 23054
rect 72896 22848 73108 22990
rect 74664 23054 74876 23060
rect 74664 22990 74670 23054
rect 74734 22990 74876 23054
rect 74664 22848 74876 22990
rect 75072 22984 75420 23060
rect 75480 23054 75692 23060
rect 75480 22990 75486 23054
rect 75550 22990 75692 23054
rect 75072 22918 75284 22984
rect 75072 22854 75078 22918
rect 75142 22854 75284 22918
rect 75072 22848 75284 22854
rect 75480 22924 75692 22990
rect 75888 23054 76780 23060
rect 75888 22990 76030 23054
rect 76094 22990 76780 23054
rect 75888 22984 76780 22990
rect 75480 22918 75828 22924
rect 75480 22854 75486 22918
rect 75550 22854 75828 22918
rect 75480 22848 75828 22854
rect 75888 22848 76100 22984
rect 76840 22848 77052 23060
rect 77248 22848 77460 23060
rect 72896 22788 72972 22848
rect 75752 22788 75828 22848
rect 76840 22788 76916 22848
rect 66368 22652 66444 22712
rect 66368 22168 66580 22652
rect 71264 22646 71476 22652
rect 71264 22582 71406 22646
rect 71470 22582 71476 22646
rect 71264 22510 71476 22582
rect 71264 22446 71270 22510
rect 71334 22446 71476 22510
rect 71264 22440 71476 22446
rect 71672 22646 71884 22652
rect 71672 22582 71814 22646
rect 71878 22582 71884 22646
rect 71672 22510 71884 22582
rect 71672 22446 71678 22510
rect 71742 22446 71884 22510
rect 71672 22440 71884 22446
rect 72080 22646 72292 22652
rect 72080 22582 72086 22646
rect 72150 22582 72292 22646
rect 72080 22516 72292 22582
rect 72488 22646 72700 22652
rect 72488 22582 72494 22646
rect 72558 22582 72700 22646
rect 72080 22440 72428 22516
rect 72488 22440 72700 22582
rect 72896 22646 73108 22788
rect 75752 22712 76916 22788
rect 72896 22582 72902 22646
rect 72966 22582 73108 22646
rect 72896 22576 73108 22582
rect 72216 22380 72292 22440
rect 24344 22108 24420 22168
rect 66504 22108 66580 22168
rect 24344 21966 24692 22108
rect 24344 21902 24350 21966
rect 24414 21902 24692 21966
rect 24344 21694 24692 21902
rect 24344 21630 24350 21694
rect 24414 21630 24486 21694
rect 24550 21630 24692 21694
rect 24344 21558 24692 21630
rect 24344 21494 24622 21558
rect 24686 21494 24692 21558
rect 24344 21488 24692 21494
rect 66368 21966 66580 22108
rect 66368 21902 66374 21966
rect 66438 21902 66580 21966
rect 66368 21694 66580 21902
rect 66368 21630 66374 21694
rect 66438 21630 66580 21694
rect 66368 21558 66580 21630
rect 71264 22238 71476 22244
rect 71264 22174 71270 22238
rect 71334 22174 71476 22238
rect 71264 22032 71476 22174
rect 71672 22238 71884 22244
rect 71672 22174 71678 22238
rect 71742 22174 71884 22238
rect 71672 22032 71884 22174
rect 72080 22102 72292 22380
rect 72352 22380 72428 22440
rect 72624 22380 72700 22440
rect 72352 22304 72700 22380
rect 72080 22038 72086 22102
rect 72150 22038 72292 22102
rect 72080 22032 72292 22038
rect 72488 22032 72700 22304
rect 72896 22374 73108 22380
rect 72896 22310 72902 22374
rect 72966 22310 73108 22374
rect 72896 22032 73108 22310
rect 89080 22292 89428 22380
rect 89080 22236 89216 22292
rect 89272 22244 89428 22292
rect 89272 22238 89836 22244
rect 89272 22236 89766 22238
rect 89080 22174 89766 22236
rect 89830 22174 89836 22238
rect 89080 22168 89836 22174
rect 71264 21972 71340 22032
rect 71672 21972 71748 22032
rect 72896 21972 72972 22032
rect 71264 21624 71476 21972
rect 71672 21624 71884 21972
rect 71400 21564 71476 21624
rect 71808 21564 71884 21624
rect 66368 21494 66510 21558
rect 66574 21494 66580 21558
rect 66368 21488 66580 21494
rect 19040 21156 19116 21216
rect 19584 21156 19660 21216
rect 17816 21150 18028 21156
rect 17816 21086 17958 21150
rect 18022 21086 18028 21150
rect 17816 21014 18028 21086
rect 17816 20950 17958 21014
rect 18022 20950 18028 21014
rect 17816 20944 18028 20950
rect 544 20878 3748 20884
rect 544 20814 550 20878
rect 614 20814 3678 20878
rect 3742 20814 3748 20878
rect 544 20808 3748 20814
rect 3128 20748 3340 20808
rect 3808 20748 4020 20884
rect 13872 20808 14900 20884
rect 13872 20748 13948 20808
rect 14824 20748 14900 20808
rect 15096 20808 15716 20884
rect 18224 20808 18436 21156
rect 18632 21150 18980 21156
rect 18632 21086 18910 21150
rect 18974 21086 18980 21150
rect 18632 20884 18980 21086
rect 19040 21014 19252 21156
rect 19040 20950 19046 21014
rect 19110 20950 19252 21014
rect 19040 20944 19252 20950
rect 19448 21014 19660 21156
rect 19448 20950 19590 21014
rect 19654 20950 19660 21014
rect 19448 20944 19660 20950
rect 24344 21286 24692 21292
rect 24344 21222 24486 21286
rect 24550 21222 24622 21286
rect 24686 21222 24692 21286
rect 24344 20944 24692 21222
rect 66368 21286 66580 21292
rect 66368 21222 66510 21286
rect 66574 21222 66580 21286
rect 66368 21150 66580 21222
rect 71264 21216 71476 21564
rect 71672 21216 71884 21564
rect 72080 21830 72292 21836
rect 72080 21766 72086 21830
rect 72150 21766 72292 21830
rect 72080 21624 72292 21766
rect 72488 21624 72700 21836
rect 72896 21830 73108 21972
rect 72896 21766 72902 21830
rect 72966 21766 73108 21830
rect 72896 21760 73108 21766
rect 74936 21624 75556 21700
rect 72080 21564 72156 21624
rect 72488 21564 72564 21624
rect 74936 21564 75012 21624
rect 75480 21564 75556 21624
rect 72080 21428 72292 21564
rect 72488 21428 72700 21564
rect 72080 21422 72700 21428
rect 72080 21358 72222 21422
rect 72286 21358 72700 21422
rect 72080 21352 72700 21358
rect 72896 21558 73108 21564
rect 72896 21494 72902 21558
rect 72966 21494 73108 21558
rect 72896 21422 73108 21494
rect 72896 21358 73038 21422
rect 73102 21358 73108 21422
rect 72896 21352 73108 21358
rect 74664 21488 75012 21564
rect 75072 21558 75284 21564
rect 75072 21494 75078 21558
rect 75142 21494 75284 21558
rect 72216 21292 72292 21352
rect 72216 21216 72564 21292
rect 74664 21286 74876 21488
rect 74664 21222 74806 21286
rect 74870 21222 74876 21286
rect 74664 21216 74876 21222
rect 75072 21292 75284 21494
rect 75480 21558 75692 21564
rect 75480 21494 75486 21558
rect 75550 21494 75692 21558
rect 75480 21422 75692 21494
rect 75480 21358 75486 21422
rect 75550 21358 75692 21422
rect 75480 21352 75692 21358
rect 75888 21422 76100 21564
rect 75888 21358 75894 21422
rect 75958 21358 76100 21422
rect 75888 21352 76100 21358
rect 75888 21292 75964 21352
rect 75072 21286 75964 21292
rect 75072 21222 75078 21286
rect 75142 21222 75964 21286
rect 75072 21216 75964 21222
rect 71400 21156 71476 21216
rect 71808 21156 71884 21216
rect 72488 21156 72564 21216
rect 66368 21086 66510 21150
rect 66574 21086 66580 21150
rect 66368 20944 66580 21086
rect 71264 21014 71476 21156
rect 71264 20950 71406 21014
rect 71470 20950 71476 21014
rect 71264 20944 71476 20950
rect 71672 21014 71884 21156
rect 71672 20950 71814 21014
rect 71878 20950 71884 21014
rect 71672 20944 71884 20950
rect 72080 21150 72292 21156
rect 72080 21086 72222 21150
rect 72286 21086 72292 21150
rect 24616 20884 24692 20944
rect 66504 20884 66580 20944
rect 18534 20878 18980 20884
rect 18496 20814 18502 20878
rect 18566 20814 18980 20878
rect 18534 20808 18980 20814
rect 15096 20748 15172 20808
rect 15640 20748 15716 20808
rect 18360 20748 18436 20808
rect 1632 20612 1844 20748
rect 1632 20556 1718 20612
rect 1774 20556 1844 20612
rect 1632 20476 1844 20556
rect 3128 20672 4020 20748
rect 3128 20536 3340 20672
rect 3808 20606 4020 20672
rect 3808 20542 3950 20606
rect 4014 20542 4020 20606
rect 3808 20536 4020 20542
rect 13600 20672 13948 20748
rect 13600 20606 13812 20672
rect 13600 20542 13606 20606
rect 13670 20542 13812 20606
rect 13600 20536 13812 20542
rect 14008 20612 14220 20748
rect 14824 20672 15172 20748
rect 14008 20606 14764 20612
rect 14008 20542 14014 20606
rect 14078 20542 14764 20606
rect 14008 20536 14764 20542
rect 14824 20536 15036 20672
rect 15232 20612 15444 20748
rect 15640 20742 15852 20748
rect 15640 20678 15782 20742
rect 15846 20678 15852 20742
rect 15232 20536 15580 20612
rect 15640 20536 15852 20678
rect 16048 20742 16260 20748
rect 16048 20678 16190 20742
rect 16254 20678 16260 20742
rect 16048 20536 16260 20678
rect 17816 20742 18028 20748
rect 17816 20678 17958 20742
rect 18022 20678 18028 20742
rect 17816 20536 18028 20678
rect 18224 20672 18980 20748
rect 18224 20612 18436 20672
rect 18224 20606 18572 20612
rect 18224 20542 18502 20606
rect 18566 20542 18572 20606
rect 18224 20536 18572 20542
rect 18632 20536 18980 20672
rect 19040 20742 19252 20748
rect 19040 20678 19046 20742
rect 19110 20678 19252 20742
rect 19040 20606 19252 20678
rect 19040 20542 19046 20606
rect 19110 20542 19252 20606
rect 19040 20536 19252 20542
rect 19448 20742 19660 20748
rect 19448 20678 19590 20742
rect 19654 20678 19660 20742
rect 19448 20606 19660 20678
rect 24344 20672 24692 20884
rect 24616 20612 24692 20672
rect 19448 20542 19454 20606
rect 19518 20542 19660 20606
rect 19448 20536 19660 20542
rect 1224 20470 1844 20476
rect 1224 20406 1230 20470
rect 1294 20406 1844 20470
rect 1224 20400 1844 20406
rect 14688 20476 14764 20536
rect 15232 20476 15308 20536
rect 14688 20400 15308 20476
rect 15504 20476 15580 20536
rect 16048 20476 16124 20536
rect 15504 20400 16124 20476
rect 24344 20400 24692 20612
rect 66368 20878 66580 20884
rect 66368 20814 66510 20878
rect 66574 20814 66580 20878
rect 66368 20672 66580 20814
rect 72080 20808 72292 21086
rect 72488 20808 72700 21156
rect 72896 21150 73108 21156
rect 72896 21086 73038 21150
rect 73102 21086 73108 21150
rect 72896 21014 73108 21086
rect 72896 20950 73038 21014
rect 73102 20950 73108 21014
rect 72896 20944 73108 20950
rect 75752 20808 76916 20884
rect 72080 20748 72156 20808
rect 72488 20748 72564 20808
rect 75752 20748 75828 20808
rect 76840 20748 76916 20808
rect 71264 20742 71476 20748
rect 71264 20678 71406 20742
rect 71470 20678 71476 20742
rect 66368 20612 66444 20672
rect 66368 20400 66580 20612
rect 71264 20536 71476 20678
rect 71672 20742 71884 20748
rect 71672 20678 71814 20742
rect 71878 20678 71884 20742
rect 71672 20536 71884 20678
rect 72080 20536 72292 20748
rect 72488 20536 72700 20748
rect 72896 20742 73108 20748
rect 72896 20678 73038 20742
rect 73102 20678 73108 20742
rect 72896 20536 73108 20678
rect 74664 20742 74876 20748
rect 74664 20678 74806 20742
rect 74870 20678 74876 20742
rect 74664 20536 74876 20678
rect 75072 20742 75284 20748
rect 75072 20678 75078 20742
rect 75142 20678 75284 20742
rect 75072 20536 75284 20678
rect 75480 20742 75828 20748
rect 75480 20678 75486 20742
rect 75550 20678 75828 20742
rect 75480 20672 75828 20678
rect 75888 20742 76100 20748
rect 75888 20678 75894 20742
rect 75958 20678 76100 20742
rect 75480 20536 75692 20672
rect 75888 20612 76100 20678
rect 76840 20612 77052 20748
rect 77248 20612 77460 20748
rect 89080 20612 89428 20748
rect 75888 20536 76780 20612
rect 76840 20606 77188 20612
rect 76840 20542 77118 20606
rect 77182 20542 77188 20606
rect 76840 20536 77188 20542
rect 77248 20606 79908 20612
rect 77248 20542 79838 20606
rect 79902 20542 79908 20606
rect 77248 20536 79908 20542
rect 89080 20556 89216 20612
rect 89272 20606 89836 20612
rect 89272 20556 89766 20606
rect 89080 20542 89766 20556
rect 89830 20542 89836 20606
rect 89080 20536 89836 20542
rect 76704 20476 76780 20536
rect 77248 20476 77324 20536
rect 76704 20400 77324 20476
rect 89080 20400 89428 20536
rect 24480 20340 24556 20400
rect 66504 20340 66580 20400
rect 24344 20204 24692 20340
rect 19448 20198 19660 20204
rect 19448 20134 19454 20198
rect 19518 20134 19660 20198
rect 19448 20068 19660 20134
rect 20264 20068 20612 20204
rect 24072 20128 24692 20204
rect 66368 20204 66580 20340
rect 79832 20334 80044 20340
rect 79832 20270 79838 20334
rect 79902 20270 80044 20334
rect 66368 20198 66988 20204
rect 66368 20134 66374 20198
rect 66438 20134 66988 20198
rect 66368 20128 66988 20134
rect 79832 20198 80044 20270
rect 79832 20134 79974 20198
rect 80038 20134 80044 20198
rect 79832 20128 80044 20134
rect 19448 19992 20612 20068
rect 19448 19932 19660 19992
rect 19214 19926 19660 19932
rect 19176 19862 19182 19926
rect 19246 19862 19660 19926
rect 19214 19856 19660 19862
rect 20264 19932 20612 19992
rect 22984 19932 23196 20068
rect 24072 19992 24284 20128
rect 66776 19992 66988 20128
rect 79288 19938 79372 19942
rect 79255 19933 79372 19938
rect 20264 19856 25236 19932
rect 79255 19877 79260 19933
rect 79316 19877 79372 19933
rect 79255 19872 79372 19877
rect 79288 19868 79372 19872
rect 25160 19796 25236 19856
rect 25160 19660 25372 19796
rect 25704 19660 25916 19796
rect 26384 19720 27820 19796
rect 26384 19660 26596 19720
rect 25160 19654 26596 19660
rect 25160 19590 25302 19654
rect 25366 19590 26526 19654
rect 26590 19590 26596 19654
rect 25160 19584 26596 19590
rect 26928 19584 27140 19720
rect 27608 19660 27820 19720
rect 28152 19660 28500 19796
rect 27608 19654 28500 19660
rect 27608 19590 28158 19654
rect 28222 19590 28500 19654
rect 27608 19584 28500 19590
rect 28832 19720 29724 19796
rect 28832 19584 29044 19720
rect 29512 19660 29724 19720
rect 30056 19660 30268 19796
rect 30736 19720 31628 19796
rect 30736 19660 30948 19720
rect 29512 19654 30268 19660
rect 30366 19654 30948 19660
rect 29512 19590 29518 19654
rect 29582 19590 29654 19654
rect 29718 19590 30268 19654
rect 30328 19590 30334 19654
rect 30398 19590 30948 19654
rect 29512 19584 30268 19590
rect 30366 19584 30948 19590
rect 31280 19654 31628 19720
rect 31280 19590 31558 19654
rect 31622 19590 31628 19654
rect 31280 19584 31628 19590
rect 31960 19660 32172 19796
rect 32640 19660 32852 19796
rect 31960 19654 32852 19660
rect 31960 19590 31966 19654
rect 32030 19590 32646 19654
rect 32710 19590 32852 19654
rect 31960 19584 32852 19590
rect 33184 19720 34076 19796
rect 33184 19654 33396 19720
rect 33184 19590 33190 19654
rect 33254 19590 33396 19654
rect 33184 19584 33396 19590
rect 33864 19660 34076 19720
rect 34408 19720 35300 19796
rect 34408 19660 34756 19720
rect 33864 19654 34756 19660
rect 33864 19590 34550 19654
rect 34614 19590 34756 19654
rect 33864 19584 34756 19590
rect 35088 19654 35300 19720
rect 35088 19590 35230 19654
rect 35294 19590 35300 19654
rect 35088 19584 35300 19590
rect 35768 19660 35980 19796
rect 36312 19660 36524 19796
rect 36992 19720 38428 19796
rect 36992 19660 37204 19720
rect 35768 19654 37204 19660
rect 35768 19590 35774 19654
rect 35838 19590 36454 19654
rect 36518 19590 37204 19654
rect 35768 19584 37204 19590
rect 37536 19584 37748 19720
rect 38216 19660 38428 19720
rect 38760 19720 40332 19796
rect 38760 19660 39108 19720
rect 38216 19654 39108 19660
rect 38216 19590 38358 19654
rect 38422 19590 39108 19654
rect 38216 19584 39108 19590
rect 39440 19584 39652 19720
rect 40120 19660 40332 19720
rect 40664 19660 40876 19796
rect 41344 19720 42780 19796
rect 41344 19660 41556 19720
rect 40120 19654 41556 19660
rect 40120 19590 40806 19654
rect 40870 19590 41486 19654
rect 41550 19590 41556 19654
rect 40120 19584 41556 19590
rect 41888 19584 42236 19720
rect 42568 19660 42780 19720
rect 43248 19720 44004 19796
rect 43248 19660 43460 19720
rect 42568 19654 43460 19660
rect 42568 19590 42710 19654
rect 42774 19590 43460 19654
rect 42568 19584 43460 19590
rect 43792 19654 44004 19720
rect 43792 19590 43934 19654
rect 43998 19590 44004 19654
rect 43792 19584 44004 19590
rect 44472 19660 44684 19796
rect 45016 19720 46588 19796
rect 45016 19660 45364 19720
rect 44472 19654 45636 19660
rect 44472 19590 44478 19654
rect 44542 19590 45566 19654
rect 45630 19590 45636 19654
rect 44472 19584 45636 19590
rect 45696 19584 45908 19720
rect 46376 19660 46588 19720
rect 46920 19660 47132 19796
rect 47600 19720 48356 19796
rect 47600 19660 47812 19720
rect 48144 19660 48356 19720
rect 46376 19654 47812 19660
rect 47910 19654 48356 19660
rect 46376 19590 46926 19654
rect 46990 19590 47812 19654
rect 47872 19590 47878 19654
rect 47942 19590 48356 19654
rect 46376 19584 47812 19590
rect 47910 19584 48356 19590
rect 48824 19660 49036 19796
rect 49368 19660 49716 19796
rect 50048 19660 50260 19796
rect 48824 19654 50260 19660
rect 48824 19590 49374 19654
rect 49438 19590 50190 19654
rect 50254 19590 50260 19654
rect 48824 19584 50260 19590
rect 50728 19660 50940 19796
rect 51272 19660 51484 19796
rect 51952 19720 52844 19796
rect 51952 19660 52164 19720
rect 50728 19654 52164 19660
rect 50728 19590 50734 19654
rect 50798 19590 51958 19654
rect 52022 19590 52164 19654
rect 50728 19584 52164 19590
rect 52496 19660 52844 19720
rect 53176 19660 53388 19796
rect 53856 19720 55292 19796
rect 53856 19660 54068 19720
rect 54400 19660 54612 19720
rect 52496 19654 54068 19660
rect 54166 19654 54612 19660
rect 52496 19590 53182 19654
rect 53246 19590 54068 19654
rect 54128 19590 54134 19654
rect 54198 19590 54612 19654
rect 52496 19584 54068 19590
rect 54166 19584 54612 19590
rect 55080 19660 55292 19720
rect 55624 19660 55972 19796
rect 56304 19720 57196 19796
rect 56304 19660 56516 19720
rect 55080 19654 56516 19660
rect 55080 19590 55766 19654
rect 55830 19590 56516 19654
rect 55080 19584 56516 19590
rect 56984 19660 57196 19720
rect 57528 19660 57740 19796
rect 56984 19654 57740 19660
rect 56984 19590 56990 19654
rect 57054 19590 57740 19654
rect 56984 19584 57740 19590
rect 58208 19720 58964 19796
rect 58208 19654 58420 19720
rect 58208 19590 58214 19654
rect 58278 19590 58420 19654
rect 58208 19584 58420 19590
rect 58752 19654 58964 19720
rect 58752 19590 58894 19654
rect 58958 19590 58964 19654
rect 58752 19584 58964 19590
rect 59432 19660 59644 19796
rect 59976 19660 60324 19796
rect 59432 19654 60324 19660
rect 59432 19590 59438 19654
rect 59502 19590 60118 19654
rect 60182 19590 60324 19654
rect 59432 19584 60324 19590
rect 60656 19720 61548 19796
rect 60656 19654 60868 19720
rect 60656 19590 60662 19654
rect 60726 19590 60868 19654
rect 60656 19584 60868 19590
rect 61336 19660 61548 19720
rect 61880 19660 62092 19796
rect 62560 19720 63996 19796
rect 62560 19660 62772 19720
rect 63104 19660 63452 19720
rect 61336 19654 62772 19660
rect 62870 19654 63452 19660
rect 61336 19590 61886 19654
rect 61950 19590 62772 19654
rect 62832 19590 62838 19654
rect 62902 19590 63452 19654
rect 61336 19584 62772 19590
rect 62870 19584 63452 19590
rect 63784 19660 63996 19720
rect 64464 19720 65900 19796
rect 64464 19660 64676 19720
rect 63784 19654 64676 19660
rect 63784 19590 63926 19654
rect 63990 19590 64676 19654
rect 63784 19584 64676 19590
rect 65008 19584 65220 19720
rect 65688 19654 65900 19720
rect 65688 19590 65694 19654
rect 65758 19590 65900 19654
rect 80240 19720 91060 19796
rect 80240 19677 80452 19720
rect 80240 19621 80342 19677
rect 80398 19621 80452 19677
rect 65688 19584 65900 19590
rect 79054 19608 79120 19611
rect 79392 19608 79458 19611
rect 79054 19606 79458 19608
rect 79054 19550 79059 19606
rect 79115 19550 79397 19606
rect 79453 19550 79458 19606
rect 80240 19584 80452 19621
rect 79054 19548 79458 19550
rect 79054 19545 79120 19548
rect 79392 19545 79458 19548
rect 3128 19312 4020 19388
rect 3128 19246 3340 19312
rect 3128 19182 3134 19246
rect 3198 19182 3340 19246
rect 3128 19176 3340 19182
rect 3808 19176 4020 19312
rect 11560 19382 13676 19388
rect 11560 19318 13606 19382
rect 13670 19318 13676 19382
rect 11560 19312 13676 19318
rect 11560 19246 11772 19312
rect 11560 19182 11566 19246
rect 11630 19182 11772 19246
rect 11560 19176 11772 19182
rect 25160 19110 25780 19116
rect 25160 19046 25302 19110
rect 25366 19046 25780 19110
rect 25160 19040 25780 19046
rect 1632 18974 3204 18980
rect 1632 18932 3134 18974
rect 1632 18876 1718 18932
rect 1774 18910 3134 18932
rect 3198 18910 3204 18974
rect 1774 18904 3204 18910
rect 25160 18904 25508 19040
rect 25568 18904 25780 19040
rect 26520 19110 27140 19116
rect 26520 19046 26526 19110
rect 26590 19046 27140 19110
rect 26520 19040 27140 19046
rect 26520 18904 26732 19040
rect 26792 18974 27140 19040
rect 26792 18910 26798 18974
rect 26862 18910 27140 18974
rect 26792 18904 27140 18910
rect 27744 18980 27956 19116
rect 28152 19110 28364 19116
rect 28152 19046 28158 19110
rect 28222 19046 28364 19110
rect 28152 18980 28364 19046
rect 28968 19110 29588 19116
rect 29686 19110 30812 19116
rect 28968 19046 29518 19110
rect 29582 19046 29588 19110
rect 29648 19046 29654 19110
rect 29718 19046 30334 19110
rect 30398 19046 30812 19110
rect 28968 19040 29588 19046
rect 29686 19040 30812 19046
rect 28968 18980 29180 19040
rect 27744 18904 29180 18980
rect 29376 18904 29588 19040
rect 30192 18904 30404 19040
rect 30600 18974 30812 19040
rect 30600 18910 30742 18974
rect 30806 18910 30812 18974
rect 30600 18904 30812 18910
rect 31416 19110 32036 19116
rect 31416 19046 31558 19110
rect 31622 19046 31966 19110
rect 32030 19046 32036 19110
rect 31416 19040 32036 19046
rect 31416 18904 31628 19040
rect 31824 18904 32036 19040
rect 32640 19110 32988 19116
rect 32640 19046 32646 19110
rect 32710 19046 32988 19110
rect 32640 18980 32988 19046
rect 33048 19110 33260 19116
rect 33048 19046 33190 19110
rect 33254 19046 33260 19110
rect 33048 18980 33260 19046
rect 32640 18904 33260 18980
rect 34000 19110 34620 19116
rect 34000 19046 34550 19110
rect 34614 19046 34620 19110
rect 34000 19040 34620 19046
rect 34000 18904 34212 19040
rect 34272 18904 34620 19040
rect 35224 19110 35844 19116
rect 35224 19046 35230 19110
rect 35294 19046 35774 19110
rect 35838 19046 35844 19110
rect 35224 19040 35844 19046
rect 35224 18904 35436 19040
rect 35632 18904 35844 19040
rect 36448 19110 36660 19116
rect 36448 19046 36454 19110
rect 36518 19046 36660 19110
rect 36448 18980 36660 19046
rect 36856 18980 37068 19116
rect 36448 18974 37068 18980
rect 36448 18910 36454 18974
rect 36518 18910 37068 18974
rect 36448 18904 37068 18910
rect 37672 19040 38292 19116
rect 38390 19110 39516 19116
rect 38352 19046 38358 19110
rect 38422 19046 39516 19110
rect 38390 19040 39516 19046
rect 37672 18904 37884 19040
rect 38080 18980 38292 19040
rect 38896 18980 39244 19040
rect 38080 18904 39244 18980
rect 39304 18904 39516 19040
rect 40256 18980 40468 19116
rect 40528 19110 40876 19116
rect 40528 19046 40806 19110
rect 40870 19046 40876 19110
rect 40528 18980 40876 19046
rect 40256 18904 40876 18980
rect 41480 19110 42100 19116
rect 41480 19046 41486 19110
rect 41550 19046 42100 19110
rect 41480 19040 42100 19046
rect 41480 18974 41692 19040
rect 41480 18910 41486 18974
rect 41550 18910 41692 18974
rect 41480 18904 41692 18910
rect 41888 18904 42100 19040
rect 42704 19110 43324 19116
rect 42704 19046 42710 19110
rect 42774 19046 43324 19110
rect 42704 19040 43324 19046
rect 42704 18904 42916 19040
rect 43112 18904 43324 19040
rect 43928 19110 44548 19116
rect 43928 19046 43934 19110
rect 43998 19046 44478 19110
rect 44542 19046 44548 19110
rect 43928 19040 44548 19046
rect 43928 18904 44140 19040
rect 44336 18904 44548 19040
rect 45152 18980 45364 19116
rect 45560 19110 45772 19116
rect 45560 19046 45566 19110
rect 45630 19046 45772 19110
rect 45560 18980 45772 19046
rect 45152 18974 45772 18980
rect 45152 18910 45702 18974
rect 45766 18910 45772 18974
rect 45152 18904 45772 18910
rect 46376 18980 46724 19116
rect 46784 19110 46996 19116
rect 46784 19046 46926 19110
rect 46990 19046 46996 19110
rect 46784 18980 46996 19046
rect 46376 18904 46996 18980
rect 47736 19110 48356 19116
rect 47736 19046 47878 19110
rect 47942 19046 48356 19110
rect 47736 19040 48356 19046
rect 47736 18904 47948 19040
rect 48008 18980 48356 19040
rect 48960 18980 49172 19116
rect 49368 19110 49580 19116
rect 49368 19046 49374 19110
rect 49438 19046 49580 19110
rect 49368 18980 49580 19046
rect 48008 18904 49580 18980
rect 50184 19110 50804 19116
rect 50184 19046 50190 19110
rect 50254 19046 50734 19110
rect 50798 19046 50804 19110
rect 50184 19040 50804 19046
rect 50184 18904 50396 19040
rect 50592 18904 50804 19040
rect 51408 19110 52028 19116
rect 51408 19046 51958 19110
rect 52022 19046 52028 19110
rect 51408 19040 52028 19046
rect 51408 18974 51620 19040
rect 51408 18910 51414 18974
rect 51478 18910 51620 18974
rect 51408 18904 51620 18910
rect 51816 18904 52028 19040
rect 52632 19110 53252 19116
rect 52632 19046 53182 19110
rect 53246 19046 53252 19110
rect 52632 19040 53252 19046
rect 52632 18904 52844 19040
rect 53040 18904 53252 19040
rect 53856 19110 54476 19116
rect 53856 19046 54134 19110
rect 54198 19046 54476 19110
rect 53856 19040 54476 19046
rect 53856 18904 54204 19040
rect 54264 18904 54476 19040
rect 55216 19110 55836 19116
rect 55216 19046 55766 19110
rect 55830 19046 55836 19110
rect 55216 19040 55836 19046
rect 55216 18904 55428 19040
rect 55488 18974 55836 19040
rect 55488 18910 55766 18974
rect 55830 18910 55836 18974
rect 55488 18904 55836 18910
rect 56440 19110 57876 19116
rect 56440 19046 56990 19110
rect 57054 19046 57876 19110
rect 56440 19040 57876 19046
rect 56440 18904 56652 19040
rect 56848 18904 57060 19040
rect 57664 18980 57876 19040
rect 58072 19110 58284 19116
rect 58072 19046 58214 19110
rect 58278 19046 58284 19110
rect 58072 18980 58284 19046
rect 57664 18904 58284 18980
rect 58888 19110 59508 19116
rect 58888 19046 58894 19110
rect 58958 19046 59438 19110
rect 59502 19046 59508 19110
rect 58888 19040 59508 19046
rect 58888 18904 59100 19040
rect 59296 18904 59508 19040
rect 60112 19110 60460 19116
rect 60112 19046 60118 19110
rect 60182 19046 60460 19110
rect 60112 18980 60460 19046
rect 60520 19110 60732 19116
rect 60520 19046 60662 19110
rect 60726 19046 60732 19110
rect 60520 18980 60732 19046
rect 60112 18904 60732 18980
rect 61472 18980 61684 19116
rect 61744 19110 62092 19116
rect 61744 19046 61886 19110
rect 61950 19046 62092 19110
rect 61744 18980 62092 19046
rect 61472 18974 62092 18980
rect 61472 18910 61478 18974
rect 61542 18910 62092 18974
rect 61472 18904 62092 18910
rect 62696 19110 63316 19116
rect 62696 19046 62838 19110
rect 62902 19046 63316 19110
rect 62696 19040 63316 19046
rect 62696 18904 62908 19040
rect 63104 18904 63316 19040
rect 63920 19110 64540 19116
rect 63920 19046 63926 19110
rect 63990 19046 64540 19110
rect 63920 19040 64540 19046
rect 63920 18904 64132 19040
rect 64328 18904 64540 19040
rect 65144 19110 65764 19116
rect 65144 19046 65694 19110
rect 65758 19046 65764 19110
rect 65144 19040 65764 19046
rect 65144 18904 65356 19040
rect 77150 18974 80044 18980
rect 77112 18910 77118 18974
rect 77182 18910 80044 18974
rect 77150 18904 80044 18910
rect 1774 18876 1844 18904
rect 1632 18844 1844 18876
rect 1224 18838 1844 18844
rect 1224 18774 1230 18838
rect 1294 18774 1844 18838
rect 1224 18768 1844 18774
rect 79832 18702 80044 18904
rect 89080 18932 89428 18980
rect 89080 18876 89216 18932
rect 89272 18876 89428 18932
rect 89080 18844 89428 18876
rect 89080 18838 89836 18844
rect 89080 18774 89766 18838
rect 89830 18774 89836 18838
rect 89080 18768 89836 18774
rect 79832 18638 79838 18702
rect 79902 18638 80044 18702
rect 79832 18632 80044 18638
rect 11669 18622 11735 18625
rect 19811 18622 19877 18625
rect 11669 18620 19877 18622
rect 11669 18564 11674 18620
rect 11730 18564 19816 18620
rect 19872 18564 19877 18620
rect 11669 18562 19877 18564
rect 11669 18559 11735 18562
rect 19811 18559 19877 18562
rect 2455 18261 2461 18325
rect 2525 18323 2531 18325
rect 2525 18263 25447 18323
rect 2525 18261 2531 18263
rect 78974 18050 79040 18053
rect 79392 18050 79458 18053
rect 78974 18048 79458 18050
rect 3128 17892 3340 18028
rect 3808 18022 4020 18028
rect 3808 17958 3950 18022
rect 4014 17958 4020 18022
rect 3808 17892 4020 17958
rect 3128 17816 4020 17892
rect 11560 18022 14084 18028
rect 11560 17958 14014 18022
rect 14078 17958 14084 18022
rect 78974 17992 78979 18048
rect 79035 17992 79397 18048
rect 79453 17992 79458 18048
rect 78974 17990 79458 17992
rect 78974 17987 79040 17990
rect 79392 17987 79458 17990
rect 11560 17952 14084 17958
rect 80240 17977 91060 18028
rect 11560 17886 11772 17952
rect 11560 17822 11702 17886
rect 11766 17822 11772 17886
rect 11560 17816 11772 17822
rect 80240 17921 80342 17977
rect 80398 17952 91060 17977
rect 80398 17921 80452 17952
rect 80240 17816 80452 17921
rect 16456 17620 16668 17756
rect 17816 17750 19116 17756
rect 17816 17686 19046 17750
rect 19110 17686 19116 17750
rect 17816 17680 19116 17686
rect 17816 17620 18028 17680
rect 16456 17614 18028 17620
rect 16456 17550 16598 17614
rect 16662 17550 18028 17614
rect 16456 17544 18028 17550
rect 25976 17484 26324 17620
rect 27336 17484 27548 17620
rect 28560 17544 29996 17620
rect 28560 17484 28772 17544
rect 25976 17478 28772 17484
rect 25976 17414 25982 17478
rect 26046 17414 28772 17478
rect 25976 17408 28772 17414
rect 29784 17484 29996 17544
rect 31008 17544 32444 17620
rect 31008 17484 31220 17544
rect 29784 17478 31220 17484
rect 29784 17414 31150 17478
rect 31214 17414 31220 17478
rect 29784 17408 31220 17414
rect 32232 17484 32444 17544
rect 33456 17544 36252 17620
rect 33456 17484 33804 17544
rect 32232 17408 33804 17484
rect 34816 17408 35028 17544
rect 36040 17484 36252 17544
rect 37264 17544 38700 17620
rect 37264 17484 37476 17544
rect 36040 17478 37476 17484
rect 36040 17414 36182 17478
rect 36246 17414 37476 17478
rect 36040 17408 37476 17414
rect 38488 17484 38700 17544
rect 39712 17544 42508 17620
rect 39712 17484 40060 17544
rect 41072 17484 41284 17544
rect 38488 17408 40060 17484
rect 40974 17478 41284 17484
rect 40936 17414 40942 17478
rect 41006 17414 41284 17478
rect 40974 17408 41284 17414
rect 42296 17484 42508 17544
rect 43520 17544 44956 17620
rect 43520 17484 43732 17544
rect 42296 17408 43732 17484
rect 44744 17484 44956 17544
rect 45968 17544 47540 17620
rect 45968 17484 46180 17544
rect 44744 17478 46180 17484
rect 44744 17414 45974 17478
rect 46038 17414 46180 17478
rect 44744 17408 46180 17414
rect 47192 17484 47540 17544
rect 48552 17484 48764 17620
rect 49776 17544 51212 17620
rect 49776 17484 49988 17544
rect 47192 17408 49988 17484
rect 51000 17484 51212 17544
rect 52224 17544 53660 17620
rect 52224 17484 52436 17544
rect 51000 17478 52436 17484
rect 51000 17414 51142 17478
rect 51206 17414 52436 17478
rect 51000 17408 52436 17414
rect 53448 17484 53660 17544
rect 54672 17484 55020 17620
rect 56032 17544 57468 17620
rect 56032 17484 56244 17544
rect 53448 17478 56244 17484
rect 53448 17414 56174 17478
rect 56238 17414 56244 17478
rect 53448 17408 56244 17414
rect 57256 17484 57468 17544
rect 58480 17544 59916 17620
rect 58480 17484 58692 17544
rect 57256 17408 58692 17484
rect 59704 17484 59916 17544
rect 60928 17544 63724 17620
rect 60928 17484 61276 17544
rect 59704 17478 61276 17484
rect 59704 17414 60934 17478
rect 60998 17414 61276 17478
rect 59704 17408 61276 17414
rect 62288 17408 62500 17544
rect 63512 17484 63724 17544
rect 64736 17614 66444 17620
rect 64736 17550 66374 17614
rect 66438 17550 66444 17614
rect 64736 17544 66444 17550
rect 64736 17484 64948 17544
rect 63512 17408 64948 17484
rect 79832 17478 80044 17484
rect 79832 17414 79974 17478
rect 80038 17414 80044 17478
rect 1632 17252 1844 17348
rect 79832 17342 80044 17414
rect 79832 17278 79974 17342
rect 80038 17278 80044 17342
rect 79832 17272 80044 17278
rect 1632 17212 1718 17252
rect 1224 17206 1718 17212
rect 1224 17142 1230 17206
rect 1294 17196 1718 17206
rect 1774 17212 1844 17252
rect 89080 17252 89428 17348
rect 1774 17206 2524 17212
rect 1774 17196 2454 17206
rect 1294 17142 2454 17196
rect 2518 17142 2524 17206
rect 1224 17136 2524 17142
rect 89080 17196 89216 17252
rect 89272 17212 89428 17252
rect 89272 17206 89836 17212
rect 89272 17196 89766 17206
rect 89080 17142 89766 17196
rect 89830 17142 89836 17206
rect 89080 17136 89836 17142
rect 80240 16864 91060 16940
rect 80240 16849 80452 16864
rect 80240 16793 80342 16849
rect 80398 16793 80452 16849
rect 78894 16780 78960 16783
rect 79392 16780 79458 16783
rect 78894 16778 79458 16780
rect 78894 16722 78899 16778
rect 78955 16722 79397 16778
rect 79453 16722 79458 16778
rect 80240 16728 80452 16793
rect 78894 16720 79458 16722
rect 78894 16717 78960 16720
rect 79392 16717 79458 16720
rect 2486 16526 3340 16532
rect 2448 16462 2454 16526
rect 2518 16462 3340 16526
rect 2486 16456 3340 16462
rect 3128 16396 3340 16456
rect 3808 16396 4020 16532
rect 11560 16526 11772 16532
rect 11560 16462 11566 16526
rect 11630 16462 11772 16526
rect 11560 16396 11772 16462
rect 3128 16320 4020 16396
rect 11424 16390 11772 16396
rect 11424 16326 11430 16390
rect 11494 16326 11772 16390
rect 11424 16320 11772 16326
rect 16456 16390 19252 16396
rect 16456 16326 19182 16390
rect 19246 16326 19252 16390
rect 16456 16320 19252 16326
rect 16456 16254 16668 16320
rect 16456 16190 16462 16254
rect 16526 16190 16668 16254
rect 16456 16184 16668 16190
rect 17816 16184 18028 16320
rect 79832 16118 80044 16124
rect 79832 16054 79838 16118
rect 79902 16054 80044 16118
rect 79832 15982 80044 16054
rect 79832 15918 79838 15982
rect 79902 15918 80044 15982
rect 79832 15912 80044 15918
rect 11669 15792 11735 15797
rect 11669 15736 11674 15792
rect 11730 15777 11735 15792
rect 11730 15772 23580 15777
rect 11730 15736 23519 15772
rect 11669 15717 23519 15736
rect 23514 15716 23519 15717
rect 23575 15716 23580 15772
rect 1224 15710 1844 15716
rect 23514 15711 23580 15716
rect 1224 15646 1230 15710
rect 1294 15646 1844 15710
rect 1224 15640 1844 15646
rect 1632 15572 1844 15640
rect 1632 15516 1718 15572
rect 1774 15516 1844 15572
rect 1632 15368 1844 15516
rect 89080 15580 89428 15716
rect 89080 15574 89836 15580
rect 89080 15572 89766 15574
rect 89080 15516 89216 15572
rect 89272 15516 89766 15572
rect 89080 15510 89766 15516
rect 89830 15510 89836 15574
rect 89080 15504 89836 15510
rect 89080 15368 89428 15504
rect 78814 15222 78880 15225
rect 79392 15222 79458 15225
rect 78814 15220 79458 15222
rect 544 15166 3340 15172
rect 544 15102 550 15166
rect 614 15102 3340 15166
rect 544 15096 3340 15102
rect 3128 15036 3340 15096
rect 3808 15036 4020 15172
rect 3128 14960 4020 15036
rect 11560 15166 11772 15172
rect 11560 15102 11702 15166
rect 11766 15102 11772 15166
rect 78814 15164 78819 15220
rect 78875 15164 79397 15220
rect 79453 15164 79458 15220
rect 78814 15162 79458 15164
rect 78814 15159 78880 15162
rect 79392 15159 79458 15162
rect 11560 15030 11772 15102
rect 80240 15149 91060 15172
rect 80240 15093 80342 15149
rect 80398 15096 91060 15149
rect 80398 15093 80452 15096
rect 25929 15036 26027 15068
rect 30921 15036 31019 15068
rect 35913 15036 36011 15068
rect 40905 15036 41003 15068
rect 45897 15036 45995 15068
rect 50889 15036 50987 15068
rect 55881 15036 55979 15068
rect 60873 15036 60971 15068
rect 11560 14966 11566 15030
rect 11630 14966 11772 15030
rect 11560 14960 11772 14966
rect 25840 15030 26150 15036
rect 30872 15030 31220 15036
rect 25840 14966 25982 15030
rect 26046 14966 26118 15030
rect 26182 14966 26188 15030
rect 30872 14966 31014 15030
rect 31078 14966 31150 15030
rect 31214 14966 31220 15030
rect 25840 14960 26150 14966
rect 30872 14960 31220 14966
rect 35904 15030 36252 15036
rect 35904 14966 36046 15030
rect 36110 14966 36182 15030
rect 36246 14966 36252 15030
rect 35904 14960 36252 14966
rect 40800 15030 41110 15036
rect 45832 15030 46044 15036
rect 40800 14966 40942 15030
rect 41006 14966 41078 15030
rect 41142 14966 41148 15030
rect 45832 14966 45838 15030
rect 45902 14966 45974 15030
rect 46038 14966 46044 15030
rect 40800 14960 41110 14966
rect 45832 14960 46044 14966
rect 50864 15030 51212 15036
rect 50864 14966 51006 15030
rect 51070 14966 51142 15030
rect 51206 14966 51212 15030
rect 50864 14960 51212 14966
rect 55760 15030 56244 15036
rect 55760 14966 56038 15030
rect 56102 14966 56174 15030
rect 56238 14966 56244 15030
rect 55760 14960 56244 14966
rect 60792 15030 61102 15036
rect 60792 14966 60934 15030
rect 60998 14966 61070 15030
rect 61134 14966 61140 15030
rect 60792 14960 61102 14966
rect 80240 14960 80452 15093
rect 16456 14894 16668 14900
rect 16456 14830 16598 14894
rect 16662 14830 16668 14894
rect 16456 14764 16668 14830
rect 17816 14764 18028 14900
rect 16456 14758 18028 14764
rect 16456 14694 16598 14758
rect 16662 14694 18028 14758
rect 16456 14688 18028 14694
rect 79832 14622 80044 14628
rect 79832 14558 79974 14622
rect 80038 14558 80044 14622
rect 79832 14486 80044 14558
rect 79832 14422 79974 14486
rect 80038 14422 80044 14486
rect 79832 14416 80044 14422
rect 11669 14380 11735 14383
rect 23762 14380 23828 14383
rect 11669 14378 23828 14380
rect 11669 14322 11674 14378
rect 11730 14322 23767 14378
rect 23823 14322 23828 14378
rect 11669 14320 23828 14322
rect 11669 14317 11735 14320
rect 23762 14317 23828 14320
rect 25840 14350 26868 14356
rect 25840 14286 26798 14350
rect 26862 14286 26868 14350
rect 25840 14280 26868 14286
rect 30736 14350 30948 14356
rect 30736 14286 30742 14350
rect 30806 14286 30948 14350
rect 25840 14214 26052 14280
rect 25840 14150 25982 14214
rect 26046 14150 26052 14214
rect 25840 14144 26052 14150
rect 30736 14214 30948 14286
rect 30736 14150 30742 14214
rect 30806 14150 30948 14214
rect 30736 14144 30948 14150
rect 35768 14350 36524 14356
rect 35768 14286 36454 14350
rect 36518 14286 36524 14350
rect 35768 14280 36524 14286
rect 40800 14350 41556 14356
rect 40800 14286 41486 14350
rect 41550 14286 41556 14350
rect 40800 14280 41556 14286
rect 45696 14350 46044 14356
rect 45696 14286 45702 14350
rect 45766 14286 46044 14350
rect 35768 14214 35980 14280
rect 35768 14150 35774 14214
rect 35838 14150 35980 14214
rect 35768 14144 35980 14150
rect 40800 14214 41012 14280
rect 40800 14150 40942 14214
rect 41006 14150 41012 14214
rect 40800 14144 41012 14150
rect 45696 14214 46044 14286
rect 45696 14150 45974 14214
rect 46038 14150 46044 14214
rect 45696 14144 46044 14150
rect 50728 14350 51484 14356
rect 50728 14286 51414 14350
rect 51478 14286 51484 14350
rect 50728 14280 51484 14286
rect 55760 14350 55972 14356
rect 55760 14286 55766 14350
rect 55830 14286 55972 14350
rect 50728 14214 50940 14280
rect 50728 14150 50734 14214
rect 50798 14150 50940 14214
rect 50728 14144 50940 14150
rect 55760 14214 55972 14286
rect 55760 14150 55766 14214
rect 55830 14150 55972 14214
rect 55760 14144 55972 14150
rect 60656 14350 61548 14356
rect 60656 14286 61478 14350
rect 61542 14286 61548 14350
rect 60656 14280 61548 14286
rect 60656 14214 61004 14280
rect 60656 14150 60798 14214
rect 60862 14150 61004 14214
rect 60656 14144 61004 14150
rect 80240 14021 91060 14084
rect 80240 13965 80342 14021
rect 80398 14008 91060 14021
rect 80398 13965 80452 14008
rect 78734 13952 78800 13955
rect 79392 13952 79458 13955
rect 78734 13950 79458 13952
rect 1632 13892 1844 13948
rect 1632 13836 1718 13892
rect 1774 13836 1844 13892
rect 78734 13894 78739 13950
rect 78795 13894 79397 13950
rect 79453 13894 79458 13950
rect 78734 13892 79458 13894
rect 78734 13889 78800 13892
rect 79392 13889 79458 13892
rect 80240 13872 80452 13965
rect 89080 13942 89836 13948
rect 89080 13892 89766 13942
rect 1632 13812 1844 13836
rect 89080 13836 89216 13892
rect 89272 13878 89766 13892
rect 89830 13878 89836 13942
rect 89272 13872 89836 13878
rect 89272 13836 89428 13872
rect 1224 13806 3340 13812
rect 1224 13742 1230 13806
rect 1294 13742 3340 13806
rect 1224 13736 3340 13742
rect 3128 13676 3340 13736
rect 3808 13676 4020 13812
rect 11462 13806 11772 13812
rect 11424 13742 11430 13806
rect 11494 13742 11772 13806
rect 11462 13736 11772 13742
rect 89080 13736 89428 13836
rect 3128 13600 4020 13676
rect 3128 13464 3340 13600
rect 3808 13464 4020 13600
rect 11560 13534 11772 13736
rect 11560 13470 11702 13534
rect 11766 13470 11772 13534
rect 11560 13464 11772 13470
rect 16456 13534 16668 13540
rect 16456 13470 16462 13534
rect 16526 13470 16668 13534
rect 16456 13404 16668 13470
rect 17816 13404 18028 13540
rect 25840 13534 26052 13540
rect 25840 13470 25982 13534
rect 26046 13470 26052 13534
rect 25840 13464 26052 13470
rect 30736 13534 31084 13540
rect 30736 13470 30742 13534
rect 30806 13470 31084 13534
rect 30736 13464 31084 13470
rect 35768 13534 35980 13540
rect 35768 13470 35774 13534
rect 35838 13470 35980 13534
rect 35768 13464 35980 13470
rect 40800 13534 41012 13540
rect 40800 13470 40942 13534
rect 41006 13470 41012 13534
rect 40800 13464 41012 13470
rect 16456 13398 18028 13404
rect 16456 13334 17958 13398
rect 18022 13334 18028 13398
rect 25859 13398 26052 13464
rect 25859 13358 25982 13398
rect 16456 13328 18028 13334
rect 25976 13334 25982 13358
rect 26046 13334 26052 13398
rect 30851 13398 31084 13464
rect 30851 13358 30878 13398
rect 25976 13328 26052 13334
rect 30872 13334 30878 13358
rect 30942 13334 31084 13398
rect 35843 13398 35980 13464
rect 35843 13358 35910 13398
rect 30872 13328 31084 13334
rect 35904 13334 35910 13358
rect 35974 13334 35980 13398
rect 40835 13398 41012 13464
rect 40835 13358 40942 13398
rect 35904 13328 35980 13334
rect 40936 13334 40942 13358
rect 41006 13334 41012 13398
rect 40936 13328 41012 13334
rect 45696 13534 46044 13540
rect 45696 13470 45974 13534
rect 46038 13470 46044 13534
rect 45696 13398 46044 13470
rect 50728 13534 50940 13540
rect 50728 13470 50734 13534
rect 50798 13470 50940 13534
rect 50728 13464 50940 13470
rect 55760 13534 55972 13540
rect 55760 13470 55766 13534
rect 55830 13470 55972 13534
rect 55760 13464 55972 13470
rect 60792 13534 61004 13540
rect 60792 13470 60798 13534
rect 60862 13470 61004 13534
rect 60792 13464 61004 13470
rect 45696 13334 45702 13398
rect 45766 13334 46044 13398
rect 50819 13398 50940 13464
rect 50819 13358 50870 13398
rect 45696 13328 46044 13334
rect 50864 13334 50870 13358
rect 50934 13334 50940 13398
rect 55811 13398 55972 13464
rect 55811 13358 55902 13398
rect 50864 13328 50940 13334
rect 55896 13334 55902 13358
rect 55966 13334 55972 13398
rect 60803 13398 61004 13464
rect 60803 13358 60934 13398
rect 55896 13328 55972 13334
rect 60928 13334 60934 13358
rect 60998 13334 61004 13398
rect 60928 13328 61004 13334
rect 25568 13132 25780 13268
rect 25976 13262 26188 13268
rect 25976 13198 26118 13262
rect 26182 13198 26188 13262
rect 25976 13192 26188 13198
rect 25976 13134 26052 13192
rect 25568 13076 25626 13132
rect 25682 13076 25780 13132
rect 25568 12996 25780 13076
rect 25859 13036 26052 13134
rect 25296 12990 25780 12996
rect 11669 12982 11735 12985
rect 23638 12982 23704 12985
rect 11669 12980 23704 12982
rect 11669 12924 11674 12980
rect 11730 12924 23643 12980
rect 23699 12924 23704 12980
rect 11669 12922 23704 12924
rect 11669 12919 11735 12922
rect 23638 12919 23704 12922
rect 25296 12926 25302 12990
rect 25366 12926 25780 12990
rect 25296 12920 25780 12926
rect 25976 12860 26052 13036
rect 30464 13153 30676 13268
rect 30872 13262 31084 13268
rect 30872 13198 31014 13262
rect 31078 13198 31084 13262
rect 30464 13132 30695 13153
rect 30872 13134 31084 13198
rect 30464 13076 30618 13132
rect 30674 13076 30695 13132
rect 30464 13055 30695 13076
rect 30464 12990 30676 13055
rect 30851 13036 31084 13134
rect 30464 12926 30470 12990
rect 30534 12926 30676 12990
rect 30464 12920 30676 12926
rect 30872 12990 31084 13036
rect 30872 12926 31014 12990
rect 31078 12926 31084 12990
rect 30872 12920 31084 12926
rect 35496 13132 35708 13268
rect 35904 13262 36116 13268
rect 35904 13198 36046 13262
rect 36110 13198 36116 13262
rect 35904 13192 36116 13198
rect 35904 13134 35980 13192
rect 35496 13076 35610 13132
rect 35666 13076 35708 13132
rect 35496 12990 35708 13076
rect 35843 13036 35980 13134
rect 35496 12926 35502 12990
rect 35566 12926 35708 12990
rect 35496 12920 35708 12926
rect 35904 12860 35980 13036
rect 40528 13132 40740 13268
rect 40936 13262 41148 13268
rect 40936 13198 41078 13262
rect 41142 13198 41148 13262
rect 40936 13192 41148 13198
rect 40936 13134 41012 13192
rect 40528 13076 40602 13132
rect 40658 13076 40740 13132
rect 40528 12990 40740 13076
rect 40835 13036 41012 13134
rect 40528 12926 40534 12990
rect 40598 12926 40740 12990
rect 40528 12920 40740 12926
rect 40936 12860 41012 13036
rect 45560 13153 45636 13268
rect 45832 13262 46044 13268
rect 45832 13198 45838 13262
rect 45902 13198 46044 13262
rect 45560 13132 45671 13153
rect 45832 13134 46044 13198
rect 45560 13076 45594 13132
rect 45650 13076 45671 13132
rect 45560 13055 45671 13076
rect 45560 12990 45636 13055
rect 45827 13036 46044 13134
rect 45560 12926 45566 12990
rect 45630 12926 45636 12990
rect 45560 12920 45636 12926
rect 45832 12990 46044 13036
rect 45832 12926 45838 12990
rect 45902 12926 46044 12990
rect 45832 12920 46044 12926
rect 50456 13132 50668 13268
rect 50864 13262 51076 13268
rect 50864 13198 51006 13262
rect 51070 13198 51076 13262
rect 50864 13192 51076 13198
rect 50864 13134 50940 13192
rect 50456 13076 50586 13132
rect 50642 13076 50668 13132
rect 50456 12990 50668 13076
rect 50819 13036 50940 13134
rect 50456 12926 50462 12990
rect 50526 12926 50668 12990
rect 50456 12920 50668 12926
rect 50864 12860 50940 13036
rect 55488 13132 55700 13268
rect 55896 13262 56108 13268
rect 55896 13198 56038 13262
rect 56102 13198 56108 13262
rect 55896 13192 56108 13198
rect 55896 13134 55972 13192
rect 55488 13076 55578 13132
rect 55634 13076 55700 13132
rect 55488 12990 55700 13076
rect 55811 13036 55972 13134
rect 55488 12926 55494 12990
rect 55558 12926 55700 12990
rect 55488 12920 55700 12926
rect 55896 12860 55972 13036
rect 60520 13132 60732 13268
rect 60928 13262 61140 13268
rect 60928 13198 61070 13262
rect 61134 13198 61140 13262
rect 60928 13192 61140 13198
rect 79832 13262 80044 13268
rect 79832 13198 79838 13262
rect 79902 13198 80044 13262
rect 60928 13134 61004 13192
rect 60520 13076 60570 13132
rect 60626 13076 60732 13132
rect 60520 12990 60732 13076
rect 60803 13036 61004 13134
rect 79832 13126 80044 13198
rect 79832 13062 79838 13126
rect 79902 13062 80044 13126
rect 79832 13056 80044 13062
rect 60520 12926 60526 12990
rect 60590 12926 60732 12990
rect 60520 12920 60732 12926
rect 60928 12860 61004 13036
rect 25878 12854 26052 12860
rect 35806 12854 35980 12860
rect 40838 12854 41012 12860
rect 50766 12854 50940 12860
rect 55798 12854 55972 12860
rect 60830 12854 61004 12860
rect 25840 12790 25846 12854
rect 25910 12790 26052 12854
rect 35768 12790 35774 12854
rect 35838 12790 35980 12854
rect 40800 12790 40806 12854
rect 40870 12790 41012 12854
rect 50728 12790 50734 12854
rect 50798 12790 50940 12854
rect 55760 12790 55766 12854
rect 55830 12790 55972 12854
rect 60792 12790 60798 12854
rect 60862 12790 61004 12854
rect 25878 12784 26052 12790
rect 35806 12784 35980 12790
rect 40838 12784 41012 12790
rect 50766 12784 50940 12790
rect 55798 12784 55972 12790
rect 60830 12784 61004 12790
rect 25704 12446 25916 12452
rect 25704 12382 25846 12446
rect 25910 12382 25916 12446
rect 1224 12310 1844 12316
rect 1224 12246 1230 12310
rect 1294 12246 1844 12310
rect 1224 12240 1844 12246
rect 1632 12212 1844 12240
rect 1632 12156 1718 12212
rect 1774 12156 1844 12212
rect 1632 12104 1844 12156
rect 11560 12310 11772 12316
rect 11560 12246 11566 12310
rect 11630 12246 11772 12310
rect 11560 12174 11772 12246
rect 25704 12310 25916 12382
rect 25704 12246 25846 12310
rect 25910 12246 25916 12310
rect 25704 12240 25916 12246
rect 30736 12446 31084 12452
rect 30736 12382 31014 12446
rect 31078 12382 31084 12446
rect 30736 12376 31084 12382
rect 35632 12446 35844 12452
rect 35632 12382 35774 12446
rect 35838 12382 35844 12446
rect 30736 12310 30948 12376
rect 30736 12246 30742 12310
rect 30806 12246 30948 12310
rect 30736 12240 30948 12246
rect 35632 12310 35844 12382
rect 35632 12246 35638 12310
rect 35702 12246 35844 12310
rect 35632 12240 35844 12246
rect 40664 12446 40876 12452
rect 40664 12382 40806 12446
rect 40870 12382 40876 12446
rect 40664 12316 40876 12382
rect 45696 12446 45908 12452
rect 45696 12382 45838 12446
rect 45902 12382 45908 12446
rect 40664 12310 41148 12316
rect 40664 12246 41078 12310
rect 41142 12246 41148 12310
rect 40664 12240 41148 12246
rect 45696 12310 45908 12382
rect 45696 12246 45838 12310
rect 45902 12246 45908 12310
rect 45696 12240 45908 12246
rect 50592 12446 50804 12452
rect 50592 12382 50734 12446
rect 50798 12382 50804 12446
rect 50592 12316 50804 12382
rect 55624 12446 55836 12452
rect 55624 12382 55766 12446
rect 55830 12382 55836 12446
rect 55624 12316 55836 12382
rect 60656 12446 60868 12452
rect 60656 12382 60798 12446
rect 60862 12382 60868 12446
rect 50592 12310 51076 12316
rect 50592 12246 51006 12310
rect 51070 12246 51076 12310
rect 50592 12240 51076 12246
rect 55624 12310 56108 12316
rect 55624 12246 56038 12310
rect 56102 12246 56108 12310
rect 55624 12240 56108 12246
rect 60656 12310 60868 12382
rect 78654 12394 78720 12397
rect 79392 12394 79458 12397
rect 78654 12392 79458 12394
rect 78654 12336 78659 12392
rect 78715 12336 79397 12392
rect 79453 12336 79458 12392
rect 78654 12334 79458 12336
rect 78654 12331 78720 12334
rect 79392 12331 79458 12334
rect 80240 12376 91060 12452
rect 60656 12246 60662 12310
rect 60726 12246 60868 12310
rect 60656 12240 60868 12246
rect 80240 12321 80452 12376
rect 80240 12265 80342 12321
rect 80398 12265 80452 12321
rect 80240 12240 80452 12265
rect 89080 12310 89836 12316
rect 89080 12246 89766 12310
rect 89830 12246 89836 12310
rect 89080 12240 89836 12246
rect 89080 12212 89428 12240
rect 11560 12110 11566 12174
rect 11630 12110 11772 12174
rect 11560 12104 11772 12110
rect 16456 12174 16668 12180
rect 16456 12110 16598 12174
rect 16662 12110 16668 12174
rect 16456 11908 16668 12110
rect 17816 11908 18028 12180
rect 89080 12156 89216 12212
rect 89272 12156 89428 12212
rect 89080 12104 89428 12156
rect 16456 11902 18028 11908
rect 16456 11838 16598 11902
rect 16662 11838 18028 11902
rect 16456 11832 18028 11838
rect 25704 11902 26052 11908
rect 25704 11838 25982 11902
rect 26046 11838 26052 11902
rect 25704 11832 26052 11838
rect 30600 11902 30948 11908
rect 30600 11838 30878 11902
rect 30942 11838 30948 11902
rect 25704 11766 25916 11832
rect 25704 11702 25710 11766
rect 25774 11702 25916 11766
rect 25704 11696 25916 11702
rect 30600 11766 30948 11838
rect 30600 11702 30878 11766
rect 30942 11702 30948 11766
rect 30600 11696 30948 11702
rect 35632 11902 35980 11908
rect 35632 11838 35910 11902
rect 35974 11838 35980 11902
rect 35632 11832 35980 11838
rect 40664 11902 41012 11908
rect 40664 11838 40942 11902
rect 41006 11838 41012 11902
rect 40664 11832 41012 11838
rect 45696 11902 45908 11908
rect 45696 11838 45702 11902
rect 45766 11838 45908 11902
rect 35632 11766 35844 11832
rect 35632 11702 35774 11766
rect 35838 11702 35844 11766
rect 35632 11696 35844 11702
rect 40664 11766 40876 11832
rect 40664 11702 40806 11766
rect 40870 11702 40876 11766
rect 40664 11696 40876 11702
rect 45696 11766 45908 11838
rect 45696 11702 45702 11766
rect 45766 11702 45908 11766
rect 45696 11696 45908 11702
rect 50592 11902 50940 11908
rect 50592 11838 50870 11902
rect 50934 11838 50940 11902
rect 50592 11832 50940 11838
rect 55624 11902 55972 11908
rect 55624 11838 55902 11902
rect 55966 11838 55972 11902
rect 55624 11832 55972 11838
rect 60656 11902 61004 11908
rect 60656 11838 60934 11902
rect 60998 11838 61004 11902
rect 60656 11832 61004 11838
rect 79832 11902 80044 11908
rect 79832 11838 79974 11902
rect 80038 11838 80044 11902
rect 50592 11766 50804 11832
rect 50592 11702 50734 11766
rect 50798 11702 50804 11766
rect 50592 11696 50804 11702
rect 55624 11766 55836 11832
rect 55624 11702 55766 11766
rect 55830 11702 55836 11766
rect 55624 11696 55836 11702
rect 60656 11766 60868 11832
rect 60656 11702 60798 11766
rect 60862 11702 60868 11766
rect 60656 11696 60868 11702
rect 25840 11630 26052 11636
rect 25840 11566 25846 11630
rect 25910 11566 26052 11630
rect 25840 11500 26052 11566
rect 30736 11630 30948 11636
rect 35670 11630 35980 11636
rect 30736 11566 30742 11630
rect 30806 11566 30948 11630
rect 35632 11566 35638 11630
rect 35702 11566 35980 11630
rect 30736 11500 30948 11566
rect 35670 11560 35980 11566
rect 35768 11500 35980 11560
rect 40800 11630 41110 11636
rect 45696 11630 46044 11636
rect 40800 11566 41078 11630
rect 41142 11566 41148 11630
rect 45696 11566 45838 11630
rect 45902 11566 46044 11630
rect 40800 11560 41110 11566
rect 40800 11500 41012 11560
rect 25704 11424 26052 11500
rect 25704 11228 25916 11424
rect 25198 11222 25916 11228
rect 25160 11158 25166 11222
rect 25230 11158 25916 11222
rect 25198 11152 25916 11158
rect 30600 11152 30948 11500
rect 35632 11424 35980 11500
rect 40664 11424 41012 11500
rect 45696 11424 46044 11566
rect 50728 11630 51038 11636
rect 55760 11630 56070 11636
rect 60694 11630 61004 11636
rect 50728 11566 51006 11630
rect 51070 11566 51076 11630
rect 55760 11566 56038 11630
rect 56102 11566 56108 11630
rect 60656 11566 60662 11630
rect 60726 11566 61004 11630
rect 50728 11560 51038 11566
rect 55760 11560 56070 11566
rect 60694 11560 61004 11566
rect 79832 11560 80044 11838
rect 50728 11500 50940 11560
rect 55760 11500 55972 11560
rect 60792 11500 61004 11560
rect 50592 11424 50940 11500
rect 55624 11424 55972 11500
rect 60656 11494 65492 11500
rect 60656 11430 65422 11494
rect 65486 11430 65492 11494
rect 60656 11424 65492 11430
rect 35632 11152 35844 11424
rect 40664 11152 40876 11424
rect 45696 11152 45908 11424
rect 50592 11152 50804 11424
rect 55624 11152 55836 11424
rect 60656 11152 60868 11424
rect 80240 11193 80452 11228
rect 80240 11137 80342 11193
rect 80398 11137 80452 11193
rect 78574 11124 78640 11127
rect 79392 11124 79458 11127
rect 78574 11122 79458 11124
rect 78574 11066 78579 11122
rect 78635 11066 79397 11122
rect 79453 11066 79458 11122
rect 78574 11064 79458 11066
rect 78574 11061 78640 11064
rect 79392 11061 79458 11064
rect 80240 11092 80452 11137
rect 80240 11016 91060 11092
rect 544 10950 2660 10956
rect 544 10886 550 10950
rect 614 10886 2660 10950
rect 544 10880 2660 10886
rect 2448 10744 2660 10880
rect 11560 10950 11772 10956
rect 25606 10950 25916 10956
rect 11560 10886 11702 10950
rect 11766 10886 11772 10950
rect 25568 10886 25574 10950
rect 25638 10886 25710 10950
rect 25774 10886 25916 10950
rect 11560 10814 11772 10886
rect 25606 10880 25916 10886
rect 30736 10950 30948 10956
rect 30736 10886 30878 10950
rect 30942 10886 30948 10950
rect 30736 10880 30948 10886
rect 35632 10950 35844 10956
rect 35632 10886 35774 10950
rect 35838 10886 35844 10950
rect 35632 10880 35844 10886
rect 40664 10950 40876 10956
rect 40664 10886 40806 10950
rect 40870 10886 40876 10950
rect 40664 10880 40876 10886
rect 45696 10950 45908 10956
rect 45696 10886 45702 10950
rect 45766 10886 45908 10950
rect 45696 10880 45908 10886
rect 50592 10950 50940 10956
rect 50592 10886 50734 10950
rect 50798 10886 50940 10950
rect 50592 10880 50940 10886
rect 55624 10950 55836 10956
rect 55624 10886 55766 10950
rect 55830 10886 55836 10950
rect 55624 10880 55836 10886
rect 60656 10950 65356 10956
rect 60656 10886 60798 10950
rect 60862 10886 65286 10950
rect 65350 10886 65356 10950
rect 60656 10880 65356 10886
rect 25754 10856 25852 10880
rect 30746 10856 30844 10880
rect 35738 10856 35836 10880
rect 40730 10856 40828 10880
rect 45722 10856 45820 10880
rect 50714 10856 50812 10880
rect 55706 10856 55804 10880
rect 60698 10856 60796 10880
rect 11560 10750 11702 10814
rect 11766 10750 11772 10814
rect 11560 10744 11772 10750
rect 1632 10548 1844 10684
rect 1224 10542 1844 10548
rect 1224 10478 1230 10542
rect 1294 10532 1844 10542
rect 1294 10478 1718 10532
rect 1224 10476 1718 10478
rect 1774 10476 1844 10532
rect 1224 10472 1844 10476
rect 16456 10678 18028 10684
rect 16456 10614 17958 10678
rect 18022 10614 18028 10678
rect 16456 10608 18028 10614
rect 16456 10542 16668 10608
rect 16456 10478 16462 10542
rect 16526 10478 16668 10542
rect 16456 10472 16668 10478
rect 17816 10472 18028 10608
rect 24072 10542 25644 10548
rect 24072 10478 25574 10542
rect 25638 10478 25644 10542
rect 24072 10472 25644 10478
rect 65280 10542 65628 10548
rect 65280 10478 65286 10542
rect 65350 10478 65628 10542
rect 1697 10455 1795 10472
rect 2584 10279 2796 10412
rect 24072 10336 24284 10472
rect 65280 10336 65628 10478
rect 89080 10532 89428 10684
rect 89080 10476 89216 10532
rect 89272 10476 89428 10532
rect 89080 10412 89428 10476
rect 79832 10406 80044 10412
rect 79832 10342 79838 10406
rect 79902 10342 80044 10406
rect 2584 10276 2678 10279
rect 0 10223 2678 10276
rect 2734 10223 2796 10279
rect 0 10200 2796 10223
rect 79832 10200 80044 10342
rect 89080 10406 89836 10412
rect 89080 10342 89766 10406
rect 89830 10342 89836 10406
rect 89080 10336 89836 10342
rect 2448 9318 2660 9460
rect 2448 9254 2454 9318
rect 2518 9254 2660 9318
rect 2448 9248 2660 9254
rect 11560 9454 11772 9460
rect 11560 9390 11566 9454
rect 11630 9390 11772 9454
rect 11560 9248 11772 9390
rect 24072 9454 25236 9460
rect 24072 9390 25166 9454
rect 25230 9390 25236 9454
rect 24072 9384 25236 9390
rect 65280 9454 65628 9460
rect 65280 9390 65422 9454
rect 65486 9390 65628 9454
rect 16456 9318 18028 9324
rect 16456 9254 16598 9318
rect 16662 9254 18028 9318
rect 16456 9248 18028 9254
rect 24072 9248 24284 9384
rect 65280 9248 65628 9390
rect 16456 9182 16668 9248
rect 16456 9118 16598 9182
rect 16662 9118 16668 9182
rect 16456 9112 16668 9118
rect 17816 9112 18028 9248
rect 1224 8910 2524 8916
rect 1224 8846 1230 8910
rect 1294 8852 2454 8910
rect 1294 8846 1718 8852
rect 1224 8840 1718 8846
rect 1697 8796 1718 8840
rect 1774 8846 2454 8852
rect 2518 8846 2524 8910
rect 1774 8840 2524 8846
rect 89080 8852 89428 8916
rect 1774 8796 1795 8840
rect 1697 8775 1795 8796
rect 89080 8796 89216 8852
rect 89272 8796 89428 8852
rect 89080 8780 89428 8796
rect 5848 8684 6060 8780
rect 89080 8774 89836 8780
rect 89080 8710 89766 8774
rect 89830 8710 89836 8774
rect 89080 8704 89836 8710
rect 5848 8644 5899 8684
rect 0 8579 2796 8644
rect 0 8568 2678 8579
rect 2584 8523 2678 8568
rect 2734 8523 2796 8579
rect 2856 8638 5899 8644
rect 2856 8574 2862 8638
rect 2926 8628 5899 8638
rect 5955 8628 6060 8684
rect 2926 8574 6060 8628
rect 2856 8568 6060 8574
rect 2584 8432 2796 8523
rect 0 8366 2894 8372
rect 0 8302 2862 8366
rect 2926 8302 2932 8366
rect 0 8296 2894 8302
rect 2448 7964 2660 8100
rect 544 7958 2660 7964
rect 544 7894 550 7958
rect 614 7894 2660 7958
rect 544 7888 2660 7894
rect 11560 8094 11772 8100
rect 11560 8030 11702 8094
rect 11766 8030 11772 8094
rect 11560 7888 11772 8030
rect 16456 7822 16668 7828
rect 16456 7758 16462 7822
rect 16526 7758 16668 7822
rect 16456 7692 16668 7758
rect 17816 7692 18028 7828
rect 16456 7686 18028 7692
rect 16456 7622 16462 7686
rect 16526 7622 18028 7686
rect 16456 7616 18028 7622
rect 1632 7172 1844 7284
rect 1632 7148 1718 7172
rect 1224 7142 1718 7148
rect 1224 7078 1230 7142
rect 1294 7116 1718 7142
rect 1774 7116 1844 7172
rect 1294 7078 1844 7116
rect 1224 7072 1844 7078
rect 89080 7278 89836 7284
rect 89080 7214 89766 7278
rect 89830 7214 89836 7278
rect 89080 7208 89836 7214
rect 89080 7172 89428 7208
rect 89080 7116 89216 7172
rect 89272 7116 89428 7172
rect 89080 7072 89428 7116
rect 16456 6462 16668 6468
rect 16456 6398 16598 6462
rect 16662 6398 16668 6462
rect 16456 6332 16668 6398
rect 17816 6332 18028 6468
rect 16456 6256 18028 6332
rect 1632 5492 1844 5516
rect 1632 5436 1718 5492
rect 1774 5436 1844 5492
rect 1632 5380 1844 5436
rect 1224 5374 1844 5380
rect 1224 5310 1230 5374
rect 1294 5310 1844 5374
rect 1224 5304 1844 5310
rect 89080 5492 89428 5516
rect 89080 5436 89216 5492
rect 89272 5436 89428 5492
rect 89080 5380 89428 5436
rect 89080 5374 89836 5380
rect 89080 5310 89766 5374
rect 89830 5310 89836 5374
rect 89080 5304 89836 5310
rect 13328 3944 14764 4020
rect 1632 3812 1844 3884
rect 1632 3756 1718 3812
rect 1774 3756 1844 3812
rect 1632 3748 1844 3756
rect 1224 3742 1844 3748
rect 1224 3678 1230 3742
rect 1294 3678 1844 3742
rect 1224 3672 1844 3678
rect 13328 3672 13540 3944
rect 14552 3748 14764 3944
rect 15640 4014 16532 4020
rect 15640 3950 16462 4014
rect 16526 3950 16532 4014
rect 15640 3944 16532 3950
rect 15640 3884 15852 3944
rect 16864 3884 17076 4020
rect 17952 3944 19388 4020
rect 17952 3884 18300 3944
rect 15640 3808 18300 3884
rect 15640 3748 15852 3808
rect 14552 3672 15852 3748
rect 16864 3672 17076 3808
rect 17952 3672 18300 3808
rect 19176 3884 19388 3944
rect 20413 3884 20511 3903
rect 21581 3884 21679 3903
rect 22749 3884 22847 3903
rect 23917 3884 24015 3903
rect 25085 3884 25183 3903
rect 26253 3884 26351 3903
rect 19176 3808 24148 3884
rect 19176 3672 19388 3808
rect 20400 3672 20612 3808
rect 21488 3672 21700 3808
rect 22712 3672 22924 3808
rect 23800 3748 24148 3808
rect 25024 3748 25236 3884
rect 26248 3748 26460 3884
rect 23800 3742 26460 3748
rect 23800 3678 25166 3742
rect 25230 3678 26460 3742
rect 23800 3672 26460 3678
rect 89080 3812 89428 3884
rect 89080 3756 89216 3812
rect 89272 3756 89428 3812
rect 89080 3748 89428 3756
rect 89080 3742 89836 3748
rect 89080 3678 89766 3742
rect 89830 3678 89836 3742
rect 89080 3672 89836 3678
rect 12920 3032 13132 3068
rect 12920 2976 13012 3032
rect 13068 2976 13132 3032
rect 12920 2926 13132 2976
rect 12920 2862 12926 2926
rect 12990 2862 13132 2926
rect 12920 2856 13132 2862
rect 14144 3032 14356 3068
rect 14144 2976 14180 3032
rect 14236 2976 14356 3032
rect 14144 2926 14356 2976
rect 14144 2862 14286 2926
rect 14350 2862 14356 2926
rect 14144 2856 14356 2862
rect 15232 3032 15444 3068
rect 15232 2976 15348 3032
rect 15404 2976 15444 3032
rect 15232 2926 15444 2976
rect 15232 2862 15374 2926
rect 15438 2862 15444 2926
rect 15232 2856 15444 2862
rect 16456 3032 16668 3068
rect 17680 3053 17892 3068
rect 18904 3053 18980 3068
rect 16456 2976 16516 3032
rect 16572 2976 16668 3032
rect 16456 2926 16668 2976
rect 17663 3032 17892 3053
rect 17663 2976 17684 3032
rect 17740 2976 17892 3032
rect 17663 2932 17892 2976
rect 18831 3032 18980 3053
rect 18831 2976 18852 3032
rect 18908 2976 18980 3032
rect 18831 2932 18980 2976
rect 16456 2862 16462 2926
rect 16526 2862 16668 2926
rect 16456 2856 16668 2862
rect 17544 2926 17892 2932
rect 17544 2862 17686 2926
rect 17750 2862 17892 2926
rect 17544 2856 17892 2862
rect 18768 2926 18980 2932
rect 18768 2862 18910 2926
rect 18974 2862 18980 2926
rect 18768 2856 18980 2862
rect 19992 3032 20204 3068
rect 21216 3053 21292 3068
rect 19992 2976 20020 3032
rect 20076 2976 20204 3032
rect 19992 2926 20204 2976
rect 21167 3032 21292 3053
rect 21167 2976 21188 3032
rect 21244 2976 21292 3032
rect 21167 2932 21292 2976
rect 19992 2862 19998 2926
rect 20062 2862 20204 2926
rect 19992 2856 20204 2862
rect 21080 2926 21292 2932
rect 21080 2862 21086 2926
rect 21150 2862 21292 2926
rect 21080 2856 21292 2862
rect 22304 3032 22516 3068
rect 23528 3053 23604 3068
rect 24752 3053 24828 3068
rect 25840 3053 26052 3068
rect 22304 2976 22356 3032
rect 22412 2976 22516 3032
rect 22304 2926 22516 2976
rect 23503 3032 23604 3053
rect 23503 2976 23524 3032
rect 23580 2976 23604 3032
rect 23503 2932 23604 2976
rect 24671 3032 24828 3053
rect 24671 2976 24692 3032
rect 24748 2976 24828 3032
rect 24671 2932 24828 2976
rect 25839 3032 26052 3053
rect 25839 2976 25860 3032
rect 25916 2976 26052 3032
rect 25839 2932 26052 2976
rect 22304 2862 22310 2926
rect 22374 2862 22516 2926
rect 22304 2856 22516 2862
rect 23392 2926 23604 2932
rect 23392 2862 23398 2926
rect 23462 2862 23604 2926
rect 23392 2856 23604 2862
rect 24616 2926 24828 2932
rect 24616 2862 24758 2926
rect 24822 2862 24828 2926
rect 24616 2856 24828 2862
rect 25704 2926 26052 2932
rect 25704 2862 25710 2926
rect 25774 2862 26052 2926
rect 25704 2856 26052 2862
rect 11753 2778 11819 2781
rect 11753 2776 14622 2778
rect 11753 2720 11758 2776
rect 11814 2720 14622 2776
rect 11753 2718 14622 2720
rect 11753 2715 11819 2718
rect 13328 2448 17076 2524
rect 13328 2382 13540 2448
rect 13328 2318 13334 2382
rect 13398 2318 13540 2382
rect 13328 2312 13540 2318
rect 14552 2312 14764 2448
rect 15640 2312 15852 2448
rect 16864 2388 17076 2448
rect 17952 2448 19388 2524
rect 17952 2388 18300 2448
rect 16864 2312 18300 2388
rect 19176 2388 19388 2448
rect 20400 2388 20612 2524
rect 21488 2388 21700 2524
rect 22712 2388 22924 2524
rect 23800 2448 26460 2524
rect 23800 2388 24148 2448
rect 19176 2312 24148 2388
rect 25024 2312 25236 2448
rect 26248 2312 26460 2448
rect 1632 2132 1844 2252
rect 1632 2076 1718 2132
rect 1774 2116 1844 2132
rect 89080 2132 89428 2252
rect 1774 2110 1980 2116
rect 1774 2076 1910 2110
rect 1632 2046 1910 2076
rect 1974 2046 1980 2110
rect 1632 2040 1980 2046
rect 89080 2076 89216 2132
rect 89272 2116 89428 2132
rect 89272 2110 89836 2116
rect 89272 2076 89766 2110
rect 89080 2046 89766 2076
rect 89830 2046 89836 2110
rect 89080 2040 89836 2046
rect 1904 1838 2252 1844
rect 1904 1774 1910 1838
rect 1974 1796 2252 1838
rect 1974 1774 2054 1796
rect 1904 1740 2054 1774
rect 2110 1740 2252 1796
rect 1904 1702 2252 1740
rect 1904 1638 1910 1702
rect 1974 1638 2252 1702
rect 1904 1632 2252 1638
rect 3672 1796 3884 1844
rect 3672 1740 3734 1796
rect 3790 1740 3884 1796
rect 3672 1702 3884 1740
rect 3672 1638 3678 1702
rect 3742 1638 3884 1702
rect 3672 1632 3884 1638
rect 5304 1796 5516 1844
rect 5304 1740 5414 1796
rect 5470 1740 5516 1796
rect 5304 1702 5516 1740
rect 5304 1638 5310 1702
rect 5374 1638 5516 1702
rect 5304 1632 5516 1638
rect 7072 1796 7284 1844
rect 7072 1740 7094 1796
rect 7150 1740 7284 1796
rect 7072 1702 7284 1740
rect 7072 1638 7078 1702
rect 7142 1638 7284 1702
rect 7072 1632 7284 1638
rect 8704 1796 8916 1844
rect 8704 1740 8774 1796
rect 8830 1740 8916 1796
rect 8704 1702 8916 1740
rect 8704 1638 8846 1702
rect 8910 1638 8916 1702
rect 8704 1632 8916 1638
rect 10336 1796 10548 1844
rect 10336 1740 10454 1796
rect 10510 1740 10548 1796
rect 10336 1702 10548 1740
rect 10336 1638 10342 1702
rect 10406 1638 10548 1702
rect 10336 1632 10548 1638
rect 12104 1796 12316 1844
rect 12104 1740 12134 1796
rect 12190 1740 12316 1796
rect 12104 1702 12316 1740
rect 12104 1638 12110 1702
rect 12174 1638 12316 1702
rect 12104 1632 12316 1638
rect 13736 1796 13948 1844
rect 13736 1740 13814 1796
rect 13870 1740 13948 1796
rect 13736 1702 13948 1740
rect 13736 1638 13878 1702
rect 13942 1638 13948 1702
rect 13736 1632 13948 1638
rect 15368 1796 15580 1844
rect 15368 1740 15494 1796
rect 15550 1740 15580 1796
rect 15368 1702 15580 1740
rect 15368 1638 15510 1702
rect 15574 1638 15580 1702
rect 15368 1632 15580 1638
rect 17136 1796 17348 1844
rect 17136 1740 17174 1796
rect 17230 1740 17348 1796
rect 17136 1702 17348 1740
rect 17136 1638 17142 1702
rect 17206 1638 17348 1702
rect 17136 1632 17348 1638
rect 18768 1796 18980 1844
rect 18768 1740 18854 1796
rect 18910 1740 18980 1796
rect 18768 1702 18980 1740
rect 18768 1638 18774 1702
rect 18838 1638 18980 1702
rect 18768 1632 18980 1638
rect 20400 1796 20612 1844
rect 20400 1740 20534 1796
rect 20590 1740 20612 1796
rect 20400 1702 20612 1740
rect 20400 1638 20406 1702
rect 20470 1638 20612 1702
rect 20400 1632 20612 1638
rect 22168 1796 22380 1844
rect 22168 1740 22214 1796
rect 22270 1740 22380 1796
rect 22168 1702 22380 1740
rect 22168 1638 22174 1702
rect 22238 1638 22380 1702
rect 22168 1632 22380 1638
rect 23800 1796 24012 1844
rect 25198 1838 25780 1844
rect 23800 1740 23894 1796
rect 23950 1740 24012 1796
rect 25160 1774 25166 1838
rect 25230 1796 25780 1838
rect 25230 1774 25574 1796
rect 25198 1768 25574 1774
rect 23800 1702 24012 1740
rect 23800 1638 23806 1702
rect 23870 1638 24012 1702
rect 23800 1632 24012 1638
rect 25432 1740 25574 1768
rect 25630 1740 25780 1796
rect 25432 1702 25780 1740
rect 25432 1638 25574 1702
rect 25638 1638 25780 1702
rect 25432 1632 25780 1638
rect 27200 1796 27412 1844
rect 27200 1740 27254 1796
rect 27310 1740 27412 1796
rect 27200 1702 27412 1740
rect 27200 1638 27342 1702
rect 27406 1638 27412 1702
rect 27200 1632 27412 1638
rect 28832 1796 29044 1844
rect 28832 1740 28934 1796
rect 28990 1740 29044 1796
rect 28832 1702 29044 1740
rect 28832 1638 28838 1702
rect 28902 1638 29044 1702
rect 28832 1632 29044 1638
rect 30464 1796 30812 1844
rect 30464 1740 30614 1796
rect 30670 1740 30812 1796
rect 30464 1702 30812 1740
rect 30464 1638 30742 1702
rect 30806 1638 30812 1702
rect 30464 1632 30812 1638
rect 32232 1796 32444 1844
rect 32232 1740 32294 1796
rect 32350 1740 32444 1796
rect 32232 1702 32444 1740
rect 32232 1638 32374 1702
rect 32438 1638 32444 1702
rect 32232 1632 32444 1638
rect 33864 1796 34076 1844
rect 33864 1740 33974 1796
rect 34030 1740 34076 1796
rect 33864 1702 34076 1740
rect 33864 1638 33870 1702
rect 33934 1638 34076 1702
rect 33864 1632 34076 1638
rect 35632 1796 35844 1844
rect 35632 1740 35654 1796
rect 35710 1740 35844 1796
rect 35632 1702 35844 1740
rect 35632 1638 35638 1702
rect 35702 1638 35844 1702
rect 35632 1632 35844 1638
rect 37264 1796 37476 1844
rect 37264 1740 37334 1796
rect 37390 1740 37476 1796
rect 37264 1702 37476 1740
rect 37264 1638 37406 1702
rect 37470 1638 37476 1702
rect 37264 1632 37476 1638
rect 38896 1796 39108 1844
rect 38896 1740 39014 1796
rect 39070 1740 39108 1796
rect 38896 1702 39108 1740
rect 38896 1638 38902 1702
rect 38966 1638 39108 1702
rect 38896 1632 39108 1638
rect 40664 1796 40876 1844
rect 40664 1740 40694 1796
rect 40750 1740 40876 1796
rect 40664 1702 40876 1740
rect 40664 1638 40806 1702
rect 40870 1638 40876 1702
rect 40664 1632 40876 1638
rect 42296 1796 42508 1844
rect 42296 1740 42374 1796
rect 42430 1740 42508 1796
rect 42296 1702 42508 1740
rect 42296 1638 42302 1702
rect 42366 1638 42508 1702
rect 42296 1632 42508 1638
rect 43928 1796 44140 1844
rect 43928 1740 44054 1796
rect 44110 1740 44140 1796
rect 43928 1702 44140 1740
rect 43928 1638 43934 1702
rect 43998 1638 44140 1702
rect 43928 1632 44140 1638
rect 45696 1796 45908 1844
rect 45696 1740 45734 1796
rect 45790 1740 45908 1796
rect 45696 1702 45908 1740
rect 45696 1638 45838 1702
rect 45902 1638 45908 1702
rect 45696 1632 45908 1638
rect 47328 1796 47540 1844
rect 47328 1740 47414 1796
rect 47470 1740 47540 1796
rect 47328 1702 47540 1740
rect 47328 1638 47334 1702
rect 47398 1638 47540 1702
rect 47328 1632 47540 1638
rect 48960 1796 49172 1844
rect 48960 1740 49094 1796
rect 49150 1740 49172 1796
rect 48960 1702 49172 1740
rect 48960 1638 49102 1702
rect 49166 1638 49172 1702
rect 48960 1632 49172 1638
rect 50728 1796 50940 1844
rect 50728 1740 50774 1796
rect 50830 1740 50940 1796
rect 50728 1702 50940 1740
rect 50728 1638 50870 1702
rect 50934 1638 50940 1702
rect 50728 1632 50940 1638
rect 52360 1796 52572 1844
rect 52360 1740 52454 1796
rect 52510 1740 52572 1796
rect 52360 1702 52572 1740
rect 52360 1638 52366 1702
rect 52430 1638 52572 1702
rect 52360 1632 52572 1638
rect 53992 1796 54340 1844
rect 53992 1740 54134 1796
rect 54190 1740 54340 1796
rect 53992 1702 54340 1740
rect 53992 1638 54134 1702
rect 54198 1638 54340 1702
rect 53992 1632 54340 1638
rect 55760 1796 55972 1844
rect 55760 1740 55814 1796
rect 55870 1740 55972 1796
rect 55760 1702 55972 1740
rect 55760 1638 55902 1702
rect 55966 1638 55972 1702
rect 55760 1632 55972 1638
rect 57392 1796 57604 1844
rect 57392 1740 57494 1796
rect 57550 1740 57604 1796
rect 57392 1702 57604 1740
rect 57392 1638 57398 1702
rect 57462 1638 57604 1702
rect 57392 1632 57604 1638
rect 59024 1796 59372 1844
rect 59024 1740 59174 1796
rect 59230 1740 59372 1796
rect 59024 1702 59372 1740
rect 59024 1638 59302 1702
rect 59366 1638 59372 1702
rect 59024 1632 59372 1638
rect 60792 1796 61004 1844
rect 60792 1740 60854 1796
rect 60910 1740 61004 1796
rect 60792 1702 61004 1740
rect 60792 1638 60798 1702
rect 60862 1638 61004 1702
rect 60792 1632 61004 1638
rect 62424 1796 62636 1844
rect 62424 1740 62534 1796
rect 62590 1740 62636 1796
rect 62424 1702 62636 1740
rect 62424 1638 62430 1702
rect 62494 1638 62636 1702
rect 62424 1632 62636 1638
rect 64192 1796 64404 1844
rect 64192 1740 64214 1796
rect 64270 1740 64404 1796
rect 64192 1702 64404 1740
rect 64192 1638 64334 1702
rect 64398 1638 64404 1702
rect 64192 1632 64404 1638
rect 65824 1796 66036 1844
rect 65824 1740 65894 1796
rect 65950 1740 66036 1796
rect 65824 1702 66036 1740
rect 65824 1638 65830 1702
rect 65894 1638 66036 1702
rect 65824 1632 66036 1638
rect 67456 1796 67668 1844
rect 67456 1740 67574 1796
rect 67630 1740 67668 1796
rect 67456 1702 67668 1740
rect 67456 1638 67598 1702
rect 67662 1638 67668 1702
rect 67456 1632 67668 1638
rect 69224 1796 69436 1844
rect 69224 1740 69254 1796
rect 69310 1740 69436 1796
rect 69224 1702 69436 1740
rect 69224 1638 69366 1702
rect 69430 1638 69436 1702
rect 69224 1632 69436 1638
rect 70856 1796 71068 1844
rect 70856 1740 70934 1796
rect 70990 1740 71068 1796
rect 70856 1702 71068 1740
rect 70856 1638 70862 1702
rect 70926 1638 71068 1702
rect 70856 1632 71068 1638
rect 72488 1796 72700 1844
rect 72488 1740 72614 1796
rect 72670 1740 72700 1796
rect 72488 1702 72700 1740
rect 72488 1638 72630 1702
rect 72694 1638 72700 1702
rect 72488 1632 72700 1638
rect 74256 1796 74468 1844
rect 74256 1740 74294 1796
rect 74350 1740 74468 1796
rect 74256 1702 74468 1740
rect 74256 1638 74398 1702
rect 74462 1638 74468 1702
rect 74256 1632 74468 1638
rect 75888 1796 76100 1844
rect 75888 1740 75974 1796
rect 76030 1740 76100 1796
rect 75888 1702 76100 1740
rect 75888 1638 75894 1702
rect 75958 1638 76100 1702
rect 75888 1632 76100 1638
rect 77520 1796 77732 1844
rect 77520 1740 77654 1796
rect 77710 1740 77732 1796
rect 77520 1702 77732 1740
rect 77520 1638 77662 1702
rect 77726 1638 77732 1702
rect 77520 1632 77732 1638
rect 79288 1796 79500 1844
rect 79288 1740 79334 1796
rect 79390 1740 79500 1796
rect 79288 1702 79500 1740
rect 79288 1638 79294 1702
rect 79358 1638 79500 1702
rect 79288 1632 79500 1638
rect 80920 1796 81132 1844
rect 80920 1740 81014 1796
rect 81070 1740 81132 1796
rect 80920 1702 81132 1740
rect 80920 1638 80926 1702
rect 80990 1638 81132 1702
rect 80920 1632 81132 1638
rect 82552 1796 82900 1844
rect 82552 1740 82694 1796
rect 82750 1740 82900 1796
rect 82552 1702 82900 1740
rect 82552 1638 82830 1702
rect 82894 1638 82900 1702
rect 82552 1632 82900 1638
rect 84320 1796 84532 1844
rect 84320 1740 84374 1796
rect 84430 1740 84532 1796
rect 84320 1702 84532 1740
rect 84320 1638 84326 1702
rect 84390 1638 84532 1702
rect 84320 1632 84532 1638
rect 85952 1796 86164 1844
rect 85952 1740 86054 1796
rect 86110 1740 86164 1796
rect 85952 1702 86164 1740
rect 85952 1638 86094 1702
rect 86158 1638 86164 1702
rect 85952 1632 86164 1638
rect 87584 1796 87932 1844
rect 87584 1740 87734 1796
rect 87790 1740 87932 1796
rect 87584 1702 87932 1740
rect 87584 1638 87590 1702
rect 87654 1638 87932 1702
rect 87584 1632 87932 1638
rect 952 1294 90108 1300
rect 952 1230 958 1294
rect 1022 1230 1094 1294
rect 1158 1230 1230 1294
rect 1294 1230 1910 1294
rect 1974 1230 3678 1294
rect 3742 1230 5310 1294
rect 5374 1230 7078 1294
rect 7142 1230 8846 1294
rect 8910 1230 10342 1294
rect 10406 1230 12110 1294
rect 12174 1230 13878 1294
rect 13942 1230 15510 1294
rect 15574 1230 17142 1294
rect 17206 1230 18774 1294
rect 18838 1230 20406 1294
rect 20470 1230 22174 1294
rect 22238 1230 23806 1294
rect 23870 1230 25574 1294
rect 25638 1230 27342 1294
rect 27406 1230 28838 1294
rect 28902 1230 30742 1294
rect 30806 1230 32374 1294
rect 32438 1230 33870 1294
rect 33934 1230 35638 1294
rect 35702 1230 37406 1294
rect 37470 1230 38902 1294
rect 38966 1230 40806 1294
rect 40870 1230 42302 1294
rect 42366 1230 43934 1294
rect 43998 1230 45838 1294
rect 45902 1230 47334 1294
rect 47398 1230 49102 1294
rect 49166 1230 50870 1294
rect 50934 1230 52366 1294
rect 52430 1230 54134 1294
rect 54198 1230 55902 1294
rect 55966 1230 57398 1294
rect 57462 1230 59302 1294
rect 59366 1230 60798 1294
rect 60862 1230 62430 1294
rect 62494 1230 64334 1294
rect 64398 1230 65830 1294
rect 65894 1230 67598 1294
rect 67662 1230 69366 1294
rect 69430 1230 70862 1294
rect 70926 1230 72630 1294
rect 72694 1230 74398 1294
rect 74462 1230 75894 1294
rect 75958 1230 77662 1294
rect 77726 1230 79294 1294
rect 79358 1230 80926 1294
rect 80990 1230 82830 1294
rect 82894 1230 84326 1294
rect 84390 1230 86094 1294
rect 86158 1230 87590 1294
rect 87654 1230 89766 1294
rect 89830 1230 89902 1294
rect 89966 1230 90038 1294
rect 90102 1230 90108 1294
rect 952 1158 90108 1230
rect 952 1094 958 1158
rect 1022 1094 1094 1158
rect 1158 1094 1230 1158
rect 1294 1094 89766 1158
rect 89830 1094 89902 1158
rect 89966 1094 90038 1158
rect 90102 1094 90108 1158
rect 952 1022 90108 1094
rect 952 958 958 1022
rect 1022 958 1094 1022
rect 1158 958 1230 1022
rect 1294 958 89766 1022
rect 89830 958 89902 1022
rect 89966 958 90038 1022
rect 90102 958 90108 1022
rect 952 952 90108 958
rect 272 614 90788 620
rect 272 550 278 614
rect 342 550 414 614
rect 478 550 550 614
rect 614 550 13334 614
rect 13398 550 90446 614
rect 90510 550 90582 614
rect 90646 550 90718 614
rect 90782 550 90788 614
rect 272 478 90788 550
rect 272 414 278 478
rect 342 414 414 478
rect 478 414 550 478
rect 614 414 90446 478
rect 90510 414 90582 478
rect 90646 414 90718 478
rect 90782 414 90788 478
rect 272 342 90788 414
rect 272 278 278 342
rect 342 278 414 342
rect 478 278 550 342
rect 614 278 90446 342
rect 90510 278 90582 342
rect 90646 278 90718 342
rect 90782 278 90788 342
rect 272 272 90788 278
<< via3 >>
rect 278 88950 342 89014
rect 414 88950 478 89014
rect 550 88950 614 89014
rect 90446 88950 90510 89014
rect 90582 88950 90646 89014
rect 90718 88950 90782 89014
rect 278 88814 342 88878
rect 414 88814 478 88878
rect 550 88814 614 88878
rect 90446 88814 90510 88878
rect 90582 88814 90646 88878
rect 90718 88814 90782 88878
rect 278 88678 342 88742
rect 414 88678 478 88742
rect 550 88678 614 88742
rect 73990 88678 74054 88742
rect 90446 88678 90510 88742
rect 90582 88678 90646 88742
rect 90718 88678 90782 88742
rect 958 88270 1022 88334
rect 1094 88270 1158 88334
rect 1230 88270 1294 88334
rect 89766 88270 89830 88334
rect 89902 88270 89966 88334
rect 90038 88270 90102 88334
rect 958 88134 1022 88198
rect 1094 88134 1158 88198
rect 1230 88134 1294 88198
rect 89766 88134 89830 88198
rect 89902 88134 89966 88198
rect 90038 88134 90102 88198
rect 958 87998 1022 88062
rect 1094 87998 1158 88062
rect 1230 87998 1294 88062
rect 2182 87998 2246 88062
rect 3814 87998 3878 88062
rect 5310 87998 5374 88062
rect 7078 87998 7142 88062
rect 8846 87998 8910 88062
rect 10342 87998 10406 88062
rect 12110 87998 12174 88062
rect 13878 87998 13942 88062
rect 15374 87998 15438 88062
rect 17278 87998 17342 88062
rect 18910 87998 18974 88062
rect 20542 87998 20606 88062
rect 22174 87998 22238 88062
rect 23942 87998 24006 88062
rect 25438 87998 25502 88062
rect 27342 87998 27406 88062
rect 28838 87998 28902 88062
rect 30470 87998 30534 88062
rect 32374 87998 32438 88062
rect 33870 87998 33934 88062
rect 35910 87998 35974 88062
rect 37406 87998 37470 88062
rect 39038 87998 39102 88062
rect 40942 87998 41006 88062
rect 42438 87998 42502 88062
rect 43934 87998 43998 88062
rect 45838 87998 45902 88062
rect 47334 87998 47398 88062
rect 49102 87998 49166 88062
rect 50870 87998 50934 88062
rect 52502 87998 52566 88062
rect 54270 87998 54334 88062
rect 55902 87998 55966 88062
rect 57398 87998 57462 88062
rect 59302 87998 59366 88062
rect 60934 87998 60998 88062
rect 62566 87998 62630 88062
rect 64334 87998 64398 88062
rect 65966 87998 66030 88062
rect 67598 87998 67662 88062
rect 69366 87998 69430 88062
rect 70862 87998 70926 88062
rect 72630 87998 72694 88062
rect 74262 87998 74326 88062
rect 76030 87998 76094 88062
rect 77662 87998 77726 88062
rect 79430 87998 79494 88062
rect 81062 87998 81126 88062
rect 82558 87998 82622 88062
rect 84326 87998 84390 88062
rect 86094 87998 86158 88062
rect 87862 87998 87926 88062
rect 89766 87998 89830 88062
rect 89902 87998 89966 88062
rect 90038 87998 90102 88062
rect 2182 87590 2246 87654
rect 3814 87590 3878 87654
rect 5310 87590 5374 87654
rect 7078 87590 7142 87654
rect 8846 87590 8910 87654
rect 10342 87590 10406 87654
rect 12110 87590 12174 87654
rect 13878 87590 13942 87654
rect 15374 87590 15438 87654
rect 17278 87590 17342 87654
rect 18910 87590 18974 87654
rect 20542 87590 20606 87654
rect 22174 87590 22238 87654
rect 23942 87590 24006 87654
rect 25438 87590 25502 87654
rect 27342 87590 27406 87654
rect 28838 87590 28902 87654
rect 30470 87590 30534 87654
rect 32374 87590 32438 87654
rect 33870 87590 33934 87654
rect 35910 87590 35974 87654
rect 37406 87590 37470 87654
rect 39038 87590 39102 87654
rect 40942 87590 41006 87654
rect 42438 87590 42502 87654
rect 43934 87590 43998 87654
rect 45838 87590 45902 87654
rect 47334 87590 47398 87654
rect 49102 87590 49166 87654
rect 50870 87590 50934 87654
rect 52502 87590 52566 87654
rect 54270 87590 54334 87654
rect 55902 87590 55966 87654
rect 57398 87590 57462 87654
rect 59302 87590 59366 87654
rect 60934 87590 60998 87654
rect 62566 87590 62630 87654
rect 64334 87590 64398 87654
rect 65966 87590 66030 87654
rect 67598 87590 67662 87654
rect 69366 87590 69430 87654
rect 70862 87590 70926 87654
rect 72630 87590 72694 87654
rect 74262 87590 74326 87654
rect 76030 87590 76094 87654
rect 77662 87590 77726 87654
rect 76302 87318 76366 87382
rect 79430 87590 79494 87654
rect 81062 87590 81126 87654
rect 82558 87590 82622 87654
rect 84326 87590 84390 87654
rect 86094 87590 86158 87654
rect 87862 87590 87926 87654
rect 73990 86910 74054 86974
rect 74262 86774 74326 86838
rect 74534 86288 74598 86294
rect 74534 86232 74558 86288
rect 74558 86232 74598 86288
rect 74534 86230 74598 86232
rect 75622 86288 75686 86294
rect 75622 86232 75670 86288
rect 75670 86232 75686 86288
rect 75622 86230 75686 86232
rect 76710 86230 76774 86294
rect 1230 85958 1294 86022
rect 89766 85958 89830 86022
rect 76302 85414 76366 85478
rect 74126 85278 74190 85342
rect 74262 84734 74326 84798
rect 74398 84598 74462 84662
rect 1230 84326 1294 84390
rect 89766 84326 89830 84390
rect 74126 83238 74190 83302
rect 74262 83102 74326 83166
rect 1230 82694 1294 82758
rect 89766 82694 89830 82758
rect 74398 81878 74462 81942
rect 74126 81742 74190 81806
rect 1230 80926 1294 80990
rect 89766 80926 89830 80990
rect 74262 80382 74326 80446
rect 74262 80246 74326 80310
rect 79294 80110 79358 80174
rect 90446 80110 90510 80174
rect 87998 79430 88062 79494
rect 1230 79294 1294 79358
rect 89086 79294 89150 79358
rect 89766 79294 89830 79358
rect 87998 79158 88062 79222
rect 74126 79022 74190 79086
rect 74126 78886 74190 78950
rect 79566 78614 79630 78678
rect 89086 78750 89150 78814
rect 25574 77934 25638 77998
rect 25982 77798 26046 77862
rect 30606 77934 30670 77998
rect 30878 77798 30942 77862
rect 35638 77934 35702 77998
rect 35910 77798 35974 77862
rect 40670 77934 40734 77998
rect 45566 77934 45630 77998
rect 41078 77798 41142 77862
rect 45974 77798 46038 77862
rect 50462 77934 50526 77998
rect 50870 77798 50934 77862
rect 55630 77934 55694 77998
rect 60662 77934 60726 77998
rect 56038 77798 56102 77862
rect 60934 77798 60998 77862
rect 1230 77662 1294 77726
rect 25846 77526 25910 77590
rect 30742 77526 30806 77590
rect 35774 77526 35838 77590
rect 40942 77526 41006 77590
rect 45838 77526 45902 77590
rect 50734 77526 50798 77590
rect 55902 77526 55966 77590
rect 60934 77526 60998 77590
rect 74262 77662 74326 77726
rect 72902 77526 72966 77590
rect 89766 77526 89830 77590
rect 79294 77390 79358 77454
rect 79294 77254 79358 77318
rect 79430 77254 79494 77318
rect 25846 76846 25910 76910
rect 30742 76846 30806 76910
rect 25846 76574 25910 76638
rect 30334 76574 30398 76638
rect 35774 76846 35838 76910
rect 40942 76846 41006 76910
rect 36862 76574 36926 76638
rect 40806 76574 40870 76638
rect 45838 76846 45902 76910
rect 45702 76574 45766 76638
rect 50734 76846 50798 76910
rect 55902 76846 55966 76910
rect 50734 76574 50798 76638
rect 55358 76574 55422 76638
rect 60934 76846 60998 76910
rect 61478 76574 61542 76638
rect 74126 76166 74190 76230
rect 79294 76166 79358 76230
rect 25982 76030 26046 76094
rect 26118 76030 26182 76094
rect 30878 76030 30942 76094
rect 31014 76030 31078 76094
rect 35910 76030 35974 76094
rect 36046 76030 36110 76094
rect 40942 76030 41006 76094
rect 41078 76030 41142 76094
rect 45974 76030 46038 76094
rect 46110 76030 46174 76094
rect 50870 76030 50934 76094
rect 51006 76030 51070 76094
rect 56038 76030 56102 76094
rect 56174 76030 56238 76094
rect 60798 76030 60862 76094
rect 60934 76030 60998 76094
rect 72630 76030 72694 76094
rect 79566 76030 79630 76094
rect 1230 75894 1294 75958
rect 89766 75894 89830 75958
rect 79294 75758 79358 75822
rect 79566 75758 79630 75822
rect 72902 74806 72966 74870
rect 79294 74806 79358 74870
rect 72766 74670 72830 74734
rect 79430 74534 79494 74598
rect 79294 74398 79358 74462
rect 89766 74398 89830 74462
rect 1230 74262 1294 74326
rect 26118 73582 26182 73646
rect 25982 73310 26046 73374
rect 31014 73582 31078 73646
rect 36046 73582 36110 73646
rect 41078 73582 41142 73646
rect 46110 73582 46174 73646
rect 51006 73582 51070 73646
rect 56174 73582 56238 73646
rect 60934 73582 60998 73646
rect 72630 73446 72694 73510
rect 66782 73310 66846 73374
rect 74126 73174 74190 73238
rect 79566 73174 79630 73238
rect 90446 73174 90510 73238
rect 1230 72630 1294 72694
rect 88465 72661 88529 72725
rect 89086 72494 89150 72558
rect 89766 72494 89830 72558
rect 25846 71950 25910 72014
rect 25574 71814 25638 71878
rect 26798 71814 26862 71878
rect 27614 71814 27678 71878
rect 27750 71814 27814 71878
rect 28974 71814 29038 71878
rect 29518 71814 29582 71878
rect 30334 71950 30398 72014
rect 30742 71814 30806 71878
rect 31422 71814 31486 71878
rect 31966 71814 32030 71878
rect 32510 71814 32574 71878
rect 33054 71814 33118 71878
rect 34006 71814 34070 71878
rect 34414 71814 34478 71878
rect 35230 71814 35294 71878
rect 35774 71814 35838 71878
rect 36862 71950 36926 72014
rect 36454 71814 36518 71878
rect 36998 71814 37062 71878
rect 37678 71814 37742 71878
rect 38222 71814 38286 71878
rect 39446 71814 39510 71878
rect 40806 71950 40870 72014
rect 40262 71814 40326 71878
rect 40670 71814 40734 71878
rect 41622 71814 41686 71878
rect 42710 71814 42774 71878
rect 43254 71814 43318 71878
rect 43934 71814 43998 71878
rect 45702 71950 45766 72014
rect 45158 71814 45222 71878
rect 45702 71814 45766 71878
rect 46926 71814 46990 71878
rect 47742 71814 47806 71878
rect 48966 71814 49030 71878
rect 49374 71814 49438 71878
rect 50734 71950 50798 72014
rect 50190 71814 50254 71878
rect 51414 71814 51478 71878
rect 51958 71814 52022 71878
rect 52638 71814 52702 71878
rect 54134 71814 54198 71878
rect 55358 71950 55422 72014
rect 55766 71814 55830 71878
rect 56446 71814 56510 71878
rect 56990 71814 57054 71878
rect 57670 71814 57734 71878
rect 58214 71814 58278 71878
rect 58894 71814 58958 71878
rect 60662 71814 60726 71878
rect 61478 71950 61542 72014
rect 61478 71814 61542 71878
rect 62022 71814 62086 71878
rect 62702 71814 62766 71878
rect 63110 71814 63174 71878
rect 63926 71814 63990 71878
rect 64470 71814 64534 71878
rect 65150 71814 65214 71878
rect 65694 71814 65758 71878
rect 79294 71678 79358 71742
rect 89086 71678 89150 71742
rect 25574 71406 25638 71470
rect 26798 71406 26862 71470
rect 27614 71406 27678 71470
rect 27750 71406 27814 71470
rect 28974 71406 29038 71470
rect 29518 71406 29582 71470
rect 30742 71406 30806 71470
rect 31422 71406 31486 71470
rect 31966 71406 32030 71470
rect 32510 71406 32574 71470
rect 33054 71406 33118 71470
rect 34006 71406 34070 71470
rect 34414 71406 34478 71470
rect 35230 71406 35294 71470
rect 35774 71406 35838 71470
rect 36454 71406 36518 71470
rect 36998 71406 37062 71470
rect 37678 71406 37742 71470
rect 38222 71406 38286 71470
rect 39446 71406 39510 71470
rect 40262 71406 40326 71470
rect 40670 71406 40734 71470
rect 42710 71406 42774 71470
rect 41622 71270 41686 71334
rect 43254 71406 43318 71470
rect 43934 71406 43998 71470
rect 45158 71406 45222 71470
rect 45702 71406 45766 71470
rect 46926 71406 46990 71470
rect 47742 71406 47806 71470
rect 48966 71406 49030 71470
rect 49374 71406 49438 71470
rect 50190 71406 50254 71470
rect 51414 71406 51478 71470
rect 51958 71406 52022 71470
rect 52638 71406 52702 71470
rect 54134 71270 54198 71334
rect 55766 71406 55830 71470
rect 56446 71406 56510 71470
rect 56990 71406 57054 71470
rect 57670 71406 57734 71470
rect 58214 71406 58278 71470
rect 58894 71406 58958 71470
rect 60662 71406 60726 71470
rect 61478 71406 61542 71470
rect 62022 71406 62086 71470
rect 62702 71406 62766 71470
rect 63110 71406 63174 71470
rect 63926 71406 63990 71470
rect 64470 71406 64534 71470
rect 65150 71406 65214 71470
rect 65694 71406 65758 71470
rect 67734 71270 67798 71334
rect 66782 71134 66846 71198
rect 1230 70998 1294 71062
rect 67734 70998 67798 71062
rect 25982 70862 26046 70926
rect 72766 70998 72830 71062
rect 71134 70862 71198 70926
rect 71406 70862 71470 70926
rect 89766 70862 89830 70926
rect 17958 70318 18022 70382
rect 18230 70318 18294 70382
rect 18910 70318 18974 70382
rect 19046 70318 19110 70382
rect 66510 70454 66574 70518
rect 71134 70454 71198 70518
rect 71406 70454 71470 70518
rect 19590 70318 19654 70382
rect 17958 70046 18022 70110
rect 17958 69910 18022 69974
rect 18230 70046 18294 70110
rect 18230 69910 18294 69974
rect 18910 70046 18974 70110
rect 19046 70046 19110 70110
rect 19182 69910 19246 69974
rect 19590 70046 19654 70110
rect 19590 69910 19654 69974
rect 71270 70318 71334 70382
rect 71678 70318 71742 70382
rect 72222 70318 72286 70382
rect 72358 70318 72422 70382
rect 74126 70454 74190 70518
rect 73038 70318 73102 70382
rect 90446 70182 90510 70246
rect 66510 70046 66574 70110
rect 71270 70046 71334 70110
rect 71406 69910 71470 69974
rect 71678 70046 71742 70110
rect 71814 69910 71878 69974
rect 72222 70046 72286 70110
rect 72358 70046 72422 70110
rect 72630 69910 72694 69974
rect 73038 70046 73102 70110
rect 72902 69910 72966 69974
rect 17958 69638 18022 69702
rect 17822 69502 17886 69566
rect 18230 69638 18294 69702
rect 18230 69502 18294 69566
rect 19182 69638 19246 69702
rect 19182 69502 19246 69566
rect 19590 69638 19654 69702
rect 19454 69502 19518 69566
rect 71406 69638 71470 69702
rect 1230 69230 1294 69294
rect 17822 69230 17886 69294
rect 17822 69094 17886 69158
rect 18230 69230 18294 69294
rect 18230 69094 18294 69158
rect 18502 69094 18566 69158
rect 19182 69230 19246 69294
rect 19046 69094 19110 69158
rect 19454 69230 19518 69294
rect 19590 69094 19654 69158
rect 71406 69502 71470 69566
rect 71814 69638 71878 69702
rect 71678 69502 71742 69566
rect 72222 69502 72286 69566
rect 72630 69638 72694 69702
rect 72902 69638 72966 69702
rect 72902 69502 72966 69566
rect 89766 69366 89830 69430
rect 71406 69230 71470 69294
rect 71270 69094 71334 69158
rect 71678 69230 71742 69294
rect 71678 69094 71742 69158
rect 72222 69230 72286 69294
rect 72358 69094 72422 69158
rect 72902 69230 72966 69294
rect 89086 69230 89150 69294
rect 73038 69094 73102 69158
rect 17822 68822 17886 68886
rect 18230 68822 18294 68886
rect 18502 68822 18566 68886
rect 18366 68686 18430 68750
rect 18502 68686 18566 68750
rect 19046 68822 19110 68886
rect 19182 68686 19246 68750
rect 19590 68822 19654 68886
rect 19454 68686 19518 68750
rect 71270 68822 71334 68886
rect 71406 68686 71470 68750
rect 71678 68822 71742 68886
rect 71814 68686 71878 68750
rect 72358 68822 72422 68886
rect 72086 68686 72150 68750
rect 72494 68686 72558 68750
rect 73038 68822 73102 68886
rect 89086 68958 89150 69022
rect 66374 68550 66438 68614
rect 18366 68414 18430 68478
rect 18502 68414 18566 68478
rect 19182 68414 19246 68478
rect 19046 68278 19110 68342
rect 19454 68414 19518 68478
rect 19590 68278 19654 68342
rect 18502 67870 18566 67934
rect 19046 68006 19110 68070
rect 19046 67870 19110 67934
rect 19590 68006 19654 68070
rect 19454 67870 19518 67934
rect 66374 68278 66438 68342
rect 66510 68278 66574 68342
rect 71406 68414 71470 68478
rect 71270 68278 71334 68342
rect 71814 68414 71878 68478
rect 71814 68278 71878 68342
rect 72086 68414 72150 68478
rect 72494 68414 72558 68478
rect 71270 68006 71334 68070
rect 1230 67734 1294 67798
rect 66510 67870 66574 67934
rect 71270 67870 71334 67934
rect 71814 68006 71878 68070
rect 71678 67870 71742 67934
rect 72358 67870 72422 67934
rect 17822 67598 17886 67662
rect 18502 67598 18566 67662
rect 17822 67326 17886 67390
rect 17822 67190 17886 67254
rect 18502 67190 18566 67254
rect 19046 67598 19110 67662
rect 19454 67598 19518 67662
rect 24350 67326 24414 67390
rect 71270 67598 71334 67662
rect 66510 67326 66574 67390
rect 24350 67054 24414 67118
rect 17822 66918 17886 66982
rect 17822 66782 17886 66846
rect 18502 66918 18566 66982
rect 17822 66510 17886 66574
rect 17958 66374 18022 66438
rect 18910 66374 18974 66438
rect 19182 66374 19246 66438
rect 24622 66918 24686 66982
rect 24622 66646 24686 66710
rect 66510 67054 66574 67118
rect 66510 66918 66574 66982
rect 66510 66646 66574 66710
rect 71678 67598 71742 67662
rect 72358 67598 72422 67662
rect 72902 67598 72966 67662
rect 89766 67734 89830 67798
rect 72086 67190 72150 67254
rect 72630 67190 72694 67254
rect 72902 67326 72966 67390
rect 87726 67326 87790 67390
rect 72902 67190 72966 67254
rect 72086 66918 72150 66982
rect 72630 66918 72694 66982
rect 72086 66646 72150 66710
rect 19454 66374 19518 66438
rect 17958 66102 18022 66166
rect 17822 65966 17886 66030
rect 18230 65966 18294 66030
rect 18910 66102 18974 66166
rect 18774 65966 18838 66030
rect 19182 66102 19246 66166
rect 19046 65966 19110 66030
rect 19454 66102 19518 66166
rect 19454 65966 19518 66030
rect 24622 66102 24686 66166
rect 71406 66374 71470 66438
rect 71814 66374 71878 66438
rect 72902 66918 72966 66982
rect 72902 66782 72966 66846
rect 72902 66510 72966 66574
rect 72902 66374 72966 66438
rect 72086 66238 72150 66302
rect 66510 66102 66574 66166
rect 71406 66102 71470 66166
rect 71270 65966 71334 66030
rect 71814 66102 71878 66166
rect 71678 65966 71742 66030
rect 72222 65966 72286 66030
rect 72358 65966 72422 66030
rect 72902 66102 72966 66166
rect 73038 65966 73102 66030
rect 1230 65830 1294 65894
rect 24622 65830 24686 65894
rect 17822 65694 17886 65758
rect 17822 65558 17886 65622
rect 18230 65694 18294 65758
rect 18774 65694 18838 65758
rect 18230 65558 18294 65622
rect 18502 65558 18566 65622
rect 19046 65694 19110 65758
rect 19046 65558 19110 65622
rect 19454 65694 19518 65758
rect 19454 65558 19518 65622
rect 66510 65830 66574 65894
rect 89766 65830 89830 65894
rect 17822 65286 17886 65350
rect 17822 65150 17886 65214
rect 18230 65286 18294 65350
rect 18502 65286 18566 65350
rect 18638 65150 18702 65214
rect 19046 65286 19110 65350
rect 19182 65150 19246 65214
rect 19454 65286 19518 65350
rect 19454 65150 19518 65214
rect 17822 64878 17886 64942
rect 18230 64742 18294 64806
rect 18638 64878 18702 64942
rect 18910 64742 18974 64806
rect 19182 64878 19246 64942
rect 19046 64742 19110 64806
rect 19454 64878 19518 64942
rect 71270 65694 71334 65758
rect 71406 65558 71470 65622
rect 71678 65694 71742 65758
rect 71678 65558 71742 65622
rect 72222 65694 72286 65758
rect 72358 65694 72422 65758
rect 72086 65558 72150 65622
rect 72494 65558 72558 65622
rect 73038 65694 73102 65758
rect 72902 65558 72966 65622
rect 71406 65286 71470 65350
rect 71406 65150 71470 65214
rect 71678 65286 71742 65350
rect 71814 65150 71878 65214
rect 72086 65286 72150 65350
rect 72494 65286 72558 65350
rect 72358 65150 72422 65214
rect 72902 65286 72966 65350
rect 73038 65150 73102 65214
rect 19590 64742 19654 64806
rect 71406 64878 71470 64942
rect 71270 64742 71334 64806
rect 71814 64878 71878 64942
rect 71678 64742 71742 64806
rect 72358 64878 72422 64942
rect 72222 64742 72286 64806
rect 72630 64742 72694 64806
rect 73038 64878 73102 64942
rect 17958 64334 18022 64398
rect 18230 64470 18294 64534
rect 18366 64334 18430 64398
rect 18910 64470 18974 64534
rect 19046 64470 19110 64534
rect 19182 64334 19246 64398
rect 19590 64470 19654 64534
rect 19590 64334 19654 64398
rect 1230 64198 1294 64262
rect 17958 64062 18022 64126
rect 18366 64062 18430 64126
rect 18910 63926 18974 63990
rect 19182 64062 19246 64126
rect 19182 63926 19246 63990
rect 19590 64062 19654 64126
rect 71270 64470 71334 64534
rect 71406 64334 71470 64398
rect 71678 64470 71742 64534
rect 71678 64334 71742 64398
rect 72222 64470 72286 64534
rect 72630 64470 72694 64534
rect 72494 64334 72558 64398
rect 87726 64606 87790 64670
rect 87590 64470 87654 64534
rect 90446 64470 90510 64534
rect 72902 64334 72966 64398
rect 89766 64198 89830 64262
rect 71406 64062 71470 64126
rect 19590 63926 19654 63990
rect 24486 63790 24550 63854
rect 71270 63926 71334 63990
rect 71678 64062 71742 64126
rect 71678 63926 71742 63990
rect 72494 64062 72558 64126
rect 72086 63926 72150 63990
rect 72358 63926 72422 63990
rect 72902 64062 72966 64126
rect 66510 63790 66574 63854
rect 17822 63654 17886 63718
rect 18910 63654 18974 63718
rect 19182 63654 19246 63718
rect 19590 63654 19654 63718
rect 17822 63382 17886 63446
rect 17958 63246 18022 63310
rect 18502 63246 18566 63310
rect 17958 62974 18022 63038
rect 17958 62838 18022 62902
rect 18502 62974 18566 63038
rect 1230 62430 1294 62494
rect 17958 62566 18022 62630
rect 17822 62430 17886 62494
rect 18366 62430 18430 62494
rect 24486 63518 24550 63582
rect 24622 63382 24686 63446
rect 66510 63518 66574 63582
rect 66374 63382 66438 63446
rect 71270 63654 71334 63718
rect 71678 63654 71742 63718
rect 72086 63654 72150 63718
rect 72358 63654 72422 63718
rect 73038 63654 73102 63718
rect 24622 63110 24686 63174
rect 24350 62974 24414 63038
rect 24350 62702 24414 62766
rect 19046 62430 19110 62494
rect 19590 62430 19654 62494
rect 17822 62158 17886 62222
rect 17822 62022 17886 62086
rect 18366 62158 18430 62222
rect 18910 62022 18974 62086
rect 19046 62158 19110 62222
rect 19182 62022 19246 62086
rect 19590 62158 19654 62222
rect 19454 62022 19518 62086
rect 66374 63110 66438 63174
rect 66374 62974 66438 63038
rect 66374 62702 66438 62766
rect 66510 62702 66574 62766
rect 72086 63246 72150 63310
rect 73038 63382 73102 63446
rect 72902 63246 72966 63310
rect 89086 63110 89150 63174
rect 72086 62974 72150 63038
rect 72902 62974 72966 63038
rect 72902 62838 72966 62902
rect 66510 62430 66574 62494
rect 71406 62430 71470 62494
rect 71678 62430 71742 62494
rect 72494 62430 72558 62494
rect 72902 62566 72966 62630
rect 72902 62430 72966 62494
rect 89086 62566 89150 62630
rect 89766 62566 89830 62630
rect 88465 62486 88529 62490
rect 88465 62430 88469 62486
rect 88469 62430 88525 62486
rect 88525 62430 88529 62486
rect 88465 62426 88529 62430
rect 71406 62158 71470 62222
rect 71406 62022 71470 62086
rect 71678 62158 71742 62222
rect 71678 62022 71742 62086
rect 72494 62158 72558 62222
rect 72086 62022 72150 62086
rect 72358 62022 72422 62086
rect 72902 62158 72966 62222
rect 72902 62022 72966 62086
rect 17822 61750 17886 61814
rect 17822 61614 17886 61678
rect 18230 61614 18294 61678
rect 18910 61750 18974 61814
rect 18774 61614 18838 61678
rect 19182 61750 19246 61814
rect 19046 61614 19110 61678
rect 19454 61750 19518 61814
rect 87726 61886 87790 61950
rect 19454 61614 19518 61678
rect 71406 61750 71470 61814
rect 71270 61614 71334 61678
rect 71678 61750 71742 61814
rect 71814 61614 71878 61678
rect 72086 61750 72150 61814
rect 72358 61750 72422 61814
rect 72222 61614 72286 61678
rect 72358 61614 72422 61678
rect 72902 61750 72966 61814
rect 73038 61614 73102 61678
rect 17822 61342 17886 61406
rect 17958 61206 18022 61270
rect 18230 61342 18294 61406
rect 18366 61206 18430 61270
rect 18774 61342 18838 61406
rect 18774 61206 18838 61270
rect 19046 61342 19110 61406
rect 19046 61206 19110 61270
rect 19454 61342 19518 61406
rect 19590 61206 19654 61270
rect 71270 61342 71334 61406
rect 71406 61206 71470 61270
rect 71814 61342 71878 61406
rect 71814 61206 71878 61270
rect 72222 61342 72286 61406
rect 72358 61342 72422 61406
rect 72086 61206 72150 61270
rect 72630 61206 72694 61270
rect 73038 61342 73102 61406
rect 73038 61206 73102 61270
rect 1230 60798 1294 60862
rect 17958 60934 18022 60998
rect 18366 60934 18430 60998
rect 18774 60934 18838 60998
rect 18638 60798 18702 60862
rect 19046 60934 19110 60998
rect 19046 60798 19110 60862
rect 19590 60934 19654 60998
rect 19454 60798 19518 60862
rect 71406 60934 71470 60998
rect 17958 60390 18022 60454
rect 18230 60390 18294 60454
rect 18638 60526 18702 60590
rect 18910 60390 18974 60454
rect 19046 60526 19110 60590
rect 19046 60390 19110 60454
rect 19454 60526 19518 60590
rect 19454 60390 19518 60454
rect 71270 60798 71334 60862
rect 71814 60934 71878 60998
rect 71678 60798 71742 60862
rect 72086 60934 72150 60998
rect 72630 60934 72694 60998
rect 73038 60934 73102 60998
rect 89766 60934 89830 60998
rect 71270 60526 71334 60590
rect 71270 60390 71334 60454
rect 71678 60526 71742 60590
rect 71678 60390 71742 60454
rect 72222 60390 72286 60454
rect 72630 60390 72694 60454
rect 73038 60390 73102 60454
rect 17958 60118 18022 60182
rect 18230 60118 18294 60182
rect 18910 60118 18974 60182
rect 18366 59982 18430 60046
rect 18502 59982 18566 60046
rect 18774 59982 18838 60046
rect 19046 60118 19110 60182
rect 19182 59982 19246 60046
rect 19454 60118 19518 60182
rect 19454 59982 19518 60046
rect 24622 59846 24686 59910
rect 17822 59710 17886 59774
rect 18366 59710 18430 59774
rect 18502 59710 18566 59774
rect 18774 59710 18838 59774
rect 19182 59710 19246 59774
rect 19182 59574 19246 59638
rect 19454 59710 19518 59774
rect 19590 59574 19654 59638
rect 24622 59574 24686 59638
rect 17822 59438 17886 59502
rect 1230 59166 1294 59230
rect 18910 59166 18974 59230
rect 19182 59302 19246 59366
rect 19590 59302 19654 59366
rect 71270 60118 71334 60182
rect 71406 59982 71470 60046
rect 71678 60118 71742 60182
rect 71678 59982 71742 60046
rect 72222 60118 72286 60182
rect 72086 59982 72150 60046
rect 72630 60118 72694 60182
rect 73038 60118 73102 60182
rect 66374 59846 66438 59910
rect 66374 59574 66438 59638
rect 66510 59574 66574 59638
rect 71406 59710 71470 59774
rect 71270 59574 71334 59638
rect 71678 59710 71742 59774
rect 71814 59574 71878 59638
rect 72086 59710 72150 59774
rect 72902 59710 72966 59774
rect 71270 59302 71334 59366
rect 17822 58894 17886 58958
rect 18910 58894 18974 58958
rect 18502 58758 18566 58822
rect 17822 58622 17886 58686
rect 17822 58486 17886 58550
rect 18502 58486 18566 58550
rect 18774 58486 18838 58550
rect 24350 58622 24414 58686
rect 66510 59166 66574 59230
rect 66374 59030 66438 59094
rect 66374 58758 66438 58822
rect 66510 58622 66574 58686
rect 71814 59302 71878 59366
rect 72358 59166 72422 59230
rect 72902 59438 72966 59502
rect 89766 59166 89830 59230
rect 72358 58894 72422 58958
rect 72902 58894 72966 58958
rect 24350 58350 24414 58414
rect 17822 58214 17886 58278
rect 17822 58078 17886 58142
rect 18774 58214 18838 58278
rect 19046 58078 19110 58142
rect 19454 58078 19518 58142
rect 66510 58350 66574 58414
rect 72086 58486 72150 58550
rect 72358 58486 72422 58550
rect 72902 58622 72966 58686
rect 73038 58486 73102 58550
rect 71270 58078 71334 58142
rect 71814 58078 71878 58142
rect 72086 58214 72150 58278
rect 72358 58214 72422 58278
rect 17822 57806 17886 57870
rect 17822 57670 17886 57734
rect 18638 57670 18702 57734
rect 19046 57806 19110 57870
rect 19182 57670 19246 57734
rect 19454 57806 19518 57870
rect 71270 57806 71334 57870
rect 19454 57670 19518 57734
rect 1230 57398 1294 57462
rect 17822 57398 17886 57462
rect 17822 57262 17886 57326
rect 18638 57398 18702 57462
rect 18230 57262 18294 57326
rect 19182 57398 19246 57462
rect 19046 57262 19110 57326
rect 19454 57398 19518 57462
rect 19590 57262 19654 57326
rect 71406 57670 71470 57734
rect 71814 57806 71878 57870
rect 71814 57670 71878 57734
rect 73038 58214 73102 58278
rect 72902 58078 72966 58142
rect 72358 57670 72422 57734
rect 72902 57806 72966 57870
rect 72902 57670 72966 57734
rect 71406 57398 71470 57462
rect 71270 57262 71334 57326
rect 71814 57398 71878 57462
rect 72358 57398 72422 57462
rect 71814 57262 71878 57326
rect 72222 57262 72286 57326
rect 72902 57398 72966 57462
rect 89766 57398 89830 57462
rect 73038 57262 73102 57326
rect 17822 56990 17886 57054
rect 17958 56854 18022 56918
rect 18230 56990 18294 57054
rect 18366 56854 18430 56918
rect 18502 56854 18566 56918
rect 19046 56990 19110 57054
rect 19182 56854 19246 56918
rect 19590 56990 19654 57054
rect 19590 56854 19654 56918
rect 17958 56582 18022 56646
rect 17822 56446 17886 56510
rect 18366 56582 18430 56646
rect 18502 56582 18566 56646
rect 18366 56446 18430 56510
rect 18502 56446 18566 56510
rect 19182 56582 19246 56646
rect 19182 56446 19246 56510
rect 19590 56582 19654 56646
rect 19590 56446 19654 56510
rect 71270 56990 71334 57054
rect 71270 56854 71334 56918
rect 71814 56990 71878 57054
rect 71678 56854 71742 56918
rect 72222 56990 72286 57054
rect 72086 56854 72150 56918
rect 72494 56854 72558 56918
rect 73038 56990 73102 57054
rect 72902 56854 72966 56918
rect 71270 56582 71334 56646
rect 71406 56446 71470 56510
rect 71678 56582 71742 56646
rect 71678 56446 71742 56510
rect 72086 56582 72150 56646
rect 72494 56582 72558 56646
rect 72358 56446 72422 56510
rect 72902 56582 72966 56646
rect 72902 56446 72966 56510
rect 17822 56174 17886 56238
rect 18366 56174 18430 56238
rect 18502 56174 18566 56238
rect 18910 56038 18974 56102
rect 19182 56174 19246 56238
rect 19046 56038 19110 56102
rect 19590 56174 19654 56238
rect 19590 56038 19654 56102
rect 1230 55766 1294 55830
rect 71406 56174 71470 56238
rect 71270 56038 71334 56102
rect 71678 56174 71742 56238
rect 71678 56038 71742 56102
rect 72358 56174 72422 56238
rect 72630 56038 72694 56102
rect 72902 56174 72966 56238
rect 18910 55766 18974 55830
rect 19046 55766 19110 55830
rect 19182 55630 19246 55694
rect 19590 55766 19654 55830
rect 19590 55630 19654 55694
rect 18638 55222 18702 55286
rect 19182 55358 19246 55422
rect 19590 55358 19654 55422
rect 71270 55766 71334 55830
rect 71406 55630 71470 55694
rect 71678 55766 71742 55830
rect 71814 55630 71878 55694
rect 72630 55766 72694 55830
rect 89766 55766 89830 55830
rect 71406 55358 71470 55422
rect 17958 54950 18022 55014
rect 18638 54950 18702 55014
rect 17958 54678 18022 54742
rect 17822 54542 17886 54606
rect 18366 54542 18430 54606
rect 18502 54542 18566 54606
rect 24622 54678 24686 54742
rect 71814 55358 71878 55422
rect 72222 55222 72286 55286
rect 72358 55222 72422 55286
rect 66510 55086 66574 55150
rect 66510 54814 66574 54878
rect 66510 54678 66574 54742
rect 72222 54950 72286 55014
rect 72358 54950 72422 55014
rect 73038 54950 73102 55014
rect 1230 54134 1294 54198
rect 17822 54270 17886 54334
rect 17958 54134 18022 54198
rect 18366 54270 18430 54334
rect 18502 54270 18566 54334
rect 17958 53862 18022 53926
rect 17822 53726 17886 53790
rect 19182 54134 19246 54198
rect 19454 54134 19518 54198
rect 24622 54406 24686 54470
rect 24350 54270 24414 54334
rect 66510 54406 66574 54470
rect 72358 54542 72422 54606
rect 73038 54678 73102 54742
rect 72902 54542 72966 54606
rect 71406 54134 71470 54198
rect 71814 54134 71878 54198
rect 72358 54270 72422 54334
rect 24350 53998 24414 54062
rect 19182 53862 19246 53926
rect 19182 53726 19246 53790
rect 19454 53862 19518 53926
rect 19454 53726 19518 53790
rect 17822 53454 17886 53518
rect 17822 53318 17886 53382
rect 18502 53318 18566 53382
rect 19182 53454 19246 53518
rect 19182 53318 19246 53382
rect 19454 53454 19518 53518
rect 19454 53318 19518 53382
rect 72902 54270 72966 54334
rect 73038 54134 73102 54198
rect 89766 54134 89830 54198
rect 71406 53862 71470 53926
rect 71406 53726 71470 53790
rect 71814 53862 71878 53926
rect 71678 53726 71742 53790
rect 72086 53726 72150 53790
rect 73038 53862 73102 53926
rect 73038 53726 73102 53790
rect 71406 53454 71470 53518
rect 71406 53318 71470 53382
rect 71678 53454 71742 53518
rect 71678 53318 71742 53382
rect 72086 53454 72150 53518
rect 72086 53318 72150 53382
rect 72358 53318 72422 53382
rect 73038 53454 73102 53518
rect 72902 53318 72966 53382
rect 17822 53046 17886 53110
rect 17822 52910 17886 52974
rect 18502 53046 18566 53110
rect 18230 52910 18294 52974
rect 18910 52910 18974 52974
rect 19182 53046 19246 53110
rect 19046 52910 19110 52974
rect 19454 53046 19518 53110
rect 19454 52910 19518 52974
rect 71406 53046 71470 53110
rect 71270 52910 71334 52974
rect 71678 53046 71742 53110
rect 71678 52910 71742 52974
rect 72086 53046 72150 53110
rect 72358 53046 72422 53110
rect 72222 52910 72286 52974
rect 72902 53046 72966 53110
rect 73038 52910 73102 52974
rect 17822 52638 17886 52702
rect 1230 52502 1294 52566
rect 17822 52502 17886 52566
rect 18230 52638 18294 52702
rect 18910 52638 18974 52702
rect 18366 52502 18430 52566
rect 18502 52502 18566 52566
rect 19046 52638 19110 52702
rect 19046 52502 19110 52566
rect 19454 52638 19518 52702
rect 19590 52502 19654 52566
rect 71270 52638 71334 52702
rect 71270 52502 71334 52566
rect 71678 52638 71742 52702
rect 71678 52502 71742 52566
rect 72222 52638 72286 52702
rect 72086 52502 72150 52566
rect 72630 52502 72694 52566
rect 73038 52638 73102 52702
rect 72902 52502 72966 52566
rect 17822 52230 17886 52294
rect 18366 52230 18430 52294
rect 18502 52230 18566 52294
rect 18910 52094 18974 52158
rect 19046 52230 19110 52294
rect 19182 52094 19246 52158
rect 19590 52230 19654 52294
rect 19454 52094 19518 52158
rect 89766 52366 89830 52430
rect 71270 52230 71334 52294
rect 18910 51822 18974 51886
rect 19182 51822 19246 51886
rect 19046 51686 19110 51750
rect 19454 51822 19518 51886
rect 19590 51686 19654 51750
rect 18502 51278 18566 51342
rect 19046 51414 19110 51478
rect 19182 51278 19246 51342
rect 19590 51414 19654 51478
rect 71270 52094 71334 52158
rect 71678 52230 71742 52294
rect 71678 52094 71742 52158
rect 72086 52230 72150 52294
rect 72630 52230 72694 52294
rect 72358 52094 72422 52158
rect 72902 52230 72966 52294
rect 71270 51822 71334 51886
rect 71270 51686 71334 51750
rect 71678 51822 71742 51886
rect 71678 51686 71742 51750
rect 72358 51822 72422 51886
rect 72494 51686 72558 51750
rect 19454 51278 19518 51342
rect 18910 51142 18974 51206
rect 24622 51142 24686 51206
rect 17822 51006 17886 51070
rect 18502 51006 18566 51070
rect 1230 50734 1294 50798
rect 19182 51006 19246 51070
rect 17822 50734 17886 50798
rect 17958 50598 18022 50662
rect 18910 50734 18974 50798
rect 18638 50598 18702 50662
rect 19454 51006 19518 51070
rect 24486 50870 24550 50934
rect 24622 50870 24686 50934
rect 71270 51414 71334 51478
rect 71406 51278 71470 51342
rect 71678 51414 71742 51478
rect 71678 51278 71742 51342
rect 72358 51414 72422 51478
rect 72494 51278 72558 51342
rect 66374 51142 66438 51206
rect 66374 50870 66438 50934
rect 71406 51006 71470 51070
rect 66374 50734 66438 50798
rect 66510 50734 66574 50798
rect 17958 50326 18022 50390
rect 17958 50190 18022 50254
rect 18638 50326 18702 50390
rect 24486 50462 24550 50526
rect 66374 50462 66438 50526
rect 71678 51006 71742 51070
rect 72494 51006 72558 51070
rect 72902 51006 72966 51070
rect 72358 50598 72422 50662
rect 72902 50734 72966 50798
rect 89766 50734 89830 50798
rect 73038 50598 73102 50662
rect 66510 50326 66574 50390
rect 17958 49918 18022 49982
rect 17958 49782 18022 49846
rect 18230 49782 18294 49846
rect 18774 49782 18838 49846
rect 19182 49782 19246 49846
rect 19590 49782 19654 49846
rect 17958 49510 18022 49574
rect 17822 49374 17886 49438
rect 18230 49510 18294 49574
rect 18774 49510 18838 49574
rect 18774 49374 18838 49438
rect 19182 49510 19246 49574
rect 19182 49374 19246 49438
rect 19590 49510 19654 49574
rect 19454 49374 19518 49438
rect 71270 49782 71334 49846
rect 71678 49782 71742 49846
rect 72358 50326 72422 50390
rect 73038 50326 73102 50390
rect 72902 50190 72966 50254
rect 72086 49782 72150 49846
rect 72630 49782 72694 49846
rect 72902 49918 72966 49982
rect 73038 49782 73102 49846
rect 71270 49510 71334 49574
rect 71270 49374 71334 49438
rect 71678 49510 71742 49574
rect 71678 49374 71742 49438
rect 72086 49510 72150 49574
rect 72630 49510 72694 49574
rect 72630 49374 72694 49438
rect 73038 49510 73102 49574
rect 73038 49374 73102 49438
rect 1230 48966 1294 49030
rect 17822 49102 17886 49166
rect 17958 48966 18022 49030
rect 18774 49102 18838 49166
rect 18638 48966 18702 49030
rect 19182 49102 19246 49166
rect 19182 48966 19246 49030
rect 19454 49102 19518 49166
rect 71270 49102 71334 49166
rect 19454 48966 19518 49030
rect 17958 48694 18022 48758
rect 17822 48558 17886 48622
rect 18230 48558 18294 48622
rect 18638 48694 18702 48758
rect 18910 48558 18974 48622
rect 19182 48694 19246 48758
rect 19046 48558 19110 48622
rect 19454 48694 19518 48758
rect 19590 48558 19654 48622
rect 71406 48966 71470 49030
rect 71678 49102 71742 49166
rect 71814 48966 71878 49030
rect 72086 48966 72150 49030
rect 72630 49102 72694 49166
rect 72494 48966 72558 49030
rect 73038 49102 73102 49166
rect 72902 48966 72966 49030
rect 89766 49102 89830 49166
rect 71406 48694 71470 48758
rect 71270 48558 71334 48622
rect 71814 48694 71878 48758
rect 71678 48558 71742 48622
rect 72086 48694 72150 48758
rect 72494 48694 72558 48758
rect 72222 48558 72286 48622
rect 72902 48694 72966 48758
rect 73038 48558 73102 48622
rect 17822 48286 17886 48350
rect 18230 48286 18294 48350
rect 18230 48150 18294 48214
rect 18910 48286 18974 48350
rect 19046 48286 19110 48350
rect 19046 48150 19110 48214
rect 19590 48286 19654 48350
rect 19454 48150 19518 48214
rect 1230 47334 1294 47398
rect 18230 47878 18294 47942
rect 19046 47878 19110 47942
rect 19182 47742 19246 47806
rect 19454 47878 19518 47942
rect 19454 47742 19518 47806
rect 71270 48286 71334 48350
rect 71270 48150 71334 48214
rect 71678 48286 71742 48350
rect 71814 48150 71878 48214
rect 72222 48286 72286 48350
rect 72086 48150 72150 48214
rect 73038 48286 73102 48350
rect 71270 47878 71334 47942
rect 71270 47742 71334 47806
rect 71814 47878 71878 47942
rect 71814 47742 71878 47806
rect 72086 47878 72150 47942
rect 19182 47470 19246 47534
rect 18910 47334 18974 47398
rect 19046 47334 19110 47398
rect 19454 47470 19518 47534
rect 19590 47334 19654 47398
rect 71270 47470 71334 47534
rect 71270 47334 71334 47398
rect 71814 47470 71878 47534
rect 71814 47334 71878 47398
rect 72222 47334 72286 47398
rect 89766 47334 89830 47398
rect 17958 47062 18022 47126
rect 18910 47062 18974 47126
rect 18502 46926 18566 46990
rect 19046 47062 19110 47126
rect 19590 47062 19654 47126
rect 17958 46790 18022 46854
rect 17822 46654 17886 46718
rect 18502 46654 18566 46718
rect 18774 46654 18838 46718
rect 24486 46790 24550 46854
rect 71270 47062 71334 47126
rect 66374 46790 66438 46854
rect 24486 46518 24550 46582
rect 17822 46382 17886 46446
rect 17958 46246 18022 46310
rect 18774 46382 18838 46446
rect 17958 45974 18022 46038
rect 17958 45838 18022 45902
rect 18366 45838 18430 45902
rect 18502 45838 18566 45902
rect 22854 46110 22918 46174
rect 24486 46110 24550 46174
rect 19182 45838 19246 45902
rect 66374 46518 66438 46582
rect 66510 46382 66574 46446
rect 66510 46110 66574 46174
rect 71814 47062 71878 47126
rect 72222 47062 72286 47126
rect 72902 47062 72966 47126
rect 72494 46654 72558 46718
rect 72902 46790 72966 46854
rect 72902 46654 72966 46718
rect 69366 45974 69430 46038
rect 19454 45838 19518 45902
rect 24486 45838 24550 45902
rect 1230 45702 1294 45766
rect 17958 45566 18022 45630
rect 17958 45430 18022 45494
rect 18366 45566 18430 45630
rect 18502 45566 18566 45630
rect 19182 45566 19246 45630
rect 19454 45566 19518 45630
rect 19046 45430 19110 45494
rect 19454 45430 19518 45494
rect 22854 45566 22918 45630
rect 24350 45566 24414 45630
rect 71406 45838 71470 45902
rect 71678 45838 71742 45902
rect 72086 45838 72150 45902
rect 72494 46382 72558 46446
rect 72902 46382 72966 46446
rect 73038 46246 73102 46310
rect 72494 45838 72558 45902
rect 73038 45974 73102 46038
rect 72902 45838 72966 45902
rect 89766 45702 89830 45766
rect 69366 45566 69430 45630
rect 71406 45566 71470 45630
rect 70726 45430 70790 45494
rect 71270 45430 71334 45494
rect 71678 45566 71742 45630
rect 71678 45430 71742 45494
rect 72086 45566 72150 45630
rect 72494 45566 72558 45630
rect 72222 45430 72286 45494
rect 72358 45430 72422 45494
rect 72902 45566 72966 45630
rect 73038 45430 73102 45494
rect 24350 45294 24414 45358
rect 17958 45158 18022 45222
rect 17822 45022 17886 45086
rect 18366 45022 18430 45086
rect 19046 45158 19110 45222
rect 19046 45022 19110 45086
rect 19454 45158 19518 45222
rect 70726 45158 70790 45222
rect 71270 45158 71334 45222
rect 19454 45022 19518 45086
rect 71270 45022 71334 45086
rect 71678 45158 71742 45222
rect 71678 45022 71742 45086
rect 72222 45158 72286 45222
rect 72358 45158 72422 45222
rect 72494 45022 72558 45086
rect 73038 45158 73102 45222
rect 73038 45022 73102 45086
rect 17822 44750 17886 44814
rect 17822 44614 17886 44678
rect 18366 44750 18430 44814
rect 18638 44614 18702 44678
rect 19046 44750 19110 44814
rect 19182 44614 19246 44678
rect 19454 44750 19518 44814
rect 19590 44614 19654 44678
rect 71270 44750 71334 44814
rect 71406 44614 71470 44678
rect 71678 44750 71742 44814
rect 71814 44614 71878 44678
rect 72494 44750 72558 44814
rect 72086 44614 72150 44678
rect 72358 44614 72422 44678
rect 73038 44750 73102 44814
rect 72902 44614 72966 44678
rect 17822 44342 17886 44406
rect 1230 44206 1294 44270
rect 18230 44206 18294 44270
rect 18638 44342 18702 44406
rect 18910 44206 18974 44270
rect 19182 44342 19246 44406
rect 19046 44206 19110 44270
rect 19590 44342 19654 44406
rect 19590 44206 19654 44270
rect 71406 44342 71470 44406
rect 71270 44206 71334 44270
rect 71814 44342 71878 44406
rect 71678 44206 71742 44270
rect 72086 44342 72150 44406
rect 72358 44342 72422 44406
rect 72222 44206 72286 44270
rect 72902 44342 72966 44406
rect 17958 43798 18022 43862
rect 18230 43934 18294 43998
rect 18366 43798 18430 43862
rect 18910 43934 18974 43998
rect 19046 43934 19110 43998
rect 19046 43798 19110 43862
rect 19590 43934 19654 43998
rect 19590 43798 19654 43862
rect 71270 43934 71334 43998
rect 71270 43798 71334 43862
rect 71678 43934 71742 43998
rect 71678 43798 71742 43862
rect 72222 43934 72286 43998
rect 72630 43798 72694 43862
rect 89766 43934 89830 43998
rect 73038 43798 73102 43862
rect 17958 43526 18022 43590
rect 18366 43526 18430 43590
rect 18910 43390 18974 43454
rect 19046 43526 19110 43590
rect 19046 43390 19110 43454
rect 19590 43526 19654 43590
rect 19454 43390 19518 43454
rect 71270 43526 71334 43590
rect 71406 43390 71470 43454
rect 71678 43526 71742 43590
rect 71814 43390 71878 43454
rect 72630 43526 72694 43590
rect 72222 43390 72286 43454
rect 72358 43390 72422 43454
rect 73038 43526 73102 43590
rect 17822 43118 17886 43182
rect 18910 43118 18974 43182
rect 19046 43118 19110 43182
rect 19046 42982 19110 43046
rect 19454 43118 19518 43182
rect 19454 42982 19518 43046
rect 17822 42846 17886 42910
rect 18366 42574 18430 42638
rect 19046 42710 19110 42774
rect 1230 42302 1294 42366
rect 17822 42302 17886 42366
rect 18366 42302 18430 42366
rect 19454 42710 19518 42774
rect 24350 42710 24414 42774
rect 24350 42438 24414 42502
rect 24622 42438 24686 42502
rect 24622 42166 24686 42230
rect 17822 42030 17886 42094
rect 17822 41894 17886 41958
rect 18230 41894 18294 41958
rect 19182 41894 19246 41958
rect 19454 41894 19518 41958
rect 71406 43118 71470 43182
rect 71270 42982 71334 43046
rect 71814 43118 71878 43182
rect 71814 42982 71878 43046
rect 72222 43118 72286 43182
rect 72358 43118 72422 43182
rect 73038 43118 73102 43182
rect 71270 42710 71334 42774
rect 66510 42438 66574 42502
rect 66374 42166 66438 42230
rect 66510 42166 66574 42230
rect 71814 42710 71878 42774
rect 72086 42574 72150 42638
rect 73038 42846 73102 42910
rect 72086 42302 72150 42366
rect 72902 42302 72966 42366
rect 89766 42302 89830 42366
rect 19046 41758 19110 41822
rect 17822 41622 17886 41686
rect 18230 41622 18294 41686
rect 17958 41486 18022 41550
rect 19182 41622 19246 41686
rect 19182 41486 19246 41550
rect 19454 41622 19518 41686
rect 19590 41486 19654 41550
rect 18502 41350 18566 41414
rect 17958 41214 18022 41278
rect 17958 41078 18022 41142
rect 18502 41078 18566 41142
rect 19046 41214 19110 41278
rect 19182 41214 19246 41278
rect 19182 41078 19246 41142
rect 19590 41214 19654 41278
rect 19454 41078 19518 41142
rect 66374 41894 66438 41958
rect 71270 41894 71334 41958
rect 71678 41894 71742 41958
rect 72630 41894 72694 41958
rect 72902 42030 72966 42094
rect 73038 41894 73102 41958
rect 66374 41622 66438 41686
rect 71270 41622 71334 41686
rect 71406 41486 71470 41550
rect 71678 41622 71742 41686
rect 71814 41486 71878 41550
rect 66374 41350 66438 41414
rect 72630 41622 72694 41686
rect 73038 41622 73102 41686
rect 72902 41486 72966 41550
rect 71406 41214 71470 41278
rect 71406 41078 71470 41142
rect 71814 41214 71878 41278
rect 71814 41078 71878 41142
rect 72086 41078 72150 41142
rect 72902 41214 72966 41278
rect 72902 41078 72966 41142
rect 1230 40670 1294 40734
rect 17958 40806 18022 40870
rect 17822 40670 17886 40734
rect 18366 40670 18430 40734
rect 18502 40670 18566 40734
rect 19182 40806 19246 40870
rect 19182 40670 19246 40734
rect 19454 40806 19518 40870
rect 19454 40670 19518 40734
rect 71406 40806 71470 40870
rect 71406 40670 71470 40734
rect 71814 40806 71878 40870
rect 71678 40670 71742 40734
rect 72086 40806 72150 40870
rect 72494 40670 72558 40734
rect 72902 40806 72966 40870
rect 72902 40670 72966 40734
rect 89766 40806 89830 40870
rect 17822 40398 17886 40462
rect 17958 40262 18022 40326
rect 18366 40398 18430 40462
rect 18502 40398 18566 40462
rect 18638 40262 18702 40326
rect 19182 40398 19246 40462
rect 19182 40262 19246 40326
rect 19454 40398 19518 40462
rect 71406 40398 71470 40462
rect 19590 40262 19654 40326
rect 17958 39990 18022 40054
rect 17822 39854 17886 39918
rect 18230 39854 18294 39918
rect 18638 39990 18702 40054
rect 18910 39854 18974 39918
rect 19182 39990 19246 40054
rect 19046 39854 19110 39918
rect 19590 39990 19654 40054
rect 19590 39854 19654 39918
rect 71406 40262 71470 40326
rect 71678 40398 71742 40462
rect 71678 40262 71742 40326
rect 72494 40398 72558 40462
rect 72086 40262 72150 40326
rect 72358 40262 72422 40326
rect 72902 40398 72966 40462
rect 72902 40262 72966 40326
rect 71406 39990 71470 40054
rect 71270 39854 71334 39918
rect 71678 39990 71742 40054
rect 71814 39854 71878 39918
rect 72086 39990 72150 40054
rect 72358 39990 72422 40054
rect 72222 39854 72286 39918
rect 72358 39854 72422 39918
rect 72902 39990 72966 40054
rect 73038 39854 73102 39918
rect 17822 39582 17886 39646
rect 18230 39582 18294 39646
rect 18910 39582 18974 39646
rect 18366 39446 18430 39510
rect 18502 39446 18566 39510
rect 18774 39446 18838 39510
rect 19046 39582 19110 39646
rect 19182 39446 19246 39510
rect 19590 39582 19654 39646
rect 19454 39446 19518 39510
rect 1230 39174 1294 39238
rect 24350 39310 24414 39374
rect 71270 39582 71334 39646
rect 71270 39446 71334 39510
rect 71814 39582 71878 39646
rect 71814 39446 71878 39510
rect 72222 39582 72286 39646
rect 72358 39582 72422 39646
rect 72086 39446 72150 39510
rect 73038 39582 73102 39646
rect 66374 39310 66438 39374
rect 18366 39174 18430 39238
rect 18502 39174 18566 39238
rect 18774 39174 18838 39238
rect 19182 39174 19246 39238
rect 19046 39038 19110 39102
rect 19454 39174 19518 39238
rect 19454 39038 19518 39102
rect 24350 39038 24414 39102
rect 18910 38630 18974 38694
rect 19046 38766 19110 38830
rect 19454 38766 19518 38830
rect 66374 39038 66438 39102
rect 71270 39174 71334 39238
rect 71270 39038 71334 39102
rect 71814 39174 71878 39238
rect 71814 39038 71878 39102
rect 72086 39174 72150 39238
rect 89766 39174 89830 39238
rect 66510 38766 66574 38830
rect 71270 38766 71334 38830
rect 17822 38358 17886 38422
rect 18910 38358 18974 38422
rect 11158 37950 11222 38014
rect 17822 38086 17886 38150
rect 17822 37950 17886 38014
rect 18502 37950 18566 38014
rect 24622 38086 24686 38150
rect 66510 38494 66574 38558
rect 71814 38766 71878 38830
rect 72222 38630 72286 38694
rect 66374 38086 66438 38150
rect 66510 38086 66574 38150
rect 17822 37678 17886 37742
rect 17958 37542 18022 37606
rect 18502 37678 18566 37742
rect 19046 37542 19110 37606
rect 19590 37542 19654 37606
rect 24622 37814 24686 37878
rect 66374 37814 66438 37878
rect 66510 37678 66574 37742
rect 72222 38358 72286 38422
rect 72902 38358 72966 38422
rect 72086 37950 72150 38014
rect 72902 38086 72966 38150
rect 72902 37950 72966 38014
rect 71270 37542 71334 37606
rect 71678 37542 71742 37606
rect 72086 37678 72150 37742
rect 72902 37678 72966 37742
rect 73038 37542 73102 37606
rect 1230 37270 1294 37334
rect 17958 37270 18022 37334
rect 17822 37134 17886 37198
rect 18366 37134 18430 37198
rect 19046 37270 19110 37334
rect 19182 37134 19246 37198
rect 19590 37270 19654 37334
rect 71270 37270 71334 37334
rect 19454 37134 19518 37198
rect 17822 36862 17886 36926
rect 17958 36726 18022 36790
rect 18366 36862 18430 36926
rect 18230 36726 18294 36790
rect 18910 36726 18974 36790
rect 19182 36862 19246 36926
rect 19182 36726 19246 36790
rect 19454 36862 19518 36926
rect 19590 36726 19654 36790
rect 24622 36862 24686 36926
rect 71406 37134 71470 37198
rect 71678 37270 71742 37334
rect 71678 37134 71742 37198
rect 72494 37134 72558 37198
rect 73038 37270 73102 37334
rect 89766 37270 89830 37334
rect 72902 37134 72966 37198
rect 66374 36862 66438 36926
rect 71406 36862 71470 36926
rect 71270 36726 71334 36790
rect 71678 36862 71742 36926
rect 71678 36726 71742 36790
rect 72494 36862 72558 36926
rect 72086 36726 72150 36790
rect 72358 36726 72422 36790
rect 72902 36862 72966 36926
rect 73038 36726 73102 36790
rect 24622 36590 24686 36654
rect 11294 36454 11358 36518
rect 17958 36454 18022 36518
rect 17822 36318 17886 36382
rect 18230 36454 18294 36518
rect 18910 36454 18974 36518
rect 19182 36454 19246 36518
rect 19046 36318 19110 36382
rect 19590 36454 19654 36518
rect 66374 36590 66438 36654
rect 19454 36318 19518 36382
rect 71270 36454 71334 36518
rect 71270 36318 71334 36382
rect 71678 36454 71742 36518
rect 71678 36318 71742 36382
rect 72086 36454 72150 36518
rect 72358 36454 72422 36518
rect 72494 36318 72558 36382
rect 73038 36454 73102 36518
rect 72902 36318 72966 36382
rect 17822 36046 17886 36110
rect 17822 35910 17886 35974
rect 18910 35910 18974 35974
rect 19046 36046 19110 36110
rect 19182 35910 19246 35974
rect 19454 36046 19518 36110
rect 19454 35910 19518 35974
rect 71270 36046 71334 36110
rect 71406 35910 71470 35974
rect 71678 36046 71742 36110
rect 71678 35910 71742 35974
rect 72494 36046 72558 36110
rect 72086 35910 72150 35974
rect 72358 35910 72422 35974
rect 72902 36046 72966 36110
rect 72902 35910 72966 35974
rect 1230 35638 1294 35702
rect 17822 35638 17886 35702
rect 18910 35638 18974 35702
rect 18502 35502 18566 35566
rect 18910 35502 18974 35566
rect 19182 35638 19246 35702
rect 19046 35502 19110 35566
rect 19454 35638 19518 35702
rect 19590 35502 19654 35566
rect 11158 35230 11222 35294
rect 11022 35094 11086 35158
rect 71406 35638 71470 35702
rect 71270 35502 71334 35566
rect 71678 35638 71742 35702
rect 71814 35502 71878 35566
rect 72086 35638 72150 35702
rect 72358 35638 72422 35702
rect 72222 35502 72286 35566
rect 72358 35502 72422 35566
rect 72902 35638 72966 35702
rect 89766 35638 89830 35702
rect 18502 35230 18566 35294
rect 18910 35230 18974 35294
rect 19046 35230 19110 35294
rect 19046 35094 19110 35158
rect 19590 35230 19654 35294
rect 19454 35094 19518 35158
rect 18638 34686 18702 34750
rect 19046 34822 19110 34886
rect 19046 34686 19110 34750
rect 19454 34822 19518 34886
rect 19454 34686 19518 34750
rect 71270 35230 71334 35294
rect 71270 35094 71334 35158
rect 71814 35230 71878 35294
rect 71814 35094 71878 35158
rect 72222 35230 72286 35294
rect 72358 35230 72422 35294
rect 24622 34550 24686 34614
rect 71270 34822 71334 34886
rect 71270 34686 71334 34750
rect 71814 34822 71878 34886
rect 71678 34686 71742 34750
rect 72222 34686 72286 34750
rect 17958 34414 18022 34478
rect 18638 34414 18702 34478
rect 19046 34414 19110 34478
rect 19454 34414 19518 34478
rect 24622 34278 24686 34342
rect 17958 34142 18022 34206
rect 1230 34006 1294 34070
rect 17822 34006 17886 34070
rect 18230 34006 18294 34070
rect 18638 34006 18702 34070
rect 11294 33870 11358 33934
rect 24622 34142 24686 34206
rect 66510 34142 66574 34206
rect 71270 34414 71334 34478
rect 71678 34414 71742 34478
rect 72222 34414 72286 34478
rect 73038 34414 73102 34478
rect 11158 33598 11222 33662
rect 17822 33734 17886 33798
rect 17822 33598 17886 33662
rect 18230 33734 18294 33798
rect 18638 33734 18702 33798
rect 18502 33598 18566 33662
rect 19182 33598 19246 33662
rect 19590 33598 19654 33662
rect 24486 33734 24550 33798
rect 24622 33734 24686 33798
rect 66510 33870 66574 33934
rect 66374 33734 66438 33798
rect 71406 33598 71470 33662
rect 72630 34006 72694 34070
rect 73038 34142 73102 34206
rect 72902 34006 72966 34070
rect 89766 34006 89830 34070
rect 71814 33598 71878 33662
rect 24486 33462 24550 33526
rect 17822 33326 17886 33390
rect 17958 33190 18022 33254
rect 18502 33326 18566 33390
rect 18638 33190 18702 33254
rect 19182 33326 19246 33390
rect 19046 33190 19110 33254
rect 19590 33326 19654 33390
rect 19590 33190 19654 33254
rect 66374 33462 66438 33526
rect 72630 33734 72694 33798
rect 72902 33734 72966 33798
rect 72902 33598 72966 33662
rect 72358 33462 72422 33526
rect 17958 32918 18022 32982
rect 17822 32782 17886 32846
rect 18366 32782 18430 32846
rect 18638 32918 18702 32982
rect 19046 32918 19110 32982
rect 19182 32782 19246 32846
rect 19590 32918 19654 32982
rect 19454 32782 19518 32846
rect 17822 32510 17886 32574
rect 1230 32238 1294 32302
rect 11022 32374 11086 32438
rect 17958 32374 18022 32438
rect 18366 32510 18430 32574
rect 18366 32374 18430 32438
rect 18774 32374 18838 32438
rect 19182 32510 19246 32574
rect 19182 32374 19246 32438
rect 19454 32510 19518 32574
rect 19590 32374 19654 32438
rect 11022 32238 11086 32302
rect 71406 33326 71470 33390
rect 71270 33190 71334 33254
rect 71814 33326 71878 33390
rect 71814 33190 71878 33254
rect 72358 33190 72422 33254
rect 72630 33190 72694 33254
rect 72902 33326 72966 33390
rect 73038 33190 73102 33254
rect 66374 32918 66438 32982
rect 71270 32918 71334 32982
rect 71406 32782 71470 32846
rect 71814 32918 71878 32982
rect 71678 32782 71742 32846
rect 72630 32918 72694 32982
rect 72358 32782 72422 32846
rect 73038 32918 73102 32982
rect 72902 32782 72966 32846
rect 66374 32646 66438 32710
rect 71406 32510 71470 32574
rect 71406 32374 71470 32438
rect 71678 32510 71742 32574
rect 71814 32374 71878 32438
rect 72358 32510 72422 32574
rect 72086 32374 72150 32438
rect 72630 32374 72694 32438
rect 72902 32510 72966 32574
rect 73038 32374 73102 32438
rect 89766 32374 89830 32438
rect 17958 32102 18022 32166
rect 17958 31966 18022 32030
rect 18366 32102 18430 32166
rect 18774 32102 18838 32166
rect 18502 31966 18566 32030
rect 19182 32102 19246 32166
rect 19046 31966 19110 32030
rect 19590 32102 19654 32166
rect 19454 31966 19518 32030
rect 71406 32102 71470 32166
rect 71406 31966 71470 32030
rect 71814 32102 71878 32166
rect 71678 31966 71742 32030
rect 72086 32102 72150 32166
rect 72630 32102 72694 32166
rect 72494 31966 72558 32030
rect 73038 32102 73102 32166
rect 73038 31966 73102 32030
rect 17958 31694 18022 31758
rect 18502 31694 18566 31758
rect 18366 31558 18430 31622
rect 19046 31694 19110 31758
rect 19182 31558 19246 31622
rect 19454 31694 19518 31758
rect 71406 31694 71470 31758
rect 19454 31558 19518 31622
rect 24486 31422 24550 31486
rect 18366 31286 18430 31350
rect 19182 31286 19246 31350
rect 19046 31150 19110 31214
rect 19454 31286 19518 31350
rect 19454 31150 19518 31214
rect 24486 31150 24550 31214
rect 11158 31014 11222 31078
rect 11158 30878 11222 30942
rect 1230 30742 1294 30806
rect 18502 30742 18566 30806
rect 19046 30878 19110 30942
rect 19182 30742 19246 30806
rect 19454 30878 19518 30942
rect 19590 30742 19654 30806
rect 71406 31558 71470 31622
rect 71678 31694 71742 31758
rect 71678 31558 71742 31622
rect 72494 31694 72558 31758
rect 72086 31558 72150 31622
rect 73038 31694 73102 31758
rect 71406 31286 71470 31350
rect 71270 31150 71334 31214
rect 71678 31286 71742 31350
rect 71814 31150 71878 31214
rect 72086 31286 72150 31350
rect 24622 30606 24686 30670
rect 71270 30878 71334 30942
rect 71406 30742 71470 30806
rect 71814 30878 71878 30942
rect 71814 30742 71878 30806
rect 72086 30742 72150 30806
rect 17822 30470 17886 30534
rect 18502 30470 18566 30534
rect 19182 30470 19246 30534
rect 17822 30198 17886 30262
rect 17822 30062 17886 30126
rect 18638 30062 18702 30126
rect 19590 30470 19654 30534
rect 24622 30334 24686 30398
rect 24486 30198 24550 30262
rect 71406 30470 71470 30534
rect 71814 30470 71878 30534
rect 66374 30198 66438 30262
rect 24486 29926 24550 29990
rect 17822 29790 17886 29854
rect 17822 29654 17886 29718
rect 11022 29518 11086 29582
rect 18638 29790 18702 29854
rect 14830 29382 14894 29446
rect 17822 29382 17886 29446
rect 17822 29246 17886 29310
rect 18774 29246 18838 29310
rect 19046 29246 19110 29310
rect 19454 29246 19518 29310
rect 1230 28838 1294 28902
rect 17822 28974 17886 29038
rect 17822 28838 17886 28902
rect 18774 28974 18838 29038
rect 18230 28838 18294 28902
rect 18502 28838 18566 28902
rect 19046 28974 19110 29038
rect 19046 28838 19110 28902
rect 19454 28974 19518 29038
rect 19590 28838 19654 28902
rect 66374 29926 66438 29990
rect 72086 30470 72150 30534
rect 89766 30606 89830 30670
rect 72902 30470 72966 30534
rect 72222 30062 72286 30126
rect 72630 30062 72694 30126
rect 72902 30198 72966 30262
rect 73038 30062 73102 30126
rect 66510 29790 66574 29854
rect 66510 29518 66574 29582
rect 71406 29246 71470 29310
rect 72222 29790 72286 29854
rect 72630 29790 72694 29854
rect 73038 29790 73102 29854
rect 73038 29654 73102 29718
rect 71814 29246 71878 29310
rect 73038 29382 73102 29446
rect 73038 29246 73102 29310
rect 66510 28974 66574 29038
rect 71406 28974 71470 29038
rect 71270 28838 71334 28902
rect 71814 28974 71878 29038
rect 71814 28838 71878 28902
rect 72494 28838 72558 28902
rect 73038 28974 73102 29038
rect 73038 28838 73102 28902
rect 89766 28974 89830 29038
rect 17822 28566 17886 28630
rect 17822 28430 17886 28494
rect 18230 28566 18294 28630
rect 18502 28566 18566 28630
rect 18366 28430 18430 28494
rect 19046 28566 19110 28630
rect 19182 28430 19246 28494
rect 19590 28566 19654 28630
rect 66510 28702 66574 28766
rect 71270 28566 71334 28630
rect 19590 28430 19654 28494
rect 11158 28158 11222 28222
rect 17822 28158 17886 28222
rect 12926 28022 12990 28086
rect 17822 28022 17886 28086
rect 18366 28158 18430 28222
rect 18230 28022 18294 28086
rect 18774 28022 18838 28086
rect 19182 28158 19246 28222
rect 19046 28022 19110 28086
rect 19590 28158 19654 28222
rect 19590 28022 19654 28086
rect 71406 28430 71470 28494
rect 71814 28566 71878 28630
rect 71678 28430 71742 28494
rect 72086 28430 72150 28494
rect 72494 28566 72558 28630
rect 72494 28430 72558 28494
rect 73038 28566 73102 28630
rect 72902 28430 72966 28494
rect 71406 28158 71470 28222
rect 71270 28022 71334 28086
rect 71678 28158 71742 28222
rect 71678 28022 71742 28086
rect 72086 28158 72150 28222
rect 72222 28022 72286 28086
rect 72494 28158 72558 28222
rect 72902 28158 72966 28222
rect 72902 28022 72966 28086
rect 14558 27614 14622 27678
rect 14830 27750 14894 27814
rect 15374 27614 15438 27678
rect 15782 27614 15846 27678
rect 17822 27750 17886 27814
rect 18230 27750 18294 27814
rect 18774 27750 18838 27814
rect 18502 27614 18566 27678
rect 18774 27614 18838 27678
rect 19046 27750 19110 27814
rect 19046 27614 19110 27678
rect 19590 27750 19654 27814
rect 19454 27614 19518 27678
rect 1230 27206 1294 27270
rect 71270 27750 71334 27814
rect 71270 27614 71334 27678
rect 71678 27750 71742 27814
rect 71678 27614 71742 27678
rect 72222 27750 72286 27814
rect 72630 27614 72694 27678
rect 72902 27750 72966 27814
rect 74806 27614 74870 27678
rect 75214 27614 75278 27678
rect 76438 27614 76502 27678
rect 17822 27206 17886 27270
rect 18502 27342 18566 27406
rect 18774 27342 18838 27406
rect 18638 27206 18702 27270
rect 19046 27342 19110 27406
rect 19182 27206 19246 27270
rect 19454 27342 19518 27406
rect 19590 27206 19654 27270
rect 14558 26934 14622 26998
rect 15374 26934 15438 26998
rect 14422 26798 14486 26862
rect 15102 26798 15166 26862
rect 15782 26934 15846 26998
rect 15646 26798 15710 26862
rect 16190 26798 16254 26862
rect 17822 26934 17886 26998
rect 18638 26934 18702 26998
rect 18502 26798 18566 26862
rect 18910 26798 18974 26862
rect 19182 26934 19246 26998
rect 19046 26798 19110 26862
rect 19590 26934 19654 26998
rect 19454 26798 19518 26862
rect 71270 27342 71334 27406
rect 71406 27206 71470 27270
rect 71678 27342 71742 27406
rect 71678 27206 71742 27270
rect 72630 27342 72694 27406
rect 72494 27206 72558 27270
rect 72902 27206 72966 27270
rect 89766 27342 89830 27406
rect 71406 26934 71470 26998
rect 71270 26798 71334 26862
rect 71678 26934 71742 26998
rect 71814 26798 71878 26862
rect 72494 26934 72558 26998
rect 72358 26798 72422 26862
rect 72902 26934 72966 26998
rect 74806 26934 74870 26998
rect 75214 26934 75278 26998
rect 75214 26798 75278 26862
rect 76030 26798 76094 26862
rect 76438 26934 76502 26998
rect 76302 26798 76366 26862
rect 17958 26526 18022 26590
rect 18502 26526 18566 26590
rect 18910 26526 18974 26590
rect 19046 26526 19110 26590
rect 19182 26390 19246 26454
rect 19454 26526 19518 26590
rect 19454 26390 19518 26454
rect 550 26254 614 26318
rect 14422 26254 14486 26318
rect 14422 25982 14486 26046
rect 15102 26254 15166 26318
rect 15918 26254 15982 26318
rect 17958 26254 18022 26318
rect 14830 25982 14894 26046
rect 15102 25982 15166 26046
rect 15646 26118 15710 26182
rect 15782 25982 15846 26046
rect 16190 26118 16254 26182
rect 16054 25982 16118 26046
rect 17686 25982 17750 26046
rect 19182 26118 19246 26182
rect 18638 25982 18702 26046
rect 19454 26118 19518 26182
rect 2461 25728 2525 25732
rect 2461 25672 2465 25728
rect 2465 25672 2521 25728
rect 2521 25672 2525 25728
rect 2461 25668 2525 25672
rect 17958 25710 18022 25774
rect 1230 25574 1294 25638
rect 2182 25574 2246 25638
rect 14830 25574 14894 25638
rect 17686 25574 17750 25638
rect 18638 25710 18702 25774
rect 12926 25438 12990 25502
rect 14422 25438 14486 25502
rect 15102 25438 15166 25502
rect 15782 25438 15846 25502
rect 15918 25438 15982 25502
rect 16054 25438 16118 25502
rect 14694 25302 14758 25366
rect 17958 25438 18022 25502
rect 17822 25302 17886 25366
rect 18230 25302 18294 25366
rect 18502 25302 18566 25366
rect 19046 25302 19110 25366
rect 71270 26526 71334 26590
rect 71270 26390 71334 26454
rect 71814 26526 71878 26590
rect 71678 26390 71742 26454
rect 72358 26526 72422 26590
rect 73038 26526 73102 26590
rect 74670 26390 74734 26454
rect 71270 26118 71334 26182
rect 24622 25846 24686 25910
rect 24622 25574 24686 25638
rect 71678 26118 71742 26182
rect 72222 25982 72286 26046
rect 73038 26254 73102 26318
rect 76030 26254 76094 26318
rect 76302 26254 76366 26318
rect 74670 26118 74734 26182
rect 74670 25982 74734 26046
rect 75214 26118 75278 26182
rect 75078 25982 75142 26046
rect 75758 25982 75822 26046
rect 76302 25982 76366 26046
rect 76438 25982 76502 26046
rect 66374 25846 66438 25910
rect 66374 25574 66438 25638
rect 19590 25302 19654 25366
rect 15238 25166 15302 25230
rect 2182 25030 2246 25094
rect 17822 25030 17886 25094
rect 17822 24894 17886 24958
rect 18230 25030 18294 25094
rect 18502 25030 18566 25094
rect 18774 24894 18838 24958
rect 19046 25030 19110 25094
rect 19182 24894 19246 24958
rect 19590 25030 19654 25094
rect 19454 24894 19518 24958
rect 24622 25030 24686 25094
rect 72222 25710 72286 25774
rect 77390 25846 77454 25910
rect 73038 25710 73102 25774
rect 76302 25574 76366 25638
rect 89766 25574 89830 25638
rect 71406 25302 71470 25366
rect 71678 25302 71742 25366
rect 72222 25302 72286 25366
rect 73038 25438 73102 25502
rect 72902 25302 72966 25366
rect 74670 25438 74734 25502
rect 75078 25438 75142 25502
rect 74670 25302 74734 25366
rect 75758 25438 75822 25502
rect 76438 25438 76502 25502
rect 77390 25438 77454 25502
rect 76302 25302 76366 25366
rect 66374 25030 66438 25094
rect 71406 25030 71470 25094
rect 71406 24894 71470 24958
rect 71678 25030 71742 25094
rect 71678 24894 71742 24958
rect 72222 25030 72286 25094
rect 72222 24894 72286 24958
rect 72902 25030 72966 25094
rect 73038 24894 73102 24958
rect 24622 24758 24686 24822
rect 17822 24622 17886 24686
rect 17958 24486 18022 24550
rect 18230 24486 18294 24550
rect 18774 24622 18838 24686
rect 18638 24486 18702 24550
rect 19182 24622 19246 24686
rect 19046 24486 19110 24550
rect 19454 24622 19518 24686
rect 19590 24486 19654 24550
rect 66374 24758 66438 24822
rect 71406 24622 71470 24686
rect 71270 24486 71334 24550
rect 71678 24622 71742 24686
rect 71678 24486 71742 24550
rect 72222 24622 72286 24686
rect 72630 24486 72694 24550
rect 73038 24622 73102 24686
rect 73038 24486 73102 24550
rect 17958 24214 18022 24278
rect 17822 24078 17886 24142
rect 18230 24214 18294 24278
rect 18638 24214 18702 24278
rect 18366 24078 18430 24142
rect 18502 24078 18566 24142
rect 19046 24214 19110 24278
rect 19182 24078 19246 24142
rect 19590 24214 19654 24278
rect 19454 24078 19518 24142
rect 71270 24214 71334 24278
rect 71406 24078 71470 24142
rect 71678 24214 71742 24278
rect 71678 24078 71742 24142
rect 72086 24078 72150 24142
rect 72630 24214 72694 24278
rect 72494 24078 72558 24142
rect 73038 24214 73102 24278
rect 72902 24078 72966 24142
rect 75078 24078 75142 24142
rect 1230 23806 1294 23870
rect 14694 23806 14758 23870
rect 15238 23806 15302 23870
rect 15238 23670 15302 23734
rect 15782 23670 15846 23734
rect 16190 23670 16254 23734
rect 17822 23806 17886 23870
rect 17822 23670 17886 23734
rect 18366 23806 18430 23870
rect 18502 23806 18566 23870
rect 18230 23670 18294 23734
rect 19182 23806 19246 23870
rect 19182 23670 19246 23734
rect 19454 23806 19518 23870
rect 71406 23806 71470 23870
rect 19454 23670 19518 23734
rect 71270 23670 71334 23734
rect 71678 23806 71742 23870
rect 71678 23670 71742 23734
rect 72086 23806 72150 23870
rect 72086 23670 72150 23734
rect 72494 23806 72558 23870
rect 72902 23806 72966 23870
rect 73038 23670 73102 23734
rect 74670 23806 74734 23870
rect 75078 23806 75142 23870
rect 74670 23670 74734 23734
rect 75486 23670 75550 23734
rect 76302 23806 76366 23870
rect 89766 23806 89830 23870
rect 76030 23670 76094 23734
rect 3678 23398 3742 23462
rect 17822 23398 17886 23462
rect 17822 23262 17886 23326
rect 18230 23398 18294 23462
rect 18502 23262 18566 23326
rect 19182 23398 19246 23462
rect 19182 23262 19246 23326
rect 19454 23398 19518 23462
rect 19590 23262 19654 23326
rect 71270 23398 71334 23462
rect 71270 23262 71334 23326
rect 71678 23398 71742 23462
rect 71678 23262 71742 23326
rect 72086 23398 72150 23462
rect 72086 23262 72150 23326
rect 73038 23398 73102 23462
rect 72902 23262 72966 23326
rect 15238 22990 15302 23054
rect 15238 22854 15302 22918
rect 15782 22990 15846 23054
rect 15646 22854 15710 22918
rect 16190 22990 16254 23054
rect 17822 22990 17886 23054
rect 18502 22990 18566 23054
rect 19182 22990 19246 23054
rect 19182 22854 19246 22918
rect 19590 22990 19654 23054
rect 71270 22990 71334 23054
rect 19590 22854 19654 22918
rect 15102 22582 15166 22646
rect 15646 22582 15710 22646
rect 17958 22582 18022 22646
rect 19182 22582 19246 22646
rect 19046 22446 19110 22510
rect 19590 22582 19654 22646
rect 19454 22446 19518 22510
rect 1230 22174 1294 22238
rect 17958 22310 18022 22374
rect 18366 22038 18430 22102
rect 18774 22038 18838 22102
rect 19046 22174 19110 22238
rect 19454 22174 19518 22238
rect 17822 21766 17886 21830
rect 18366 21766 18430 21830
rect 18774 21766 18838 21830
rect 15102 21494 15166 21558
rect 15238 21494 15302 21558
rect 15782 21222 15846 21286
rect 17822 21494 17886 21558
rect 17958 21358 18022 21422
rect 18910 21358 18974 21422
rect 16190 21222 16254 21286
rect 71406 22854 71470 22918
rect 71678 22990 71742 23054
rect 71814 22854 71878 22918
rect 72086 22990 72150 23054
rect 72086 22854 72150 22918
rect 72494 22854 72558 22918
rect 72902 22990 72966 23054
rect 74670 22990 74734 23054
rect 75486 22990 75550 23054
rect 75078 22854 75142 22918
rect 76030 22990 76094 23054
rect 75486 22854 75550 22918
rect 71406 22582 71470 22646
rect 71270 22446 71334 22510
rect 71814 22582 71878 22646
rect 71678 22446 71742 22510
rect 72086 22582 72150 22646
rect 72494 22582 72558 22646
rect 72902 22582 72966 22646
rect 24350 21902 24414 21966
rect 24350 21630 24414 21694
rect 24486 21630 24550 21694
rect 24622 21494 24686 21558
rect 66374 21902 66438 21966
rect 66374 21630 66438 21694
rect 71270 22174 71334 22238
rect 71678 22174 71742 22238
rect 72086 22038 72150 22102
rect 72902 22310 72966 22374
rect 89766 22174 89830 22238
rect 66510 21494 66574 21558
rect 17958 21086 18022 21150
rect 17958 20950 18022 21014
rect 550 20814 614 20878
rect 3678 20814 3742 20878
rect 18910 21086 18974 21150
rect 19046 20950 19110 21014
rect 19590 20950 19654 21014
rect 24486 21222 24550 21286
rect 24622 21222 24686 21286
rect 66510 21222 66574 21286
rect 72086 21766 72150 21830
rect 72902 21766 72966 21830
rect 72222 21358 72286 21422
rect 72902 21494 72966 21558
rect 73038 21358 73102 21422
rect 75078 21494 75142 21558
rect 74806 21222 74870 21286
rect 75486 21494 75550 21558
rect 75486 21358 75550 21422
rect 75894 21358 75958 21422
rect 75078 21222 75142 21286
rect 66510 21086 66574 21150
rect 71406 20950 71470 21014
rect 71814 20950 71878 21014
rect 72222 21086 72286 21150
rect 18502 20814 18566 20878
rect 3950 20542 4014 20606
rect 13606 20542 13670 20606
rect 14014 20542 14078 20606
rect 15782 20678 15846 20742
rect 16190 20678 16254 20742
rect 17958 20678 18022 20742
rect 18502 20542 18566 20606
rect 19046 20678 19110 20742
rect 19046 20542 19110 20606
rect 19590 20678 19654 20742
rect 19454 20542 19518 20606
rect 1230 20406 1294 20470
rect 66510 20814 66574 20878
rect 73038 21086 73102 21150
rect 73038 20950 73102 21014
rect 71406 20678 71470 20742
rect 71814 20678 71878 20742
rect 73038 20678 73102 20742
rect 74806 20678 74870 20742
rect 75078 20678 75142 20742
rect 75486 20678 75550 20742
rect 75894 20678 75958 20742
rect 77118 20542 77182 20606
rect 79838 20542 79902 20606
rect 89766 20542 89830 20606
rect 19454 20134 19518 20198
rect 79838 20270 79902 20334
rect 66374 20134 66438 20198
rect 79974 20134 80038 20198
rect 19182 19862 19246 19926
rect 25302 19590 25366 19654
rect 26526 19590 26590 19654
rect 28158 19590 28222 19654
rect 29518 19590 29582 19654
rect 29654 19590 29718 19654
rect 30334 19590 30398 19654
rect 31558 19590 31622 19654
rect 31966 19590 32030 19654
rect 32646 19590 32710 19654
rect 33190 19590 33254 19654
rect 34550 19590 34614 19654
rect 35230 19590 35294 19654
rect 35774 19590 35838 19654
rect 36454 19590 36518 19654
rect 38358 19590 38422 19654
rect 40806 19590 40870 19654
rect 41486 19590 41550 19654
rect 42710 19590 42774 19654
rect 43934 19590 43998 19654
rect 44478 19590 44542 19654
rect 45566 19590 45630 19654
rect 46926 19590 46990 19654
rect 47878 19590 47942 19654
rect 49374 19590 49438 19654
rect 50190 19590 50254 19654
rect 50734 19590 50798 19654
rect 51958 19590 52022 19654
rect 53182 19590 53246 19654
rect 54134 19590 54198 19654
rect 55766 19590 55830 19654
rect 56990 19590 57054 19654
rect 58214 19590 58278 19654
rect 58894 19590 58958 19654
rect 59438 19590 59502 19654
rect 60118 19590 60182 19654
rect 60662 19590 60726 19654
rect 61886 19590 61950 19654
rect 62838 19590 62902 19654
rect 63926 19590 63990 19654
rect 65694 19590 65758 19654
rect 3134 19182 3198 19246
rect 13606 19318 13670 19382
rect 11566 19182 11630 19246
rect 25302 19046 25366 19110
rect 3134 18910 3198 18974
rect 26526 19046 26590 19110
rect 26798 18910 26862 18974
rect 28158 19046 28222 19110
rect 29518 19046 29582 19110
rect 29654 19046 29718 19110
rect 30334 19046 30398 19110
rect 30742 18910 30806 18974
rect 31558 19046 31622 19110
rect 31966 19046 32030 19110
rect 32646 19046 32710 19110
rect 33190 19046 33254 19110
rect 34550 19046 34614 19110
rect 35230 19046 35294 19110
rect 35774 19046 35838 19110
rect 36454 19046 36518 19110
rect 36454 18910 36518 18974
rect 38358 19046 38422 19110
rect 40806 19046 40870 19110
rect 41486 19046 41550 19110
rect 41486 18910 41550 18974
rect 42710 19046 42774 19110
rect 43934 19046 43998 19110
rect 44478 19046 44542 19110
rect 45566 19046 45630 19110
rect 45702 18910 45766 18974
rect 46926 19046 46990 19110
rect 47878 19046 47942 19110
rect 49374 19046 49438 19110
rect 50190 19046 50254 19110
rect 50734 19046 50798 19110
rect 51958 19046 52022 19110
rect 51414 18910 51478 18974
rect 53182 19046 53246 19110
rect 54134 19046 54198 19110
rect 55766 19046 55830 19110
rect 55766 18910 55830 18974
rect 56990 19046 57054 19110
rect 58214 19046 58278 19110
rect 58894 19046 58958 19110
rect 59438 19046 59502 19110
rect 60118 19046 60182 19110
rect 60662 19046 60726 19110
rect 61886 19046 61950 19110
rect 61478 18910 61542 18974
rect 62838 19046 62902 19110
rect 63926 19046 63990 19110
rect 65694 19046 65758 19110
rect 77118 18910 77182 18974
rect 1230 18774 1294 18838
rect 89766 18774 89830 18838
rect 79838 18638 79902 18702
rect 2461 18261 2525 18325
rect 3950 17958 4014 18022
rect 14014 17958 14078 18022
rect 11702 17822 11766 17886
rect 19046 17686 19110 17750
rect 16598 17550 16662 17614
rect 25982 17414 26046 17478
rect 31150 17414 31214 17478
rect 36182 17414 36246 17478
rect 40942 17414 41006 17478
rect 45974 17414 46038 17478
rect 51142 17414 51206 17478
rect 56174 17414 56238 17478
rect 60934 17414 60998 17478
rect 66374 17550 66438 17614
rect 79974 17414 80038 17478
rect 79974 17278 80038 17342
rect 1230 17142 1294 17206
rect 2454 17142 2518 17206
rect 89766 17142 89830 17206
rect 2454 16462 2518 16526
rect 11566 16462 11630 16526
rect 11430 16326 11494 16390
rect 19182 16326 19246 16390
rect 16462 16190 16526 16254
rect 79838 16054 79902 16118
rect 79838 15918 79902 15982
rect 1230 15646 1294 15710
rect 89766 15510 89830 15574
rect 550 15102 614 15166
rect 11702 15102 11766 15166
rect 11566 14966 11630 15030
rect 25982 14966 26046 15030
rect 26118 14966 26182 15030
rect 31014 14966 31078 15030
rect 31150 14966 31214 15030
rect 36046 14966 36110 15030
rect 36182 14966 36246 15030
rect 40942 14966 41006 15030
rect 41078 14966 41142 15030
rect 45838 14966 45902 15030
rect 45974 14966 46038 15030
rect 51006 14966 51070 15030
rect 51142 14966 51206 15030
rect 56038 14966 56102 15030
rect 56174 14966 56238 15030
rect 60934 14966 60998 15030
rect 61070 14966 61134 15030
rect 16598 14830 16662 14894
rect 16598 14694 16662 14758
rect 79974 14558 80038 14622
rect 79974 14422 80038 14486
rect 26798 14286 26862 14350
rect 30742 14286 30806 14350
rect 25982 14150 26046 14214
rect 30742 14150 30806 14214
rect 36454 14286 36518 14350
rect 41486 14286 41550 14350
rect 45702 14286 45766 14350
rect 35774 14150 35838 14214
rect 40942 14150 41006 14214
rect 45974 14150 46038 14214
rect 51414 14286 51478 14350
rect 55766 14286 55830 14350
rect 50734 14150 50798 14214
rect 55766 14150 55830 14214
rect 61478 14286 61542 14350
rect 60798 14150 60862 14214
rect 89766 13878 89830 13942
rect 1230 13742 1294 13806
rect 11430 13742 11494 13806
rect 11702 13470 11766 13534
rect 16462 13470 16526 13534
rect 25982 13470 26046 13534
rect 30742 13470 30806 13534
rect 35774 13470 35838 13534
rect 40942 13470 41006 13534
rect 17958 13334 18022 13398
rect 25982 13334 26046 13398
rect 30878 13334 30942 13398
rect 35910 13334 35974 13398
rect 40942 13334 41006 13398
rect 45974 13470 46038 13534
rect 50734 13470 50798 13534
rect 55766 13470 55830 13534
rect 60798 13470 60862 13534
rect 45702 13334 45766 13398
rect 50870 13334 50934 13398
rect 55902 13334 55966 13398
rect 60934 13334 60998 13398
rect 26118 13198 26182 13262
rect 25302 12926 25366 12990
rect 31014 13198 31078 13262
rect 30470 12926 30534 12990
rect 31014 12926 31078 12990
rect 36046 13198 36110 13262
rect 35502 12926 35566 12990
rect 41078 13198 41142 13262
rect 40534 12926 40598 12990
rect 45838 13198 45902 13262
rect 45566 12926 45630 12990
rect 45838 12926 45902 12990
rect 51006 13198 51070 13262
rect 50462 12926 50526 12990
rect 56038 13198 56102 13262
rect 55494 12926 55558 12990
rect 61070 13198 61134 13262
rect 79838 13198 79902 13262
rect 79838 13062 79902 13126
rect 60526 12926 60590 12990
rect 25846 12790 25910 12854
rect 35774 12790 35838 12854
rect 40806 12790 40870 12854
rect 50734 12790 50798 12854
rect 55766 12790 55830 12854
rect 60798 12790 60862 12854
rect 25846 12382 25910 12446
rect 1230 12246 1294 12310
rect 11566 12246 11630 12310
rect 25846 12246 25910 12310
rect 31014 12382 31078 12446
rect 35774 12382 35838 12446
rect 30742 12246 30806 12310
rect 35638 12246 35702 12310
rect 40806 12382 40870 12446
rect 45838 12382 45902 12446
rect 41078 12246 41142 12310
rect 45838 12246 45902 12310
rect 50734 12382 50798 12446
rect 55766 12382 55830 12446
rect 60798 12382 60862 12446
rect 51006 12246 51070 12310
rect 56038 12246 56102 12310
rect 60662 12246 60726 12310
rect 89766 12246 89830 12310
rect 11566 12110 11630 12174
rect 16598 12110 16662 12174
rect 16598 11838 16662 11902
rect 25982 11838 26046 11902
rect 30878 11838 30942 11902
rect 25710 11702 25774 11766
rect 30878 11702 30942 11766
rect 35910 11838 35974 11902
rect 40942 11838 41006 11902
rect 45702 11838 45766 11902
rect 35774 11702 35838 11766
rect 40806 11702 40870 11766
rect 45702 11702 45766 11766
rect 50870 11838 50934 11902
rect 55902 11838 55966 11902
rect 60934 11838 60998 11902
rect 79974 11838 80038 11902
rect 50734 11702 50798 11766
rect 55766 11702 55830 11766
rect 60798 11702 60862 11766
rect 25846 11566 25910 11630
rect 30742 11566 30806 11630
rect 35638 11566 35702 11630
rect 41078 11566 41142 11630
rect 45838 11566 45902 11630
rect 25166 11158 25230 11222
rect 51006 11566 51070 11630
rect 56038 11566 56102 11630
rect 60662 11566 60726 11630
rect 65422 11430 65486 11494
rect 550 10886 614 10950
rect 11702 10886 11766 10950
rect 25574 10886 25638 10950
rect 25710 10886 25774 10950
rect 30878 10886 30942 10950
rect 35774 10886 35838 10950
rect 40806 10886 40870 10950
rect 45702 10886 45766 10950
rect 50734 10886 50798 10950
rect 55766 10886 55830 10950
rect 60798 10886 60862 10950
rect 65286 10886 65350 10950
rect 11702 10750 11766 10814
rect 1230 10478 1294 10542
rect 17958 10614 18022 10678
rect 16462 10478 16526 10542
rect 25574 10478 25638 10542
rect 65286 10478 65350 10542
rect 79838 10342 79902 10406
rect 89766 10342 89830 10406
rect 2454 9254 2518 9318
rect 11566 9390 11630 9454
rect 25166 9390 25230 9454
rect 65422 9390 65486 9454
rect 16598 9254 16662 9318
rect 16598 9118 16662 9182
rect 1230 8846 1294 8910
rect 2454 8846 2518 8910
rect 89766 8710 89830 8774
rect 2862 8574 2926 8638
rect 2862 8302 2926 8366
rect 550 7894 614 7958
rect 11702 8030 11766 8094
rect 16462 7758 16526 7822
rect 16462 7622 16526 7686
rect 1230 7078 1294 7142
rect 89766 7214 89830 7278
rect 16598 6398 16662 6462
rect 1230 5310 1294 5374
rect 89766 5310 89830 5374
rect 1230 3678 1294 3742
rect 16462 3950 16526 4014
rect 25166 3678 25230 3742
rect 89766 3678 89830 3742
rect 12926 2862 12990 2926
rect 14286 2862 14350 2926
rect 15374 2862 15438 2926
rect 16462 2862 16526 2926
rect 17686 2862 17750 2926
rect 18910 2862 18974 2926
rect 19998 2862 20062 2926
rect 21086 2862 21150 2926
rect 22310 2862 22374 2926
rect 23398 2862 23462 2926
rect 24758 2862 24822 2926
rect 25710 2862 25774 2926
rect 13334 2318 13398 2382
rect 1910 2046 1974 2110
rect 89766 2046 89830 2110
rect 1910 1774 1974 1838
rect 1910 1638 1974 1702
rect 3678 1638 3742 1702
rect 5310 1638 5374 1702
rect 7078 1638 7142 1702
rect 8846 1638 8910 1702
rect 10342 1638 10406 1702
rect 12110 1638 12174 1702
rect 13878 1638 13942 1702
rect 15510 1638 15574 1702
rect 17142 1638 17206 1702
rect 18774 1638 18838 1702
rect 20406 1638 20470 1702
rect 22174 1638 22238 1702
rect 25166 1774 25230 1838
rect 23806 1638 23870 1702
rect 25574 1638 25638 1702
rect 27342 1638 27406 1702
rect 28838 1638 28902 1702
rect 30742 1638 30806 1702
rect 32374 1638 32438 1702
rect 33870 1638 33934 1702
rect 35638 1638 35702 1702
rect 37406 1638 37470 1702
rect 38902 1638 38966 1702
rect 40806 1638 40870 1702
rect 42302 1638 42366 1702
rect 43934 1638 43998 1702
rect 45838 1638 45902 1702
rect 47334 1638 47398 1702
rect 49102 1638 49166 1702
rect 50870 1638 50934 1702
rect 52366 1638 52430 1702
rect 54134 1638 54198 1702
rect 55902 1638 55966 1702
rect 57398 1638 57462 1702
rect 59302 1638 59366 1702
rect 60798 1638 60862 1702
rect 62430 1638 62494 1702
rect 64334 1638 64398 1702
rect 65830 1638 65894 1702
rect 67598 1638 67662 1702
rect 69366 1638 69430 1702
rect 70862 1638 70926 1702
rect 72630 1638 72694 1702
rect 74398 1638 74462 1702
rect 75894 1638 75958 1702
rect 77662 1638 77726 1702
rect 79294 1638 79358 1702
rect 80926 1638 80990 1702
rect 82830 1638 82894 1702
rect 84326 1638 84390 1702
rect 86094 1638 86158 1702
rect 87590 1638 87654 1702
rect 958 1230 1022 1294
rect 1094 1230 1158 1294
rect 1230 1230 1294 1294
rect 1910 1230 1974 1294
rect 3678 1230 3742 1294
rect 5310 1230 5374 1294
rect 7078 1230 7142 1294
rect 8846 1230 8910 1294
rect 10342 1230 10406 1294
rect 12110 1230 12174 1294
rect 13878 1230 13942 1294
rect 15510 1230 15574 1294
rect 17142 1230 17206 1294
rect 18774 1230 18838 1294
rect 20406 1230 20470 1294
rect 22174 1230 22238 1294
rect 23806 1230 23870 1294
rect 25574 1230 25638 1294
rect 27342 1230 27406 1294
rect 28838 1230 28902 1294
rect 30742 1230 30806 1294
rect 32374 1230 32438 1294
rect 33870 1230 33934 1294
rect 35638 1230 35702 1294
rect 37406 1230 37470 1294
rect 38902 1230 38966 1294
rect 40806 1230 40870 1294
rect 42302 1230 42366 1294
rect 43934 1230 43998 1294
rect 45838 1230 45902 1294
rect 47334 1230 47398 1294
rect 49102 1230 49166 1294
rect 50870 1230 50934 1294
rect 52366 1230 52430 1294
rect 54134 1230 54198 1294
rect 55902 1230 55966 1294
rect 57398 1230 57462 1294
rect 59302 1230 59366 1294
rect 60798 1230 60862 1294
rect 62430 1230 62494 1294
rect 64334 1230 64398 1294
rect 65830 1230 65894 1294
rect 67598 1230 67662 1294
rect 69366 1230 69430 1294
rect 70862 1230 70926 1294
rect 72630 1230 72694 1294
rect 74398 1230 74462 1294
rect 75894 1230 75958 1294
rect 77662 1230 77726 1294
rect 79294 1230 79358 1294
rect 80926 1230 80990 1294
rect 82830 1230 82894 1294
rect 84326 1230 84390 1294
rect 86094 1230 86158 1294
rect 87590 1230 87654 1294
rect 89766 1230 89830 1294
rect 89902 1230 89966 1294
rect 90038 1230 90102 1294
rect 958 1094 1022 1158
rect 1094 1094 1158 1158
rect 1230 1094 1294 1158
rect 89766 1094 89830 1158
rect 89902 1094 89966 1158
rect 90038 1094 90102 1158
rect 958 958 1022 1022
rect 1094 958 1158 1022
rect 1230 958 1294 1022
rect 89766 958 89830 1022
rect 89902 958 89966 1022
rect 90038 958 90102 1022
rect 278 550 342 614
rect 414 550 478 614
rect 550 550 614 614
rect 13334 550 13398 614
rect 90446 550 90510 614
rect 90582 550 90646 614
rect 90718 550 90782 614
rect 278 414 342 478
rect 414 414 478 478
rect 550 414 614 478
rect 90446 414 90510 478
rect 90582 414 90646 478
rect 90718 414 90782 478
rect 278 278 342 342
rect 414 278 478 342
rect 550 278 614 342
rect 90446 278 90510 342
rect 90582 278 90646 342
rect 90718 278 90782 342
<< metal4 >>
rect 272 89014 620 89020
rect 272 88950 278 89014
rect 342 88950 414 89014
rect 478 88950 550 89014
rect 614 88950 620 89014
rect 272 88878 620 88950
rect 272 88814 278 88878
rect 342 88814 414 88878
rect 478 88814 550 88878
rect 614 88814 620 88878
rect 272 88742 620 88814
rect 272 88678 278 88742
rect 342 88678 414 88742
rect 478 88678 550 88742
rect 614 88678 620 88742
rect 272 26318 620 88678
rect 272 26254 550 26318
rect 614 26254 620 26318
rect 272 20878 620 26254
rect 272 20814 550 20878
rect 614 20814 620 20878
rect 272 15166 620 20814
rect 272 15102 550 15166
rect 614 15102 620 15166
rect 272 10950 620 15102
rect 272 10886 550 10950
rect 614 10886 620 10950
rect 272 7958 620 10886
rect 272 7894 550 7958
rect 614 7894 620 7958
rect 272 614 620 7894
rect 952 88334 1300 88340
rect 952 88270 958 88334
rect 1022 88270 1094 88334
rect 1158 88270 1230 88334
rect 1294 88270 1300 88334
rect 952 88198 1300 88270
rect 952 88134 958 88198
rect 1022 88134 1094 88198
rect 1158 88134 1230 88198
rect 1294 88134 1300 88198
rect 952 88062 1300 88134
rect 952 87998 958 88062
rect 1022 87998 1094 88062
rect 1158 87998 1230 88062
rect 1294 87998 1300 88062
rect 952 86022 1300 87998
rect 2176 88062 2252 88068
rect 2176 87998 2182 88062
rect 2246 87998 2252 88062
rect 2176 87654 2252 87998
rect 2176 87622 2182 87654
rect 2181 87590 2182 87622
rect 2246 87622 2252 87654
rect 3808 88062 3884 88068
rect 3808 87998 3814 88062
rect 3878 87998 3884 88062
rect 3808 87654 3884 87998
rect 3808 87622 3814 87654
rect 2246 87590 2247 87622
rect 2181 87589 2247 87590
rect 3813 87590 3814 87622
rect 3878 87622 3884 87654
rect 5304 88062 5380 88068
rect 5304 87998 5310 88062
rect 5374 87998 5380 88062
rect 5304 87654 5380 87998
rect 5304 87622 5310 87654
rect 3878 87590 3879 87622
rect 3813 87589 3879 87590
rect 5309 87590 5310 87622
rect 5374 87622 5380 87654
rect 7072 88062 7148 88068
rect 7072 87998 7078 88062
rect 7142 87998 7148 88062
rect 7072 87654 7148 87998
rect 7072 87622 7078 87654
rect 5374 87590 5375 87622
rect 5309 87589 5375 87590
rect 7077 87590 7078 87622
rect 7142 87622 7148 87654
rect 8840 88062 8916 88068
rect 8840 87998 8846 88062
rect 8910 87998 8916 88062
rect 8840 87654 8916 87998
rect 8840 87622 8846 87654
rect 7142 87590 7143 87622
rect 7077 87589 7143 87590
rect 8845 87590 8846 87622
rect 8910 87622 8916 87654
rect 10336 88062 10412 88068
rect 10336 87998 10342 88062
rect 10406 87998 10412 88062
rect 10336 87654 10412 87998
rect 10336 87622 10342 87654
rect 8910 87590 8911 87622
rect 8845 87589 8911 87590
rect 10341 87590 10342 87622
rect 10406 87622 10412 87654
rect 12104 88062 12180 88068
rect 12104 87998 12110 88062
rect 12174 87998 12180 88062
rect 12104 87654 12180 87998
rect 12104 87622 12110 87654
rect 10406 87590 10407 87622
rect 10341 87589 10407 87590
rect 12109 87590 12110 87622
rect 12174 87622 12180 87654
rect 13872 88062 13948 88068
rect 13872 87998 13878 88062
rect 13942 87998 13948 88062
rect 13872 87654 13948 87998
rect 13872 87622 13878 87654
rect 12174 87590 12175 87622
rect 12109 87589 12175 87590
rect 13877 87590 13878 87622
rect 13942 87622 13948 87654
rect 15368 88062 15444 88068
rect 15368 87998 15374 88062
rect 15438 87998 15444 88062
rect 15368 87654 15444 87998
rect 15368 87622 15374 87654
rect 13942 87590 13943 87622
rect 13877 87589 13943 87590
rect 15373 87590 15374 87622
rect 15438 87622 15444 87654
rect 17272 88062 17348 88068
rect 17272 87998 17278 88062
rect 17342 87998 17348 88062
rect 17272 87654 17348 87998
rect 17272 87622 17278 87654
rect 15438 87590 15439 87622
rect 15373 87589 15439 87590
rect 17277 87590 17278 87622
rect 17342 87622 17348 87654
rect 18904 88062 18980 88068
rect 18904 87998 18910 88062
rect 18974 87998 18980 88062
rect 18904 87654 18980 87998
rect 18904 87622 18910 87654
rect 17342 87590 17343 87622
rect 17277 87589 17343 87590
rect 18909 87590 18910 87622
rect 18974 87622 18980 87654
rect 20536 88062 20612 88068
rect 20536 87998 20542 88062
rect 20606 87998 20612 88062
rect 20536 87654 20612 87998
rect 20536 87622 20542 87654
rect 18974 87590 18975 87622
rect 18909 87589 18975 87590
rect 20541 87590 20542 87622
rect 20606 87622 20612 87654
rect 22168 88062 22244 88068
rect 22168 87998 22174 88062
rect 22238 87998 22244 88062
rect 22168 87654 22244 87998
rect 22168 87622 22174 87654
rect 20606 87590 20607 87622
rect 20541 87589 20607 87590
rect 22173 87590 22174 87622
rect 22238 87622 22244 87654
rect 23936 88062 24012 88068
rect 23936 87998 23942 88062
rect 24006 87998 24012 88062
rect 23936 87654 24012 87998
rect 23936 87622 23942 87654
rect 22238 87590 22239 87622
rect 22173 87589 22239 87590
rect 23941 87590 23942 87622
rect 24006 87622 24012 87654
rect 25432 88062 25508 88068
rect 25432 87998 25438 88062
rect 25502 87998 25508 88062
rect 25432 87654 25508 87998
rect 25432 87622 25438 87654
rect 24006 87590 24007 87622
rect 23941 87589 24007 87590
rect 25437 87590 25438 87622
rect 25502 87622 25508 87654
rect 25502 87590 25503 87622
rect 25437 87589 25503 87590
rect 952 85958 1230 86022
rect 1294 85958 1300 86022
rect 952 84390 1300 85958
rect 952 84326 1230 84390
rect 1294 84326 1300 84390
rect 952 82758 1300 84326
rect 952 82694 1230 82758
rect 1294 82694 1300 82758
rect 952 80990 1300 82694
rect 952 80926 1230 80990
rect 1294 80926 1300 80990
rect 952 79358 1300 80926
rect 952 79294 1230 79358
rect 1294 79294 1300 79358
rect 952 77726 1300 79294
rect 25568 77998 25644 89292
rect 27336 88062 27412 88068
rect 27336 87998 27342 88062
rect 27406 87998 27412 88062
rect 27336 87654 27412 87998
rect 27336 87622 27342 87654
rect 27341 87590 27342 87622
rect 27406 87622 27412 87654
rect 28832 88062 28908 88068
rect 28832 87998 28838 88062
rect 28902 87998 28908 88062
rect 28832 87654 28908 87998
rect 28832 87622 28838 87654
rect 27406 87590 27407 87622
rect 27341 87589 27407 87590
rect 28837 87590 28838 87622
rect 28902 87622 28908 87654
rect 30464 88062 30540 88068
rect 30464 87998 30470 88062
rect 30534 87998 30540 88062
rect 30464 87654 30540 87998
rect 30464 87622 30470 87654
rect 28902 87590 28903 87622
rect 28837 87589 28903 87590
rect 30469 87590 30470 87622
rect 30534 87622 30540 87654
rect 30534 87590 30535 87622
rect 30469 87589 30535 87590
rect 25568 77966 25574 77998
rect 25573 77934 25574 77966
rect 25638 77966 25644 77998
rect 30600 77998 30676 89292
rect 32368 88062 32444 88068
rect 32368 87998 32374 88062
rect 32438 87998 32444 88062
rect 32368 87654 32444 87998
rect 32368 87622 32374 87654
rect 32373 87590 32374 87622
rect 32438 87622 32444 87654
rect 33864 88062 33940 88068
rect 33864 87998 33870 88062
rect 33934 87998 33940 88062
rect 33864 87654 33940 87998
rect 33864 87622 33870 87654
rect 32438 87590 32439 87622
rect 32373 87589 32439 87590
rect 33869 87590 33870 87622
rect 33934 87622 33940 87654
rect 33934 87590 33935 87622
rect 33869 87589 33935 87590
rect 30600 77966 30606 77998
rect 25638 77934 25639 77966
rect 25573 77933 25639 77934
rect 30605 77934 30606 77966
rect 30670 77966 30676 77998
rect 35632 77998 35708 89292
rect 35904 88062 35980 88068
rect 35904 87998 35910 88062
rect 35974 87998 35980 88062
rect 35904 87654 35980 87998
rect 35904 87622 35910 87654
rect 35909 87590 35910 87622
rect 35974 87622 35980 87654
rect 37400 88062 37476 88068
rect 37400 87998 37406 88062
rect 37470 87998 37476 88062
rect 37400 87654 37476 87998
rect 37400 87622 37406 87654
rect 35974 87590 35975 87622
rect 35909 87589 35975 87590
rect 37405 87590 37406 87622
rect 37470 87622 37476 87654
rect 39032 88062 39108 88068
rect 39032 87998 39038 88062
rect 39102 87998 39108 88062
rect 39032 87654 39108 87998
rect 39032 87622 39038 87654
rect 37470 87590 37471 87622
rect 37405 87589 37471 87590
rect 39037 87590 39038 87622
rect 39102 87622 39108 87654
rect 39102 87590 39103 87622
rect 39037 87589 39103 87590
rect 35632 77966 35638 77998
rect 30670 77934 30671 77966
rect 30605 77933 30671 77934
rect 35637 77934 35638 77966
rect 35702 77966 35708 77998
rect 40664 77998 40740 89292
rect 40936 88062 41012 88068
rect 40936 87998 40942 88062
rect 41006 87998 41012 88062
rect 40936 87654 41012 87998
rect 40936 87622 40942 87654
rect 40941 87590 40942 87622
rect 41006 87622 41012 87654
rect 42432 88062 42508 88068
rect 42432 87998 42438 88062
rect 42502 87998 42508 88062
rect 42432 87654 42508 87998
rect 42432 87622 42438 87654
rect 41006 87590 41007 87622
rect 40941 87589 41007 87590
rect 42437 87590 42438 87622
rect 42502 87622 42508 87654
rect 43928 88062 44004 88068
rect 43928 87998 43934 88062
rect 43998 87998 44004 88062
rect 43928 87654 44004 87998
rect 43928 87622 43934 87654
rect 42502 87590 42503 87622
rect 42437 87589 42503 87590
rect 43933 87590 43934 87622
rect 43998 87622 44004 87654
rect 43998 87590 43999 87622
rect 43933 87589 43999 87590
rect 40664 77966 40670 77998
rect 35702 77934 35703 77966
rect 35637 77933 35703 77934
rect 40669 77934 40670 77966
rect 40734 77966 40740 77998
rect 45560 77998 45636 89292
rect 45832 88062 45908 88068
rect 45832 87998 45838 88062
rect 45902 87998 45908 88062
rect 45832 87654 45908 87998
rect 45832 87622 45838 87654
rect 45837 87590 45838 87622
rect 45902 87622 45908 87654
rect 47328 88062 47404 88068
rect 47328 87998 47334 88062
rect 47398 87998 47404 88062
rect 47328 87654 47404 87998
rect 47328 87622 47334 87654
rect 45902 87590 45903 87622
rect 45837 87589 45903 87590
rect 47333 87590 47334 87622
rect 47398 87622 47404 87654
rect 49096 88062 49172 88068
rect 49096 87998 49102 88062
rect 49166 87998 49172 88062
rect 49096 87654 49172 87998
rect 49096 87622 49102 87654
rect 47398 87590 47399 87622
rect 47333 87589 47399 87590
rect 49101 87590 49102 87622
rect 49166 87622 49172 87654
rect 49166 87590 49167 87622
rect 49101 87589 49167 87590
rect 45560 77966 45566 77998
rect 40734 77934 40735 77966
rect 40669 77933 40735 77934
rect 45565 77934 45566 77966
rect 45630 77966 45636 77998
rect 50456 77998 50532 89292
rect 50864 88062 50940 88068
rect 50864 87998 50870 88062
rect 50934 87998 50940 88062
rect 50864 87654 50940 87998
rect 50864 87622 50870 87654
rect 50869 87590 50870 87622
rect 50934 87622 50940 87654
rect 52496 88062 52572 88068
rect 52496 87998 52502 88062
rect 52566 87998 52572 88062
rect 52496 87654 52572 87998
rect 52496 87622 52502 87654
rect 50934 87590 50935 87622
rect 50869 87589 50935 87590
rect 52501 87590 52502 87622
rect 52566 87622 52572 87654
rect 54264 88062 54340 88068
rect 54264 87998 54270 88062
rect 54334 87998 54340 88062
rect 54264 87654 54340 87998
rect 54264 87622 54270 87654
rect 52566 87590 52567 87622
rect 52501 87589 52567 87590
rect 54269 87590 54270 87622
rect 54334 87622 54340 87654
rect 54334 87590 54335 87622
rect 54269 87589 54335 87590
rect 50456 77966 50462 77998
rect 45630 77934 45631 77966
rect 45565 77933 45631 77934
rect 50461 77934 50462 77966
rect 50526 77966 50532 77998
rect 55624 77998 55700 89292
rect 55896 88062 55972 88068
rect 55896 87998 55902 88062
rect 55966 87998 55972 88062
rect 55896 87654 55972 87998
rect 55896 87622 55902 87654
rect 55901 87590 55902 87622
rect 55966 87622 55972 87654
rect 57392 88062 57468 88068
rect 57392 87998 57398 88062
rect 57462 87998 57468 88062
rect 57392 87654 57468 87998
rect 57392 87622 57398 87654
rect 55966 87590 55967 87622
rect 55901 87589 55967 87590
rect 57397 87590 57398 87622
rect 57462 87622 57468 87654
rect 59296 88062 59372 88068
rect 59296 87998 59302 88062
rect 59366 87998 59372 88062
rect 59296 87654 59372 87998
rect 59296 87622 59302 87654
rect 57462 87590 57463 87622
rect 57397 87589 57463 87590
rect 59301 87590 59302 87622
rect 59366 87622 59372 87654
rect 59366 87590 59367 87622
rect 59301 87589 59367 87590
rect 55624 77966 55630 77998
rect 50526 77934 50527 77966
rect 50461 77933 50527 77934
rect 55629 77934 55630 77966
rect 55694 77966 55700 77998
rect 60656 77998 60732 89292
rect 73984 88742 74060 88748
rect 73984 88678 73990 88742
rect 74054 88678 74060 88742
rect 60928 88062 61004 88068
rect 60928 87998 60934 88062
rect 60998 87998 61004 88062
rect 60928 87654 61004 87998
rect 60928 87622 60934 87654
rect 60933 87590 60934 87622
rect 60998 87622 61004 87654
rect 62560 88062 62636 88068
rect 62560 87998 62566 88062
rect 62630 87998 62636 88062
rect 62560 87654 62636 87998
rect 62560 87622 62566 87654
rect 60998 87590 60999 87622
rect 60933 87589 60999 87590
rect 62565 87590 62566 87622
rect 62630 87622 62636 87654
rect 64328 88062 64404 88068
rect 64328 87998 64334 88062
rect 64398 87998 64404 88062
rect 64328 87654 64404 87998
rect 64328 87622 64334 87654
rect 62630 87590 62631 87622
rect 62565 87589 62631 87590
rect 64333 87590 64334 87622
rect 64398 87622 64404 87654
rect 65960 88062 66036 88068
rect 65960 87998 65966 88062
rect 66030 87998 66036 88062
rect 65960 87654 66036 87998
rect 65960 87622 65966 87654
rect 64398 87590 64399 87622
rect 64333 87589 64399 87590
rect 65965 87590 65966 87622
rect 66030 87622 66036 87654
rect 67592 88062 67668 88068
rect 67592 87998 67598 88062
rect 67662 87998 67668 88062
rect 67592 87654 67668 87998
rect 67592 87622 67598 87654
rect 66030 87590 66031 87622
rect 65965 87589 66031 87590
rect 67597 87590 67598 87622
rect 67662 87622 67668 87654
rect 69360 88062 69436 88068
rect 69360 87998 69366 88062
rect 69430 87998 69436 88062
rect 69360 87654 69436 87998
rect 69360 87622 69366 87654
rect 67662 87590 67663 87622
rect 67597 87589 67663 87590
rect 69365 87590 69366 87622
rect 69430 87622 69436 87654
rect 70856 88062 70932 88068
rect 70856 87998 70862 88062
rect 70926 87998 70932 88062
rect 70856 87654 70932 87998
rect 70856 87622 70862 87654
rect 69430 87590 69431 87622
rect 69365 87589 69431 87590
rect 70861 87590 70862 87622
rect 70926 87622 70932 87654
rect 72624 88062 72700 88068
rect 72624 87998 72630 88062
rect 72694 87998 72700 88062
rect 72624 87654 72700 87998
rect 72624 87622 72630 87654
rect 70926 87590 70927 87622
rect 70861 87589 70927 87590
rect 72629 87590 72630 87622
rect 72694 87622 72700 87654
rect 72694 87590 72695 87622
rect 72629 87589 72695 87590
rect 73984 86974 74060 88678
rect 74256 88062 74332 88068
rect 74256 87998 74262 88062
rect 74326 87998 74332 88062
rect 74256 87654 74332 87998
rect 74256 87622 74262 87654
rect 74261 87590 74262 87622
rect 74326 87622 74332 87654
rect 74326 87590 74327 87622
rect 74261 87589 74327 87590
rect 73984 86942 73990 86974
rect 73989 86910 73990 86942
rect 74054 86942 74060 86974
rect 74054 86910 74055 86942
rect 73989 86909 74055 86910
rect 74261 86838 74327 86839
rect 74261 86806 74262 86838
rect 74256 86774 74262 86806
rect 74326 86806 74327 86838
rect 74326 86774 74332 86806
rect 74125 85342 74191 85343
rect 74125 85310 74126 85342
rect 74120 85278 74126 85310
rect 74190 85310 74191 85342
rect 74190 85278 74196 85310
rect 74120 83302 74196 85278
rect 74256 84798 74332 86774
rect 74528 86294 74604 89292
rect 74528 86262 74534 86294
rect 74533 86230 74534 86262
rect 74598 86262 74604 86294
rect 75616 86294 75692 89292
rect 76024 88062 76100 88068
rect 76024 87998 76030 88062
rect 76094 87998 76100 88062
rect 76024 87654 76100 87998
rect 76024 87622 76030 87654
rect 76029 87590 76030 87622
rect 76094 87622 76100 87654
rect 76094 87590 76095 87622
rect 76029 87589 76095 87590
rect 76301 87382 76367 87383
rect 76301 87350 76302 87382
rect 75616 86262 75622 86294
rect 74598 86230 74599 86262
rect 74533 86229 74599 86230
rect 75621 86230 75622 86262
rect 75686 86262 75692 86294
rect 76296 87318 76302 87350
rect 76366 87350 76367 87382
rect 76366 87318 76372 87350
rect 75686 86230 75687 86262
rect 75621 86229 75687 86230
rect 76296 85478 76372 87318
rect 76704 86294 76780 89292
rect 90440 89014 90788 89020
rect 90440 88950 90446 89014
rect 90510 88950 90582 89014
rect 90646 88950 90718 89014
rect 90782 88950 90788 89014
rect 90440 88878 90788 88950
rect 90440 88814 90446 88878
rect 90510 88814 90582 88878
rect 90646 88814 90718 88878
rect 90782 88814 90788 88878
rect 90440 88742 90788 88814
rect 90440 88678 90446 88742
rect 90510 88678 90582 88742
rect 90646 88678 90718 88742
rect 90782 88678 90788 88742
rect 89760 88334 90108 88340
rect 89760 88270 89766 88334
rect 89830 88270 89902 88334
rect 89966 88270 90038 88334
rect 90102 88270 90108 88334
rect 89760 88198 90108 88270
rect 89760 88134 89766 88198
rect 89830 88134 89902 88198
rect 89966 88134 90038 88198
rect 90102 88134 90108 88198
rect 77656 88062 77732 88068
rect 77656 87998 77662 88062
rect 77726 87998 77732 88062
rect 77656 87654 77732 87998
rect 77656 87622 77662 87654
rect 77661 87590 77662 87622
rect 77726 87622 77732 87654
rect 79424 88062 79500 88068
rect 79424 87998 79430 88062
rect 79494 87998 79500 88062
rect 79424 87654 79500 87998
rect 79424 87622 79430 87654
rect 77726 87590 77727 87622
rect 77661 87589 77727 87590
rect 79429 87590 79430 87622
rect 79494 87622 79500 87654
rect 81056 88062 81132 88068
rect 81056 87998 81062 88062
rect 81126 87998 81132 88062
rect 81056 87654 81132 87998
rect 81056 87622 81062 87654
rect 79494 87590 79495 87622
rect 79429 87589 79495 87590
rect 81061 87590 81062 87622
rect 81126 87622 81132 87654
rect 82552 88062 82628 88068
rect 82552 87998 82558 88062
rect 82622 87998 82628 88062
rect 82552 87654 82628 87998
rect 82552 87622 82558 87654
rect 81126 87590 81127 87622
rect 81061 87589 81127 87590
rect 82557 87590 82558 87622
rect 82622 87622 82628 87654
rect 84320 88062 84396 88068
rect 84320 87998 84326 88062
rect 84390 87998 84396 88062
rect 84320 87654 84396 87998
rect 84320 87622 84326 87654
rect 82622 87590 82623 87622
rect 82557 87589 82623 87590
rect 84325 87590 84326 87622
rect 84390 87622 84396 87654
rect 86088 88062 86164 88068
rect 86088 87998 86094 88062
rect 86158 87998 86164 88062
rect 86088 87654 86164 87998
rect 86088 87622 86094 87654
rect 84390 87590 84391 87622
rect 84325 87589 84391 87590
rect 86093 87590 86094 87622
rect 86158 87622 86164 87654
rect 87856 88062 87932 88068
rect 87856 87998 87862 88062
rect 87926 87998 87932 88062
rect 87856 87654 87932 87998
rect 87856 87622 87862 87654
rect 86158 87590 86159 87622
rect 86093 87589 86159 87590
rect 87861 87590 87862 87622
rect 87926 87622 87932 87654
rect 89760 88062 90108 88134
rect 89760 87998 89766 88062
rect 89830 87998 89902 88062
rect 89966 87998 90038 88062
rect 90102 87998 90108 88062
rect 87926 87590 87927 87622
rect 87861 87589 87927 87590
rect 76704 86262 76710 86294
rect 76709 86230 76710 86262
rect 76774 86262 76780 86294
rect 76774 86230 76775 86262
rect 76709 86229 76775 86230
rect 76296 85414 76302 85478
rect 76366 85414 76372 85478
rect 76296 85408 76372 85414
rect 89760 86022 90108 87998
rect 89760 85958 89766 86022
rect 89830 85958 90108 86022
rect 74256 84734 74262 84798
rect 74326 84734 74332 84798
rect 74256 84728 74332 84734
rect 74120 83238 74126 83302
rect 74190 83238 74196 83302
rect 74120 83232 74196 83238
rect 74392 84662 74468 84668
rect 74392 84598 74398 84662
rect 74462 84598 74468 84662
rect 74256 83166 74332 83172
rect 74256 83102 74262 83166
rect 74326 83102 74332 83166
rect 74120 81806 74196 81812
rect 74120 81742 74126 81806
rect 74190 81742 74196 81806
rect 74120 79086 74196 81742
rect 74256 80446 74332 83102
rect 74392 81942 74468 84598
rect 74392 81910 74398 81942
rect 74397 81878 74398 81910
rect 74462 81910 74468 81942
rect 89760 84390 90108 85958
rect 89760 84326 89766 84390
rect 89830 84326 90108 84390
rect 89760 82758 90108 84326
rect 89760 82694 89766 82758
rect 89830 82694 90108 82758
rect 74462 81878 74463 81910
rect 74397 81877 74463 81878
rect 74256 80414 74262 80446
rect 74261 80382 74262 80414
rect 74326 80414 74332 80446
rect 89760 80990 90108 82694
rect 89760 80926 89766 80990
rect 89830 80926 90108 80990
rect 74326 80382 74327 80414
rect 74261 80381 74327 80382
rect 74261 80310 74327 80311
rect 74261 80278 74262 80310
rect 74120 79054 74126 79086
rect 74125 79022 74126 79054
rect 74190 79054 74196 79086
rect 74256 80246 74262 80278
rect 74326 80278 74327 80310
rect 74326 80246 74332 80278
rect 74190 79022 74191 79054
rect 74125 79021 74191 79022
rect 60656 77966 60662 77998
rect 55694 77934 55695 77966
rect 55629 77933 55695 77934
rect 60661 77934 60662 77966
rect 60726 77966 60732 77998
rect 74120 78950 74196 78956
rect 74120 78886 74126 78950
rect 74190 78886 74196 78950
rect 60726 77934 60727 77966
rect 60661 77933 60727 77934
rect 25981 77862 26047 77863
rect 25981 77830 25982 77862
rect 952 77662 1230 77726
rect 1294 77662 1300 77726
rect 952 75958 1300 77662
rect 25976 77798 25982 77830
rect 26046 77830 26047 77862
rect 30877 77862 30943 77863
rect 30877 77830 30878 77862
rect 26046 77798 26052 77830
rect 25840 77590 25916 77596
rect 25840 77526 25846 77590
rect 25910 77526 25916 77590
rect 25840 76910 25916 77526
rect 25840 76878 25846 76910
rect 25845 76846 25846 76878
rect 25910 76878 25916 76910
rect 25910 76846 25911 76878
rect 25845 76845 25911 76846
rect 952 75894 1230 75958
rect 1294 75894 1300 75958
rect 952 74326 1300 75894
rect 952 74262 1230 74326
rect 1294 74262 1300 74326
rect 952 72694 1300 74262
rect 952 72630 1230 72694
rect 1294 72630 1300 72694
rect 952 71062 1300 72630
rect 25840 76638 25916 76644
rect 25840 76574 25846 76638
rect 25910 76574 25916 76638
rect 25840 72014 25916 76574
rect 25976 76094 26052 77798
rect 30872 77798 30878 77830
rect 30942 77830 30943 77862
rect 35909 77862 35975 77863
rect 35909 77830 35910 77862
rect 30942 77798 30948 77830
rect 30736 77590 30812 77596
rect 30736 77526 30742 77590
rect 30806 77526 30812 77590
rect 30736 76910 30812 77526
rect 30736 76878 30742 76910
rect 30741 76846 30742 76878
rect 30806 76878 30812 76910
rect 30806 76846 30807 76878
rect 30741 76845 30807 76846
rect 30328 76638 30404 76644
rect 30328 76574 30334 76638
rect 30398 76574 30404 76638
rect 25976 76030 25982 76094
rect 26046 76030 26052 76094
rect 26117 76094 26183 76095
rect 26117 76062 26118 76094
rect 25976 76024 26052 76030
rect 26112 76030 26118 76062
rect 26182 76062 26183 76094
rect 26182 76030 26188 76062
rect 26112 73646 26188 76030
rect 26112 73582 26118 73646
rect 26182 73582 26188 73646
rect 26112 73576 26188 73582
rect 25840 71982 25846 72014
rect 25845 71950 25846 71982
rect 25910 71982 25916 72014
rect 25976 73374 26052 73380
rect 25976 73310 25982 73374
rect 26046 73310 26052 73374
rect 25910 71950 25911 71982
rect 25845 71949 25911 71950
rect 25568 71878 25644 71884
rect 25568 71814 25574 71878
rect 25638 71814 25644 71878
rect 25568 71470 25644 71814
rect 25568 71438 25574 71470
rect 25573 71406 25574 71438
rect 25638 71438 25644 71470
rect 25638 71406 25639 71438
rect 25573 71405 25639 71406
rect 952 70998 1230 71062
rect 1294 70998 1300 71062
rect 952 69294 1300 70998
rect 25976 70926 26052 73310
rect 30328 72014 30404 76574
rect 30872 76094 30948 77798
rect 35904 77798 35910 77830
rect 35974 77830 35975 77862
rect 41077 77862 41143 77863
rect 41077 77830 41078 77862
rect 35974 77798 35980 77830
rect 35768 77590 35844 77596
rect 35768 77526 35774 77590
rect 35838 77526 35844 77590
rect 35768 76910 35844 77526
rect 35768 76878 35774 76910
rect 35773 76846 35774 76878
rect 35838 76878 35844 76910
rect 35838 76846 35839 76878
rect 35773 76845 35839 76846
rect 30872 76030 30878 76094
rect 30942 76030 30948 76094
rect 31013 76094 31079 76095
rect 31013 76062 31014 76094
rect 30872 76024 30948 76030
rect 31008 76030 31014 76062
rect 31078 76062 31079 76094
rect 35904 76094 35980 77798
rect 41072 77798 41078 77830
rect 41142 77830 41143 77862
rect 45973 77862 46039 77863
rect 45973 77830 45974 77862
rect 41142 77798 41148 77830
rect 40936 77590 41012 77596
rect 40936 77526 40942 77590
rect 41006 77526 41012 77590
rect 40936 76910 41012 77526
rect 40936 76878 40942 76910
rect 40941 76846 40942 76878
rect 41006 76878 41012 76910
rect 41006 76846 41007 76878
rect 40941 76845 41007 76846
rect 36861 76638 36927 76639
rect 36861 76606 36862 76638
rect 36856 76574 36862 76606
rect 36926 76606 36927 76638
rect 40800 76638 40876 76644
rect 36926 76574 36932 76606
rect 31078 76030 31084 76062
rect 31008 73646 31084 76030
rect 35904 76030 35910 76094
rect 35974 76030 35980 76094
rect 36045 76094 36111 76095
rect 36045 76062 36046 76094
rect 35904 76024 35980 76030
rect 36040 76030 36046 76062
rect 36110 76062 36111 76094
rect 36110 76030 36116 76062
rect 31008 73582 31014 73646
rect 31078 73582 31084 73646
rect 31008 73576 31084 73582
rect 36040 73646 36116 76030
rect 36040 73582 36046 73646
rect 36110 73582 36116 73646
rect 36040 73576 36116 73582
rect 30328 71982 30334 72014
rect 30333 71950 30334 71982
rect 30398 71982 30404 72014
rect 36856 72014 36932 76574
rect 30398 71950 30399 71982
rect 30333 71949 30399 71950
rect 36856 71950 36862 72014
rect 36926 71950 36932 72014
rect 40800 76574 40806 76638
rect 40870 76574 40876 76638
rect 40800 72014 40876 76574
rect 40941 76094 41007 76095
rect 40941 76062 40942 76094
rect 40936 76030 40942 76062
rect 41006 76062 41007 76094
rect 41072 76094 41148 77798
rect 45968 77798 45974 77830
rect 46038 77830 46039 77862
rect 50869 77862 50935 77863
rect 50869 77830 50870 77862
rect 46038 77798 46044 77830
rect 45832 77590 45908 77596
rect 45832 77526 45838 77590
rect 45902 77526 45908 77590
rect 45832 76910 45908 77526
rect 45832 76878 45838 76910
rect 45837 76846 45838 76878
rect 45902 76878 45908 76910
rect 45902 76846 45903 76878
rect 45837 76845 45903 76846
rect 41006 76030 41012 76062
rect 40936 73652 41012 76030
rect 41072 76030 41078 76094
rect 41142 76030 41148 76094
rect 41072 76024 41148 76030
rect 45696 76638 45772 76644
rect 45696 76574 45702 76638
rect 45766 76574 45772 76638
rect 40936 73646 41148 73652
rect 40936 73582 41078 73646
rect 41142 73582 41148 73646
rect 40936 73576 41148 73582
rect 40800 71982 40806 72014
rect 36856 71944 36932 71950
rect 40805 71950 40806 71982
rect 40870 71982 40876 72014
rect 45696 72014 45772 76574
rect 45968 76094 46044 77798
rect 50864 77798 50870 77830
rect 50934 77830 50935 77862
rect 56037 77862 56103 77863
rect 56037 77830 56038 77862
rect 50934 77798 50940 77830
rect 50728 77590 50804 77596
rect 50728 77526 50734 77590
rect 50798 77526 50804 77590
rect 50728 76910 50804 77526
rect 50728 76878 50734 76910
rect 50733 76846 50734 76878
rect 50798 76878 50804 76910
rect 50798 76846 50799 76878
rect 50733 76845 50799 76846
rect 50728 76638 50804 76644
rect 50728 76574 50734 76638
rect 50798 76574 50804 76638
rect 45968 76030 45974 76094
rect 46038 76030 46044 76094
rect 46109 76094 46175 76095
rect 46109 76062 46110 76094
rect 45968 76024 46044 76030
rect 46104 76030 46110 76062
rect 46174 76062 46175 76094
rect 46174 76030 46180 76062
rect 46104 73646 46180 76030
rect 46104 73582 46110 73646
rect 46174 73582 46180 73646
rect 46104 73576 46180 73582
rect 45696 71982 45702 72014
rect 40870 71950 40871 71982
rect 40805 71949 40871 71950
rect 45701 71950 45702 71982
rect 45766 71982 45772 72014
rect 50728 72014 50804 76574
rect 50864 76094 50940 77798
rect 56032 77798 56038 77830
rect 56102 77830 56103 77862
rect 60933 77862 60999 77863
rect 60933 77830 60934 77862
rect 56102 77798 56108 77830
rect 55896 77590 55972 77596
rect 55896 77526 55902 77590
rect 55966 77526 55972 77590
rect 55896 76910 55972 77526
rect 55896 76878 55902 76910
rect 55901 76846 55902 76878
rect 55966 76878 55972 76910
rect 55966 76846 55967 76878
rect 55901 76845 55967 76846
rect 55352 76638 55428 76644
rect 55352 76574 55358 76638
rect 55422 76574 55428 76638
rect 50864 76030 50870 76094
rect 50934 76030 50940 76094
rect 51005 76094 51071 76095
rect 51005 76062 51006 76094
rect 50864 76024 50940 76030
rect 51000 76030 51006 76062
rect 51070 76062 51071 76094
rect 51070 76030 51076 76062
rect 51000 73646 51076 76030
rect 51000 73582 51006 73646
rect 51070 73582 51076 73646
rect 51000 73576 51076 73582
rect 50728 71982 50734 72014
rect 45766 71950 45767 71982
rect 45701 71949 45767 71950
rect 50733 71950 50734 71982
rect 50798 71982 50804 72014
rect 55352 72014 55428 76574
rect 56032 76094 56108 77798
rect 60928 77798 60934 77830
rect 60998 77830 60999 77862
rect 60998 77798 61004 77830
rect 60928 77732 61004 77798
rect 60792 77656 61004 77732
rect 56032 76030 56038 76094
rect 56102 76030 56108 76094
rect 56173 76094 56239 76095
rect 56173 76062 56174 76094
rect 56032 76024 56108 76030
rect 56168 76030 56174 76062
rect 56238 76062 56239 76094
rect 60792 76094 60868 77656
rect 60928 77590 61004 77596
rect 60928 77526 60934 77590
rect 60998 77526 61004 77590
rect 72901 77590 72967 77591
rect 72901 77558 72902 77590
rect 60928 76910 61004 77526
rect 60928 76878 60934 76910
rect 60933 76846 60934 76878
rect 60998 76878 61004 76910
rect 72896 77526 72902 77558
rect 72966 77558 72967 77590
rect 72966 77526 72972 77558
rect 60998 76846 60999 76878
rect 60933 76845 60999 76846
rect 61477 76638 61543 76639
rect 61477 76606 61478 76638
rect 61472 76574 61478 76606
rect 61542 76606 61543 76638
rect 61542 76574 61548 76606
rect 56238 76030 56244 76062
rect 56168 73646 56244 76030
rect 60792 76030 60798 76094
rect 60862 76030 60868 76094
rect 60933 76094 60999 76095
rect 60933 76062 60934 76094
rect 60792 76024 60868 76030
rect 60928 76030 60934 76062
rect 60998 76062 60999 76094
rect 60998 76030 61004 76062
rect 56168 73582 56174 73646
rect 56238 73582 56244 73646
rect 56168 73576 56244 73582
rect 60928 73646 61004 76030
rect 60928 73582 60934 73646
rect 60998 73582 61004 73646
rect 60928 73576 61004 73582
rect 55352 71982 55358 72014
rect 50798 71950 50799 71982
rect 50733 71949 50799 71950
rect 55357 71950 55358 71982
rect 55422 71982 55428 72014
rect 61472 72014 61548 76574
rect 72629 76094 72695 76095
rect 72629 76062 72630 76094
rect 72624 76030 72630 76062
rect 72694 76062 72695 76094
rect 72694 76030 72700 76062
rect 72624 73510 72700 76030
rect 72896 74870 72972 77526
rect 74120 76230 74196 78886
rect 74256 77726 74332 80246
rect 79293 80174 79359 80175
rect 79293 80142 79294 80174
rect 74256 77662 74262 77726
rect 74326 77662 74332 77726
rect 74256 77656 74332 77662
rect 79288 80110 79294 80142
rect 79358 80142 79359 80174
rect 79358 80110 79364 80142
rect 79288 77454 79364 80110
rect 87997 79494 88063 79495
rect 87997 79462 87998 79494
rect 87992 79430 87998 79462
rect 88062 79462 88063 79494
rect 88062 79430 88068 79462
rect 87992 79222 88068 79430
rect 87992 79158 87998 79222
rect 88062 79158 88068 79222
rect 87992 79152 88068 79158
rect 89080 79358 89156 79364
rect 89080 79294 89086 79358
rect 89150 79294 89156 79358
rect 89080 78814 89156 79294
rect 89080 78782 89086 78814
rect 89085 78750 89086 78782
rect 89150 78782 89156 78814
rect 89760 79358 90108 80926
rect 89760 79294 89766 79358
rect 89830 79294 90108 79358
rect 89150 78750 89151 78782
rect 89085 78749 89151 78750
rect 79565 78678 79631 78679
rect 79565 78646 79566 78678
rect 79288 77390 79294 77454
rect 79358 77390 79364 77454
rect 79288 77384 79364 77390
rect 79560 78614 79566 78646
rect 79630 78646 79631 78678
rect 79630 78614 79636 78646
rect 74120 76198 74126 76230
rect 74125 76166 74126 76198
rect 74190 76198 74196 76230
rect 79288 77318 79364 77324
rect 79288 77254 79294 77318
rect 79358 77254 79364 77318
rect 79288 76230 79364 77254
rect 79288 76198 79294 76230
rect 74190 76166 74191 76198
rect 74125 76165 74191 76166
rect 79293 76166 79294 76198
rect 79358 76198 79364 76230
rect 79424 77318 79500 77324
rect 79424 77254 79430 77318
rect 79494 77254 79500 77318
rect 79358 76166 79359 76198
rect 79293 76165 79359 76166
rect 72896 74806 72902 74870
rect 72966 74806 72972 74870
rect 79288 75822 79364 75828
rect 79288 75758 79294 75822
rect 79358 75758 79364 75822
rect 79288 74870 79364 75758
rect 79288 74838 79294 74870
rect 72896 74800 72972 74806
rect 79293 74806 79294 74838
rect 79358 74838 79364 74870
rect 79358 74806 79359 74838
rect 79293 74805 79359 74806
rect 72624 73446 72630 73510
rect 72694 73446 72700 73510
rect 72624 73440 72700 73446
rect 72760 74734 72836 74740
rect 72760 74670 72766 74734
rect 72830 74670 72836 74734
rect 66781 73374 66847 73375
rect 66781 73342 66782 73374
rect 55422 71950 55423 71982
rect 55357 71949 55423 71950
rect 61472 71950 61478 72014
rect 61542 71950 61548 72014
rect 61472 71944 61548 71950
rect 66776 73310 66782 73342
rect 66846 73342 66847 73374
rect 66846 73310 66852 73342
rect 26792 71878 26868 71884
rect 26792 71814 26798 71878
rect 26862 71814 26868 71878
rect 27613 71878 27679 71879
rect 27613 71846 27614 71878
rect 26792 71470 26868 71814
rect 26792 71438 26798 71470
rect 26797 71406 26798 71438
rect 26862 71438 26868 71470
rect 27608 71814 27614 71846
rect 27678 71846 27679 71878
rect 27744 71878 27820 71884
rect 27678 71814 27684 71846
rect 27608 71470 27684 71814
rect 26862 71406 26863 71438
rect 26797 71405 26863 71406
rect 27608 71406 27614 71470
rect 27678 71406 27684 71470
rect 27744 71814 27750 71878
rect 27814 71814 27820 71878
rect 27744 71470 27820 71814
rect 27744 71438 27750 71470
rect 27608 71400 27684 71406
rect 27749 71406 27750 71438
rect 27814 71438 27820 71470
rect 28968 71878 29044 71884
rect 28968 71814 28974 71878
rect 29038 71814 29044 71878
rect 29517 71878 29583 71879
rect 29517 71846 29518 71878
rect 28968 71470 29044 71814
rect 28968 71438 28974 71470
rect 27814 71406 27815 71438
rect 27749 71405 27815 71406
rect 28973 71406 28974 71438
rect 29038 71438 29044 71470
rect 29512 71814 29518 71846
rect 29582 71846 29583 71878
rect 30741 71878 30807 71879
rect 30741 71846 30742 71878
rect 29582 71814 29588 71846
rect 29512 71470 29588 71814
rect 29038 71406 29039 71438
rect 28973 71405 29039 71406
rect 29512 71406 29518 71470
rect 29582 71406 29588 71470
rect 29512 71400 29588 71406
rect 30736 71814 30742 71846
rect 30806 71846 30807 71878
rect 31416 71878 31492 71884
rect 30806 71814 30812 71846
rect 30736 71470 30812 71814
rect 30736 71406 30742 71470
rect 30806 71406 30812 71470
rect 31416 71814 31422 71878
rect 31486 71814 31492 71878
rect 31965 71878 32031 71879
rect 31965 71846 31966 71878
rect 31416 71470 31492 71814
rect 31416 71438 31422 71470
rect 30736 71400 30812 71406
rect 31421 71406 31422 71438
rect 31486 71438 31492 71470
rect 31960 71814 31966 71846
rect 32030 71846 32031 71878
rect 32504 71878 32580 71884
rect 32030 71814 32036 71846
rect 31960 71470 32036 71814
rect 31486 71406 31487 71438
rect 31421 71405 31487 71406
rect 31960 71406 31966 71470
rect 32030 71406 32036 71470
rect 32504 71814 32510 71878
rect 32574 71814 32580 71878
rect 32504 71470 32580 71814
rect 32504 71438 32510 71470
rect 31960 71400 32036 71406
rect 32509 71406 32510 71438
rect 32574 71438 32580 71470
rect 33048 71878 33124 71884
rect 33048 71814 33054 71878
rect 33118 71814 33124 71878
rect 33048 71470 33124 71814
rect 33048 71438 33054 71470
rect 32574 71406 32575 71438
rect 32509 71405 32575 71406
rect 33053 71406 33054 71438
rect 33118 71438 33124 71470
rect 34000 71878 34076 71884
rect 34000 71814 34006 71878
rect 34070 71814 34076 71878
rect 34413 71878 34479 71879
rect 34413 71846 34414 71878
rect 34000 71470 34076 71814
rect 34000 71438 34006 71470
rect 33118 71406 33119 71438
rect 33053 71405 33119 71406
rect 34005 71406 34006 71438
rect 34070 71438 34076 71470
rect 34408 71814 34414 71846
rect 34478 71846 34479 71878
rect 35224 71878 35300 71884
rect 34478 71814 34484 71846
rect 34408 71470 34484 71814
rect 34070 71406 34071 71438
rect 34005 71405 34071 71406
rect 34408 71406 34414 71470
rect 34478 71406 34484 71470
rect 35224 71814 35230 71878
rect 35294 71814 35300 71878
rect 35773 71878 35839 71879
rect 35773 71846 35774 71878
rect 35224 71470 35300 71814
rect 35224 71438 35230 71470
rect 34408 71400 34484 71406
rect 35229 71406 35230 71438
rect 35294 71438 35300 71470
rect 35768 71814 35774 71846
rect 35838 71846 35839 71878
rect 36448 71878 36524 71884
rect 35838 71814 35844 71846
rect 35768 71470 35844 71814
rect 35294 71406 35295 71438
rect 35229 71405 35295 71406
rect 35768 71406 35774 71470
rect 35838 71406 35844 71470
rect 36448 71814 36454 71878
rect 36518 71814 36524 71878
rect 36997 71878 37063 71879
rect 36997 71846 36998 71878
rect 36448 71470 36524 71814
rect 36448 71438 36454 71470
rect 35768 71400 35844 71406
rect 36453 71406 36454 71438
rect 36518 71438 36524 71470
rect 36992 71814 36998 71846
rect 37062 71846 37063 71878
rect 37672 71878 37748 71884
rect 37062 71814 37068 71846
rect 36992 71470 37068 71814
rect 36518 71406 36519 71438
rect 36453 71405 36519 71406
rect 36992 71406 36998 71470
rect 37062 71406 37068 71470
rect 37672 71814 37678 71878
rect 37742 71814 37748 71878
rect 38221 71878 38287 71879
rect 38221 71846 38222 71878
rect 37672 71470 37748 71814
rect 37672 71438 37678 71470
rect 36992 71400 37068 71406
rect 37677 71406 37678 71438
rect 37742 71438 37748 71470
rect 38216 71814 38222 71846
rect 38286 71846 38287 71878
rect 39445 71878 39511 71879
rect 39445 71846 39446 71878
rect 38286 71814 38292 71846
rect 38216 71470 38292 71814
rect 37742 71406 37743 71438
rect 37677 71405 37743 71406
rect 38216 71406 38222 71470
rect 38286 71406 38292 71470
rect 38216 71400 38292 71406
rect 39440 71814 39446 71846
rect 39510 71846 39511 71878
rect 40256 71878 40332 71884
rect 39510 71814 39516 71846
rect 39440 71470 39516 71814
rect 39440 71406 39446 71470
rect 39510 71406 39516 71470
rect 40256 71814 40262 71878
rect 40326 71814 40332 71878
rect 40669 71878 40735 71879
rect 40669 71846 40670 71878
rect 40256 71470 40332 71814
rect 40256 71438 40262 71470
rect 39440 71400 39516 71406
rect 40261 71406 40262 71438
rect 40326 71438 40332 71470
rect 40664 71814 40670 71846
rect 40734 71846 40735 71878
rect 41621 71878 41687 71879
rect 41621 71846 41622 71878
rect 40734 71814 40740 71846
rect 40664 71470 40740 71814
rect 40326 71406 40327 71438
rect 40261 71405 40327 71406
rect 40664 71406 40670 71470
rect 40734 71406 40740 71470
rect 40664 71400 40740 71406
rect 41616 71814 41622 71846
rect 41686 71846 41687 71878
rect 42704 71878 42780 71884
rect 41686 71814 41692 71846
rect 41616 71334 41692 71814
rect 42704 71814 42710 71878
rect 42774 71814 42780 71878
rect 43253 71878 43319 71879
rect 43253 71846 43254 71878
rect 42704 71470 42780 71814
rect 42704 71438 42710 71470
rect 42709 71406 42710 71438
rect 42774 71438 42780 71470
rect 43248 71814 43254 71846
rect 43318 71846 43319 71878
rect 43928 71878 44004 71884
rect 43318 71814 43324 71846
rect 43248 71470 43324 71814
rect 42774 71406 42775 71438
rect 42709 71405 42775 71406
rect 43248 71406 43254 71470
rect 43318 71406 43324 71470
rect 43928 71814 43934 71878
rect 43998 71814 44004 71878
rect 43928 71470 44004 71814
rect 43928 71438 43934 71470
rect 43248 71400 43324 71406
rect 43933 71406 43934 71438
rect 43998 71438 44004 71470
rect 45152 71878 45228 71884
rect 45152 71814 45158 71878
rect 45222 71814 45228 71878
rect 45701 71878 45767 71879
rect 45701 71846 45702 71878
rect 45152 71470 45228 71814
rect 45152 71438 45158 71470
rect 43998 71406 43999 71438
rect 43933 71405 43999 71406
rect 45157 71406 45158 71438
rect 45222 71438 45228 71470
rect 45696 71814 45702 71846
rect 45766 71846 45767 71878
rect 46925 71878 46991 71879
rect 46925 71846 46926 71878
rect 45766 71814 45772 71846
rect 45696 71470 45772 71814
rect 45222 71406 45223 71438
rect 45157 71405 45223 71406
rect 45696 71406 45702 71470
rect 45766 71406 45772 71470
rect 45696 71400 45772 71406
rect 46920 71814 46926 71846
rect 46990 71846 46991 71878
rect 47736 71878 47812 71884
rect 46990 71814 46996 71846
rect 46920 71470 46996 71814
rect 46920 71406 46926 71470
rect 46990 71406 46996 71470
rect 47736 71814 47742 71878
rect 47806 71814 47812 71878
rect 47736 71470 47812 71814
rect 47736 71438 47742 71470
rect 46920 71400 46996 71406
rect 47741 71406 47742 71438
rect 47806 71438 47812 71470
rect 48960 71878 49036 71884
rect 48960 71814 48966 71878
rect 49030 71814 49036 71878
rect 49373 71878 49439 71879
rect 49373 71846 49374 71878
rect 48960 71470 49036 71814
rect 48960 71438 48966 71470
rect 47806 71406 47807 71438
rect 47741 71405 47807 71406
rect 48965 71406 48966 71438
rect 49030 71438 49036 71470
rect 49368 71814 49374 71846
rect 49438 71846 49439 71878
rect 50184 71878 50260 71884
rect 49438 71814 49444 71846
rect 49368 71470 49444 71814
rect 49030 71406 49031 71438
rect 48965 71405 49031 71406
rect 49368 71406 49374 71470
rect 49438 71406 49444 71470
rect 50184 71814 50190 71878
rect 50254 71814 50260 71878
rect 50184 71470 50260 71814
rect 50184 71438 50190 71470
rect 49368 71400 49444 71406
rect 50189 71406 50190 71438
rect 50254 71438 50260 71470
rect 51408 71878 51484 71884
rect 51408 71814 51414 71878
rect 51478 71814 51484 71878
rect 51957 71878 52023 71879
rect 51957 71846 51958 71878
rect 51408 71470 51484 71814
rect 51408 71438 51414 71470
rect 50254 71406 50255 71438
rect 50189 71405 50255 71406
rect 51413 71406 51414 71438
rect 51478 71438 51484 71470
rect 51952 71814 51958 71846
rect 52022 71846 52023 71878
rect 52632 71878 52708 71884
rect 52022 71814 52028 71846
rect 51952 71470 52028 71814
rect 51478 71406 51479 71438
rect 51413 71405 51479 71406
rect 51952 71406 51958 71470
rect 52022 71406 52028 71470
rect 52632 71814 52638 71878
rect 52702 71814 52708 71878
rect 54133 71878 54199 71879
rect 54133 71846 54134 71878
rect 52632 71470 52708 71814
rect 52632 71438 52638 71470
rect 51952 71400 52028 71406
rect 52637 71406 52638 71438
rect 52702 71438 52708 71470
rect 54128 71814 54134 71846
rect 54198 71846 54199 71878
rect 55765 71878 55831 71879
rect 55765 71846 55766 71878
rect 54198 71814 54204 71846
rect 52702 71406 52703 71438
rect 52637 71405 52703 71406
rect 41616 71270 41622 71334
rect 41686 71270 41692 71334
rect 41616 71264 41692 71270
rect 54128 71334 54204 71814
rect 55760 71814 55766 71846
rect 55830 71846 55831 71878
rect 56440 71878 56516 71884
rect 55830 71814 55836 71846
rect 55760 71470 55836 71814
rect 55760 71406 55766 71470
rect 55830 71406 55836 71470
rect 56440 71814 56446 71878
rect 56510 71814 56516 71878
rect 56989 71878 57055 71879
rect 56989 71846 56990 71878
rect 56440 71470 56516 71814
rect 56440 71438 56446 71470
rect 55760 71400 55836 71406
rect 56445 71406 56446 71438
rect 56510 71438 56516 71470
rect 56984 71814 56990 71846
rect 57054 71846 57055 71878
rect 57664 71878 57740 71884
rect 57054 71814 57060 71846
rect 56984 71470 57060 71814
rect 56510 71406 56511 71438
rect 56445 71405 56511 71406
rect 56984 71406 56990 71470
rect 57054 71406 57060 71470
rect 57664 71814 57670 71878
rect 57734 71814 57740 71878
rect 58213 71878 58279 71879
rect 58213 71846 58214 71878
rect 57664 71470 57740 71814
rect 57664 71438 57670 71470
rect 56984 71400 57060 71406
rect 57669 71406 57670 71438
rect 57734 71438 57740 71470
rect 58208 71814 58214 71846
rect 58278 71846 58279 71878
rect 58888 71878 58964 71884
rect 58278 71814 58284 71846
rect 58208 71470 58284 71814
rect 57734 71406 57735 71438
rect 57669 71405 57735 71406
rect 58208 71406 58214 71470
rect 58278 71406 58284 71470
rect 58888 71814 58894 71878
rect 58958 71814 58964 71878
rect 60661 71878 60727 71879
rect 60661 71846 60662 71878
rect 58888 71470 58964 71814
rect 58888 71438 58894 71470
rect 58208 71400 58284 71406
rect 58893 71406 58894 71438
rect 58958 71438 58964 71470
rect 60656 71814 60662 71846
rect 60726 71846 60727 71878
rect 61472 71878 61548 71884
rect 60726 71814 60732 71846
rect 60656 71470 60732 71814
rect 58958 71406 58959 71438
rect 58893 71405 58959 71406
rect 60656 71406 60662 71470
rect 60726 71406 60732 71470
rect 61472 71814 61478 71878
rect 61542 71814 61548 71878
rect 62021 71878 62087 71879
rect 62021 71846 62022 71878
rect 61472 71470 61548 71814
rect 61472 71438 61478 71470
rect 60656 71400 60732 71406
rect 61477 71406 61478 71438
rect 61542 71438 61548 71470
rect 62016 71814 62022 71846
rect 62086 71846 62087 71878
rect 62696 71878 62772 71884
rect 62086 71814 62092 71846
rect 62016 71470 62092 71814
rect 61542 71406 61543 71438
rect 61477 71405 61543 71406
rect 62016 71406 62022 71470
rect 62086 71406 62092 71470
rect 62696 71814 62702 71878
rect 62766 71814 62772 71878
rect 63109 71878 63175 71879
rect 63109 71846 63110 71878
rect 62696 71470 62772 71814
rect 62696 71438 62702 71470
rect 62016 71400 62092 71406
rect 62701 71406 62702 71438
rect 62766 71438 62772 71470
rect 63104 71814 63110 71846
rect 63174 71846 63175 71878
rect 63920 71878 63996 71884
rect 63174 71814 63180 71846
rect 63104 71470 63180 71814
rect 62766 71406 62767 71438
rect 62701 71405 62767 71406
rect 63104 71406 63110 71470
rect 63174 71406 63180 71470
rect 63920 71814 63926 71878
rect 63990 71814 63996 71878
rect 64469 71878 64535 71879
rect 64469 71846 64470 71878
rect 63920 71470 63996 71814
rect 63920 71438 63926 71470
rect 63104 71400 63180 71406
rect 63925 71406 63926 71438
rect 63990 71438 63996 71470
rect 64464 71814 64470 71846
rect 64534 71846 64535 71878
rect 65144 71878 65220 71884
rect 64534 71814 64540 71846
rect 64464 71470 64540 71814
rect 63990 71406 63991 71438
rect 63925 71405 63991 71406
rect 64464 71406 64470 71470
rect 64534 71406 64540 71470
rect 65144 71814 65150 71878
rect 65214 71814 65220 71878
rect 65693 71878 65759 71879
rect 65693 71846 65694 71878
rect 65144 71470 65220 71814
rect 65144 71438 65150 71470
rect 64464 71400 64540 71406
rect 65149 71406 65150 71438
rect 65214 71438 65220 71470
rect 65688 71814 65694 71846
rect 65758 71846 65759 71878
rect 65758 71814 65764 71846
rect 65688 71470 65764 71814
rect 65214 71406 65215 71438
rect 65149 71405 65215 71406
rect 65688 71406 65694 71470
rect 65758 71406 65764 71470
rect 65688 71400 65764 71406
rect 54128 71270 54134 71334
rect 54198 71270 54204 71334
rect 54128 71264 54204 71270
rect 66776 71198 66852 73310
rect 67733 71334 67799 71335
rect 67733 71302 67734 71334
rect 66776 71134 66782 71198
rect 66846 71134 66852 71198
rect 66776 71128 66852 71134
rect 67728 71270 67734 71302
rect 67798 71302 67799 71334
rect 67798 71270 67804 71302
rect 67728 71062 67804 71270
rect 67728 70998 67734 71062
rect 67798 70998 67804 71062
rect 72760 71062 72836 74670
rect 79424 74598 79500 77254
rect 79560 76094 79636 78614
rect 79560 76030 79566 76094
rect 79630 76030 79636 76094
rect 79560 76024 79636 76030
rect 89760 77590 90108 79294
rect 89760 77526 89766 77590
rect 89830 77526 90108 77590
rect 89760 75958 90108 77526
rect 89760 75894 89766 75958
rect 89830 75894 90108 75958
rect 79424 74566 79430 74598
rect 79429 74534 79430 74566
rect 79494 74566 79500 74598
rect 79560 75822 79636 75828
rect 79560 75758 79566 75822
rect 79630 75758 79636 75822
rect 79494 74534 79495 74566
rect 79429 74533 79495 74534
rect 79288 74462 79364 74468
rect 79288 74398 79294 74462
rect 79358 74398 79364 74462
rect 72760 71030 72766 71062
rect 67728 70992 67804 70998
rect 72765 70998 72766 71030
rect 72830 71030 72836 71062
rect 74120 73238 74196 73244
rect 74120 73174 74126 73238
rect 74190 73174 74196 73238
rect 72830 70998 72831 71030
rect 72765 70997 72831 70998
rect 25976 70894 25982 70926
rect 25981 70862 25982 70894
rect 26046 70894 26052 70926
rect 71133 70926 71199 70927
rect 71133 70894 71134 70926
rect 26046 70862 26047 70894
rect 25981 70861 26047 70862
rect 71128 70862 71134 70894
rect 71198 70894 71199 70926
rect 71405 70926 71471 70927
rect 71405 70894 71406 70926
rect 71198 70862 71204 70894
rect 66504 70518 66580 70524
rect 66504 70454 66510 70518
rect 66574 70454 66580 70518
rect 17952 70382 18028 70388
rect 17952 70318 17958 70382
rect 18022 70318 18028 70382
rect 18229 70382 18295 70383
rect 18229 70350 18230 70382
rect 17952 70110 18028 70318
rect 17952 70078 17958 70110
rect 17957 70046 17958 70078
rect 18022 70078 18028 70110
rect 18224 70318 18230 70350
rect 18294 70350 18295 70382
rect 18909 70382 18975 70383
rect 18909 70350 18910 70382
rect 18294 70318 18300 70350
rect 18224 70110 18300 70318
rect 18022 70046 18023 70078
rect 17957 70045 18023 70046
rect 18224 70046 18230 70110
rect 18294 70046 18300 70110
rect 18224 70040 18300 70046
rect 18904 70318 18910 70350
rect 18974 70350 18975 70382
rect 19040 70382 19116 70388
rect 18974 70318 18980 70350
rect 18904 70110 18980 70318
rect 18904 70046 18910 70110
rect 18974 70046 18980 70110
rect 19040 70318 19046 70382
rect 19110 70318 19116 70382
rect 19040 70110 19116 70318
rect 19040 70078 19046 70110
rect 18904 70040 18980 70046
rect 19045 70046 19046 70078
rect 19110 70078 19116 70110
rect 19584 70382 19660 70388
rect 19584 70318 19590 70382
rect 19654 70318 19660 70382
rect 19584 70110 19660 70318
rect 19584 70078 19590 70110
rect 19110 70046 19111 70078
rect 19045 70045 19111 70046
rect 19589 70046 19590 70078
rect 19654 70078 19660 70110
rect 66504 70110 66580 70454
rect 71128 70518 71204 70862
rect 71128 70454 71134 70518
rect 71198 70454 71204 70518
rect 71128 70448 71204 70454
rect 71400 70862 71406 70894
rect 71470 70894 71471 70926
rect 71470 70862 71476 70894
rect 71400 70518 71476 70862
rect 71400 70454 71406 70518
rect 71470 70454 71476 70518
rect 74120 70518 74196 73174
rect 79288 71742 79364 74398
rect 79560 73238 79636 75758
rect 79560 73206 79566 73238
rect 79565 73174 79566 73206
rect 79630 73206 79636 73238
rect 89760 74462 90108 75894
rect 89760 74398 89766 74462
rect 89830 74398 90108 74462
rect 79630 73174 79631 73206
rect 79565 73173 79631 73174
rect 88464 72725 88530 72726
rect 88464 72661 88465 72725
rect 88529 72661 88530 72725
rect 88464 72660 88530 72661
rect 79288 71710 79294 71742
rect 79293 71678 79294 71710
rect 79358 71710 79364 71742
rect 79358 71678 79359 71710
rect 79293 71677 79359 71678
rect 74120 70486 74126 70518
rect 71400 70448 71476 70454
rect 74125 70454 74126 70486
rect 74190 70486 74196 70518
rect 74190 70454 74191 70486
rect 74125 70453 74191 70454
rect 66504 70078 66510 70110
rect 19654 70046 19655 70078
rect 19589 70045 19655 70046
rect 66509 70046 66510 70078
rect 66574 70078 66580 70110
rect 71264 70382 71340 70388
rect 71264 70318 71270 70382
rect 71334 70318 71340 70382
rect 71677 70382 71743 70383
rect 71677 70350 71678 70382
rect 71264 70110 71340 70318
rect 71264 70078 71270 70110
rect 66574 70046 66575 70078
rect 66509 70045 66575 70046
rect 71269 70046 71270 70078
rect 71334 70078 71340 70110
rect 71672 70318 71678 70350
rect 71742 70350 71743 70382
rect 72216 70382 72292 70388
rect 71742 70318 71748 70350
rect 71672 70110 71748 70318
rect 71334 70046 71335 70078
rect 71269 70045 71335 70046
rect 71672 70046 71678 70110
rect 71742 70046 71748 70110
rect 72216 70318 72222 70382
rect 72286 70318 72292 70382
rect 72216 70110 72292 70318
rect 72216 70078 72222 70110
rect 71672 70040 71748 70046
rect 72221 70046 72222 70078
rect 72286 70078 72292 70110
rect 72352 70382 72428 70388
rect 72352 70318 72358 70382
rect 72422 70318 72428 70382
rect 73037 70382 73103 70383
rect 73037 70350 73038 70382
rect 72352 70110 72428 70318
rect 72352 70078 72358 70110
rect 72286 70046 72287 70078
rect 72221 70045 72287 70046
rect 72357 70046 72358 70078
rect 72422 70078 72428 70110
rect 73032 70318 73038 70350
rect 73102 70350 73103 70382
rect 73102 70318 73108 70350
rect 73032 70110 73108 70318
rect 72422 70046 72423 70078
rect 72357 70045 72423 70046
rect 73032 70046 73038 70110
rect 73102 70046 73108 70110
rect 73032 70040 73108 70046
rect 17957 69974 18023 69975
rect 17957 69942 17958 69974
rect 17952 69910 17958 69942
rect 18022 69942 18023 69974
rect 18229 69974 18295 69975
rect 18229 69942 18230 69974
rect 18022 69910 18028 69942
rect 17952 69702 18028 69910
rect 17952 69638 17958 69702
rect 18022 69638 18028 69702
rect 17952 69632 18028 69638
rect 18224 69910 18230 69942
rect 18294 69942 18295 69974
rect 19176 69974 19252 69980
rect 18294 69910 18300 69942
rect 18224 69702 18300 69910
rect 18224 69638 18230 69702
rect 18294 69638 18300 69702
rect 19176 69910 19182 69974
rect 19246 69910 19252 69974
rect 19589 69974 19655 69975
rect 19589 69942 19590 69974
rect 19176 69702 19252 69910
rect 19176 69670 19182 69702
rect 18224 69632 18300 69638
rect 19181 69638 19182 69670
rect 19246 69670 19252 69702
rect 19584 69910 19590 69942
rect 19654 69942 19655 69974
rect 71400 69974 71476 69980
rect 19654 69910 19660 69942
rect 19584 69702 19660 69910
rect 19246 69638 19247 69670
rect 19181 69637 19247 69638
rect 19584 69638 19590 69702
rect 19654 69638 19660 69702
rect 71400 69910 71406 69974
rect 71470 69910 71476 69974
rect 71813 69974 71879 69975
rect 71813 69942 71814 69974
rect 71400 69702 71476 69910
rect 71400 69670 71406 69702
rect 19584 69632 19660 69638
rect 71405 69638 71406 69670
rect 71470 69670 71476 69702
rect 71808 69910 71814 69942
rect 71878 69942 71879 69974
rect 72629 69974 72695 69975
rect 72629 69942 72630 69974
rect 71878 69910 71884 69942
rect 71808 69702 71884 69910
rect 71470 69638 71471 69670
rect 71405 69637 71471 69638
rect 71808 69638 71814 69702
rect 71878 69638 71884 69702
rect 71808 69632 71884 69638
rect 72624 69910 72630 69942
rect 72694 69942 72695 69974
rect 72896 69974 72972 69980
rect 72694 69910 72700 69942
rect 72624 69702 72700 69910
rect 72624 69638 72630 69702
rect 72694 69638 72700 69702
rect 72896 69910 72902 69974
rect 72966 69910 72972 69974
rect 72896 69702 72972 69910
rect 72896 69670 72902 69702
rect 72624 69632 72700 69638
rect 72901 69638 72902 69670
rect 72966 69670 72972 69702
rect 72966 69638 72967 69670
rect 72901 69637 72967 69638
rect 952 69230 1230 69294
rect 1294 69230 1300 69294
rect 17816 69566 17892 69572
rect 17816 69502 17822 69566
rect 17886 69502 17892 69566
rect 17816 69294 17892 69502
rect 17816 69262 17822 69294
rect 952 67798 1300 69230
rect 17821 69230 17822 69262
rect 17886 69262 17892 69294
rect 18224 69566 18300 69572
rect 18224 69502 18230 69566
rect 18294 69502 18300 69566
rect 19181 69566 19247 69567
rect 19181 69534 19182 69566
rect 18224 69294 18300 69502
rect 18224 69262 18230 69294
rect 17886 69230 17887 69262
rect 17821 69229 17887 69230
rect 18229 69230 18230 69262
rect 18294 69262 18300 69294
rect 19176 69502 19182 69534
rect 19246 69534 19247 69566
rect 19453 69566 19519 69567
rect 19453 69534 19454 69566
rect 19246 69502 19252 69534
rect 19176 69294 19252 69502
rect 18294 69230 18295 69262
rect 18229 69229 18295 69230
rect 19176 69230 19182 69294
rect 19246 69230 19252 69294
rect 19176 69224 19252 69230
rect 19448 69502 19454 69534
rect 19518 69534 19519 69566
rect 71405 69566 71471 69567
rect 71405 69534 71406 69566
rect 19518 69502 19524 69534
rect 19448 69294 19524 69502
rect 19448 69230 19454 69294
rect 19518 69230 19524 69294
rect 19448 69224 19524 69230
rect 71400 69502 71406 69534
rect 71470 69534 71471 69566
rect 71672 69566 71748 69572
rect 71470 69502 71476 69534
rect 71400 69294 71476 69502
rect 71400 69230 71406 69294
rect 71470 69230 71476 69294
rect 71672 69502 71678 69566
rect 71742 69502 71748 69566
rect 71672 69294 71748 69502
rect 71672 69262 71678 69294
rect 71400 69224 71476 69230
rect 71677 69230 71678 69262
rect 71742 69262 71748 69294
rect 72216 69566 72292 69572
rect 72216 69502 72222 69566
rect 72286 69502 72292 69566
rect 72901 69566 72967 69567
rect 72901 69534 72902 69566
rect 72216 69294 72292 69502
rect 72216 69262 72222 69294
rect 71742 69230 71743 69262
rect 71677 69229 71743 69230
rect 72221 69230 72222 69262
rect 72286 69262 72292 69294
rect 72896 69502 72902 69534
rect 72966 69534 72967 69566
rect 72966 69502 72972 69534
rect 72896 69294 72972 69502
rect 72286 69230 72287 69262
rect 72221 69229 72287 69230
rect 72896 69230 72902 69294
rect 72966 69230 72972 69294
rect 72896 69224 72972 69230
rect 17821 69158 17887 69159
rect 17821 69126 17822 69158
rect 17816 69094 17822 69126
rect 17886 69126 17887 69158
rect 18229 69158 18295 69159
rect 18229 69126 18230 69158
rect 17886 69094 17892 69126
rect 17816 68886 17892 69094
rect 17816 68822 17822 68886
rect 17886 68822 17892 68886
rect 17816 68816 17892 68822
rect 18224 69094 18230 69126
rect 18294 69126 18295 69158
rect 18496 69158 18572 69164
rect 18294 69094 18300 69126
rect 18224 68886 18300 69094
rect 18224 68822 18230 68886
rect 18294 68822 18300 68886
rect 18496 69094 18502 69158
rect 18566 69094 18572 69158
rect 18496 68886 18572 69094
rect 18496 68854 18502 68886
rect 18224 68816 18300 68822
rect 18501 68822 18502 68854
rect 18566 68854 18572 68886
rect 19040 69158 19116 69164
rect 19040 69094 19046 69158
rect 19110 69094 19116 69158
rect 19040 68886 19116 69094
rect 19040 68854 19046 68886
rect 18566 68822 18567 68854
rect 18501 68821 18567 68822
rect 19045 68822 19046 68854
rect 19110 68854 19116 68886
rect 19584 69158 19660 69164
rect 19584 69094 19590 69158
rect 19654 69094 19660 69158
rect 19584 68886 19660 69094
rect 19584 68854 19590 68886
rect 19110 68822 19111 68854
rect 19045 68821 19111 68822
rect 19589 68822 19590 68854
rect 19654 68854 19660 68886
rect 71264 69158 71340 69164
rect 71264 69094 71270 69158
rect 71334 69094 71340 69158
rect 71677 69158 71743 69159
rect 71677 69126 71678 69158
rect 71264 68886 71340 69094
rect 71264 68854 71270 68886
rect 19654 68822 19655 68854
rect 19589 68821 19655 68822
rect 71269 68822 71270 68854
rect 71334 68854 71340 68886
rect 71672 69094 71678 69126
rect 71742 69126 71743 69158
rect 72357 69158 72423 69159
rect 72357 69126 72358 69158
rect 71742 69094 71748 69126
rect 71672 68886 71748 69094
rect 71334 68822 71335 68854
rect 71269 68821 71335 68822
rect 71672 68822 71678 68886
rect 71742 68822 71748 68886
rect 71672 68816 71748 68822
rect 72352 69094 72358 69126
rect 72422 69126 72423 69158
rect 73032 69158 73108 69164
rect 72422 69094 72428 69126
rect 72352 68886 72428 69094
rect 72352 68822 72358 68886
rect 72422 68822 72428 68886
rect 73032 69094 73038 69158
rect 73102 69094 73108 69158
rect 73032 68886 73108 69094
rect 73032 68854 73038 68886
rect 72352 68816 72428 68822
rect 73037 68822 73038 68854
rect 73102 68854 73108 68886
rect 73102 68822 73103 68854
rect 73037 68821 73103 68822
rect 18360 68750 18436 68756
rect 18360 68686 18366 68750
rect 18430 68686 18436 68750
rect 18360 68478 18436 68686
rect 18360 68446 18366 68478
rect 18365 68414 18366 68446
rect 18430 68446 18436 68478
rect 18496 68750 18572 68756
rect 18496 68686 18502 68750
rect 18566 68686 18572 68750
rect 19181 68750 19247 68751
rect 19181 68718 19182 68750
rect 18496 68478 18572 68686
rect 18496 68446 18502 68478
rect 18430 68414 18431 68446
rect 18365 68413 18431 68414
rect 18501 68414 18502 68446
rect 18566 68446 18572 68478
rect 19176 68686 19182 68718
rect 19246 68718 19247 68750
rect 19453 68750 19519 68751
rect 19453 68718 19454 68750
rect 19246 68686 19252 68718
rect 19176 68478 19252 68686
rect 18566 68414 18567 68446
rect 18501 68413 18567 68414
rect 19176 68414 19182 68478
rect 19246 68414 19252 68478
rect 19176 68408 19252 68414
rect 19448 68686 19454 68718
rect 19518 68718 19519 68750
rect 71405 68750 71471 68751
rect 71405 68718 71406 68750
rect 19518 68686 19524 68718
rect 19448 68478 19524 68686
rect 71400 68686 71406 68718
rect 71470 68718 71471 68750
rect 71808 68750 71884 68756
rect 71470 68686 71476 68718
rect 66373 68614 66439 68615
rect 66373 68582 66374 68614
rect 19448 68414 19454 68478
rect 19518 68414 19524 68478
rect 19448 68408 19524 68414
rect 66368 68550 66374 68582
rect 66438 68582 66439 68614
rect 66438 68550 66444 68582
rect 19040 68342 19116 68348
rect 19040 68278 19046 68342
rect 19110 68278 19116 68342
rect 19589 68342 19655 68343
rect 19589 68310 19590 68342
rect 19040 68070 19116 68278
rect 19040 68038 19046 68070
rect 19045 68006 19046 68038
rect 19110 68038 19116 68070
rect 19584 68278 19590 68310
rect 19654 68310 19655 68342
rect 66368 68342 66444 68550
rect 71400 68478 71476 68686
rect 71400 68414 71406 68478
rect 71470 68414 71476 68478
rect 71808 68686 71814 68750
rect 71878 68686 71884 68750
rect 72085 68750 72151 68751
rect 72085 68718 72086 68750
rect 71808 68478 71884 68686
rect 71808 68446 71814 68478
rect 71400 68408 71476 68414
rect 71813 68414 71814 68446
rect 71878 68446 71884 68478
rect 72080 68686 72086 68718
rect 72150 68718 72151 68750
rect 72493 68750 72559 68751
rect 72493 68718 72494 68750
rect 72150 68686 72156 68718
rect 72080 68478 72156 68686
rect 71878 68414 71879 68446
rect 71813 68413 71879 68414
rect 72080 68414 72086 68478
rect 72150 68414 72156 68478
rect 72080 68408 72156 68414
rect 72488 68686 72494 68718
rect 72558 68718 72559 68750
rect 72558 68686 72564 68718
rect 72488 68478 72564 68686
rect 72488 68414 72494 68478
rect 72558 68414 72564 68478
rect 72488 68408 72564 68414
rect 19654 68278 19660 68310
rect 19584 68070 19660 68278
rect 66368 68278 66374 68342
rect 66438 68278 66444 68342
rect 66509 68342 66575 68343
rect 66509 68310 66510 68342
rect 66368 68272 66444 68278
rect 66504 68278 66510 68310
rect 66574 68310 66575 68342
rect 71264 68342 71340 68348
rect 66574 68278 66580 68310
rect 19110 68006 19111 68038
rect 19045 68005 19111 68006
rect 19584 68006 19590 68070
rect 19654 68006 19660 68070
rect 19584 68000 19660 68006
rect 952 67734 1230 67798
rect 1294 67734 1300 67798
rect 952 65894 1300 67734
rect 18496 67934 18572 67940
rect 18496 67870 18502 67934
rect 18566 67870 18572 67934
rect 19045 67934 19111 67935
rect 19045 67902 19046 67934
rect 17821 67662 17887 67663
rect 17821 67630 17822 67662
rect 17816 67598 17822 67630
rect 17886 67630 17887 67662
rect 18496 67662 18572 67870
rect 18496 67630 18502 67662
rect 17886 67598 17892 67630
rect 17816 67390 17892 67598
rect 18501 67598 18502 67630
rect 18566 67630 18572 67662
rect 19040 67870 19046 67902
rect 19110 67902 19111 67934
rect 19448 67934 19524 67940
rect 19110 67870 19116 67902
rect 19040 67662 19116 67870
rect 18566 67598 18567 67630
rect 18501 67597 18567 67598
rect 19040 67598 19046 67662
rect 19110 67598 19116 67662
rect 19448 67870 19454 67934
rect 19518 67870 19524 67934
rect 19448 67662 19524 67870
rect 66504 67934 66580 68278
rect 71264 68278 71270 68342
rect 71334 68278 71340 68342
rect 71813 68342 71879 68343
rect 71813 68310 71814 68342
rect 71264 68070 71340 68278
rect 71264 68038 71270 68070
rect 71269 68006 71270 68038
rect 71334 68038 71340 68070
rect 71808 68278 71814 68310
rect 71878 68310 71879 68342
rect 71878 68278 71884 68310
rect 71808 68070 71884 68278
rect 71334 68006 71335 68038
rect 71269 68005 71335 68006
rect 71808 68006 71814 68070
rect 71878 68006 71884 68070
rect 71808 68000 71884 68006
rect 66504 67870 66510 67934
rect 66574 67870 66580 67934
rect 71269 67934 71335 67935
rect 71269 67902 71270 67934
rect 66504 67864 66580 67870
rect 71264 67870 71270 67902
rect 71334 67902 71335 67934
rect 71672 67934 71748 67940
rect 71334 67870 71340 67902
rect 19448 67630 19454 67662
rect 19040 67592 19116 67598
rect 19453 67598 19454 67630
rect 19518 67630 19524 67662
rect 71264 67662 71340 67870
rect 19518 67598 19519 67630
rect 19453 67597 19519 67598
rect 71264 67598 71270 67662
rect 71334 67598 71340 67662
rect 71672 67870 71678 67934
rect 71742 67870 71748 67934
rect 72357 67934 72423 67935
rect 72357 67902 72358 67934
rect 71672 67662 71748 67870
rect 71672 67630 71678 67662
rect 71264 67592 71340 67598
rect 71677 67598 71678 67630
rect 71742 67630 71748 67662
rect 72352 67870 72358 67902
rect 72422 67902 72423 67934
rect 72422 67870 72428 67902
rect 72352 67662 72428 67870
rect 71742 67598 71743 67630
rect 71677 67597 71743 67598
rect 72352 67598 72358 67662
rect 72422 67598 72428 67662
rect 72352 67592 72428 67598
rect 72896 67662 72972 67668
rect 72896 67598 72902 67662
rect 72966 67598 72972 67662
rect 17816 67326 17822 67390
rect 17886 67326 17892 67390
rect 17816 67320 17892 67326
rect 24344 67390 24420 67396
rect 24344 67326 24350 67390
rect 24414 67326 24420 67390
rect 17816 67254 17892 67260
rect 17816 67190 17822 67254
rect 17886 67190 17892 67254
rect 18501 67254 18567 67255
rect 18501 67222 18502 67254
rect 17816 66982 17892 67190
rect 17816 66950 17822 66982
rect 17821 66918 17822 66950
rect 17886 66950 17892 66982
rect 18496 67190 18502 67222
rect 18566 67222 18567 67254
rect 18566 67190 18572 67222
rect 18496 66982 18572 67190
rect 24344 67118 24420 67326
rect 24344 67086 24350 67118
rect 24349 67054 24350 67086
rect 24414 67086 24420 67118
rect 66504 67390 66580 67396
rect 66504 67326 66510 67390
rect 66574 67326 66580 67390
rect 72896 67390 72972 67598
rect 72896 67358 72902 67390
rect 66504 67118 66580 67326
rect 72901 67326 72902 67358
rect 72966 67358 72972 67390
rect 87725 67390 87791 67391
rect 87725 67358 87726 67390
rect 72966 67326 72967 67358
rect 72901 67325 72967 67326
rect 87720 67326 87726 67358
rect 87790 67358 87791 67390
rect 87790 67326 87796 67358
rect 72085 67254 72151 67255
rect 72085 67222 72086 67254
rect 66504 67086 66510 67118
rect 24414 67054 24415 67086
rect 24349 67053 24415 67054
rect 66509 67054 66510 67086
rect 66574 67086 66580 67118
rect 72080 67190 72086 67222
rect 72150 67222 72151 67254
rect 72624 67254 72700 67260
rect 72150 67190 72156 67222
rect 66574 67054 66575 67086
rect 66509 67053 66575 67054
rect 17886 66918 17887 66950
rect 17821 66917 17887 66918
rect 18496 66918 18502 66982
rect 18566 66918 18572 66982
rect 24621 66982 24687 66983
rect 24621 66950 24622 66982
rect 18496 66912 18572 66918
rect 24616 66918 24622 66950
rect 24686 66950 24687 66982
rect 66509 66982 66575 66983
rect 66509 66950 66510 66982
rect 24686 66918 24692 66950
rect 17821 66846 17887 66847
rect 17821 66814 17822 66846
rect 17816 66782 17822 66814
rect 17886 66814 17887 66846
rect 17886 66782 17892 66814
rect 17816 66574 17892 66782
rect 24616 66710 24692 66918
rect 24616 66646 24622 66710
rect 24686 66646 24692 66710
rect 24616 66640 24692 66646
rect 66504 66918 66510 66950
rect 66574 66950 66575 66982
rect 72080 66982 72156 67190
rect 66574 66918 66580 66950
rect 66504 66710 66580 66918
rect 72080 66918 72086 66982
rect 72150 66918 72156 66982
rect 72624 67190 72630 67254
rect 72694 67190 72700 67254
rect 72901 67254 72967 67255
rect 72901 67222 72902 67254
rect 72624 66982 72700 67190
rect 72624 66950 72630 66982
rect 72080 66912 72156 66918
rect 72629 66918 72630 66950
rect 72694 66950 72700 66982
rect 72896 67190 72902 67222
rect 72966 67222 72967 67254
rect 72966 67190 72972 67222
rect 72896 66982 72972 67190
rect 72694 66918 72695 66950
rect 72629 66917 72695 66918
rect 72896 66918 72902 66982
rect 72966 66918 72972 66982
rect 72896 66912 72972 66918
rect 72896 66846 72972 66852
rect 72896 66782 72902 66846
rect 72966 66782 72972 66846
rect 66504 66646 66510 66710
rect 66574 66646 66580 66710
rect 66504 66640 66580 66646
rect 72080 66710 72156 66716
rect 72080 66646 72086 66710
rect 72150 66646 72156 66710
rect 17816 66510 17822 66574
rect 17886 66510 17892 66574
rect 17816 66504 17892 66510
rect 17952 66438 18028 66444
rect 17952 66374 17958 66438
rect 18022 66374 18028 66438
rect 18909 66438 18975 66439
rect 18909 66406 18910 66438
rect 17952 66166 18028 66374
rect 17952 66134 17958 66166
rect 17957 66102 17958 66134
rect 18022 66134 18028 66166
rect 18904 66374 18910 66406
rect 18974 66406 18975 66438
rect 19176 66438 19252 66444
rect 18974 66374 18980 66406
rect 18904 66166 18980 66374
rect 18022 66102 18023 66134
rect 17957 66101 18023 66102
rect 18904 66102 18910 66166
rect 18974 66102 18980 66166
rect 19176 66374 19182 66438
rect 19246 66374 19252 66438
rect 19453 66438 19519 66439
rect 19453 66406 19454 66438
rect 19176 66166 19252 66374
rect 19176 66134 19182 66166
rect 18904 66096 18980 66102
rect 19181 66102 19182 66134
rect 19246 66134 19252 66166
rect 19448 66374 19454 66406
rect 19518 66406 19519 66438
rect 71405 66438 71471 66439
rect 71405 66406 71406 66438
rect 19518 66374 19524 66406
rect 19448 66166 19524 66374
rect 71400 66374 71406 66406
rect 71470 66406 71471 66438
rect 71808 66438 71884 66444
rect 71470 66374 71476 66406
rect 19246 66102 19247 66134
rect 19181 66101 19247 66102
rect 19448 66102 19454 66166
rect 19518 66102 19524 66166
rect 24621 66166 24687 66167
rect 24621 66134 24622 66166
rect 19448 66096 19524 66102
rect 24616 66102 24622 66134
rect 24686 66134 24687 66166
rect 66509 66166 66575 66167
rect 66509 66134 66510 66166
rect 24686 66102 24692 66134
rect 17821 66030 17887 66031
rect 17821 65998 17822 66030
rect 952 65830 1230 65894
rect 1294 65830 1300 65894
rect 952 64262 1300 65830
rect 17816 65966 17822 65998
rect 17886 65998 17887 66030
rect 18229 66030 18295 66031
rect 18229 65998 18230 66030
rect 17886 65966 17892 65998
rect 17816 65758 17892 65966
rect 17816 65694 17822 65758
rect 17886 65694 17892 65758
rect 17816 65688 17892 65694
rect 18224 65966 18230 65998
rect 18294 65998 18295 66030
rect 18768 66030 18844 66036
rect 18294 65966 18300 65998
rect 18224 65758 18300 65966
rect 18224 65694 18230 65758
rect 18294 65694 18300 65758
rect 18768 65966 18774 66030
rect 18838 65966 18844 66030
rect 18768 65758 18844 65966
rect 18768 65726 18774 65758
rect 18224 65688 18300 65694
rect 18773 65694 18774 65726
rect 18838 65726 18844 65758
rect 19040 66030 19116 66036
rect 19040 65966 19046 66030
rect 19110 65966 19116 66030
rect 19453 66030 19519 66031
rect 19453 65998 19454 66030
rect 19040 65758 19116 65966
rect 19040 65726 19046 65758
rect 18838 65694 18839 65726
rect 18773 65693 18839 65694
rect 19045 65694 19046 65726
rect 19110 65726 19116 65758
rect 19448 65966 19454 65998
rect 19518 65998 19519 66030
rect 19518 65966 19524 65998
rect 19448 65758 19524 65966
rect 24616 65894 24692 66102
rect 24616 65830 24622 65894
rect 24686 65830 24692 65894
rect 24616 65824 24692 65830
rect 66504 66102 66510 66134
rect 66574 66134 66575 66166
rect 71400 66166 71476 66374
rect 66574 66102 66580 66134
rect 66504 65894 66580 66102
rect 71400 66102 71406 66166
rect 71470 66102 71476 66166
rect 71808 66374 71814 66438
rect 71878 66374 71884 66438
rect 71808 66166 71884 66374
rect 72080 66302 72156 66646
rect 72896 66574 72972 66782
rect 72896 66542 72902 66574
rect 72901 66510 72902 66542
rect 72966 66542 72972 66574
rect 72966 66510 72967 66542
rect 72901 66509 72967 66510
rect 72901 66438 72967 66439
rect 72901 66406 72902 66438
rect 72080 66270 72086 66302
rect 72085 66238 72086 66270
rect 72150 66270 72156 66302
rect 72896 66374 72902 66406
rect 72966 66406 72967 66438
rect 72966 66374 72972 66406
rect 72150 66238 72151 66270
rect 72085 66237 72151 66238
rect 71808 66134 71814 66166
rect 71400 66096 71476 66102
rect 71813 66102 71814 66134
rect 71878 66134 71884 66166
rect 72896 66166 72972 66374
rect 71878 66102 71879 66134
rect 71813 66101 71879 66102
rect 72896 66102 72902 66166
rect 72966 66102 72972 66166
rect 72896 66096 72972 66102
rect 71269 66030 71335 66031
rect 71269 65998 71270 66030
rect 66504 65830 66510 65894
rect 66574 65830 66580 65894
rect 66504 65824 66580 65830
rect 71264 65966 71270 65998
rect 71334 65998 71335 66030
rect 71677 66030 71743 66031
rect 71677 65998 71678 66030
rect 71334 65966 71340 65998
rect 19110 65694 19111 65726
rect 19045 65693 19111 65694
rect 19448 65694 19454 65758
rect 19518 65694 19524 65758
rect 19448 65688 19524 65694
rect 71264 65758 71340 65966
rect 71264 65694 71270 65758
rect 71334 65694 71340 65758
rect 71264 65688 71340 65694
rect 71672 65966 71678 65998
rect 71742 65998 71743 66030
rect 72216 66030 72292 66036
rect 71742 65966 71748 65998
rect 71672 65758 71748 65966
rect 71672 65694 71678 65758
rect 71742 65694 71748 65758
rect 72216 65966 72222 66030
rect 72286 65966 72292 66030
rect 72357 66030 72423 66031
rect 72357 65998 72358 66030
rect 72216 65758 72292 65966
rect 72216 65726 72222 65758
rect 71672 65688 71748 65694
rect 72221 65694 72222 65726
rect 72286 65726 72292 65758
rect 72352 65966 72358 65998
rect 72422 65998 72423 66030
rect 73032 66030 73108 66036
rect 72422 65966 72428 65998
rect 72352 65758 72428 65966
rect 72286 65694 72287 65726
rect 72221 65693 72287 65694
rect 72352 65694 72358 65758
rect 72422 65694 72428 65758
rect 73032 65966 73038 66030
rect 73102 65966 73108 66030
rect 73032 65758 73108 65966
rect 73032 65726 73038 65758
rect 72352 65688 72428 65694
rect 73037 65694 73038 65726
rect 73102 65726 73108 65758
rect 73102 65694 73103 65726
rect 73037 65693 73103 65694
rect 17816 65622 17892 65628
rect 17816 65558 17822 65622
rect 17886 65558 17892 65622
rect 18229 65622 18295 65623
rect 18229 65590 18230 65622
rect 17816 65350 17892 65558
rect 17816 65318 17822 65350
rect 17821 65286 17822 65318
rect 17886 65318 17892 65350
rect 18224 65558 18230 65590
rect 18294 65590 18295 65622
rect 18496 65622 18572 65628
rect 18294 65558 18300 65590
rect 18224 65350 18300 65558
rect 17886 65286 17887 65318
rect 17821 65285 17887 65286
rect 18224 65286 18230 65350
rect 18294 65286 18300 65350
rect 18496 65558 18502 65622
rect 18566 65558 18572 65622
rect 19045 65622 19111 65623
rect 19045 65590 19046 65622
rect 18496 65350 18572 65558
rect 18496 65318 18502 65350
rect 18224 65280 18300 65286
rect 18501 65286 18502 65318
rect 18566 65318 18572 65350
rect 19040 65558 19046 65590
rect 19110 65590 19111 65622
rect 19448 65622 19524 65628
rect 19110 65558 19116 65590
rect 19040 65350 19116 65558
rect 18566 65286 18567 65318
rect 18501 65285 18567 65286
rect 19040 65286 19046 65350
rect 19110 65286 19116 65350
rect 19448 65558 19454 65622
rect 19518 65558 19524 65622
rect 19448 65350 19524 65558
rect 19448 65318 19454 65350
rect 19040 65280 19116 65286
rect 19453 65286 19454 65318
rect 19518 65318 19524 65350
rect 71400 65622 71476 65628
rect 71400 65558 71406 65622
rect 71470 65558 71476 65622
rect 71400 65350 71476 65558
rect 71400 65318 71406 65350
rect 19518 65286 19519 65318
rect 19453 65285 19519 65286
rect 71405 65286 71406 65318
rect 71470 65318 71476 65350
rect 71672 65622 71748 65628
rect 71672 65558 71678 65622
rect 71742 65558 71748 65622
rect 71672 65350 71748 65558
rect 71672 65318 71678 65350
rect 71470 65286 71471 65318
rect 71405 65285 71471 65286
rect 71677 65286 71678 65318
rect 71742 65318 71748 65350
rect 72080 65622 72156 65628
rect 72080 65558 72086 65622
rect 72150 65558 72156 65622
rect 72080 65350 72156 65558
rect 72080 65318 72086 65350
rect 71742 65286 71743 65318
rect 71677 65285 71743 65286
rect 72085 65286 72086 65318
rect 72150 65318 72156 65350
rect 72488 65622 72564 65628
rect 72488 65558 72494 65622
rect 72558 65558 72564 65622
rect 72488 65350 72564 65558
rect 72488 65318 72494 65350
rect 72150 65286 72151 65318
rect 72085 65285 72151 65286
rect 72493 65286 72494 65318
rect 72558 65318 72564 65350
rect 72896 65622 72972 65628
rect 72896 65558 72902 65622
rect 72966 65558 72972 65622
rect 72896 65350 72972 65558
rect 72896 65318 72902 65350
rect 72558 65286 72559 65318
rect 72493 65285 72559 65286
rect 72901 65286 72902 65318
rect 72966 65318 72972 65350
rect 72966 65286 72967 65318
rect 72901 65285 72967 65286
rect 17816 65214 17892 65220
rect 17816 65150 17822 65214
rect 17886 65150 17892 65214
rect 18637 65214 18703 65215
rect 18637 65182 18638 65214
rect 17816 64942 17892 65150
rect 17816 64910 17822 64942
rect 17821 64878 17822 64910
rect 17886 64910 17892 64942
rect 18632 65150 18638 65182
rect 18702 65182 18703 65214
rect 19181 65214 19247 65215
rect 19181 65182 19182 65214
rect 18702 65150 18708 65182
rect 18632 64942 18708 65150
rect 17886 64878 17887 64910
rect 17821 64877 17887 64878
rect 18632 64878 18638 64942
rect 18702 64878 18708 64942
rect 18632 64872 18708 64878
rect 19176 65150 19182 65182
rect 19246 65182 19247 65214
rect 19453 65214 19519 65215
rect 19453 65182 19454 65214
rect 19246 65150 19252 65182
rect 19176 64942 19252 65150
rect 19176 64878 19182 64942
rect 19246 64878 19252 64942
rect 19176 64872 19252 64878
rect 19448 65150 19454 65182
rect 19518 65182 19519 65214
rect 71405 65214 71471 65215
rect 71405 65182 71406 65214
rect 19518 65150 19524 65182
rect 19448 64942 19524 65150
rect 19448 64878 19454 64942
rect 19518 64878 19524 64942
rect 19448 64872 19524 64878
rect 71400 65150 71406 65182
rect 71470 65182 71471 65214
rect 71813 65214 71879 65215
rect 71813 65182 71814 65214
rect 71470 65150 71476 65182
rect 71400 64942 71476 65150
rect 71400 64878 71406 64942
rect 71470 64878 71476 64942
rect 71400 64872 71476 64878
rect 71808 65150 71814 65182
rect 71878 65182 71879 65214
rect 72352 65214 72428 65220
rect 71878 65150 71884 65182
rect 71808 64942 71884 65150
rect 71808 64878 71814 64942
rect 71878 64878 71884 64942
rect 72352 65150 72358 65214
rect 72422 65150 72428 65214
rect 72352 64942 72428 65150
rect 72352 64910 72358 64942
rect 71808 64872 71884 64878
rect 72357 64878 72358 64910
rect 72422 64910 72428 64942
rect 73032 65214 73108 65220
rect 73032 65150 73038 65214
rect 73102 65150 73108 65214
rect 73032 64942 73108 65150
rect 73032 64910 73038 64942
rect 72422 64878 72423 64910
rect 72357 64877 72423 64878
rect 73037 64878 73038 64910
rect 73102 64910 73108 64942
rect 73102 64878 73103 64910
rect 73037 64877 73103 64878
rect 18229 64806 18295 64807
rect 18229 64774 18230 64806
rect 18224 64742 18230 64774
rect 18294 64774 18295 64806
rect 18909 64806 18975 64807
rect 18909 64774 18910 64806
rect 18294 64742 18300 64774
rect 18224 64534 18300 64742
rect 18224 64470 18230 64534
rect 18294 64470 18300 64534
rect 18224 64464 18300 64470
rect 18904 64742 18910 64774
rect 18974 64774 18975 64806
rect 19040 64806 19116 64812
rect 18974 64742 18980 64774
rect 18904 64534 18980 64742
rect 18904 64470 18910 64534
rect 18974 64470 18980 64534
rect 19040 64742 19046 64806
rect 19110 64742 19116 64806
rect 19040 64534 19116 64742
rect 19040 64502 19046 64534
rect 18904 64464 18980 64470
rect 19045 64470 19046 64502
rect 19110 64502 19116 64534
rect 19584 64806 19660 64812
rect 19584 64742 19590 64806
rect 19654 64742 19660 64806
rect 19584 64534 19660 64742
rect 19584 64502 19590 64534
rect 19110 64470 19111 64502
rect 19045 64469 19111 64470
rect 19589 64470 19590 64502
rect 19654 64502 19660 64534
rect 71264 64806 71340 64812
rect 71264 64742 71270 64806
rect 71334 64742 71340 64806
rect 71677 64806 71743 64807
rect 71677 64774 71678 64806
rect 71264 64534 71340 64742
rect 71264 64502 71270 64534
rect 19654 64470 19655 64502
rect 19589 64469 19655 64470
rect 71269 64470 71270 64502
rect 71334 64502 71340 64534
rect 71672 64742 71678 64774
rect 71742 64774 71743 64806
rect 72216 64806 72292 64812
rect 71742 64742 71748 64774
rect 71672 64534 71748 64742
rect 71334 64470 71335 64502
rect 71269 64469 71335 64470
rect 71672 64470 71678 64534
rect 71742 64470 71748 64534
rect 72216 64742 72222 64806
rect 72286 64742 72292 64806
rect 72216 64534 72292 64742
rect 72216 64502 72222 64534
rect 71672 64464 71748 64470
rect 72221 64470 72222 64502
rect 72286 64502 72292 64534
rect 72624 64806 72700 64812
rect 72624 64742 72630 64806
rect 72694 64742 72700 64806
rect 72624 64534 72700 64742
rect 87720 64670 87796 67326
rect 87720 64606 87726 64670
rect 87790 64606 87796 64670
rect 87720 64600 87796 64606
rect 72624 64502 72630 64534
rect 72286 64470 72287 64502
rect 72221 64469 72287 64470
rect 72629 64470 72630 64502
rect 72694 64502 72700 64534
rect 87589 64534 87655 64535
rect 87589 64502 87590 64534
rect 72694 64470 72695 64502
rect 72629 64469 72695 64470
rect 87584 64470 87590 64502
rect 87654 64502 87655 64534
rect 87654 64470 87660 64502
rect 952 64198 1230 64262
rect 1294 64198 1300 64262
rect 952 62494 1300 64198
rect 17952 64398 18028 64404
rect 17952 64334 17958 64398
rect 18022 64334 18028 64398
rect 17952 64126 18028 64334
rect 17952 64094 17958 64126
rect 17957 64062 17958 64094
rect 18022 64094 18028 64126
rect 18360 64398 18436 64404
rect 18360 64334 18366 64398
rect 18430 64334 18436 64398
rect 19181 64398 19247 64399
rect 19181 64366 19182 64398
rect 18360 64126 18436 64334
rect 18360 64094 18366 64126
rect 18022 64062 18023 64094
rect 17957 64061 18023 64062
rect 18365 64062 18366 64094
rect 18430 64094 18436 64126
rect 19176 64334 19182 64366
rect 19246 64366 19247 64398
rect 19584 64398 19660 64404
rect 19246 64334 19252 64366
rect 19176 64126 19252 64334
rect 18430 64062 18431 64094
rect 18365 64061 18431 64062
rect 19176 64062 19182 64126
rect 19246 64062 19252 64126
rect 19584 64334 19590 64398
rect 19654 64334 19660 64398
rect 19584 64126 19660 64334
rect 19584 64094 19590 64126
rect 19176 64056 19252 64062
rect 19589 64062 19590 64094
rect 19654 64094 19660 64126
rect 71400 64398 71476 64404
rect 71400 64334 71406 64398
rect 71470 64334 71476 64398
rect 71677 64398 71743 64399
rect 71677 64366 71678 64398
rect 71400 64126 71476 64334
rect 71400 64094 71406 64126
rect 19654 64062 19655 64094
rect 19589 64061 19655 64062
rect 71405 64062 71406 64094
rect 71470 64094 71476 64126
rect 71672 64334 71678 64366
rect 71742 64366 71743 64398
rect 72493 64398 72559 64399
rect 72493 64366 72494 64398
rect 71742 64334 71748 64366
rect 71672 64126 71748 64334
rect 71470 64062 71471 64094
rect 71405 64061 71471 64062
rect 71672 64062 71678 64126
rect 71742 64062 71748 64126
rect 71672 64056 71748 64062
rect 72488 64334 72494 64366
rect 72558 64366 72559 64398
rect 72896 64398 72972 64404
rect 72558 64334 72564 64366
rect 72488 64126 72564 64334
rect 72488 64062 72494 64126
rect 72558 64062 72564 64126
rect 72896 64334 72902 64398
rect 72966 64334 72972 64398
rect 72896 64126 72972 64334
rect 72896 64094 72902 64126
rect 72488 64056 72564 64062
rect 72901 64062 72902 64094
rect 72966 64094 72972 64126
rect 72966 64062 72967 64094
rect 72901 64061 72967 64062
rect 18909 63990 18975 63991
rect 18909 63958 18910 63990
rect 18904 63926 18910 63958
rect 18974 63958 18975 63990
rect 19181 63990 19247 63991
rect 19181 63958 19182 63990
rect 18974 63926 18980 63958
rect 17821 63718 17887 63719
rect 17821 63686 17822 63718
rect 17816 63654 17822 63686
rect 17886 63686 17887 63718
rect 18904 63718 18980 63926
rect 17886 63654 17892 63686
rect 17816 63446 17892 63654
rect 18904 63654 18910 63718
rect 18974 63654 18980 63718
rect 18904 63648 18980 63654
rect 19176 63926 19182 63958
rect 19246 63958 19247 63990
rect 19589 63990 19655 63991
rect 19589 63958 19590 63990
rect 19246 63926 19252 63958
rect 19176 63718 19252 63926
rect 19176 63654 19182 63718
rect 19246 63654 19252 63718
rect 19176 63648 19252 63654
rect 19584 63926 19590 63958
rect 19654 63958 19655 63990
rect 71264 63990 71340 63996
rect 19654 63926 19660 63958
rect 19584 63718 19660 63926
rect 71264 63926 71270 63990
rect 71334 63926 71340 63990
rect 19584 63654 19590 63718
rect 19654 63654 19660 63718
rect 19584 63648 19660 63654
rect 24480 63854 24556 63860
rect 24480 63790 24486 63854
rect 24550 63790 24556 63854
rect 66509 63854 66575 63855
rect 66509 63822 66510 63854
rect 24480 63582 24556 63790
rect 24480 63550 24486 63582
rect 24485 63518 24486 63550
rect 24550 63550 24556 63582
rect 66504 63790 66510 63822
rect 66574 63822 66575 63854
rect 66574 63790 66580 63822
rect 66504 63582 66580 63790
rect 71264 63718 71340 63926
rect 71264 63686 71270 63718
rect 71269 63654 71270 63686
rect 71334 63686 71340 63718
rect 71672 63990 71748 63996
rect 71672 63926 71678 63990
rect 71742 63926 71748 63990
rect 72085 63990 72151 63991
rect 72085 63958 72086 63990
rect 71672 63718 71748 63926
rect 71672 63686 71678 63718
rect 71334 63654 71335 63686
rect 71269 63653 71335 63654
rect 71677 63654 71678 63686
rect 71742 63686 71748 63718
rect 72080 63926 72086 63958
rect 72150 63958 72151 63990
rect 72352 63990 72428 63996
rect 72150 63926 72156 63958
rect 72080 63718 72156 63926
rect 71742 63654 71743 63686
rect 71677 63653 71743 63654
rect 72080 63654 72086 63718
rect 72150 63654 72156 63718
rect 72352 63926 72358 63990
rect 72422 63926 72428 63990
rect 72352 63718 72428 63926
rect 72352 63686 72358 63718
rect 72080 63648 72156 63654
rect 72357 63654 72358 63686
rect 72422 63686 72428 63718
rect 73037 63718 73103 63719
rect 73037 63686 73038 63718
rect 72422 63654 72423 63686
rect 72357 63653 72423 63654
rect 73032 63654 73038 63686
rect 73102 63686 73103 63718
rect 73102 63654 73108 63686
rect 24550 63518 24551 63550
rect 24485 63517 24551 63518
rect 66504 63518 66510 63582
rect 66574 63518 66580 63582
rect 66504 63512 66580 63518
rect 17816 63382 17822 63446
rect 17886 63382 17892 63446
rect 17816 63376 17892 63382
rect 24616 63446 24692 63452
rect 24616 63382 24622 63446
rect 24686 63382 24692 63446
rect 17952 63310 18028 63316
rect 17952 63246 17958 63310
rect 18022 63246 18028 63310
rect 18501 63310 18567 63311
rect 18501 63278 18502 63310
rect 17952 63038 18028 63246
rect 17952 63006 17958 63038
rect 17957 62974 17958 63006
rect 18022 63006 18028 63038
rect 18496 63246 18502 63278
rect 18566 63278 18567 63310
rect 18566 63246 18572 63278
rect 18496 63038 18572 63246
rect 24616 63174 24692 63382
rect 24616 63142 24622 63174
rect 24621 63110 24622 63142
rect 24686 63142 24692 63174
rect 66368 63446 66444 63452
rect 66368 63382 66374 63446
rect 66438 63382 66444 63446
rect 66368 63174 66444 63382
rect 73032 63446 73108 63654
rect 73032 63382 73038 63446
rect 73102 63382 73108 63446
rect 73032 63376 73108 63382
rect 72085 63310 72151 63311
rect 72085 63278 72086 63310
rect 66368 63142 66374 63174
rect 24686 63110 24687 63142
rect 24621 63109 24687 63110
rect 66373 63110 66374 63142
rect 66438 63142 66444 63174
rect 72080 63246 72086 63278
rect 72150 63278 72151 63310
rect 72896 63310 72972 63316
rect 72150 63246 72156 63278
rect 66438 63110 66439 63142
rect 66373 63109 66439 63110
rect 18022 62974 18023 63006
rect 17957 62973 18023 62974
rect 18496 62974 18502 63038
rect 18566 62974 18572 63038
rect 18496 62968 18572 62974
rect 24344 63038 24420 63044
rect 24344 62974 24350 63038
rect 24414 62974 24420 63038
rect 66373 63038 66439 63039
rect 66373 63006 66374 63038
rect 17957 62902 18023 62903
rect 17957 62870 17958 62902
rect 17952 62838 17958 62870
rect 18022 62870 18023 62902
rect 18022 62838 18028 62870
rect 17952 62630 18028 62838
rect 24344 62766 24420 62974
rect 24344 62734 24350 62766
rect 24349 62702 24350 62734
rect 24414 62734 24420 62766
rect 66368 62974 66374 63006
rect 66438 63006 66439 63038
rect 72080 63038 72156 63246
rect 66438 62974 66444 63006
rect 66368 62766 66444 62974
rect 72080 62974 72086 63038
rect 72150 62974 72156 63038
rect 72896 63246 72902 63310
rect 72966 63246 72972 63310
rect 72896 63038 72972 63246
rect 72896 63006 72902 63038
rect 72080 62968 72156 62974
rect 72901 62974 72902 63006
rect 72966 63006 72972 63038
rect 72966 62974 72967 63006
rect 72901 62973 72967 62974
rect 72901 62902 72967 62903
rect 72901 62870 72902 62902
rect 72896 62838 72902 62870
rect 72966 62870 72967 62902
rect 72966 62838 72972 62870
rect 24414 62702 24415 62734
rect 24349 62701 24415 62702
rect 66368 62702 66374 62766
rect 66438 62702 66444 62766
rect 66368 62696 66444 62702
rect 66504 62766 66580 62772
rect 66504 62702 66510 62766
rect 66574 62702 66580 62766
rect 17952 62566 17958 62630
rect 18022 62566 18028 62630
rect 17952 62560 18028 62566
rect 952 62430 1230 62494
rect 1294 62430 1300 62494
rect 952 60862 1300 62430
rect 17816 62494 17892 62500
rect 17816 62430 17822 62494
rect 17886 62430 17892 62494
rect 17816 62222 17892 62430
rect 17816 62190 17822 62222
rect 17821 62158 17822 62190
rect 17886 62190 17892 62222
rect 18360 62494 18436 62500
rect 18360 62430 18366 62494
rect 18430 62430 18436 62494
rect 19045 62494 19111 62495
rect 19045 62462 19046 62494
rect 18360 62222 18436 62430
rect 18360 62190 18366 62222
rect 17886 62158 17887 62190
rect 17821 62157 17887 62158
rect 18365 62158 18366 62190
rect 18430 62190 18436 62222
rect 19040 62430 19046 62462
rect 19110 62462 19111 62494
rect 19589 62494 19655 62495
rect 19589 62462 19590 62494
rect 19110 62430 19116 62462
rect 19040 62222 19116 62430
rect 18430 62158 18431 62190
rect 18365 62157 18431 62158
rect 19040 62158 19046 62222
rect 19110 62158 19116 62222
rect 19040 62152 19116 62158
rect 19584 62430 19590 62462
rect 19654 62462 19655 62494
rect 66504 62494 66580 62702
rect 72896 62630 72972 62838
rect 72896 62566 72902 62630
rect 72966 62566 72972 62630
rect 72896 62560 72972 62566
rect 66504 62462 66510 62494
rect 19654 62430 19660 62462
rect 19584 62222 19660 62430
rect 66509 62430 66510 62462
rect 66574 62462 66580 62494
rect 71400 62494 71476 62500
rect 66574 62430 66575 62462
rect 66509 62429 66575 62430
rect 71400 62430 71406 62494
rect 71470 62430 71476 62494
rect 71677 62494 71743 62495
rect 71677 62462 71678 62494
rect 19584 62158 19590 62222
rect 19654 62158 19660 62222
rect 71400 62222 71476 62430
rect 71400 62190 71406 62222
rect 19584 62152 19660 62158
rect 71405 62158 71406 62190
rect 71470 62190 71476 62222
rect 71672 62430 71678 62462
rect 71742 62462 71743 62494
rect 72488 62494 72564 62500
rect 71742 62430 71748 62462
rect 71672 62222 71748 62430
rect 71470 62158 71471 62190
rect 71405 62157 71471 62158
rect 71672 62158 71678 62222
rect 71742 62158 71748 62222
rect 72488 62430 72494 62494
rect 72558 62430 72564 62494
rect 72488 62222 72564 62430
rect 72488 62190 72494 62222
rect 71672 62152 71748 62158
rect 72493 62158 72494 62190
rect 72558 62190 72564 62222
rect 72896 62494 72972 62500
rect 72896 62430 72902 62494
rect 72966 62430 72972 62494
rect 72896 62222 72972 62430
rect 72896 62190 72902 62222
rect 72558 62158 72559 62190
rect 72493 62157 72559 62158
rect 72901 62158 72902 62190
rect 72966 62190 72972 62222
rect 72966 62158 72967 62190
rect 72901 62157 72967 62158
rect 17821 62086 17887 62087
rect 17821 62054 17822 62086
rect 17816 62022 17822 62054
rect 17886 62054 17887 62086
rect 18909 62086 18975 62087
rect 18909 62054 18910 62086
rect 17886 62022 17892 62054
rect 17816 61814 17892 62022
rect 17816 61750 17822 61814
rect 17886 61750 17892 61814
rect 17816 61744 17892 61750
rect 18904 62022 18910 62054
rect 18974 62054 18975 62086
rect 19176 62086 19252 62092
rect 18974 62022 18980 62054
rect 18904 61814 18980 62022
rect 18904 61750 18910 61814
rect 18974 61750 18980 61814
rect 19176 62022 19182 62086
rect 19246 62022 19252 62086
rect 19453 62086 19519 62087
rect 19453 62054 19454 62086
rect 19176 61814 19252 62022
rect 19176 61782 19182 61814
rect 18904 61744 18980 61750
rect 19181 61750 19182 61782
rect 19246 61782 19252 61814
rect 19448 62022 19454 62054
rect 19518 62054 19519 62086
rect 71400 62086 71476 62092
rect 19518 62022 19524 62054
rect 19448 61814 19524 62022
rect 19246 61750 19247 61782
rect 19181 61749 19247 61750
rect 19448 61750 19454 61814
rect 19518 61750 19524 61814
rect 71400 62022 71406 62086
rect 71470 62022 71476 62086
rect 71677 62086 71743 62087
rect 71677 62054 71678 62086
rect 71400 61814 71476 62022
rect 71400 61782 71406 61814
rect 19448 61744 19524 61750
rect 71405 61750 71406 61782
rect 71470 61782 71476 61814
rect 71672 62022 71678 62054
rect 71742 62054 71743 62086
rect 72085 62086 72151 62087
rect 72085 62054 72086 62086
rect 71742 62022 71748 62054
rect 71672 61814 71748 62022
rect 71470 61750 71471 61782
rect 71405 61749 71471 61750
rect 71672 61750 71678 61814
rect 71742 61750 71748 61814
rect 71672 61744 71748 61750
rect 72080 62022 72086 62054
rect 72150 62054 72151 62086
rect 72352 62086 72428 62092
rect 72150 62022 72156 62054
rect 72080 61814 72156 62022
rect 72080 61750 72086 61814
rect 72150 61750 72156 61814
rect 72352 62022 72358 62086
rect 72422 62022 72428 62086
rect 72901 62086 72967 62087
rect 72901 62054 72902 62086
rect 72352 61814 72428 62022
rect 72352 61782 72358 61814
rect 72080 61744 72156 61750
rect 72357 61750 72358 61782
rect 72422 61782 72428 61814
rect 72896 62022 72902 62054
rect 72966 62054 72967 62086
rect 72966 62022 72972 62054
rect 72896 61814 72972 62022
rect 87584 61956 87660 64470
rect 88467 62491 88527 72660
rect 89080 72558 89156 72564
rect 89080 72494 89086 72558
rect 89150 72494 89156 72558
rect 89080 71742 89156 72494
rect 89080 71710 89086 71742
rect 89085 71678 89086 71710
rect 89150 71710 89156 71742
rect 89760 72558 90108 74398
rect 89760 72494 89766 72558
rect 89830 72494 90108 72558
rect 89150 71678 89151 71710
rect 89085 71677 89151 71678
rect 89760 70926 90108 72494
rect 89760 70862 89766 70926
rect 89830 70862 90108 70926
rect 89760 69430 90108 70862
rect 89760 69366 89766 69430
rect 89830 69366 90108 69430
rect 89080 69294 89156 69300
rect 89080 69230 89086 69294
rect 89150 69230 89156 69294
rect 89080 69022 89156 69230
rect 89080 68990 89086 69022
rect 89085 68958 89086 68990
rect 89150 68990 89156 69022
rect 89150 68958 89151 68990
rect 89085 68957 89151 68958
rect 89760 67798 90108 69366
rect 89760 67734 89766 67798
rect 89830 67734 90108 67798
rect 89760 65894 90108 67734
rect 89760 65830 89766 65894
rect 89830 65830 90108 65894
rect 89760 64262 90108 65830
rect 89760 64198 89766 64262
rect 89830 64198 90108 64262
rect 89085 63174 89151 63175
rect 89085 63142 89086 63174
rect 89080 63110 89086 63142
rect 89150 63142 89151 63174
rect 89150 63110 89156 63142
rect 89080 62630 89156 63110
rect 89080 62566 89086 62630
rect 89150 62566 89156 62630
rect 89080 62560 89156 62566
rect 89760 62630 90108 64198
rect 89760 62566 89766 62630
rect 89830 62566 90108 62630
rect 88464 62490 88530 62491
rect 88464 62426 88465 62490
rect 88529 62426 88530 62490
rect 88464 62425 88530 62426
rect 87584 61950 87796 61956
rect 87584 61886 87726 61950
rect 87790 61886 87796 61950
rect 87584 61880 87796 61886
rect 72422 61750 72423 61782
rect 72357 61749 72423 61750
rect 72896 61750 72902 61814
rect 72966 61750 72972 61814
rect 72896 61744 72972 61750
rect 17821 61678 17887 61679
rect 17821 61646 17822 61678
rect 17816 61614 17822 61646
rect 17886 61646 17887 61678
rect 18229 61678 18295 61679
rect 18229 61646 18230 61678
rect 17886 61614 17892 61646
rect 17816 61406 17892 61614
rect 17816 61342 17822 61406
rect 17886 61342 17892 61406
rect 17816 61336 17892 61342
rect 18224 61614 18230 61646
rect 18294 61646 18295 61678
rect 18768 61678 18844 61684
rect 18294 61614 18300 61646
rect 18224 61406 18300 61614
rect 18224 61342 18230 61406
rect 18294 61342 18300 61406
rect 18768 61614 18774 61678
rect 18838 61614 18844 61678
rect 18768 61406 18844 61614
rect 18768 61374 18774 61406
rect 18224 61336 18300 61342
rect 18773 61342 18774 61374
rect 18838 61374 18844 61406
rect 19040 61678 19116 61684
rect 19040 61614 19046 61678
rect 19110 61614 19116 61678
rect 19453 61678 19519 61679
rect 19453 61646 19454 61678
rect 19040 61406 19116 61614
rect 19040 61374 19046 61406
rect 18838 61342 18839 61374
rect 18773 61341 18839 61342
rect 19045 61342 19046 61374
rect 19110 61374 19116 61406
rect 19448 61614 19454 61646
rect 19518 61646 19519 61678
rect 71269 61678 71335 61679
rect 71269 61646 71270 61678
rect 19518 61614 19524 61646
rect 19448 61406 19524 61614
rect 19110 61342 19111 61374
rect 19045 61341 19111 61342
rect 19448 61342 19454 61406
rect 19518 61342 19524 61406
rect 19448 61336 19524 61342
rect 71264 61614 71270 61646
rect 71334 61646 71335 61678
rect 71808 61678 71884 61684
rect 71334 61614 71340 61646
rect 71264 61406 71340 61614
rect 71264 61342 71270 61406
rect 71334 61342 71340 61406
rect 71808 61614 71814 61678
rect 71878 61614 71884 61678
rect 72221 61678 72287 61679
rect 72221 61646 72222 61678
rect 71808 61406 71884 61614
rect 71808 61374 71814 61406
rect 71264 61336 71340 61342
rect 71813 61342 71814 61374
rect 71878 61374 71884 61406
rect 72216 61614 72222 61646
rect 72286 61646 72287 61678
rect 72357 61678 72423 61679
rect 72357 61646 72358 61678
rect 72286 61614 72292 61646
rect 72216 61406 72292 61614
rect 71878 61342 71879 61374
rect 71813 61341 71879 61342
rect 72216 61342 72222 61406
rect 72286 61342 72292 61406
rect 72216 61336 72292 61342
rect 72352 61614 72358 61646
rect 72422 61646 72423 61678
rect 73032 61678 73108 61684
rect 72422 61614 72428 61646
rect 72352 61406 72428 61614
rect 72352 61342 72358 61406
rect 72422 61342 72428 61406
rect 73032 61614 73038 61678
rect 73102 61614 73108 61678
rect 73032 61406 73108 61614
rect 73032 61374 73038 61406
rect 72352 61336 72428 61342
rect 73037 61342 73038 61374
rect 73102 61374 73108 61406
rect 73102 61342 73103 61374
rect 73037 61341 73103 61342
rect 17952 61270 18028 61276
rect 17952 61206 17958 61270
rect 18022 61206 18028 61270
rect 17952 60998 18028 61206
rect 17952 60966 17958 60998
rect 17957 60934 17958 60966
rect 18022 60966 18028 60998
rect 18360 61270 18436 61276
rect 18360 61206 18366 61270
rect 18430 61206 18436 61270
rect 18360 60998 18436 61206
rect 18360 60966 18366 60998
rect 18022 60934 18023 60966
rect 17957 60933 18023 60934
rect 18365 60934 18366 60966
rect 18430 60966 18436 60998
rect 18768 61270 18844 61276
rect 18768 61206 18774 61270
rect 18838 61206 18844 61270
rect 19045 61270 19111 61271
rect 19045 61238 19046 61270
rect 18768 60998 18844 61206
rect 18768 60966 18774 60998
rect 18430 60934 18431 60966
rect 18365 60933 18431 60934
rect 18773 60934 18774 60966
rect 18838 60966 18844 60998
rect 19040 61206 19046 61238
rect 19110 61238 19111 61270
rect 19589 61270 19655 61271
rect 19589 61238 19590 61270
rect 19110 61206 19116 61238
rect 19040 60998 19116 61206
rect 18838 60934 18839 60966
rect 18773 60933 18839 60934
rect 19040 60934 19046 60998
rect 19110 60934 19116 60998
rect 19040 60928 19116 60934
rect 19584 61206 19590 61238
rect 19654 61238 19655 61270
rect 71400 61270 71476 61276
rect 19654 61206 19660 61238
rect 19584 60998 19660 61206
rect 19584 60934 19590 60998
rect 19654 60934 19660 60998
rect 71400 61206 71406 61270
rect 71470 61206 71476 61270
rect 71813 61270 71879 61271
rect 71813 61238 71814 61270
rect 71400 60998 71476 61206
rect 71400 60966 71406 60998
rect 19584 60928 19660 60934
rect 71405 60934 71406 60966
rect 71470 60966 71476 60998
rect 71808 61206 71814 61238
rect 71878 61238 71879 61270
rect 72080 61270 72156 61276
rect 71878 61206 71884 61238
rect 71808 60998 71884 61206
rect 71470 60934 71471 60966
rect 71405 60933 71471 60934
rect 71808 60934 71814 60998
rect 71878 60934 71884 60998
rect 72080 61206 72086 61270
rect 72150 61206 72156 61270
rect 72629 61270 72695 61271
rect 72629 61238 72630 61270
rect 72080 60998 72156 61206
rect 72080 60966 72086 60998
rect 71808 60928 71884 60934
rect 72085 60934 72086 60966
rect 72150 60966 72156 60998
rect 72624 61206 72630 61238
rect 72694 61238 72695 61270
rect 73037 61270 73103 61271
rect 73037 61238 73038 61270
rect 72694 61206 72700 61238
rect 72624 60998 72700 61206
rect 72150 60934 72151 60966
rect 72085 60933 72151 60934
rect 72624 60934 72630 60998
rect 72694 60934 72700 60998
rect 72624 60928 72700 60934
rect 73032 61206 73038 61238
rect 73102 61238 73103 61270
rect 73102 61206 73108 61238
rect 73032 60998 73108 61206
rect 73032 60934 73038 60998
rect 73102 60934 73108 60998
rect 73032 60928 73108 60934
rect 89760 60998 90108 62566
rect 89760 60934 89766 60998
rect 89830 60934 90108 60998
rect 952 60798 1230 60862
rect 1294 60798 1300 60862
rect 18637 60862 18703 60863
rect 18637 60830 18638 60862
rect 952 59230 1300 60798
rect 18632 60798 18638 60830
rect 18702 60830 18703 60862
rect 19040 60862 19116 60868
rect 18702 60798 18708 60830
rect 18632 60590 18708 60798
rect 18632 60526 18638 60590
rect 18702 60526 18708 60590
rect 19040 60798 19046 60862
rect 19110 60798 19116 60862
rect 19040 60590 19116 60798
rect 19040 60558 19046 60590
rect 18632 60520 18708 60526
rect 19045 60526 19046 60558
rect 19110 60558 19116 60590
rect 19448 60862 19524 60868
rect 19448 60798 19454 60862
rect 19518 60798 19524 60862
rect 19448 60590 19524 60798
rect 19448 60558 19454 60590
rect 19110 60526 19111 60558
rect 19045 60525 19111 60526
rect 19453 60526 19454 60558
rect 19518 60558 19524 60590
rect 71264 60862 71340 60868
rect 71264 60798 71270 60862
rect 71334 60798 71340 60862
rect 71264 60590 71340 60798
rect 71264 60558 71270 60590
rect 19518 60526 19519 60558
rect 19453 60525 19519 60526
rect 71269 60526 71270 60558
rect 71334 60558 71340 60590
rect 71672 60862 71748 60868
rect 71672 60798 71678 60862
rect 71742 60798 71748 60862
rect 71672 60590 71748 60798
rect 71672 60558 71678 60590
rect 71334 60526 71335 60558
rect 71269 60525 71335 60526
rect 71677 60526 71678 60558
rect 71742 60558 71748 60590
rect 71742 60526 71743 60558
rect 71677 60525 71743 60526
rect 17952 60454 18028 60460
rect 17952 60390 17958 60454
rect 18022 60390 18028 60454
rect 18229 60454 18295 60455
rect 18229 60422 18230 60454
rect 17952 60182 18028 60390
rect 17952 60150 17958 60182
rect 17957 60118 17958 60150
rect 18022 60150 18028 60182
rect 18224 60390 18230 60422
rect 18294 60422 18295 60454
rect 18904 60454 18980 60460
rect 18294 60390 18300 60422
rect 18224 60182 18300 60390
rect 18022 60118 18023 60150
rect 17957 60117 18023 60118
rect 18224 60118 18230 60182
rect 18294 60118 18300 60182
rect 18904 60390 18910 60454
rect 18974 60390 18980 60454
rect 18904 60182 18980 60390
rect 18904 60150 18910 60182
rect 18224 60112 18300 60118
rect 18909 60118 18910 60150
rect 18974 60150 18980 60182
rect 19040 60454 19116 60460
rect 19040 60390 19046 60454
rect 19110 60390 19116 60454
rect 19453 60454 19519 60455
rect 19453 60422 19454 60454
rect 19040 60182 19116 60390
rect 19040 60150 19046 60182
rect 18974 60118 18975 60150
rect 18909 60117 18975 60118
rect 19045 60118 19046 60150
rect 19110 60150 19116 60182
rect 19448 60390 19454 60422
rect 19518 60422 19519 60454
rect 71269 60454 71335 60455
rect 71269 60422 71270 60454
rect 19518 60390 19524 60422
rect 19448 60182 19524 60390
rect 19110 60118 19111 60150
rect 19045 60117 19111 60118
rect 19448 60118 19454 60182
rect 19518 60118 19524 60182
rect 19448 60112 19524 60118
rect 71264 60390 71270 60422
rect 71334 60422 71335 60454
rect 71677 60454 71743 60455
rect 71677 60422 71678 60454
rect 71334 60390 71340 60422
rect 71264 60182 71340 60390
rect 71264 60118 71270 60182
rect 71334 60118 71340 60182
rect 71264 60112 71340 60118
rect 71672 60390 71678 60422
rect 71742 60422 71743 60454
rect 72221 60454 72287 60455
rect 72221 60422 72222 60454
rect 71742 60390 71748 60422
rect 71672 60182 71748 60390
rect 71672 60118 71678 60182
rect 71742 60118 71748 60182
rect 71672 60112 71748 60118
rect 72216 60390 72222 60422
rect 72286 60422 72287 60454
rect 72629 60454 72695 60455
rect 72629 60422 72630 60454
rect 72286 60390 72292 60422
rect 72216 60182 72292 60390
rect 72216 60118 72222 60182
rect 72286 60118 72292 60182
rect 72216 60112 72292 60118
rect 72624 60390 72630 60422
rect 72694 60422 72695 60454
rect 73032 60454 73108 60460
rect 72694 60390 72700 60422
rect 72624 60182 72700 60390
rect 72624 60118 72630 60182
rect 72694 60118 72700 60182
rect 73032 60390 73038 60454
rect 73102 60390 73108 60454
rect 73032 60182 73108 60390
rect 73032 60150 73038 60182
rect 72624 60112 72700 60118
rect 73037 60118 73038 60150
rect 73102 60150 73108 60182
rect 73102 60118 73103 60150
rect 73037 60117 73103 60118
rect 18365 60046 18431 60047
rect 18365 60014 18366 60046
rect 18360 59982 18366 60014
rect 18430 60014 18431 60046
rect 18501 60046 18567 60047
rect 18501 60014 18502 60046
rect 18430 59982 18436 60014
rect 17821 59774 17887 59775
rect 17821 59742 17822 59774
rect 17816 59710 17822 59742
rect 17886 59742 17887 59774
rect 18360 59774 18436 59982
rect 17886 59710 17892 59742
rect 17816 59502 17892 59710
rect 18360 59710 18366 59774
rect 18430 59710 18436 59774
rect 18360 59704 18436 59710
rect 18496 59982 18502 60014
rect 18566 60014 18567 60046
rect 18768 60046 18844 60052
rect 18566 59982 18572 60014
rect 18496 59774 18572 59982
rect 18496 59710 18502 59774
rect 18566 59710 18572 59774
rect 18768 59982 18774 60046
rect 18838 59982 18844 60046
rect 19181 60046 19247 60047
rect 19181 60014 19182 60046
rect 18768 59774 18844 59982
rect 18768 59742 18774 59774
rect 18496 59704 18572 59710
rect 18773 59710 18774 59742
rect 18838 59742 18844 59774
rect 19176 59982 19182 60014
rect 19246 60014 19247 60046
rect 19453 60046 19519 60047
rect 19453 60014 19454 60046
rect 19246 59982 19252 60014
rect 19176 59774 19252 59982
rect 18838 59710 18839 59742
rect 18773 59709 18839 59710
rect 19176 59710 19182 59774
rect 19246 59710 19252 59774
rect 19176 59704 19252 59710
rect 19448 59982 19454 60014
rect 19518 60014 19519 60046
rect 71405 60046 71471 60047
rect 71405 60014 71406 60046
rect 19518 59982 19524 60014
rect 19448 59774 19524 59982
rect 71400 59982 71406 60014
rect 71470 60014 71471 60046
rect 71677 60046 71743 60047
rect 71677 60014 71678 60046
rect 71470 59982 71476 60014
rect 24621 59910 24687 59911
rect 24621 59878 24622 59910
rect 19448 59710 19454 59774
rect 19518 59710 19524 59774
rect 19448 59704 19524 59710
rect 24616 59846 24622 59878
rect 24686 59878 24687 59910
rect 66373 59910 66439 59911
rect 66373 59878 66374 59910
rect 24686 59846 24692 59878
rect 19181 59638 19247 59639
rect 19181 59606 19182 59638
rect 17816 59438 17822 59502
rect 17886 59438 17892 59502
rect 17816 59432 17892 59438
rect 19176 59574 19182 59606
rect 19246 59606 19247 59638
rect 19584 59638 19660 59644
rect 19246 59574 19252 59606
rect 19176 59366 19252 59574
rect 19176 59302 19182 59366
rect 19246 59302 19252 59366
rect 19584 59574 19590 59638
rect 19654 59574 19660 59638
rect 19584 59366 19660 59574
rect 24616 59638 24692 59846
rect 24616 59574 24622 59638
rect 24686 59574 24692 59638
rect 24616 59568 24692 59574
rect 66368 59846 66374 59878
rect 66438 59878 66439 59910
rect 66438 59846 66444 59878
rect 66368 59638 66444 59846
rect 71400 59774 71476 59982
rect 71400 59710 71406 59774
rect 71470 59710 71476 59774
rect 71400 59704 71476 59710
rect 71672 59982 71678 60014
rect 71742 60014 71743 60046
rect 72085 60046 72151 60047
rect 72085 60014 72086 60046
rect 71742 59982 71748 60014
rect 71672 59774 71748 59982
rect 71672 59710 71678 59774
rect 71742 59710 71748 59774
rect 71672 59704 71748 59710
rect 72080 59982 72086 60014
rect 72150 60014 72151 60046
rect 72150 59982 72156 60014
rect 72080 59774 72156 59982
rect 72080 59710 72086 59774
rect 72150 59710 72156 59774
rect 72080 59704 72156 59710
rect 72896 59774 72972 59780
rect 72896 59710 72902 59774
rect 72966 59710 72972 59774
rect 66368 59574 66374 59638
rect 66438 59574 66444 59638
rect 66509 59638 66575 59639
rect 66509 59606 66510 59638
rect 66368 59568 66444 59574
rect 66504 59574 66510 59606
rect 66574 59606 66575 59638
rect 71264 59638 71340 59644
rect 66574 59574 66580 59606
rect 19584 59334 19590 59366
rect 19176 59296 19252 59302
rect 19589 59302 19590 59334
rect 19654 59334 19660 59366
rect 19654 59302 19655 59334
rect 19589 59301 19655 59302
rect 952 59166 1230 59230
rect 1294 59166 1300 59230
rect 18909 59230 18975 59231
rect 18909 59198 18910 59230
rect 952 57462 1300 59166
rect 18904 59166 18910 59198
rect 18974 59198 18975 59230
rect 66504 59230 66580 59574
rect 71264 59574 71270 59638
rect 71334 59574 71340 59638
rect 71264 59366 71340 59574
rect 71264 59334 71270 59366
rect 71269 59302 71270 59334
rect 71334 59334 71340 59366
rect 71808 59638 71884 59644
rect 71808 59574 71814 59638
rect 71878 59574 71884 59638
rect 71808 59366 71884 59574
rect 72896 59502 72972 59710
rect 72896 59470 72902 59502
rect 72901 59438 72902 59470
rect 72966 59470 72972 59502
rect 72966 59438 72967 59470
rect 72901 59437 72967 59438
rect 71808 59334 71814 59366
rect 71334 59302 71335 59334
rect 71269 59301 71335 59302
rect 71813 59302 71814 59334
rect 71878 59334 71884 59366
rect 71878 59302 71879 59334
rect 71813 59301 71879 59302
rect 18974 59166 18980 59198
rect 17821 58958 17887 58959
rect 17821 58926 17822 58958
rect 17816 58894 17822 58926
rect 17886 58926 17887 58958
rect 18904 58958 18980 59166
rect 66504 59166 66510 59230
rect 66574 59166 66580 59230
rect 72357 59230 72423 59231
rect 72357 59198 72358 59230
rect 66504 59160 66580 59166
rect 72352 59166 72358 59198
rect 72422 59198 72423 59230
rect 89760 59230 90108 60934
rect 72422 59166 72428 59198
rect 17886 58894 17892 58926
rect 17816 58686 17892 58894
rect 18904 58894 18910 58958
rect 18974 58894 18980 58958
rect 18904 58888 18980 58894
rect 66368 59094 66444 59100
rect 66368 59030 66374 59094
rect 66438 59030 66444 59094
rect 17816 58622 17822 58686
rect 17886 58622 17892 58686
rect 17816 58616 17892 58622
rect 18496 58822 18572 58828
rect 18496 58758 18502 58822
rect 18566 58758 18572 58822
rect 66368 58822 66444 59030
rect 72352 58958 72428 59166
rect 89760 59166 89766 59230
rect 89830 59166 90108 59230
rect 72352 58894 72358 58958
rect 72422 58894 72428 58958
rect 72352 58888 72428 58894
rect 72896 58958 72972 58964
rect 72896 58894 72902 58958
rect 72966 58894 72972 58958
rect 66368 58790 66374 58822
rect 17816 58550 17892 58556
rect 17816 58486 17822 58550
rect 17886 58486 17892 58550
rect 18496 58550 18572 58758
rect 66373 58758 66374 58790
rect 66438 58790 66444 58822
rect 66438 58758 66439 58790
rect 66373 58757 66439 58758
rect 24344 58686 24420 58692
rect 24344 58622 24350 58686
rect 24414 58622 24420 58686
rect 18496 58518 18502 58550
rect 17816 58278 17892 58486
rect 18501 58486 18502 58518
rect 18566 58518 18572 58550
rect 18773 58550 18839 58551
rect 18773 58518 18774 58550
rect 18566 58486 18567 58518
rect 18501 58485 18567 58486
rect 18768 58486 18774 58518
rect 18838 58518 18839 58550
rect 18838 58486 18844 58518
rect 17816 58246 17822 58278
rect 17821 58214 17822 58246
rect 17886 58246 17892 58278
rect 18768 58278 18844 58486
rect 24344 58414 24420 58622
rect 24344 58382 24350 58414
rect 24349 58350 24350 58382
rect 24414 58382 24420 58414
rect 66504 58686 66580 58692
rect 66504 58622 66510 58686
rect 66574 58622 66580 58686
rect 72896 58686 72972 58894
rect 72896 58654 72902 58686
rect 66504 58414 66580 58622
rect 72901 58622 72902 58654
rect 72966 58654 72972 58686
rect 72966 58622 72967 58654
rect 72901 58621 72967 58622
rect 72085 58550 72151 58551
rect 72085 58518 72086 58550
rect 66504 58382 66510 58414
rect 24414 58350 24415 58382
rect 24349 58349 24415 58350
rect 66509 58350 66510 58382
rect 66574 58382 66580 58414
rect 72080 58486 72086 58518
rect 72150 58518 72151 58550
rect 72352 58550 72428 58556
rect 72150 58486 72156 58518
rect 66574 58350 66575 58382
rect 66509 58349 66575 58350
rect 17886 58214 17887 58246
rect 17821 58213 17887 58214
rect 18768 58214 18774 58278
rect 18838 58214 18844 58278
rect 18768 58208 18844 58214
rect 72080 58278 72156 58486
rect 72080 58214 72086 58278
rect 72150 58214 72156 58278
rect 72352 58486 72358 58550
rect 72422 58486 72428 58550
rect 72352 58278 72428 58486
rect 72352 58246 72358 58278
rect 72080 58208 72156 58214
rect 72357 58214 72358 58246
rect 72422 58246 72428 58278
rect 73032 58550 73108 58556
rect 73032 58486 73038 58550
rect 73102 58486 73108 58550
rect 73032 58278 73108 58486
rect 73032 58246 73038 58278
rect 72422 58214 72423 58246
rect 72357 58213 72423 58214
rect 73037 58214 73038 58246
rect 73102 58246 73108 58278
rect 73102 58214 73103 58246
rect 73037 58213 73103 58214
rect 17816 58142 17892 58148
rect 17816 58078 17822 58142
rect 17886 58078 17892 58142
rect 19045 58142 19111 58143
rect 19045 58110 19046 58142
rect 17816 57870 17892 58078
rect 17816 57838 17822 57870
rect 17821 57806 17822 57838
rect 17886 57838 17892 57870
rect 19040 58078 19046 58110
rect 19110 58110 19111 58142
rect 19448 58142 19524 58148
rect 19110 58078 19116 58110
rect 19040 57870 19116 58078
rect 17886 57806 17887 57838
rect 17821 57805 17887 57806
rect 19040 57806 19046 57870
rect 19110 57806 19116 57870
rect 19448 58078 19454 58142
rect 19518 58078 19524 58142
rect 71269 58142 71335 58143
rect 71269 58110 71270 58142
rect 19448 57870 19524 58078
rect 19448 57838 19454 57870
rect 19040 57800 19116 57806
rect 19453 57806 19454 57838
rect 19518 57838 19524 57870
rect 71264 58078 71270 58110
rect 71334 58110 71335 58142
rect 71813 58142 71879 58143
rect 71813 58110 71814 58142
rect 71334 58078 71340 58110
rect 71264 57870 71340 58078
rect 19518 57806 19519 57838
rect 19453 57805 19519 57806
rect 71264 57806 71270 57870
rect 71334 57806 71340 57870
rect 71264 57800 71340 57806
rect 71808 58078 71814 58110
rect 71878 58110 71879 58142
rect 72896 58142 72972 58148
rect 71878 58078 71884 58110
rect 71808 57870 71884 58078
rect 71808 57806 71814 57870
rect 71878 57806 71884 57870
rect 72896 58078 72902 58142
rect 72966 58078 72972 58142
rect 72896 57870 72972 58078
rect 72896 57838 72902 57870
rect 71808 57800 71884 57806
rect 72901 57806 72902 57838
rect 72966 57838 72972 57870
rect 72966 57806 72967 57838
rect 72901 57805 72967 57806
rect 17821 57734 17887 57735
rect 17821 57702 17822 57734
rect 952 57398 1230 57462
rect 1294 57398 1300 57462
rect 952 55830 1300 57398
rect 17816 57670 17822 57702
rect 17886 57702 17887 57734
rect 18632 57734 18708 57740
rect 17886 57670 17892 57702
rect 17816 57462 17892 57670
rect 17816 57398 17822 57462
rect 17886 57398 17892 57462
rect 18632 57670 18638 57734
rect 18702 57670 18708 57734
rect 18632 57462 18708 57670
rect 18632 57430 18638 57462
rect 17816 57392 17892 57398
rect 18637 57398 18638 57430
rect 18702 57430 18708 57462
rect 19176 57734 19252 57740
rect 19176 57670 19182 57734
rect 19246 57670 19252 57734
rect 19453 57734 19519 57735
rect 19453 57702 19454 57734
rect 19176 57462 19252 57670
rect 19176 57430 19182 57462
rect 18702 57398 18703 57430
rect 18637 57397 18703 57398
rect 19181 57398 19182 57430
rect 19246 57430 19252 57462
rect 19448 57670 19454 57702
rect 19518 57702 19519 57734
rect 71405 57734 71471 57735
rect 71405 57702 71406 57734
rect 19518 57670 19524 57702
rect 19448 57462 19524 57670
rect 19246 57398 19247 57430
rect 19181 57397 19247 57398
rect 19448 57398 19454 57462
rect 19518 57398 19524 57462
rect 19448 57392 19524 57398
rect 71400 57670 71406 57702
rect 71470 57702 71471 57734
rect 71808 57734 71884 57740
rect 71470 57670 71476 57702
rect 71400 57462 71476 57670
rect 71400 57398 71406 57462
rect 71470 57398 71476 57462
rect 71808 57670 71814 57734
rect 71878 57670 71884 57734
rect 71808 57462 71884 57670
rect 71808 57430 71814 57462
rect 71400 57392 71476 57398
rect 71813 57398 71814 57430
rect 71878 57430 71884 57462
rect 72352 57734 72428 57740
rect 72352 57670 72358 57734
rect 72422 57670 72428 57734
rect 72901 57734 72967 57735
rect 72901 57702 72902 57734
rect 72352 57462 72428 57670
rect 72352 57430 72358 57462
rect 71878 57398 71879 57430
rect 71813 57397 71879 57398
rect 72357 57398 72358 57430
rect 72422 57430 72428 57462
rect 72896 57670 72902 57702
rect 72966 57702 72967 57734
rect 72966 57670 72972 57702
rect 72896 57462 72972 57670
rect 72422 57398 72423 57430
rect 72357 57397 72423 57398
rect 72896 57398 72902 57462
rect 72966 57398 72972 57462
rect 72896 57392 72972 57398
rect 89760 57462 90108 59166
rect 89760 57398 89766 57462
rect 89830 57398 90108 57462
rect 17821 57326 17887 57327
rect 17821 57294 17822 57326
rect 17816 57262 17822 57294
rect 17886 57294 17887 57326
rect 18229 57326 18295 57327
rect 18229 57294 18230 57326
rect 17886 57262 17892 57294
rect 17816 57054 17892 57262
rect 17816 56990 17822 57054
rect 17886 56990 17892 57054
rect 17816 56984 17892 56990
rect 18224 57262 18230 57294
rect 18294 57294 18295 57326
rect 19045 57326 19111 57327
rect 19045 57294 19046 57326
rect 18294 57262 18300 57294
rect 18224 57054 18300 57262
rect 18224 56990 18230 57054
rect 18294 56990 18300 57054
rect 18224 56984 18300 56990
rect 19040 57262 19046 57294
rect 19110 57294 19111 57326
rect 19584 57326 19660 57332
rect 19110 57262 19116 57294
rect 19040 57054 19116 57262
rect 19040 56990 19046 57054
rect 19110 56990 19116 57054
rect 19584 57262 19590 57326
rect 19654 57262 19660 57326
rect 19584 57054 19660 57262
rect 19584 57022 19590 57054
rect 19040 56984 19116 56990
rect 19589 56990 19590 57022
rect 19654 57022 19660 57054
rect 71264 57326 71340 57332
rect 71264 57262 71270 57326
rect 71334 57262 71340 57326
rect 71264 57054 71340 57262
rect 71264 57022 71270 57054
rect 19654 56990 19655 57022
rect 19589 56989 19655 56990
rect 71269 56990 71270 57022
rect 71334 57022 71340 57054
rect 71808 57326 71884 57332
rect 71808 57262 71814 57326
rect 71878 57262 71884 57326
rect 71808 57054 71884 57262
rect 71808 57022 71814 57054
rect 71334 56990 71335 57022
rect 71269 56989 71335 56990
rect 71813 56990 71814 57022
rect 71878 57022 71884 57054
rect 72216 57326 72292 57332
rect 72216 57262 72222 57326
rect 72286 57262 72292 57326
rect 73037 57326 73103 57327
rect 73037 57294 73038 57326
rect 72216 57054 72292 57262
rect 72216 57022 72222 57054
rect 71878 56990 71879 57022
rect 71813 56989 71879 56990
rect 72221 56990 72222 57022
rect 72286 57022 72292 57054
rect 73032 57262 73038 57294
rect 73102 57294 73103 57326
rect 73102 57262 73108 57294
rect 73032 57054 73108 57262
rect 72286 56990 72287 57022
rect 72221 56989 72287 56990
rect 73032 56990 73038 57054
rect 73102 56990 73108 57054
rect 73032 56984 73108 56990
rect 17957 56918 18023 56919
rect 17957 56886 17958 56918
rect 17952 56854 17958 56886
rect 18022 56886 18023 56918
rect 18360 56918 18436 56924
rect 18022 56854 18028 56886
rect 17952 56646 18028 56854
rect 17952 56582 17958 56646
rect 18022 56582 18028 56646
rect 18360 56854 18366 56918
rect 18430 56854 18436 56918
rect 18360 56646 18436 56854
rect 18360 56614 18366 56646
rect 17952 56576 18028 56582
rect 18365 56582 18366 56614
rect 18430 56614 18436 56646
rect 18496 56918 18572 56924
rect 18496 56854 18502 56918
rect 18566 56854 18572 56918
rect 18496 56646 18572 56854
rect 18496 56614 18502 56646
rect 18430 56582 18431 56614
rect 18365 56581 18431 56582
rect 18501 56582 18502 56614
rect 18566 56614 18572 56646
rect 19176 56918 19252 56924
rect 19176 56854 19182 56918
rect 19246 56854 19252 56918
rect 19589 56918 19655 56919
rect 19589 56886 19590 56918
rect 19176 56646 19252 56854
rect 19176 56614 19182 56646
rect 18566 56582 18567 56614
rect 18501 56581 18567 56582
rect 19181 56582 19182 56614
rect 19246 56614 19252 56646
rect 19584 56854 19590 56886
rect 19654 56886 19655 56918
rect 71269 56918 71335 56919
rect 71269 56886 71270 56918
rect 19654 56854 19660 56886
rect 19584 56646 19660 56854
rect 19246 56582 19247 56614
rect 19181 56581 19247 56582
rect 19584 56582 19590 56646
rect 19654 56582 19660 56646
rect 19584 56576 19660 56582
rect 71264 56854 71270 56886
rect 71334 56886 71335 56918
rect 71672 56918 71748 56924
rect 71334 56854 71340 56886
rect 71264 56646 71340 56854
rect 71264 56582 71270 56646
rect 71334 56582 71340 56646
rect 71672 56854 71678 56918
rect 71742 56854 71748 56918
rect 71672 56646 71748 56854
rect 71672 56614 71678 56646
rect 71264 56576 71340 56582
rect 71677 56582 71678 56614
rect 71742 56614 71748 56646
rect 72080 56918 72156 56924
rect 72080 56854 72086 56918
rect 72150 56854 72156 56918
rect 72080 56646 72156 56854
rect 72080 56614 72086 56646
rect 71742 56582 71743 56614
rect 71677 56581 71743 56582
rect 72085 56582 72086 56614
rect 72150 56614 72156 56646
rect 72488 56918 72564 56924
rect 72488 56854 72494 56918
rect 72558 56854 72564 56918
rect 72488 56646 72564 56854
rect 72488 56614 72494 56646
rect 72150 56582 72151 56614
rect 72085 56581 72151 56582
rect 72493 56582 72494 56614
rect 72558 56614 72564 56646
rect 72896 56918 72972 56924
rect 72896 56854 72902 56918
rect 72966 56854 72972 56918
rect 72896 56646 72972 56854
rect 72896 56614 72902 56646
rect 72558 56582 72559 56614
rect 72493 56581 72559 56582
rect 72901 56582 72902 56614
rect 72966 56614 72972 56646
rect 72966 56582 72967 56614
rect 72901 56581 72967 56582
rect 17816 56510 17892 56516
rect 17816 56446 17822 56510
rect 17886 56446 17892 56510
rect 18365 56510 18431 56511
rect 18365 56478 18366 56510
rect 17816 56238 17892 56446
rect 17816 56206 17822 56238
rect 17821 56174 17822 56206
rect 17886 56206 17892 56238
rect 18360 56446 18366 56478
rect 18430 56478 18431 56510
rect 18501 56510 18567 56511
rect 18501 56478 18502 56510
rect 18430 56446 18436 56478
rect 18360 56238 18436 56446
rect 17886 56174 17887 56206
rect 17821 56173 17887 56174
rect 18360 56174 18366 56238
rect 18430 56174 18436 56238
rect 18360 56168 18436 56174
rect 18496 56446 18502 56478
rect 18566 56478 18567 56510
rect 19181 56510 19247 56511
rect 19181 56478 19182 56510
rect 18566 56446 18572 56478
rect 18496 56238 18572 56446
rect 18496 56174 18502 56238
rect 18566 56174 18572 56238
rect 18496 56168 18572 56174
rect 19176 56446 19182 56478
rect 19246 56478 19247 56510
rect 19589 56510 19655 56511
rect 19589 56478 19590 56510
rect 19246 56446 19252 56478
rect 19176 56238 19252 56446
rect 19176 56174 19182 56238
rect 19246 56174 19252 56238
rect 19176 56168 19252 56174
rect 19584 56446 19590 56478
rect 19654 56478 19655 56510
rect 71405 56510 71471 56511
rect 71405 56478 71406 56510
rect 19654 56446 19660 56478
rect 19584 56238 19660 56446
rect 19584 56174 19590 56238
rect 19654 56174 19660 56238
rect 19584 56168 19660 56174
rect 71400 56446 71406 56478
rect 71470 56478 71471 56510
rect 71677 56510 71743 56511
rect 71677 56478 71678 56510
rect 71470 56446 71476 56478
rect 71400 56238 71476 56446
rect 71400 56174 71406 56238
rect 71470 56174 71476 56238
rect 71400 56168 71476 56174
rect 71672 56446 71678 56478
rect 71742 56478 71743 56510
rect 72352 56510 72428 56516
rect 71742 56446 71748 56478
rect 71672 56238 71748 56446
rect 71672 56174 71678 56238
rect 71742 56174 71748 56238
rect 72352 56446 72358 56510
rect 72422 56446 72428 56510
rect 72901 56510 72967 56511
rect 72901 56478 72902 56510
rect 72352 56238 72428 56446
rect 72352 56206 72358 56238
rect 71672 56168 71748 56174
rect 72357 56174 72358 56206
rect 72422 56206 72428 56238
rect 72896 56446 72902 56478
rect 72966 56478 72967 56510
rect 72966 56446 72972 56478
rect 72896 56238 72972 56446
rect 72422 56174 72423 56206
rect 72357 56173 72423 56174
rect 72896 56174 72902 56238
rect 72966 56174 72972 56238
rect 72896 56168 72972 56174
rect 18909 56102 18975 56103
rect 18909 56070 18910 56102
rect 952 55766 1230 55830
rect 1294 55766 1300 55830
rect 952 54198 1300 55766
rect 18904 56038 18910 56070
rect 18974 56070 18975 56102
rect 19040 56102 19116 56108
rect 18974 56038 18980 56070
rect 18904 55830 18980 56038
rect 18904 55766 18910 55830
rect 18974 55766 18980 55830
rect 19040 56038 19046 56102
rect 19110 56038 19116 56102
rect 19040 55830 19116 56038
rect 19040 55798 19046 55830
rect 18904 55760 18980 55766
rect 19045 55766 19046 55798
rect 19110 55798 19116 55830
rect 19584 56102 19660 56108
rect 19584 56038 19590 56102
rect 19654 56038 19660 56102
rect 19584 55830 19660 56038
rect 19584 55798 19590 55830
rect 19110 55766 19111 55798
rect 19045 55765 19111 55766
rect 19589 55766 19590 55798
rect 19654 55798 19660 55830
rect 71264 56102 71340 56108
rect 71264 56038 71270 56102
rect 71334 56038 71340 56102
rect 71677 56102 71743 56103
rect 71677 56070 71678 56102
rect 71264 55830 71340 56038
rect 71264 55798 71270 55830
rect 19654 55766 19655 55798
rect 19589 55765 19655 55766
rect 71269 55766 71270 55798
rect 71334 55798 71340 55830
rect 71672 56038 71678 56070
rect 71742 56070 71743 56102
rect 72629 56102 72695 56103
rect 72629 56070 72630 56102
rect 71742 56038 71748 56070
rect 71672 55830 71748 56038
rect 71334 55766 71335 55798
rect 71269 55765 71335 55766
rect 71672 55766 71678 55830
rect 71742 55766 71748 55830
rect 71672 55760 71748 55766
rect 72624 56038 72630 56070
rect 72694 56070 72695 56102
rect 72694 56038 72700 56070
rect 72624 55830 72700 56038
rect 72624 55766 72630 55830
rect 72694 55766 72700 55830
rect 72624 55760 72700 55766
rect 89760 55830 90108 57398
rect 89760 55766 89766 55830
rect 89830 55766 90108 55830
rect 19176 55694 19252 55700
rect 19176 55630 19182 55694
rect 19246 55630 19252 55694
rect 19176 55422 19252 55630
rect 19176 55390 19182 55422
rect 19181 55358 19182 55390
rect 19246 55390 19252 55422
rect 19584 55694 19660 55700
rect 19584 55630 19590 55694
rect 19654 55630 19660 55694
rect 71405 55694 71471 55695
rect 71405 55662 71406 55694
rect 19584 55422 19660 55630
rect 19584 55390 19590 55422
rect 19246 55358 19247 55390
rect 19181 55357 19247 55358
rect 19589 55358 19590 55390
rect 19654 55390 19660 55422
rect 71400 55630 71406 55662
rect 71470 55662 71471 55694
rect 71808 55694 71884 55700
rect 71470 55630 71476 55662
rect 71400 55422 71476 55630
rect 19654 55358 19655 55390
rect 19589 55357 19655 55358
rect 71400 55358 71406 55422
rect 71470 55358 71476 55422
rect 71808 55630 71814 55694
rect 71878 55630 71884 55694
rect 71808 55422 71884 55630
rect 71808 55390 71814 55422
rect 71400 55352 71476 55358
rect 71813 55358 71814 55390
rect 71878 55390 71884 55422
rect 71878 55358 71879 55390
rect 71813 55357 71879 55358
rect 18632 55286 18708 55292
rect 18632 55222 18638 55286
rect 18702 55222 18708 55286
rect 17952 55014 18028 55020
rect 17952 54950 17958 55014
rect 18022 54950 18028 55014
rect 18632 55014 18708 55222
rect 72216 55286 72292 55292
rect 72216 55222 72222 55286
rect 72286 55222 72292 55286
rect 18632 54982 18638 55014
rect 17952 54742 18028 54950
rect 18637 54950 18638 54982
rect 18702 54982 18708 55014
rect 66504 55150 66580 55156
rect 66504 55086 66510 55150
rect 66574 55086 66580 55150
rect 18702 54950 18703 54982
rect 18637 54949 18703 54950
rect 66504 54878 66580 55086
rect 72216 55014 72292 55222
rect 72216 54982 72222 55014
rect 72221 54950 72222 54982
rect 72286 54982 72292 55014
rect 72352 55286 72428 55292
rect 72352 55222 72358 55286
rect 72422 55222 72428 55286
rect 72352 55014 72428 55222
rect 72352 54982 72358 55014
rect 72286 54950 72287 54982
rect 72221 54949 72287 54950
rect 72357 54950 72358 54982
rect 72422 54982 72428 55014
rect 73032 55014 73108 55020
rect 72422 54950 72423 54982
rect 72357 54949 72423 54950
rect 73032 54950 73038 55014
rect 73102 54950 73108 55014
rect 66504 54846 66510 54878
rect 66509 54814 66510 54846
rect 66574 54846 66580 54878
rect 66574 54814 66575 54846
rect 66509 54813 66575 54814
rect 17952 54710 17958 54742
rect 17957 54678 17958 54710
rect 18022 54710 18028 54742
rect 24616 54742 24692 54748
rect 18022 54678 18023 54710
rect 17957 54677 18023 54678
rect 24616 54678 24622 54742
rect 24686 54678 24692 54742
rect 66509 54742 66575 54743
rect 66509 54710 66510 54742
rect 17821 54606 17887 54607
rect 17821 54574 17822 54606
rect 17816 54542 17822 54574
rect 17886 54574 17887 54606
rect 18365 54606 18431 54607
rect 18365 54574 18366 54606
rect 17886 54542 17892 54574
rect 17816 54334 17892 54542
rect 17816 54270 17822 54334
rect 17886 54270 17892 54334
rect 17816 54264 17892 54270
rect 18360 54542 18366 54574
rect 18430 54574 18431 54606
rect 18501 54606 18567 54607
rect 18501 54574 18502 54606
rect 18430 54542 18436 54574
rect 18360 54334 18436 54542
rect 18360 54270 18366 54334
rect 18430 54270 18436 54334
rect 18360 54264 18436 54270
rect 18496 54542 18502 54574
rect 18566 54574 18567 54606
rect 18566 54542 18572 54574
rect 18496 54334 18572 54542
rect 24616 54470 24692 54678
rect 24616 54438 24622 54470
rect 24621 54406 24622 54438
rect 24686 54438 24692 54470
rect 66504 54678 66510 54710
rect 66574 54710 66575 54742
rect 73032 54742 73108 54950
rect 73032 54710 73038 54742
rect 66574 54678 66580 54710
rect 66504 54470 66580 54678
rect 73037 54678 73038 54710
rect 73102 54710 73108 54742
rect 73102 54678 73103 54710
rect 73037 54677 73103 54678
rect 72357 54606 72423 54607
rect 72357 54574 72358 54606
rect 24686 54406 24687 54438
rect 24621 54405 24687 54406
rect 66504 54406 66510 54470
rect 66574 54406 66580 54470
rect 66504 54400 66580 54406
rect 72352 54542 72358 54574
rect 72422 54574 72423 54606
rect 72901 54606 72967 54607
rect 72901 54574 72902 54606
rect 72422 54542 72428 54574
rect 18496 54270 18502 54334
rect 18566 54270 18572 54334
rect 18496 54264 18572 54270
rect 24344 54334 24420 54340
rect 24344 54270 24350 54334
rect 24414 54270 24420 54334
rect 952 54134 1230 54198
rect 1294 54134 1300 54198
rect 17957 54198 18023 54199
rect 17957 54166 17958 54198
rect 952 52566 1300 54134
rect 17952 54134 17958 54166
rect 18022 54166 18023 54198
rect 19181 54198 19247 54199
rect 19181 54166 19182 54198
rect 18022 54134 18028 54166
rect 17952 53926 18028 54134
rect 17952 53862 17958 53926
rect 18022 53862 18028 53926
rect 17952 53856 18028 53862
rect 19176 54134 19182 54166
rect 19246 54166 19247 54198
rect 19448 54198 19524 54204
rect 19246 54134 19252 54166
rect 19176 53926 19252 54134
rect 19176 53862 19182 53926
rect 19246 53862 19252 53926
rect 19448 54134 19454 54198
rect 19518 54134 19524 54198
rect 19448 53926 19524 54134
rect 24344 54062 24420 54270
rect 72352 54334 72428 54542
rect 72352 54270 72358 54334
rect 72422 54270 72428 54334
rect 72352 54264 72428 54270
rect 72896 54542 72902 54574
rect 72966 54574 72967 54606
rect 72966 54542 72972 54574
rect 72896 54334 72972 54542
rect 72896 54270 72902 54334
rect 72966 54270 72972 54334
rect 72896 54264 72972 54270
rect 71405 54198 71471 54199
rect 71405 54166 71406 54198
rect 24344 54030 24350 54062
rect 24349 53998 24350 54030
rect 24414 54030 24420 54062
rect 71400 54134 71406 54166
rect 71470 54166 71471 54198
rect 71813 54198 71879 54199
rect 71813 54166 71814 54198
rect 71470 54134 71476 54166
rect 24414 53998 24415 54030
rect 24349 53997 24415 53998
rect 19448 53894 19454 53926
rect 19176 53856 19252 53862
rect 19453 53862 19454 53894
rect 19518 53894 19524 53926
rect 71400 53926 71476 54134
rect 19518 53862 19519 53894
rect 19453 53861 19519 53862
rect 71400 53862 71406 53926
rect 71470 53862 71476 53926
rect 71400 53856 71476 53862
rect 71808 54134 71814 54166
rect 71878 54166 71879 54198
rect 73032 54198 73108 54204
rect 71878 54134 71884 54166
rect 71808 53926 71884 54134
rect 71808 53862 71814 53926
rect 71878 53862 71884 53926
rect 73032 54134 73038 54198
rect 73102 54134 73108 54198
rect 73032 53926 73108 54134
rect 73032 53894 73038 53926
rect 71808 53856 71884 53862
rect 73037 53862 73038 53894
rect 73102 53894 73108 53926
rect 89760 54198 90108 55766
rect 89760 54134 89766 54198
rect 89830 54134 90108 54198
rect 73102 53862 73103 53894
rect 73037 53861 73103 53862
rect 17816 53790 17892 53796
rect 17816 53726 17822 53790
rect 17886 53726 17892 53790
rect 17816 53518 17892 53726
rect 17816 53486 17822 53518
rect 17821 53454 17822 53486
rect 17886 53486 17892 53518
rect 19176 53790 19252 53796
rect 19176 53726 19182 53790
rect 19246 53726 19252 53790
rect 19176 53518 19252 53726
rect 19176 53486 19182 53518
rect 17886 53454 17887 53486
rect 17821 53453 17887 53454
rect 19181 53454 19182 53486
rect 19246 53486 19252 53518
rect 19448 53790 19524 53796
rect 19448 53726 19454 53790
rect 19518 53726 19524 53790
rect 19448 53518 19524 53726
rect 19448 53486 19454 53518
rect 19246 53454 19247 53486
rect 19181 53453 19247 53454
rect 19453 53454 19454 53486
rect 19518 53486 19524 53518
rect 71400 53790 71476 53796
rect 71400 53726 71406 53790
rect 71470 53726 71476 53790
rect 71400 53518 71476 53726
rect 71400 53486 71406 53518
rect 19518 53454 19519 53486
rect 19453 53453 19519 53454
rect 71405 53454 71406 53486
rect 71470 53486 71476 53518
rect 71672 53790 71748 53796
rect 71672 53726 71678 53790
rect 71742 53726 71748 53790
rect 71672 53518 71748 53726
rect 71672 53486 71678 53518
rect 71470 53454 71471 53486
rect 71405 53453 71471 53454
rect 71677 53454 71678 53486
rect 71742 53486 71748 53518
rect 72080 53790 72156 53796
rect 72080 53726 72086 53790
rect 72150 53726 72156 53790
rect 73037 53790 73103 53791
rect 73037 53758 73038 53790
rect 72080 53518 72156 53726
rect 72080 53486 72086 53518
rect 71742 53454 71743 53486
rect 71677 53453 71743 53454
rect 72085 53454 72086 53486
rect 72150 53486 72156 53518
rect 73032 53726 73038 53758
rect 73102 53758 73103 53790
rect 73102 53726 73108 53758
rect 73032 53518 73108 53726
rect 72150 53454 72151 53486
rect 72085 53453 72151 53454
rect 73032 53454 73038 53518
rect 73102 53454 73108 53518
rect 73032 53448 73108 53454
rect 17821 53382 17887 53383
rect 17821 53350 17822 53382
rect 17816 53318 17822 53350
rect 17886 53350 17887 53382
rect 18501 53382 18567 53383
rect 18501 53350 18502 53382
rect 17886 53318 17892 53350
rect 17816 53110 17892 53318
rect 17816 53046 17822 53110
rect 17886 53046 17892 53110
rect 17816 53040 17892 53046
rect 18496 53318 18502 53350
rect 18566 53350 18567 53382
rect 19176 53382 19252 53388
rect 18566 53318 18572 53350
rect 18496 53110 18572 53318
rect 18496 53046 18502 53110
rect 18566 53046 18572 53110
rect 19176 53318 19182 53382
rect 19246 53318 19252 53382
rect 19453 53382 19519 53383
rect 19453 53350 19454 53382
rect 19176 53110 19252 53318
rect 19176 53078 19182 53110
rect 18496 53040 18572 53046
rect 19181 53046 19182 53078
rect 19246 53078 19252 53110
rect 19448 53318 19454 53350
rect 19518 53350 19519 53382
rect 71405 53382 71471 53383
rect 71405 53350 71406 53382
rect 19518 53318 19524 53350
rect 19448 53110 19524 53318
rect 19246 53046 19247 53078
rect 19181 53045 19247 53046
rect 19448 53046 19454 53110
rect 19518 53046 19524 53110
rect 19448 53040 19524 53046
rect 71400 53318 71406 53350
rect 71470 53350 71471 53382
rect 71677 53382 71743 53383
rect 71677 53350 71678 53382
rect 71470 53318 71476 53350
rect 71400 53110 71476 53318
rect 71400 53046 71406 53110
rect 71470 53046 71476 53110
rect 71400 53040 71476 53046
rect 71672 53318 71678 53350
rect 71742 53350 71743 53382
rect 72080 53382 72156 53388
rect 71742 53318 71748 53350
rect 71672 53110 71748 53318
rect 71672 53046 71678 53110
rect 71742 53046 71748 53110
rect 72080 53318 72086 53382
rect 72150 53318 72156 53382
rect 72080 53110 72156 53318
rect 72080 53078 72086 53110
rect 71672 53040 71748 53046
rect 72085 53046 72086 53078
rect 72150 53078 72156 53110
rect 72352 53382 72428 53388
rect 72352 53318 72358 53382
rect 72422 53318 72428 53382
rect 72901 53382 72967 53383
rect 72901 53350 72902 53382
rect 72352 53110 72428 53318
rect 72352 53078 72358 53110
rect 72150 53046 72151 53078
rect 72085 53045 72151 53046
rect 72357 53046 72358 53078
rect 72422 53078 72428 53110
rect 72896 53318 72902 53350
rect 72966 53350 72967 53382
rect 72966 53318 72972 53350
rect 72896 53110 72972 53318
rect 72422 53046 72423 53078
rect 72357 53045 72423 53046
rect 72896 53046 72902 53110
rect 72966 53046 72972 53110
rect 72896 53040 72972 53046
rect 17821 52974 17887 52975
rect 17821 52942 17822 52974
rect 17816 52910 17822 52942
rect 17886 52942 17887 52974
rect 18229 52974 18295 52975
rect 18229 52942 18230 52974
rect 17886 52910 17892 52942
rect 17816 52702 17892 52910
rect 17816 52638 17822 52702
rect 17886 52638 17892 52702
rect 17816 52632 17892 52638
rect 18224 52910 18230 52942
rect 18294 52942 18295 52974
rect 18909 52974 18975 52975
rect 18909 52942 18910 52974
rect 18294 52910 18300 52942
rect 18224 52702 18300 52910
rect 18224 52638 18230 52702
rect 18294 52638 18300 52702
rect 18224 52632 18300 52638
rect 18904 52910 18910 52942
rect 18974 52942 18975 52974
rect 19045 52974 19111 52975
rect 19045 52942 19046 52974
rect 18974 52910 18980 52942
rect 18904 52702 18980 52910
rect 18904 52638 18910 52702
rect 18974 52638 18980 52702
rect 18904 52632 18980 52638
rect 19040 52910 19046 52942
rect 19110 52942 19111 52974
rect 19453 52974 19519 52975
rect 19453 52942 19454 52974
rect 19110 52910 19116 52942
rect 19040 52702 19116 52910
rect 19040 52638 19046 52702
rect 19110 52638 19116 52702
rect 19040 52632 19116 52638
rect 19448 52910 19454 52942
rect 19518 52942 19519 52974
rect 71264 52974 71340 52980
rect 19518 52910 19524 52942
rect 19448 52702 19524 52910
rect 19448 52638 19454 52702
rect 19518 52638 19524 52702
rect 71264 52910 71270 52974
rect 71334 52910 71340 52974
rect 71677 52974 71743 52975
rect 71677 52942 71678 52974
rect 71264 52702 71340 52910
rect 71264 52670 71270 52702
rect 19448 52632 19524 52638
rect 71269 52638 71270 52670
rect 71334 52670 71340 52702
rect 71672 52910 71678 52942
rect 71742 52942 71743 52974
rect 72221 52974 72287 52975
rect 72221 52942 72222 52974
rect 71742 52910 71748 52942
rect 71672 52702 71748 52910
rect 71334 52638 71335 52670
rect 71269 52637 71335 52638
rect 71672 52638 71678 52702
rect 71742 52638 71748 52702
rect 71672 52632 71748 52638
rect 72216 52910 72222 52942
rect 72286 52942 72287 52974
rect 73032 52974 73108 52980
rect 72286 52910 72292 52942
rect 72216 52702 72292 52910
rect 72216 52638 72222 52702
rect 72286 52638 72292 52702
rect 73032 52910 73038 52974
rect 73102 52910 73108 52974
rect 73032 52702 73108 52910
rect 73032 52670 73038 52702
rect 72216 52632 72292 52638
rect 73037 52638 73038 52670
rect 73102 52670 73108 52702
rect 73102 52638 73103 52670
rect 73037 52637 73103 52638
rect 952 52502 1230 52566
rect 1294 52502 1300 52566
rect 952 50798 1300 52502
rect 17816 52566 17892 52572
rect 17816 52502 17822 52566
rect 17886 52502 17892 52566
rect 17816 52294 17892 52502
rect 17816 52262 17822 52294
rect 17821 52230 17822 52262
rect 17886 52262 17892 52294
rect 18360 52566 18436 52572
rect 18360 52502 18366 52566
rect 18430 52502 18436 52566
rect 18360 52294 18436 52502
rect 18360 52262 18366 52294
rect 17886 52230 17887 52262
rect 17821 52229 17887 52230
rect 18365 52230 18366 52262
rect 18430 52262 18436 52294
rect 18496 52566 18572 52572
rect 18496 52502 18502 52566
rect 18566 52502 18572 52566
rect 19045 52566 19111 52567
rect 19045 52534 19046 52566
rect 18496 52294 18572 52502
rect 18496 52262 18502 52294
rect 18430 52230 18431 52262
rect 18365 52229 18431 52230
rect 18501 52230 18502 52262
rect 18566 52262 18572 52294
rect 19040 52502 19046 52534
rect 19110 52534 19111 52566
rect 19589 52566 19655 52567
rect 19589 52534 19590 52566
rect 19110 52502 19116 52534
rect 19040 52294 19116 52502
rect 18566 52230 18567 52262
rect 18501 52229 18567 52230
rect 19040 52230 19046 52294
rect 19110 52230 19116 52294
rect 19040 52224 19116 52230
rect 19584 52502 19590 52534
rect 19654 52534 19655 52566
rect 71269 52566 71335 52567
rect 71269 52534 71270 52566
rect 19654 52502 19660 52534
rect 19584 52294 19660 52502
rect 19584 52230 19590 52294
rect 19654 52230 19660 52294
rect 19584 52224 19660 52230
rect 71264 52502 71270 52534
rect 71334 52534 71335 52566
rect 71672 52566 71748 52572
rect 71334 52502 71340 52534
rect 71264 52294 71340 52502
rect 71264 52230 71270 52294
rect 71334 52230 71340 52294
rect 71672 52502 71678 52566
rect 71742 52502 71748 52566
rect 71672 52294 71748 52502
rect 71672 52262 71678 52294
rect 71264 52224 71340 52230
rect 71677 52230 71678 52262
rect 71742 52262 71748 52294
rect 72080 52566 72156 52572
rect 72080 52502 72086 52566
rect 72150 52502 72156 52566
rect 72629 52566 72695 52567
rect 72629 52534 72630 52566
rect 72080 52294 72156 52502
rect 72080 52262 72086 52294
rect 71742 52230 71743 52262
rect 71677 52229 71743 52230
rect 72085 52230 72086 52262
rect 72150 52262 72156 52294
rect 72624 52502 72630 52534
rect 72694 52534 72695 52566
rect 72896 52566 72972 52572
rect 72694 52502 72700 52534
rect 72624 52294 72700 52502
rect 72150 52230 72151 52262
rect 72085 52229 72151 52230
rect 72624 52230 72630 52294
rect 72694 52230 72700 52294
rect 72896 52502 72902 52566
rect 72966 52502 72972 52566
rect 72896 52294 72972 52502
rect 72896 52262 72902 52294
rect 72624 52224 72700 52230
rect 72901 52230 72902 52262
rect 72966 52262 72972 52294
rect 89760 52430 90108 54134
rect 89760 52366 89766 52430
rect 89830 52366 90108 52430
rect 72966 52230 72967 52262
rect 72901 52229 72967 52230
rect 18904 52158 18980 52164
rect 18904 52094 18910 52158
rect 18974 52094 18980 52158
rect 19181 52158 19247 52159
rect 19181 52126 19182 52158
rect 18904 51886 18980 52094
rect 18904 51854 18910 51886
rect 18909 51822 18910 51854
rect 18974 51854 18980 51886
rect 19176 52094 19182 52126
rect 19246 52126 19247 52158
rect 19448 52158 19524 52164
rect 19246 52094 19252 52126
rect 19176 51886 19252 52094
rect 18974 51822 18975 51854
rect 18909 51821 18975 51822
rect 19176 51822 19182 51886
rect 19246 51822 19252 51886
rect 19448 52094 19454 52158
rect 19518 52094 19524 52158
rect 19448 51886 19524 52094
rect 19448 51854 19454 51886
rect 19176 51816 19252 51822
rect 19453 51822 19454 51854
rect 19518 51854 19524 51886
rect 71264 52158 71340 52164
rect 71264 52094 71270 52158
rect 71334 52094 71340 52158
rect 71264 51886 71340 52094
rect 71264 51854 71270 51886
rect 19518 51822 19519 51854
rect 19453 51821 19519 51822
rect 71269 51822 71270 51854
rect 71334 51854 71340 51886
rect 71672 52158 71748 52164
rect 71672 52094 71678 52158
rect 71742 52094 71748 52158
rect 71672 51886 71748 52094
rect 71672 51854 71678 51886
rect 71334 51822 71335 51854
rect 71269 51821 71335 51822
rect 71677 51822 71678 51854
rect 71742 51854 71748 51886
rect 72352 52158 72428 52164
rect 72352 52094 72358 52158
rect 72422 52094 72428 52158
rect 72352 51886 72428 52094
rect 72352 51854 72358 51886
rect 71742 51822 71743 51854
rect 71677 51821 71743 51822
rect 72357 51822 72358 51854
rect 72422 51854 72428 51886
rect 72422 51822 72423 51854
rect 72357 51821 72423 51822
rect 19040 51750 19116 51756
rect 19040 51686 19046 51750
rect 19110 51686 19116 51750
rect 19040 51478 19116 51686
rect 19040 51446 19046 51478
rect 19045 51414 19046 51446
rect 19110 51446 19116 51478
rect 19584 51750 19660 51756
rect 19584 51686 19590 51750
rect 19654 51686 19660 51750
rect 71269 51750 71335 51751
rect 71269 51718 71270 51750
rect 19584 51478 19660 51686
rect 19584 51446 19590 51478
rect 19110 51414 19111 51446
rect 19045 51413 19111 51414
rect 19589 51414 19590 51446
rect 19654 51446 19660 51478
rect 71264 51686 71270 51718
rect 71334 51718 71335 51750
rect 71677 51750 71743 51751
rect 71677 51718 71678 51750
rect 71334 51686 71340 51718
rect 71264 51478 71340 51686
rect 19654 51414 19655 51446
rect 19589 51413 19655 51414
rect 71264 51414 71270 51478
rect 71334 51414 71340 51478
rect 71264 51408 71340 51414
rect 71672 51686 71678 51718
rect 71742 51718 71743 51750
rect 72352 51750 72564 51756
rect 71742 51686 71748 51718
rect 71672 51478 71748 51686
rect 71672 51414 71678 51478
rect 71742 51414 71748 51478
rect 72352 51686 72494 51750
rect 72558 51686 72564 51750
rect 72352 51680 72564 51686
rect 72352 51478 72428 51680
rect 72352 51446 72358 51478
rect 71672 51408 71748 51414
rect 72357 51414 72358 51446
rect 72422 51446 72428 51478
rect 72422 51414 72423 51446
rect 72357 51413 72423 51414
rect 18501 51342 18567 51343
rect 18501 51310 18502 51342
rect 18496 51278 18502 51310
rect 18566 51310 18567 51342
rect 19176 51342 19252 51348
rect 18566 51278 18572 51310
rect 952 50734 1230 50798
rect 1294 50734 1300 50798
rect 17816 51070 17892 51076
rect 17816 51006 17822 51070
rect 17886 51006 17892 51070
rect 17816 50798 17892 51006
rect 18496 51070 18572 51278
rect 19176 51278 19182 51342
rect 19246 51278 19252 51342
rect 19453 51342 19519 51343
rect 19453 51310 19454 51342
rect 18496 51006 18502 51070
rect 18566 51006 18572 51070
rect 18496 51000 18572 51006
rect 18904 51206 18980 51212
rect 18904 51142 18910 51206
rect 18974 51142 18980 51206
rect 17816 50766 17822 50798
rect 952 49030 1300 50734
rect 17821 50734 17822 50766
rect 17886 50766 17892 50798
rect 18904 50798 18980 51142
rect 19176 51070 19252 51278
rect 19176 51038 19182 51070
rect 19181 51006 19182 51038
rect 19246 51038 19252 51070
rect 19448 51278 19454 51310
rect 19518 51310 19519 51342
rect 71405 51342 71471 51343
rect 71405 51310 71406 51342
rect 19518 51278 19524 51310
rect 19448 51070 19524 51278
rect 71400 51278 71406 51310
rect 71470 51310 71471 51342
rect 71677 51342 71743 51343
rect 71677 51310 71678 51342
rect 71470 51278 71476 51310
rect 24621 51206 24687 51207
rect 24621 51174 24622 51206
rect 19246 51006 19247 51038
rect 19181 51005 19247 51006
rect 19448 51006 19454 51070
rect 19518 51006 19524 51070
rect 19448 51000 19524 51006
rect 24616 51142 24622 51174
rect 24686 51174 24687 51206
rect 66368 51206 66444 51212
rect 24686 51142 24692 51174
rect 18904 50766 18910 50798
rect 17886 50734 17887 50766
rect 17821 50733 17887 50734
rect 18909 50734 18910 50766
rect 18974 50766 18980 50798
rect 24480 50934 24556 50940
rect 24480 50870 24486 50934
rect 24550 50870 24556 50934
rect 18974 50734 18975 50766
rect 18909 50733 18975 50734
rect 17952 50662 18028 50668
rect 17952 50598 17958 50662
rect 18022 50598 18028 50662
rect 18637 50662 18703 50663
rect 18637 50630 18638 50662
rect 17952 50390 18028 50598
rect 17952 50358 17958 50390
rect 17957 50326 17958 50358
rect 18022 50358 18028 50390
rect 18632 50598 18638 50630
rect 18702 50630 18703 50662
rect 18702 50598 18708 50630
rect 18632 50390 18708 50598
rect 24480 50526 24556 50870
rect 24616 50934 24692 51142
rect 24616 50870 24622 50934
rect 24686 50870 24692 50934
rect 66368 51142 66374 51206
rect 66438 51142 66444 51206
rect 66368 50934 66444 51142
rect 71400 51070 71476 51278
rect 71400 51006 71406 51070
rect 71470 51006 71476 51070
rect 71400 51000 71476 51006
rect 71672 51278 71678 51310
rect 71742 51310 71743 51342
rect 72488 51342 72564 51348
rect 71742 51278 71748 51310
rect 71672 51070 71748 51278
rect 71672 51006 71678 51070
rect 71742 51006 71748 51070
rect 72488 51278 72494 51342
rect 72558 51278 72564 51342
rect 72488 51070 72564 51278
rect 72488 51038 72494 51070
rect 71672 51000 71748 51006
rect 72493 51006 72494 51038
rect 72558 51038 72564 51070
rect 72901 51070 72967 51071
rect 72901 51038 72902 51070
rect 72558 51006 72559 51038
rect 72493 51005 72559 51006
rect 72896 51006 72902 51038
rect 72966 51038 72967 51070
rect 72966 51006 72972 51038
rect 66368 50902 66374 50934
rect 24616 50864 24692 50870
rect 66373 50870 66374 50902
rect 66438 50902 66444 50934
rect 66438 50870 66439 50902
rect 66373 50869 66439 50870
rect 24480 50494 24486 50526
rect 24485 50462 24486 50494
rect 24550 50494 24556 50526
rect 66368 50798 66444 50804
rect 66368 50734 66374 50798
rect 66438 50734 66444 50798
rect 66368 50526 66444 50734
rect 66368 50494 66374 50526
rect 24550 50462 24551 50494
rect 24485 50461 24551 50462
rect 66373 50462 66374 50494
rect 66438 50494 66444 50526
rect 66504 50798 66580 50804
rect 66504 50734 66510 50798
rect 66574 50734 66580 50798
rect 66438 50462 66439 50494
rect 66373 50461 66439 50462
rect 18022 50326 18023 50358
rect 17957 50325 18023 50326
rect 18632 50326 18638 50390
rect 18702 50326 18708 50390
rect 66504 50390 66580 50734
rect 72896 50798 72972 51006
rect 72896 50734 72902 50798
rect 72966 50734 72972 50798
rect 72896 50728 72972 50734
rect 89760 50798 90108 52366
rect 89760 50734 89766 50798
rect 89830 50734 90108 50798
rect 72357 50662 72423 50663
rect 72357 50630 72358 50662
rect 66504 50358 66510 50390
rect 18632 50320 18708 50326
rect 66509 50326 66510 50358
rect 66574 50358 66580 50390
rect 72352 50598 72358 50630
rect 72422 50630 72423 50662
rect 73032 50662 73108 50668
rect 72422 50598 72428 50630
rect 72352 50390 72428 50598
rect 66574 50326 66575 50358
rect 66509 50325 66575 50326
rect 72352 50326 72358 50390
rect 72422 50326 72428 50390
rect 73032 50598 73038 50662
rect 73102 50598 73108 50662
rect 73032 50390 73108 50598
rect 73032 50358 73038 50390
rect 72352 50320 72428 50326
rect 73037 50326 73038 50358
rect 73102 50358 73108 50390
rect 73102 50326 73103 50358
rect 73037 50325 73103 50326
rect 17952 50254 18028 50260
rect 17952 50190 17958 50254
rect 18022 50190 18028 50254
rect 72901 50254 72967 50255
rect 72901 50222 72902 50254
rect 17952 49982 18028 50190
rect 17952 49950 17958 49982
rect 17957 49918 17958 49950
rect 18022 49950 18028 49982
rect 72896 50190 72902 50222
rect 72966 50222 72967 50254
rect 72966 50190 72972 50222
rect 72896 49982 72972 50190
rect 18022 49918 18023 49950
rect 17957 49917 18023 49918
rect 72896 49918 72902 49982
rect 72966 49918 72972 49982
rect 72896 49912 72972 49918
rect 17957 49846 18023 49847
rect 17957 49814 17958 49846
rect 17952 49782 17958 49814
rect 18022 49814 18023 49846
rect 18224 49846 18300 49852
rect 18022 49782 18028 49814
rect 17952 49574 18028 49782
rect 17952 49510 17958 49574
rect 18022 49510 18028 49574
rect 18224 49782 18230 49846
rect 18294 49782 18300 49846
rect 18773 49846 18839 49847
rect 18773 49814 18774 49846
rect 18224 49574 18300 49782
rect 18224 49542 18230 49574
rect 17952 49504 18028 49510
rect 18229 49510 18230 49542
rect 18294 49542 18300 49574
rect 18768 49782 18774 49814
rect 18838 49814 18839 49846
rect 19181 49846 19247 49847
rect 19181 49814 19182 49846
rect 18838 49782 18844 49814
rect 18768 49574 18844 49782
rect 18294 49510 18295 49542
rect 18229 49509 18295 49510
rect 18768 49510 18774 49574
rect 18838 49510 18844 49574
rect 18768 49504 18844 49510
rect 19176 49782 19182 49814
rect 19246 49814 19247 49846
rect 19584 49846 19660 49852
rect 19246 49782 19252 49814
rect 19176 49574 19252 49782
rect 19176 49510 19182 49574
rect 19246 49510 19252 49574
rect 19584 49782 19590 49846
rect 19654 49782 19660 49846
rect 19584 49574 19660 49782
rect 19584 49542 19590 49574
rect 19176 49504 19252 49510
rect 19589 49510 19590 49542
rect 19654 49542 19660 49574
rect 71264 49846 71340 49852
rect 71264 49782 71270 49846
rect 71334 49782 71340 49846
rect 71264 49574 71340 49782
rect 71264 49542 71270 49574
rect 19654 49510 19655 49542
rect 19589 49509 19655 49510
rect 71269 49510 71270 49542
rect 71334 49542 71340 49574
rect 71672 49846 71748 49852
rect 71672 49782 71678 49846
rect 71742 49782 71748 49846
rect 72085 49846 72151 49847
rect 72085 49814 72086 49846
rect 71672 49574 71748 49782
rect 71672 49542 71678 49574
rect 71334 49510 71335 49542
rect 71269 49509 71335 49510
rect 71677 49510 71678 49542
rect 71742 49542 71748 49574
rect 72080 49782 72086 49814
rect 72150 49814 72151 49846
rect 72624 49846 72700 49852
rect 72150 49782 72156 49814
rect 72080 49574 72156 49782
rect 71742 49510 71743 49542
rect 71677 49509 71743 49510
rect 72080 49510 72086 49574
rect 72150 49510 72156 49574
rect 72624 49782 72630 49846
rect 72694 49782 72700 49846
rect 72624 49574 72700 49782
rect 72624 49542 72630 49574
rect 72080 49504 72156 49510
rect 72629 49510 72630 49542
rect 72694 49542 72700 49574
rect 73032 49846 73108 49852
rect 73032 49782 73038 49846
rect 73102 49782 73108 49846
rect 73032 49574 73108 49782
rect 73032 49542 73038 49574
rect 72694 49510 72695 49542
rect 72629 49509 72695 49510
rect 73037 49510 73038 49542
rect 73102 49542 73108 49574
rect 73102 49510 73103 49542
rect 73037 49509 73103 49510
rect 17816 49438 17892 49444
rect 17816 49374 17822 49438
rect 17886 49374 17892 49438
rect 17816 49166 17892 49374
rect 17816 49134 17822 49166
rect 17821 49102 17822 49134
rect 17886 49134 17892 49166
rect 18768 49438 18844 49444
rect 18768 49374 18774 49438
rect 18838 49374 18844 49438
rect 18768 49166 18844 49374
rect 18768 49134 18774 49166
rect 17886 49102 17887 49134
rect 17821 49101 17887 49102
rect 18773 49102 18774 49134
rect 18838 49134 18844 49166
rect 19176 49438 19252 49444
rect 19176 49374 19182 49438
rect 19246 49374 19252 49438
rect 19176 49166 19252 49374
rect 19176 49134 19182 49166
rect 18838 49102 18839 49134
rect 18773 49101 18839 49102
rect 19181 49102 19182 49134
rect 19246 49134 19252 49166
rect 19448 49438 19524 49444
rect 19448 49374 19454 49438
rect 19518 49374 19524 49438
rect 71269 49438 71335 49439
rect 71269 49406 71270 49438
rect 19448 49166 19524 49374
rect 19448 49134 19454 49166
rect 19246 49102 19247 49134
rect 19181 49101 19247 49102
rect 19453 49102 19454 49134
rect 19518 49134 19524 49166
rect 71264 49374 71270 49406
rect 71334 49406 71335 49438
rect 71677 49438 71743 49439
rect 71677 49406 71678 49438
rect 71334 49374 71340 49406
rect 71264 49166 71340 49374
rect 19518 49102 19519 49134
rect 19453 49101 19519 49102
rect 71264 49102 71270 49166
rect 71334 49102 71340 49166
rect 71264 49096 71340 49102
rect 71672 49374 71678 49406
rect 71742 49406 71743 49438
rect 72629 49438 72695 49439
rect 72629 49406 72630 49438
rect 71742 49374 71748 49406
rect 71672 49166 71748 49374
rect 71672 49102 71678 49166
rect 71742 49102 71748 49166
rect 71672 49096 71748 49102
rect 72624 49374 72630 49406
rect 72694 49406 72695 49438
rect 73037 49438 73103 49439
rect 73037 49406 73038 49438
rect 72694 49374 72700 49406
rect 72624 49166 72700 49374
rect 72624 49102 72630 49166
rect 72694 49102 72700 49166
rect 72624 49096 72700 49102
rect 73032 49374 73038 49406
rect 73102 49406 73103 49438
rect 73102 49374 73108 49406
rect 73032 49166 73108 49374
rect 73032 49102 73038 49166
rect 73102 49102 73108 49166
rect 73032 49096 73108 49102
rect 89760 49166 90108 50734
rect 89760 49102 89766 49166
rect 89830 49102 90108 49166
rect 952 48966 1230 49030
rect 1294 48966 1300 49030
rect 952 47398 1300 48966
rect 17952 49030 18028 49036
rect 17952 48966 17958 49030
rect 18022 48966 18028 49030
rect 17952 48758 18028 48966
rect 17952 48726 17958 48758
rect 17957 48694 17958 48726
rect 18022 48726 18028 48758
rect 18632 49030 18708 49036
rect 18632 48966 18638 49030
rect 18702 48966 18708 49030
rect 19181 49030 19247 49031
rect 19181 48998 19182 49030
rect 18632 48758 18708 48966
rect 18632 48726 18638 48758
rect 18022 48694 18023 48726
rect 17957 48693 18023 48694
rect 18637 48694 18638 48726
rect 18702 48726 18708 48758
rect 19176 48966 19182 48998
rect 19246 48998 19247 49030
rect 19453 49030 19519 49031
rect 19453 48998 19454 49030
rect 19246 48966 19252 48998
rect 19176 48758 19252 48966
rect 18702 48694 18703 48726
rect 18637 48693 18703 48694
rect 19176 48694 19182 48758
rect 19246 48694 19252 48758
rect 19176 48688 19252 48694
rect 19448 48966 19454 48998
rect 19518 48998 19519 49030
rect 71400 49030 71476 49036
rect 19518 48966 19524 48998
rect 19448 48758 19524 48966
rect 19448 48694 19454 48758
rect 19518 48694 19524 48758
rect 71400 48966 71406 49030
rect 71470 48966 71476 49030
rect 71400 48758 71476 48966
rect 71400 48726 71406 48758
rect 19448 48688 19524 48694
rect 71405 48694 71406 48726
rect 71470 48726 71476 48758
rect 71808 49030 71884 49036
rect 71808 48966 71814 49030
rect 71878 48966 71884 49030
rect 72085 49030 72151 49031
rect 72085 48998 72086 49030
rect 71808 48758 71884 48966
rect 71808 48726 71814 48758
rect 71470 48694 71471 48726
rect 71405 48693 71471 48694
rect 71813 48694 71814 48726
rect 71878 48726 71884 48758
rect 72080 48966 72086 48998
rect 72150 48998 72151 49030
rect 72488 49030 72564 49036
rect 72150 48966 72156 48998
rect 72080 48758 72156 48966
rect 71878 48694 71879 48726
rect 71813 48693 71879 48694
rect 72080 48694 72086 48758
rect 72150 48694 72156 48758
rect 72488 48966 72494 49030
rect 72558 48966 72564 49030
rect 72901 49030 72967 49031
rect 72901 48998 72902 49030
rect 72488 48758 72564 48966
rect 72488 48726 72494 48758
rect 72080 48688 72156 48694
rect 72493 48694 72494 48726
rect 72558 48726 72564 48758
rect 72896 48966 72902 48998
rect 72966 48998 72967 49030
rect 72966 48966 72972 48998
rect 72896 48758 72972 48966
rect 72558 48694 72559 48726
rect 72493 48693 72559 48694
rect 72896 48694 72902 48758
rect 72966 48694 72972 48758
rect 72896 48688 72972 48694
rect 17821 48622 17887 48623
rect 17821 48590 17822 48622
rect 17816 48558 17822 48590
rect 17886 48590 17887 48622
rect 18229 48622 18295 48623
rect 18229 48590 18230 48622
rect 17886 48558 17892 48590
rect 17816 48350 17892 48558
rect 17816 48286 17822 48350
rect 17886 48286 17892 48350
rect 17816 48280 17892 48286
rect 18224 48558 18230 48590
rect 18294 48590 18295 48622
rect 18909 48622 18975 48623
rect 18909 48590 18910 48622
rect 18294 48558 18300 48590
rect 18224 48350 18300 48558
rect 18224 48286 18230 48350
rect 18294 48286 18300 48350
rect 18224 48280 18300 48286
rect 18904 48558 18910 48590
rect 18974 48590 18975 48622
rect 19040 48622 19116 48628
rect 18974 48558 18980 48590
rect 18904 48350 18980 48558
rect 18904 48286 18910 48350
rect 18974 48286 18980 48350
rect 19040 48558 19046 48622
rect 19110 48558 19116 48622
rect 19040 48350 19116 48558
rect 19040 48318 19046 48350
rect 18904 48280 18980 48286
rect 19045 48286 19046 48318
rect 19110 48318 19116 48350
rect 19584 48622 19660 48628
rect 19584 48558 19590 48622
rect 19654 48558 19660 48622
rect 71269 48622 71335 48623
rect 71269 48590 71270 48622
rect 19584 48350 19660 48558
rect 19584 48318 19590 48350
rect 19110 48286 19111 48318
rect 19045 48285 19111 48286
rect 19589 48286 19590 48318
rect 19654 48318 19660 48350
rect 71264 48558 71270 48590
rect 71334 48590 71335 48622
rect 71677 48622 71743 48623
rect 71677 48590 71678 48622
rect 71334 48558 71340 48590
rect 71264 48350 71340 48558
rect 19654 48286 19655 48318
rect 19589 48285 19655 48286
rect 71264 48286 71270 48350
rect 71334 48286 71340 48350
rect 71264 48280 71340 48286
rect 71672 48558 71678 48590
rect 71742 48590 71743 48622
rect 72221 48622 72287 48623
rect 72221 48590 72222 48622
rect 71742 48558 71748 48590
rect 71672 48350 71748 48558
rect 71672 48286 71678 48350
rect 71742 48286 71748 48350
rect 71672 48280 71748 48286
rect 72216 48558 72222 48590
rect 72286 48590 72287 48622
rect 73037 48622 73103 48623
rect 73037 48590 73038 48622
rect 72286 48558 72292 48590
rect 72216 48350 72292 48558
rect 72216 48286 72222 48350
rect 72286 48286 72292 48350
rect 72216 48280 72292 48286
rect 73032 48558 73038 48590
rect 73102 48590 73103 48622
rect 73102 48558 73108 48590
rect 73032 48350 73108 48558
rect 73032 48286 73038 48350
rect 73102 48286 73108 48350
rect 73032 48280 73108 48286
rect 18229 48214 18295 48215
rect 18229 48182 18230 48214
rect 18224 48150 18230 48182
rect 18294 48182 18295 48214
rect 19045 48214 19111 48215
rect 19045 48182 19046 48214
rect 18294 48150 18300 48182
rect 18224 47942 18300 48150
rect 18224 47878 18230 47942
rect 18294 47878 18300 47942
rect 18224 47872 18300 47878
rect 19040 48150 19046 48182
rect 19110 48182 19111 48214
rect 19448 48214 19524 48220
rect 19110 48150 19116 48182
rect 19040 47942 19116 48150
rect 19040 47878 19046 47942
rect 19110 47878 19116 47942
rect 19448 48150 19454 48214
rect 19518 48150 19524 48214
rect 71269 48214 71335 48215
rect 71269 48182 71270 48214
rect 19448 47942 19524 48150
rect 19448 47910 19454 47942
rect 19040 47872 19116 47878
rect 19453 47878 19454 47910
rect 19518 47910 19524 47942
rect 71264 48150 71270 48182
rect 71334 48182 71335 48214
rect 71813 48214 71879 48215
rect 71813 48182 71814 48214
rect 71334 48150 71340 48182
rect 71264 47942 71340 48150
rect 19518 47878 19519 47910
rect 19453 47877 19519 47878
rect 71264 47878 71270 47942
rect 71334 47878 71340 47942
rect 71264 47872 71340 47878
rect 71808 48150 71814 48182
rect 71878 48182 71879 48214
rect 72080 48214 72156 48220
rect 71878 48150 71884 48182
rect 71808 47942 71884 48150
rect 71808 47878 71814 47942
rect 71878 47878 71884 47942
rect 72080 48150 72086 48214
rect 72150 48150 72156 48214
rect 72080 47942 72156 48150
rect 72080 47910 72086 47942
rect 71808 47872 71884 47878
rect 72085 47878 72086 47910
rect 72150 47910 72156 47942
rect 72150 47878 72151 47910
rect 72085 47877 72151 47878
rect 19181 47806 19247 47807
rect 19181 47774 19182 47806
rect 19176 47742 19182 47774
rect 19246 47774 19247 47806
rect 19453 47806 19519 47807
rect 19453 47774 19454 47806
rect 19246 47742 19252 47774
rect 19176 47534 19252 47742
rect 19176 47470 19182 47534
rect 19246 47470 19252 47534
rect 19176 47464 19252 47470
rect 19448 47742 19454 47774
rect 19518 47774 19519 47806
rect 71264 47806 71340 47812
rect 19518 47742 19524 47774
rect 19448 47534 19524 47742
rect 19448 47470 19454 47534
rect 19518 47470 19524 47534
rect 71264 47742 71270 47806
rect 71334 47742 71340 47806
rect 71813 47806 71879 47807
rect 71813 47774 71814 47806
rect 71264 47534 71340 47742
rect 71264 47502 71270 47534
rect 19448 47464 19524 47470
rect 71269 47470 71270 47502
rect 71334 47502 71340 47534
rect 71808 47742 71814 47774
rect 71878 47774 71879 47806
rect 71878 47742 71884 47774
rect 71808 47534 71884 47742
rect 71334 47470 71335 47502
rect 71269 47469 71335 47470
rect 71808 47470 71814 47534
rect 71878 47470 71884 47534
rect 71808 47464 71884 47470
rect 952 47334 1230 47398
rect 1294 47334 1300 47398
rect 18909 47398 18975 47399
rect 18909 47366 18910 47398
rect 952 45766 1300 47334
rect 18904 47334 18910 47366
rect 18974 47366 18975 47398
rect 19045 47398 19111 47399
rect 19045 47366 19046 47398
rect 18974 47334 18980 47366
rect 17957 47126 18023 47127
rect 17957 47094 17958 47126
rect 17952 47062 17958 47094
rect 18022 47094 18023 47126
rect 18904 47126 18980 47334
rect 18022 47062 18028 47094
rect 17952 46854 18028 47062
rect 18904 47062 18910 47126
rect 18974 47062 18980 47126
rect 18904 47056 18980 47062
rect 19040 47334 19046 47366
rect 19110 47366 19111 47398
rect 19584 47398 19660 47404
rect 19110 47334 19116 47366
rect 19040 47126 19116 47334
rect 19040 47062 19046 47126
rect 19110 47062 19116 47126
rect 19584 47334 19590 47398
rect 19654 47334 19660 47398
rect 19584 47126 19660 47334
rect 19584 47094 19590 47126
rect 19040 47056 19116 47062
rect 19589 47062 19590 47094
rect 19654 47094 19660 47126
rect 71264 47398 71340 47404
rect 71264 47334 71270 47398
rect 71334 47334 71340 47398
rect 71264 47126 71340 47334
rect 71264 47094 71270 47126
rect 19654 47062 19655 47094
rect 19589 47061 19655 47062
rect 71269 47062 71270 47094
rect 71334 47094 71340 47126
rect 71808 47398 71884 47404
rect 71808 47334 71814 47398
rect 71878 47334 71884 47398
rect 72221 47398 72287 47399
rect 72221 47366 72222 47398
rect 71808 47126 71884 47334
rect 71808 47094 71814 47126
rect 71334 47062 71335 47094
rect 71269 47061 71335 47062
rect 71813 47062 71814 47094
rect 71878 47094 71884 47126
rect 72216 47334 72222 47366
rect 72286 47366 72287 47398
rect 89760 47398 90108 49102
rect 72286 47334 72292 47366
rect 72216 47126 72292 47334
rect 89760 47334 89766 47398
rect 89830 47334 90108 47398
rect 71878 47062 71879 47094
rect 71813 47061 71879 47062
rect 72216 47062 72222 47126
rect 72286 47062 72292 47126
rect 72216 47056 72292 47062
rect 72896 47126 72972 47132
rect 72896 47062 72902 47126
rect 72966 47062 72972 47126
rect 17952 46790 17958 46854
rect 18022 46790 18028 46854
rect 17952 46784 18028 46790
rect 18496 46990 18572 46996
rect 18496 46926 18502 46990
rect 18566 46926 18572 46990
rect 17816 46718 17892 46724
rect 17816 46654 17822 46718
rect 17886 46654 17892 46718
rect 18496 46718 18572 46926
rect 24480 46854 24556 46860
rect 24480 46790 24486 46854
rect 24550 46790 24556 46854
rect 66373 46854 66439 46855
rect 66373 46822 66374 46854
rect 18496 46686 18502 46718
rect 17816 46446 17892 46654
rect 18501 46654 18502 46686
rect 18566 46686 18572 46718
rect 18773 46718 18839 46719
rect 18773 46686 18774 46718
rect 18566 46654 18567 46686
rect 18501 46653 18567 46654
rect 18768 46654 18774 46686
rect 18838 46686 18839 46718
rect 18838 46654 18844 46686
rect 17816 46414 17822 46446
rect 17821 46382 17822 46414
rect 17886 46414 17892 46446
rect 18768 46446 18844 46654
rect 24480 46582 24556 46790
rect 24480 46550 24486 46582
rect 24485 46518 24486 46550
rect 24550 46550 24556 46582
rect 66368 46790 66374 46822
rect 66438 46822 66439 46854
rect 72896 46854 72972 47062
rect 72896 46822 72902 46854
rect 66438 46790 66444 46822
rect 66368 46582 66444 46790
rect 72901 46790 72902 46822
rect 72966 46822 72972 46854
rect 72966 46790 72967 46822
rect 72901 46789 72967 46790
rect 24550 46518 24551 46550
rect 24485 46517 24551 46518
rect 66368 46518 66374 46582
rect 66438 46518 66444 46582
rect 66368 46512 66444 46518
rect 72488 46718 72564 46724
rect 72488 46654 72494 46718
rect 72558 46654 72564 46718
rect 72901 46718 72967 46719
rect 72901 46686 72902 46718
rect 17886 46382 17887 46414
rect 17821 46381 17887 46382
rect 18768 46382 18774 46446
rect 18838 46382 18844 46446
rect 18768 46376 18844 46382
rect 66504 46446 66580 46452
rect 66504 46382 66510 46446
rect 66574 46382 66580 46446
rect 72488 46446 72564 46654
rect 72488 46414 72494 46446
rect 17952 46310 18028 46316
rect 17952 46246 17958 46310
rect 18022 46246 18028 46310
rect 17952 46038 18028 46246
rect 17952 46006 17958 46038
rect 17957 45974 17958 46006
rect 18022 46006 18028 46038
rect 22848 46174 22924 46180
rect 22848 46110 22854 46174
rect 22918 46110 22924 46174
rect 24485 46174 24551 46175
rect 24485 46142 24486 46174
rect 18022 45974 18023 46006
rect 17957 45973 18023 45974
rect 952 45702 1230 45766
rect 1294 45702 1300 45766
rect 952 44270 1300 45702
rect 17952 45902 18028 45908
rect 17952 45838 17958 45902
rect 18022 45838 18028 45902
rect 18365 45902 18431 45903
rect 18365 45870 18366 45902
rect 17952 45630 18028 45838
rect 17952 45598 17958 45630
rect 17957 45566 17958 45598
rect 18022 45598 18028 45630
rect 18360 45838 18366 45870
rect 18430 45870 18431 45902
rect 18496 45902 18572 45908
rect 18430 45838 18436 45870
rect 18360 45630 18436 45838
rect 18022 45566 18023 45598
rect 17957 45565 18023 45566
rect 18360 45566 18366 45630
rect 18430 45566 18436 45630
rect 18496 45838 18502 45902
rect 18566 45838 18572 45902
rect 18496 45630 18572 45838
rect 18496 45598 18502 45630
rect 18360 45560 18436 45566
rect 18501 45566 18502 45598
rect 18566 45598 18572 45630
rect 19176 45902 19252 45908
rect 19176 45838 19182 45902
rect 19246 45838 19252 45902
rect 19453 45902 19519 45903
rect 19453 45870 19454 45902
rect 19176 45630 19252 45838
rect 19176 45598 19182 45630
rect 18566 45566 18567 45598
rect 18501 45565 18567 45566
rect 19181 45566 19182 45598
rect 19246 45598 19252 45630
rect 19448 45838 19454 45870
rect 19518 45870 19519 45902
rect 19518 45838 19524 45870
rect 19448 45630 19524 45838
rect 19246 45566 19247 45598
rect 19181 45565 19247 45566
rect 19448 45566 19454 45630
rect 19518 45566 19524 45630
rect 22848 45630 22924 46110
rect 24480 46110 24486 46142
rect 24550 46142 24551 46174
rect 66504 46174 66580 46382
rect 72493 46382 72494 46414
rect 72558 46414 72564 46446
rect 72896 46654 72902 46686
rect 72966 46686 72967 46718
rect 72966 46654 72972 46686
rect 72896 46446 72972 46654
rect 72558 46382 72559 46414
rect 72493 46381 72559 46382
rect 72896 46382 72902 46446
rect 72966 46382 72972 46446
rect 72896 46376 72972 46382
rect 66504 46142 66510 46174
rect 24550 46110 24556 46142
rect 24480 45902 24556 46110
rect 66509 46110 66510 46142
rect 66574 46142 66580 46174
rect 73032 46310 73108 46316
rect 73032 46246 73038 46310
rect 73102 46246 73108 46310
rect 66574 46110 66575 46142
rect 66509 46109 66575 46110
rect 69365 46038 69431 46039
rect 69365 46006 69366 46038
rect 24480 45838 24486 45902
rect 24550 45838 24556 45902
rect 24480 45832 24556 45838
rect 69360 45974 69366 46006
rect 69430 46006 69431 46038
rect 73032 46038 73108 46246
rect 73032 46006 73038 46038
rect 69430 45974 69436 46006
rect 22848 45598 22854 45630
rect 19448 45560 19524 45566
rect 22853 45566 22854 45598
rect 22918 45598 22924 45630
rect 24344 45630 24420 45636
rect 22918 45566 22919 45598
rect 22853 45565 22919 45566
rect 24344 45566 24350 45630
rect 24414 45566 24420 45630
rect 17957 45494 18023 45495
rect 17957 45462 17958 45494
rect 17952 45430 17958 45462
rect 18022 45462 18023 45494
rect 19040 45494 19116 45500
rect 18022 45430 18028 45462
rect 17952 45222 18028 45430
rect 17952 45158 17958 45222
rect 18022 45158 18028 45222
rect 19040 45430 19046 45494
rect 19110 45430 19116 45494
rect 19040 45222 19116 45430
rect 19040 45190 19046 45222
rect 17952 45152 18028 45158
rect 19045 45158 19046 45190
rect 19110 45190 19116 45222
rect 19448 45494 19524 45500
rect 19448 45430 19454 45494
rect 19518 45430 19524 45494
rect 19448 45222 19524 45430
rect 24344 45358 24420 45566
rect 69360 45630 69436 45974
rect 73037 45974 73038 46006
rect 73102 46006 73108 46038
rect 73102 45974 73103 46006
rect 73037 45973 73103 45974
rect 69360 45566 69366 45630
rect 69430 45566 69436 45630
rect 71400 45902 71476 45908
rect 71400 45838 71406 45902
rect 71470 45838 71476 45902
rect 71677 45902 71743 45903
rect 71677 45870 71678 45902
rect 71400 45630 71476 45838
rect 71400 45598 71406 45630
rect 69360 45560 69436 45566
rect 71405 45566 71406 45598
rect 71470 45598 71476 45630
rect 71672 45838 71678 45870
rect 71742 45870 71743 45902
rect 72085 45902 72151 45903
rect 72085 45870 72086 45902
rect 71742 45838 71748 45870
rect 71672 45630 71748 45838
rect 71470 45566 71471 45598
rect 71405 45565 71471 45566
rect 71672 45566 71678 45630
rect 71742 45566 71748 45630
rect 71672 45560 71748 45566
rect 72080 45838 72086 45870
rect 72150 45870 72151 45902
rect 72493 45902 72559 45903
rect 72493 45870 72494 45902
rect 72150 45838 72156 45870
rect 72080 45630 72156 45838
rect 72080 45566 72086 45630
rect 72150 45566 72156 45630
rect 72080 45560 72156 45566
rect 72488 45838 72494 45870
rect 72558 45870 72559 45902
rect 72896 45902 72972 45908
rect 72558 45838 72564 45870
rect 72488 45630 72564 45838
rect 72488 45566 72494 45630
rect 72558 45566 72564 45630
rect 72896 45838 72902 45902
rect 72966 45838 72972 45902
rect 72896 45630 72972 45838
rect 72896 45598 72902 45630
rect 72488 45560 72564 45566
rect 72901 45566 72902 45598
rect 72966 45598 72972 45630
rect 89760 45766 90108 47334
rect 89760 45702 89766 45766
rect 89830 45702 90108 45766
rect 72966 45566 72967 45598
rect 72901 45565 72967 45566
rect 70725 45494 70791 45495
rect 70725 45462 70726 45494
rect 24344 45326 24350 45358
rect 24349 45294 24350 45326
rect 24414 45326 24420 45358
rect 70720 45430 70726 45462
rect 70790 45462 70791 45494
rect 71264 45494 71340 45500
rect 70790 45430 70796 45462
rect 24414 45294 24415 45326
rect 24349 45293 24415 45294
rect 19448 45190 19454 45222
rect 19110 45158 19111 45190
rect 19045 45157 19111 45158
rect 19453 45158 19454 45190
rect 19518 45190 19524 45222
rect 70720 45222 70796 45430
rect 19518 45158 19519 45190
rect 19453 45157 19519 45158
rect 70720 45158 70726 45222
rect 70790 45158 70796 45222
rect 71264 45430 71270 45494
rect 71334 45430 71340 45494
rect 71264 45222 71340 45430
rect 71264 45190 71270 45222
rect 70720 45152 70796 45158
rect 71269 45158 71270 45190
rect 71334 45190 71340 45222
rect 71672 45494 71748 45500
rect 71672 45430 71678 45494
rect 71742 45430 71748 45494
rect 71672 45222 71748 45430
rect 71672 45190 71678 45222
rect 71334 45158 71335 45190
rect 71269 45157 71335 45158
rect 71677 45158 71678 45190
rect 71742 45190 71748 45222
rect 72216 45494 72292 45500
rect 72216 45430 72222 45494
rect 72286 45430 72292 45494
rect 72216 45222 72292 45430
rect 72216 45190 72222 45222
rect 71742 45158 71743 45190
rect 71677 45157 71743 45158
rect 72221 45158 72222 45190
rect 72286 45190 72292 45222
rect 72352 45494 72428 45500
rect 72352 45430 72358 45494
rect 72422 45430 72428 45494
rect 72352 45222 72428 45430
rect 72352 45190 72358 45222
rect 72286 45158 72287 45190
rect 72221 45157 72287 45158
rect 72357 45158 72358 45190
rect 72422 45190 72428 45222
rect 73032 45494 73108 45500
rect 73032 45430 73038 45494
rect 73102 45430 73108 45494
rect 73032 45222 73108 45430
rect 73032 45190 73038 45222
rect 72422 45158 72423 45190
rect 72357 45157 72423 45158
rect 73037 45158 73038 45190
rect 73102 45190 73108 45222
rect 73102 45158 73103 45190
rect 73037 45157 73103 45158
rect 17821 45086 17887 45087
rect 17821 45054 17822 45086
rect 17816 45022 17822 45054
rect 17886 45054 17887 45086
rect 18360 45086 18436 45092
rect 17886 45022 17892 45054
rect 17816 44814 17892 45022
rect 17816 44750 17822 44814
rect 17886 44750 17892 44814
rect 18360 45022 18366 45086
rect 18430 45022 18436 45086
rect 19045 45086 19111 45087
rect 19045 45054 19046 45086
rect 18360 44814 18436 45022
rect 18360 44782 18366 44814
rect 17816 44744 17892 44750
rect 18365 44750 18366 44782
rect 18430 44782 18436 44814
rect 19040 45022 19046 45054
rect 19110 45054 19111 45086
rect 19448 45086 19524 45092
rect 19110 45022 19116 45054
rect 19040 44814 19116 45022
rect 18430 44750 18431 44782
rect 18365 44749 18431 44750
rect 19040 44750 19046 44814
rect 19110 44750 19116 44814
rect 19448 45022 19454 45086
rect 19518 45022 19524 45086
rect 71269 45086 71335 45087
rect 71269 45054 71270 45086
rect 19448 44814 19524 45022
rect 19448 44782 19454 44814
rect 19040 44744 19116 44750
rect 19453 44750 19454 44782
rect 19518 44782 19524 44814
rect 71264 45022 71270 45054
rect 71334 45054 71335 45086
rect 71672 45086 71748 45092
rect 71334 45022 71340 45054
rect 71264 44814 71340 45022
rect 19518 44750 19519 44782
rect 19453 44749 19519 44750
rect 71264 44750 71270 44814
rect 71334 44750 71340 44814
rect 71672 45022 71678 45086
rect 71742 45022 71748 45086
rect 71672 44814 71748 45022
rect 71672 44782 71678 44814
rect 71264 44744 71340 44750
rect 71677 44750 71678 44782
rect 71742 44782 71748 44814
rect 72488 45086 72564 45092
rect 72488 45022 72494 45086
rect 72558 45022 72564 45086
rect 73037 45086 73103 45087
rect 73037 45054 73038 45086
rect 72488 44814 72564 45022
rect 72488 44782 72494 44814
rect 71742 44750 71743 44782
rect 71677 44749 71743 44750
rect 72493 44750 72494 44782
rect 72558 44782 72564 44814
rect 73032 45022 73038 45054
rect 73102 45054 73103 45086
rect 73102 45022 73108 45054
rect 73032 44814 73108 45022
rect 72558 44750 72559 44782
rect 72493 44749 72559 44750
rect 73032 44750 73038 44814
rect 73102 44750 73108 44814
rect 73032 44744 73108 44750
rect 17821 44678 17887 44679
rect 17821 44646 17822 44678
rect 17816 44614 17822 44646
rect 17886 44646 17887 44678
rect 18632 44678 18708 44684
rect 17886 44614 17892 44646
rect 17816 44406 17892 44614
rect 17816 44342 17822 44406
rect 17886 44342 17892 44406
rect 18632 44614 18638 44678
rect 18702 44614 18708 44678
rect 18632 44406 18708 44614
rect 18632 44374 18638 44406
rect 17816 44336 17892 44342
rect 18637 44342 18638 44374
rect 18702 44374 18708 44406
rect 19176 44678 19252 44684
rect 19176 44614 19182 44678
rect 19246 44614 19252 44678
rect 19176 44406 19252 44614
rect 19176 44374 19182 44406
rect 18702 44342 18703 44374
rect 18637 44341 18703 44342
rect 19181 44342 19182 44374
rect 19246 44374 19252 44406
rect 19584 44678 19660 44684
rect 19584 44614 19590 44678
rect 19654 44614 19660 44678
rect 19584 44406 19660 44614
rect 19584 44374 19590 44406
rect 19246 44342 19247 44374
rect 19181 44341 19247 44342
rect 19589 44342 19590 44374
rect 19654 44374 19660 44406
rect 71400 44678 71476 44684
rect 71400 44614 71406 44678
rect 71470 44614 71476 44678
rect 71400 44406 71476 44614
rect 71400 44374 71406 44406
rect 19654 44342 19655 44374
rect 19589 44341 19655 44342
rect 71405 44342 71406 44374
rect 71470 44374 71476 44406
rect 71808 44678 71884 44684
rect 71808 44614 71814 44678
rect 71878 44614 71884 44678
rect 72085 44678 72151 44679
rect 72085 44646 72086 44678
rect 71808 44406 71884 44614
rect 71808 44374 71814 44406
rect 71470 44342 71471 44374
rect 71405 44341 71471 44342
rect 71813 44342 71814 44374
rect 71878 44374 71884 44406
rect 72080 44614 72086 44646
rect 72150 44646 72151 44678
rect 72352 44678 72428 44684
rect 72150 44614 72156 44646
rect 72080 44406 72156 44614
rect 71878 44342 71879 44374
rect 71813 44341 71879 44342
rect 72080 44342 72086 44406
rect 72150 44342 72156 44406
rect 72352 44614 72358 44678
rect 72422 44614 72428 44678
rect 72901 44678 72967 44679
rect 72901 44646 72902 44678
rect 72352 44406 72428 44614
rect 72352 44374 72358 44406
rect 72080 44336 72156 44342
rect 72357 44342 72358 44374
rect 72422 44374 72428 44406
rect 72896 44614 72902 44646
rect 72966 44646 72967 44678
rect 72966 44614 72972 44646
rect 72896 44406 72972 44614
rect 72422 44342 72423 44374
rect 72357 44341 72423 44342
rect 72896 44342 72902 44406
rect 72966 44342 72972 44406
rect 72896 44336 72972 44342
rect 952 44206 1230 44270
rect 1294 44206 1300 44270
rect 952 42366 1300 44206
rect 18224 44270 18300 44276
rect 18224 44206 18230 44270
rect 18294 44206 18300 44270
rect 18909 44270 18975 44271
rect 18909 44238 18910 44270
rect 18224 43998 18300 44206
rect 18224 43966 18230 43998
rect 18229 43934 18230 43966
rect 18294 43966 18300 43998
rect 18904 44206 18910 44238
rect 18974 44238 18975 44270
rect 19040 44270 19116 44276
rect 18974 44206 18980 44238
rect 18904 43998 18980 44206
rect 18294 43934 18295 43966
rect 18229 43933 18295 43934
rect 18904 43934 18910 43998
rect 18974 43934 18980 43998
rect 19040 44206 19046 44270
rect 19110 44206 19116 44270
rect 19040 43998 19116 44206
rect 19040 43966 19046 43998
rect 18904 43928 18980 43934
rect 19045 43934 19046 43966
rect 19110 43966 19116 43998
rect 19584 44270 19660 44276
rect 19584 44206 19590 44270
rect 19654 44206 19660 44270
rect 71269 44270 71335 44271
rect 71269 44238 71270 44270
rect 19584 43998 19660 44206
rect 19584 43966 19590 43998
rect 19110 43934 19111 43966
rect 19045 43933 19111 43934
rect 19589 43934 19590 43966
rect 19654 43966 19660 43998
rect 71264 44206 71270 44238
rect 71334 44238 71335 44270
rect 71677 44270 71743 44271
rect 71677 44238 71678 44270
rect 71334 44206 71340 44238
rect 71264 43998 71340 44206
rect 19654 43934 19655 43966
rect 19589 43933 19655 43934
rect 71264 43934 71270 43998
rect 71334 43934 71340 43998
rect 71264 43928 71340 43934
rect 71672 44206 71678 44238
rect 71742 44238 71743 44270
rect 72216 44270 72292 44276
rect 71742 44206 71748 44238
rect 71672 43998 71748 44206
rect 71672 43934 71678 43998
rect 71742 43934 71748 43998
rect 72216 44206 72222 44270
rect 72286 44206 72292 44270
rect 72216 43998 72292 44206
rect 72216 43966 72222 43998
rect 71672 43928 71748 43934
rect 72221 43934 72222 43966
rect 72286 43966 72292 43998
rect 89760 43998 90108 45702
rect 72286 43934 72287 43966
rect 72221 43933 72287 43934
rect 89760 43934 89766 43998
rect 89830 43934 90108 43998
rect 17957 43862 18023 43863
rect 17957 43830 17958 43862
rect 17952 43798 17958 43830
rect 18022 43830 18023 43862
rect 18360 43862 18436 43868
rect 18022 43798 18028 43830
rect 17952 43590 18028 43798
rect 17952 43526 17958 43590
rect 18022 43526 18028 43590
rect 18360 43798 18366 43862
rect 18430 43798 18436 43862
rect 19045 43862 19111 43863
rect 19045 43830 19046 43862
rect 18360 43590 18436 43798
rect 18360 43558 18366 43590
rect 17952 43520 18028 43526
rect 18365 43526 18366 43558
rect 18430 43558 18436 43590
rect 19040 43798 19046 43830
rect 19110 43830 19111 43862
rect 19589 43862 19655 43863
rect 19589 43830 19590 43862
rect 19110 43798 19116 43830
rect 19040 43590 19116 43798
rect 18430 43526 18431 43558
rect 18365 43525 18431 43526
rect 19040 43526 19046 43590
rect 19110 43526 19116 43590
rect 19040 43520 19116 43526
rect 19584 43798 19590 43830
rect 19654 43830 19655 43862
rect 71269 43862 71335 43863
rect 71269 43830 71270 43862
rect 19654 43798 19660 43830
rect 19584 43590 19660 43798
rect 19584 43526 19590 43590
rect 19654 43526 19660 43590
rect 19584 43520 19660 43526
rect 71264 43798 71270 43830
rect 71334 43830 71335 43862
rect 71672 43862 71748 43868
rect 71334 43798 71340 43830
rect 71264 43590 71340 43798
rect 71264 43526 71270 43590
rect 71334 43526 71340 43590
rect 71672 43798 71678 43862
rect 71742 43798 71748 43862
rect 72629 43862 72695 43863
rect 72629 43830 72630 43862
rect 71672 43590 71748 43798
rect 71672 43558 71678 43590
rect 71264 43520 71340 43526
rect 71677 43526 71678 43558
rect 71742 43558 71748 43590
rect 72624 43798 72630 43830
rect 72694 43830 72695 43862
rect 73037 43862 73103 43863
rect 73037 43830 73038 43862
rect 72694 43798 72700 43830
rect 72624 43590 72700 43798
rect 71742 43526 71743 43558
rect 71677 43525 71743 43526
rect 72624 43526 72630 43590
rect 72694 43526 72700 43590
rect 72624 43520 72700 43526
rect 73032 43798 73038 43830
rect 73102 43830 73103 43862
rect 73102 43798 73108 43830
rect 73032 43590 73108 43798
rect 73032 43526 73038 43590
rect 73102 43526 73108 43590
rect 73032 43520 73108 43526
rect 18904 43454 18980 43460
rect 18904 43390 18910 43454
rect 18974 43390 18980 43454
rect 17816 43182 17892 43188
rect 17816 43118 17822 43182
rect 17886 43118 17892 43182
rect 18904 43182 18980 43390
rect 18904 43150 18910 43182
rect 17816 42910 17892 43118
rect 18909 43118 18910 43150
rect 18974 43150 18980 43182
rect 19040 43454 19116 43460
rect 19040 43390 19046 43454
rect 19110 43390 19116 43454
rect 19040 43182 19116 43390
rect 19040 43150 19046 43182
rect 18974 43118 18975 43150
rect 18909 43117 18975 43118
rect 19045 43118 19046 43150
rect 19110 43150 19116 43182
rect 19448 43454 19524 43460
rect 19448 43390 19454 43454
rect 19518 43390 19524 43454
rect 71405 43454 71471 43455
rect 71405 43422 71406 43454
rect 19448 43182 19524 43390
rect 19448 43150 19454 43182
rect 19110 43118 19111 43150
rect 19045 43117 19111 43118
rect 19453 43118 19454 43150
rect 19518 43150 19524 43182
rect 71400 43390 71406 43422
rect 71470 43422 71471 43454
rect 71813 43454 71879 43455
rect 71813 43422 71814 43454
rect 71470 43390 71476 43422
rect 71400 43182 71476 43390
rect 19518 43118 19519 43150
rect 19453 43117 19519 43118
rect 71400 43118 71406 43182
rect 71470 43118 71476 43182
rect 71400 43112 71476 43118
rect 71808 43390 71814 43422
rect 71878 43422 71879 43454
rect 72216 43454 72292 43460
rect 71878 43390 71884 43422
rect 71808 43182 71884 43390
rect 71808 43118 71814 43182
rect 71878 43118 71884 43182
rect 72216 43390 72222 43454
rect 72286 43390 72292 43454
rect 72216 43182 72292 43390
rect 72216 43150 72222 43182
rect 71808 43112 71884 43118
rect 72221 43118 72222 43150
rect 72286 43150 72292 43182
rect 72352 43454 72428 43460
rect 72352 43390 72358 43454
rect 72422 43390 72428 43454
rect 72352 43182 72428 43390
rect 72352 43150 72358 43182
rect 72286 43118 72287 43150
rect 72221 43117 72287 43118
rect 72357 43118 72358 43150
rect 72422 43150 72428 43182
rect 73037 43182 73103 43183
rect 73037 43150 73038 43182
rect 72422 43118 72423 43150
rect 72357 43117 72423 43118
rect 73032 43118 73038 43150
rect 73102 43150 73103 43182
rect 73102 43118 73108 43150
rect 19045 43046 19111 43047
rect 19045 43014 19046 43046
rect 17816 42878 17822 42910
rect 17821 42846 17822 42878
rect 17886 42878 17892 42910
rect 19040 42982 19046 43014
rect 19110 43014 19111 43046
rect 19453 43046 19519 43047
rect 19453 43014 19454 43046
rect 19110 42982 19116 43014
rect 17886 42846 17887 42878
rect 17821 42845 17887 42846
rect 19040 42774 19116 42982
rect 19040 42710 19046 42774
rect 19110 42710 19116 42774
rect 19040 42704 19116 42710
rect 19448 42982 19454 43014
rect 19518 43014 19519 43046
rect 71264 43046 71340 43052
rect 19518 42982 19524 43014
rect 19448 42774 19524 42982
rect 71264 42982 71270 43046
rect 71334 42982 71340 43046
rect 19448 42710 19454 42774
rect 19518 42710 19524 42774
rect 19448 42704 19524 42710
rect 24344 42774 24420 42780
rect 24344 42710 24350 42774
rect 24414 42710 24420 42774
rect 71264 42774 71340 42982
rect 71264 42742 71270 42774
rect 18360 42638 18436 42644
rect 18360 42574 18366 42638
rect 18430 42574 18436 42638
rect 952 42302 1230 42366
rect 1294 42302 1300 42366
rect 952 40734 1300 42302
rect 17816 42366 17892 42372
rect 17816 42302 17822 42366
rect 17886 42302 17892 42366
rect 18360 42366 18436 42574
rect 24344 42502 24420 42710
rect 71269 42710 71270 42742
rect 71334 42742 71340 42774
rect 71808 43046 71884 43052
rect 71808 42982 71814 43046
rect 71878 42982 71884 43046
rect 71808 42774 71884 42982
rect 73032 42910 73108 43118
rect 73032 42846 73038 42910
rect 73102 42846 73108 42910
rect 73032 42840 73108 42846
rect 71808 42742 71814 42774
rect 71334 42710 71335 42742
rect 71269 42709 71335 42710
rect 71813 42710 71814 42742
rect 71878 42742 71884 42774
rect 71878 42710 71879 42742
rect 71813 42709 71879 42710
rect 72080 42638 72156 42644
rect 72080 42574 72086 42638
rect 72150 42574 72156 42638
rect 24344 42470 24350 42502
rect 24349 42438 24350 42470
rect 24414 42470 24420 42502
rect 24621 42502 24687 42503
rect 24621 42470 24622 42502
rect 24414 42438 24415 42470
rect 24349 42437 24415 42438
rect 24616 42438 24622 42470
rect 24686 42470 24687 42502
rect 66509 42502 66575 42503
rect 66509 42470 66510 42502
rect 24686 42438 24692 42470
rect 18360 42334 18366 42366
rect 17816 42094 17892 42302
rect 18365 42302 18366 42334
rect 18430 42334 18436 42366
rect 18430 42302 18431 42334
rect 18365 42301 18431 42302
rect 24616 42230 24692 42438
rect 66504 42438 66510 42470
rect 66574 42470 66575 42502
rect 66574 42438 66580 42470
rect 24616 42166 24622 42230
rect 24686 42166 24692 42230
rect 66373 42230 66439 42231
rect 66373 42198 66374 42230
rect 24616 42160 24692 42166
rect 66368 42166 66374 42198
rect 66438 42198 66439 42230
rect 66504 42230 66580 42438
rect 72080 42366 72156 42574
rect 72080 42334 72086 42366
rect 72085 42302 72086 42334
rect 72150 42334 72156 42366
rect 72901 42366 72967 42367
rect 72901 42334 72902 42366
rect 72150 42302 72151 42334
rect 72085 42301 72151 42302
rect 72896 42302 72902 42334
rect 72966 42334 72967 42366
rect 89760 42366 90108 43934
rect 72966 42302 72972 42334
rect 66438 42166 66444 42198
rect 17816 42062 17822 42094
rect 17821 42030 17822 42062
rect 17886 42062 17892 42094
rect 17886 42030 17887 42062
rect 17821 42029 17887 42030
rect 17821 41958 17887 41959
rect 17821 41926 17822 41958
rect 17816 41894 17822 41926
rect 17886 41926 17887 41958
rect 18229 41958 18295 41959
rect 18229 41926 18230 41958
rect 17886 41894 17892 41926
rect 17816 41686 17892 41894
rect 17816 41622 17822 41686
rect 17886 41622 17892 41686
rect 17816 41616 17892 41622
rect 18224 41894 18230 41926
rect 18294 41926 18295 41958
rect 19176 41958 19252 41964
rect 18294 41894 18300 41926
rect 18224 41686 18300 41894
rect 19176 41894 19182 41958
rect 19246 41894 19252 41958
rect 19453 41958 19519 41959
rect 19453 41926 19454 41958
rect 19045 41822 19111 41823
rect 19045 41790 19046 41822
rect 18224 41622 18230 41686
rect 18294 41622 18300 41686
rect 18224 41616 18300 41622
rect 19040 41758 19046 41790
rect 19110 41790 19111 41822
rect 19110 41758 19116 41790
rect 17952 41550 18028 41556
rect 17952 41486 17958 41550
rect 18022 41486 18028 41550
rect 17952 41278 18028 41486
rect 17952 41246 17958 41278
rect 17957 41214 17958 41246
rect 18022 41246 18028 41278
rect 18496 41414 18572 41420
rect 18496 41350 18502 41414
rect 18566 41350 18572 41414
rect 18022 41214 18023 41246
rect 17957 41213 18023 41214
rect 17957 41142 18023 41143
rect 17957 41110 17958 41142
rect 17952 41078 17958 41110
rect 18022 41110 18023 41142
rect 18496 41142 18572 41350
rect 19040 41278 19116 41758
rect 19176 41686 19252 41894
rect 19176 41654 19182 41686
rect 19181 41622 19182 41654
rect 19246 41654 19252 41686
rect 19448 41894 19454 41926
rect 19518 41926 19519 41958
rect 66368 41958 66444 42166
rect 66504 42166 66510 42230
rect 66574 42166 66580 42230
rect 66504 42160 66580 42166
rect 72896 42094 72972 42302
rect 72896 42030 72902 42094
rect 72966 42030 72972 42094
rect 72896 42024 72972 42030
rect 89760 42302 89766 42366
rect 89830 42302 90108 42366
rect 19518 41894 19524 41926
rect 19448 41686 19524 41894
rect 66368 41894 66374 41958
rect 66438 41894 66444 41958
rect 71269 41958 71335 41959
rect 71269 41926 71270 41958
rect 66368 41888 66444 41894
rect 71264 41894 71270 41926
rect 71334 41926 71335 41958
rect 71677 41958 71743 41959
rect 71677 41926 71678 41958
rect 71334 41894 71340 41926
rect 19246 41622 19247 41654
rect 19181 41621 19247 41622
rect 19448 41622 19454 41686
rect 19518 41622 19524 41686
rect 19448 41616 19524 41622
rect 66368 41686 66444 41692
rect 66368 41622 66374 41686
rect 66438 41622 66444 41686
rect 19040 41214 19046 41278
rect 19110 41214 19116 41278
rect 19176 41550 19252 41556
rect 19176 41486 19182 41550
rect 19246 41486 19252 41550
rect 19176 41278 19252 41486
rect 19176 41246 19182 41278
rect 19040 41208 19116 41214
rect 19181 41214 19182 41246
rect 19246 41246 19252 41278
rect 19584 41550 19660 41556
rect 19584 41486 19590 41550
rect 19654 41486 19660 41550
rect 19584 41278 19660 41486
rect 66368 41414 66444 41622
rect 71264 41686 71340 41894
rect 71264 41622 71270 41686
rect 71334 41622 71340 41686
rect 71264 41616 71340 41622
rect 71672 41894 71678 41926
rect 71742 41926 71743 41958
rect 72629 41958 72695 41959
rect 72629 41926 72630 41958
rect 71742 41894 71748 41926
rect 71672 41686 71748 41894
rect 71672 41622 71678 41686
rect 71742 41622 71748 41686
rect 71672 41616 71748 41622
rect 72624 41894 72630 41926
rect 72694 41926 72695 41958
rect 73032 41958 73108 41964
rect 72694 41894 72700 41926
rect 72624 41686 72700 41894
rect 72624 41622 72630 41686
rect 72694 41622 72700 41686
rect 73032 41894 73038 41958
rect 73102 41894 73108 41958
rect 73032 41686 73108 41894
rect 73032 41654 73038 41686
rect 72624 41616 72700 41622
rect 73037 41622 73038 41654
rect 73102 41654 73108 41686
rect 73102 41622 73103 41654
rect 73037 41621 73103 41622
rect 66368 41382 66374 41414
rect 66373 41350 66374 41382
rect 66438 41382 66444 41414
rect 71400 41550 71476 41556
rect 71400 41486 71406 41550
rect 71470 41486 71476 41550
rect 66438 41350 66439 41382
rect 66373 41349 66439 41350
rect 19584 41246 19590 41278
rect 19246 41214 19247 41246
rect 19181 41213 19247 41214
rect 19589 41214 19590 41246
rect 19654 41246 19660 41278
rect 71400 41278 71476 41486
rect 71400 41246 71406 41278
rect 19654 41214 19655 41246
rect 19589 41213 19655 41214
rect 71405 41214 71406 41246
rect 71470 41246 71476 41278
rect 71808 41550 71884 41556
rect 71808 41486 71814 41550
rect 71878 41486 71884 41550
rect 72901 41550 72967 41551
rect 72901 41518 72902 41550
rect 71808 41278 71884 41486
rect 71808 41246 71814 41278
rect 71470 41214 71471 41246
rect 71405 41213 71471 41214
rect 71813 41214 71814 41246
rect 71878 41246 71884 41278
rect 72896 41486 72902 41518
rect 72966 41518 72967 41550
rect 72966 41486 72972 41518
rect 72896 41278 72972 41486
rect 71878 41214 71879 41246
rect 71813 41213 71879 41214
rect 72896 41214 72902 41278
rect 72966 41214 72972 41278
rect 72896 41208 72972 41214
rect 18496 41110 18502 41142
rect 18022 41078 18028 41110
rect 17952 40870 18028 41078
rect 18501 41078 18502 41110
rect 18566 41110 18572 41142
rect 19181 41142 19247 41143
rect 19181 41110 19182 41142
rect 18566 41078 18567 41110
rect 18501 41077 18567 41078
rect 19176 41078 19182 41110
rect 19246 41110 19247 41142
rect 19448 41142 19524 41148
rect 19246 41078 19252 41110
rect 17952 40806 17958 40870
rect 18022 40806 18028 40870
rect 17952 40800 18028 40806
rect 19176 40870 19252 41078
rect 19176 40806 19182 40870
rect 19246 40806 19252 40870
rect 19448 41078 19454 41142
rect 19518 41078 19524 41142
rect 71405 41142 71471 41143
rect 71405 41110 71406 41142
rect 19448 40870 19524 41078
rect 19448 40838 19454 40870
rect 19176 40800 19252 40806
rect 19453 40806 19454 40838
rect 19518 40838 19524 40870
rect 71400 41078 71406 41110
rect 71470 41110 71471 41142
rect 71813 41142 71879 41143
rect 71813 41110 71814 41142
rect 71470 41078 71476 41110
rect 71400 40870 71476 41078
rect 19518 40806 19519 40838
rect 19453 40805 19519 40806
rect 71400 40806 71406 40870
rect 71470 40806 71476 40870
rect 71400 40800 71476 40806
rect 71808 41078 71814 41110
rect 71878 41110 71879 41142
rect 72085 41142 72151 41143
rect 72085 41110 72086 41142
rect 71878 41078 71884 41110
rect 71808 40870 71884 41078
rect 71808 40806 71814 40870
rect 71878 40806 71884 40870
rect 71808 40800 71884 40806
rect 72080 41078 72086 41110
rect 72150 41110 72151 41142
rect 72901 41142 72967 41143
rect 72901 41110 72902 41142
rect 72150 41078 72156 41110
rect 72080 40870 72156 41078
rect 72080 40806 72086 40870
rect 72150 40806 72156 40870
rect 72080 40800 72156 40806
rect 72896 41078 72902 41110
rect 72966 41110 72967 41142
rect 72966 41078 72972 41110
rect 72896 40870 72972 41078
rect 72896 40806 72902 40870
rect 72966 40806 72972 40870
rect 72896 40800 72972 40806
rect 89760 40870 90108 42302
rect 89760 40806 89766 40870
rect 89830 40806 90108 40870
rect 952 40670 1230 40734
rect 1294 40670 1300 40734
rect 17821 40734 17887 40735
rect 17821 40702 17822 40734
rect 952 39238 1300 40670
rect 17816 40670 17822 40702
rect 17886 40702 17887 40734
rect 18360 40734 18436 40740
rect 17886 40670 17892 40702
rect 17816 40462 17892 40670
rect 17816 40398 17822 40462
rect 17886 40398 17892 40462
rect 18360 40670 18366 40734
rect 18430 40670 18436 40734
rect 18360 40462 18436 40670
rect 18360 40430 18366 40462
rect 17816 40392 17892 40398
rect 18365 40398 18366 40430
rect 18430 40430 18436 40462
rect 18496 40734 18572 40740
rect 18496 40670 18502 40734
rect 18566 40670 18572 40734
rect 18496 40462 18572 40670
rect 18496 40430 18502 40462
rect 18430 40398 18431 40430
rect 18365 40397 18431 40398
rect 18501 40398 18502 40430
rect 18566 40430 18572 40462
rect 19176 40734 19252 40740
rect 19176 40670 19182 40734
rect 19246 40670 19252 40734
rect 19453 40734 19519 40735
rect 19453 40702 19454 40734
rect 19176 40462 19252 40670
rect 19176 40430 19182 40462
rect 18566 40398 18567 40430
rect 18501 40397 18567 40398
rect 19181 40398 19182 40430
rect 19246 40430 19252 40462
rect 19448 40670 19454 40702
rect 19518 40702 19519 40734
rect 71400 40734 71476 40740
rect 19518 40670 19524 40702
rect 19448 40462 19524 40670
rect 19246 40398 19247 40430
rect 19181 40397 19247 40398
rect 19448 40398 19454 40462
rect 19518 40398 19524 40462
rect 71400 40670 71406 40734
rect 71470 40670 71476 40734
rect 71677 40734 71743 40735
rect 71677 40702 71678 40734
rect 71400 40462 71476 40670
rect 71400 40430 71406 40462
rect 19448 40392 19524 40398
rect 71405 40398 71406 40430
rect 71470 40430 71476 40462
rect 71672 40670 71678 40702
rect 71742 40702 71743 40734
rect 72488 40734 72564 40740
rect 71742 40670 71748 40702
rect 71672 40462 71748 40670
rect 71470 40398 71471 40430
rect 71405 40397 71471 40398
rect 71672 40398 71678 40462
rect 71742 40398 71748 40462
rect 72488 40670 72494 40734
rect 72558 40670 72564 40734
rect 72488 40462 72564 40670
rect 72488 40430 72494 40462
rect 71672 40392 71748 40398
rect 72493 40398 72494 40430
rect 72558 40430 72564 40462
rect 72896 40734 72972 40740
rect 72896 40670 72902 40734
rect 72966 40670 72972 40734
rect 72896 40462 72972 40670
rect 72896 40430 72902 40462
rect 72558 40398 72559 40430
rect 72493 40397 72559 40398
rect 72901 40398 72902 40430
rect 72966 40430 72972 40462
rect 72966 40398 72967 40430
rect 72901 40397 72967 40398
rect 17952 40326 18028 40332
rect 17952 40262 17958 40326
rect 18022 40262 18028 40326
rect 17952 40054 18028 40262
rect 17952 40022 17958 40054
rect 17957 39990 17958 40022
rect 18022 40022 18028 40054
rect 18632 40326 18708 40332
rect 18632 40262 18638 40326
rect 18702 40262 18708 40326
rect 19181 40326 19247 40327
rect 19181 40294 19182 40326
rect 18632 40054 18708 40262
rect 18632 40022 18638 40054
rect 18022 39990 18023 40022
rect 17957 39989 18023 39990
rect 18637 39990 18638 40022
rect 18702 40022 18708 40054
rect 19176 40262 19182 40294
rect 19246 40294 19247 40326
rect 19584 40326 19660 40332
rect 19246 40262 19252 40294
rect 19176 40054 19252 40262
rect 18702 39990 18703 40022
rect 18637 39989 18703 39990
rect 19176 39990 19182 40054
rect 19246 39990 19252 40054
rect 19584 40262 19590 40326
rect 19654 40262 19660 40326
rect 71405 40326 71471 40327
rect 71405 40294 71406 40326
rect 19584 40054 19660 40262
rect 19584 40022 19590 40054
rect 19176 39984 19252 39990
rect 19589 39990 19590 40022
rect 19654 40022 19660 40054
rect 71400 40262 71406 40294
rect 71470 40294 71471 40326
rect 71677 40326 71743 40327
rect 71677 40294 71678 40326
rect 71470 40262 71476 40294
rect 71400 40054 71476 40262
rect 19654 39990 19655 40022
rect 19589 39989 19655 39990
rect 71400 39990 71406 40054
rect 71470 39990 71476 40054
rect 71400 39984 71476 39990
rect 71672 40262 71678 40294
rect 71742 40294 71743 40326
rect 72085 40326 72151 40327
rect 72085 40294 72086 40326
rect 71742 40262 71748 40294
rect 71672 40054 71748 40262
rect 71672 39990 71678 40054
rect 71742 39990 71748 40054
rect 71672 39984 71748 39990
rect 72080 40262 72086 40294
rect 72150 40294 72151 40326
rect 72352 40326 72428 40332
rect 72150 40262 72156 40294
rect 72080 40054 72156 40262
rect 72080 39990 72086 40054
rect 72150 39990 72156 40054
rect 72352 40262 72358 40326
rect 72422 40262 72428 40326
rect 72901 40326 72967 40327
rect 72901 40294 72902 40326
rect 72352 40054 72428 40262
rect 72352 40022 72358 40054
rect 72080 39984 72156 39990
rect 72357 39990 72358 40022
rect 72422 40022 72428 40054
rect 72896 40262 72902 40294
rect 72966 40294 72967 40326
rect 72966 40262 72972 40294
rect 72896 40054 72972 40262
rect 72422 39990 72423 40022
rect 72357 39989 72423 39990
rect 72896 39990 72902 40054
rect 72966 39990 72972 40054
rect 72896 39984 72972 39990
rect 17821 39918 17887 39919
rect 17821 39886 17822 39918
rect 17816 39854 17822 39886
rect 17886 39886 17887 39918
rect 18229 39918 18295 39919
rect 18229 39886 18230 39918
rect 17886 39854 17892 39886
rect 17816 39646 17892 39854
rect 17816 39582 17822 39646
rect 17886 39582 17892 39646
rect 17816 39576 17892 39582
rect 18224 39854 18230 39886
rect 18294 39886 18295 39918
rect 18909 39918 18975 39919
rect 18909 39886 18910 39918
rect 18294 39854 18300 39886
rect 18224 39646 18300 39854
rect 18224 39582 18230 39646
rect 18294 39582 18300 39646
rect 18224 39576 18300 39582
rect 18904 39854 18910 39886
rect 18974 39886 18975 39918
rect 19045 39918 19111 39919
rect 19045 39886 19046 39918
rect 18974 39854 18980 39886
rect 18904 39646 18980 39854
rect 18904 39582 18910 39646
rect 18974 39582 18980 39646
rect 18904 39576 18980 39582
rect 19040 39854 19046 39886
rect 19110 39886 19111 39918
rect 19584 39918 19660 39924
rect 19110 39854 19116 39886
rect 19040 39646 19116 39854
rect 19040 39582 19046 39646
rect 19110 39582 19116 39646
rect 19584 39854 19590 39918
rect 19654 39854 19660 39918
rect 71269 39918 71335 39919
rect 71269 39886 71270 39918
rect 19584 39646 19660 39854
rect 19584 39614 19590 39646
rect 19040 39576 19116 39582
rect 19589 39582 19590 39614
rect 19654 39614 19660 39646
rect 71264 39854 71270 39886
rect 71334 39886 71335 39918
rect 71808 39918 71884 39924
rect 71334 39854 71340 39886
rect 71264 39646 71340 39854
rect 19654 39582 19655 39614
rect 19589 39581 19655 39582
rect 71264 39582 71270 39646
rect 71334 39582 71340 39646
rect 71808 39854 71814 39918
rect 71878 39854 71884 39918
rect 72221 39918 72287 39919
rect 72221 39886 72222 39918
rect 71808 39646 71884 39854
rect 71808 39614 71814 39646
rect 71264 39576 71340 39582
rect 71813 39582 71814 39614
rect 71878 39614 71884 39646
rect 72216 39854 72222 39886
rect 72286 39886 72287 39918
rect 72357 39918 72423 39919
rect 72357 39886 72358 39918
rect 72286 39854 72292 39886
rect 72216 39646 72292 39854
rect 71878 39582 71879 39614
rect 71813 39581 71879 39582
rect 72216 39582 72222 39646
rect 72286 39582 72292 39646
rect 72216 39576 72292 39582
rect 72352 39854 72358 39886
rect 72422 39886 72423 39918
rect 73032 39918 73108 39924
rect 72422 39854 72428 39886
rect 72352 39646 72428 39854
rect 72352 39582 72358 39646
rect 72422 39582 72428 39646
rect 73032 39854 73038 39918
rect 73102 39854 73108 39918
rect 73032 39646 73108 39854
rect 73032 39614 73038 39646
rect 72352 39576 72428 39582
rect 73037 39582 73038 39614
rect 73102 39614 73108 39646
rect 73102 39582 73103 39614
rect 73037 39581 73103 39582
rect 952 39174 1230 39238
rect 1294 39174 1300 39238
rect 18360 39510 18436 39516
rect 18360 39446 18366 39510
rect 18430 39446 18436 39510
rect 18360 39238 18436 39446
rect 18360 39206 18366 39238
rect 952 37334 1300 39174
rect 18365 39174 18366 39206
rect 18430 39206 18436 39238
rect 18496 39510 18572 39516
rect 18496 39446 18502 39510
rect 18566 39446 18572 39510
rect 18496 39238 18572 39446
rect 18496 39206 18502 39238
rect 18430 39174 18431 39206
rect 18365 39173 18431 39174
rect 18501 39174 18502 39206
rect 18566 39206 18572 39238
rect 18768 39510 18844 39516
rect 18768 39446 18774 39510
rect 18838 39446 18844 39510
rect 18768 39238 18844 39446
rect 18768 39206 18774 39238
rect 18566 39174 18567 39206
rect 18501 39173 18567 39174
rect 18773 39174 18774 39206
rect 18838 39206 18844 39238
rect 19176 39510 19252 39516
rect 19176 39446 19182 39510
rect 19246 39446 19252 39510
rect 19176 39238 19252 39446
rect 19176 39206 19182 39238
rect 18838 39174 18839 39206
rect 18773 39173 18839 39174
rect 19181 39174 19182 39206
rect 19246 39206 19252 39238
rect 19448 39510 19524 39516
rect 19448 39446 19454 39510
rect 19518 39446 19524 39510
rect 71269 39510 71335 39511
rect 71269 39478 71270 39510
rect 19448 39238 19524 39446
rect 71264 39446 71270 39478
rect 71334 39478 71335 39510
rect 71808 39510 71884 39516
rect 71334 39446 71340 39478
rect 19448 39206 19454 39238
rect 19246 39174 19247 39206
rect 19181 39173 19247 39174
rect 19453 39174 19454 39206
rect 19518 39206 19524 39238
rect 24344 39374 24420 39380
rect 24344 39310 24350 39374
rect 24414 39310 24420 39374
rect 19518 39174 19519 39206
rect 19453 39173 19519 39174
rect 19040 39102 19116 39108
rect 19040 39038 19046 39102
rect 19110 39038 19116 39102
rect 19453 39102 19519 39103
rect 19453 39070 19454 39102
rect 19040 38830 19116 39038
rect 19040 38798 19046 38830
rect 19045 38766 19046 38798
rect 19110 38798 19116 38830
rect 19448 39038 19454 39070
rect 19518 39070 19519 39102
rect 24344 39102 24420 39310
rect 24344 39070 24350 39102
rect 19518 39038 19524 39070
rect 19448 38830 19524 39038
rect 24349 39038 24350 39070
rect 24414 39070 24420 39102
rect 66368 39374 66444 39380
rect 66368 39310 66374 39374
rect 66438 39310 66444 39374
rect 66368 39102 66444 39310
rect 71264 39238 71340 39446
rect 71264 39174 71270 39238
rect 71334 39174 71340 39238
rect 71808 39446 71814 39510
rect 71878 39446 71884 39510
rect 71808 39238 71884 39446
rect 71808 39206 71814 39238
rect 71264 39168 71340 39174
rect 71813 39174 71814 39206
rect 71878 39206 71884 39238
rect 72080 39510 72156 39516
rect 72080 39446 72086 39510
rect 72150 39446 72156 39510
rect 72080 39238 72156 39446
rect 72080 39206 72086 39238
rect 71878 39174 71879 39206
rect 71813 39173 71879 39174
rect 72085 39174 72086 39206
rect 72150 39206 72156 39238
rect 89760 39238 90108 40806
rect 72150 39174 72151 39206
rect 72085 39173 72151 39174
rect 89760 39174 89766 39238
rect 89830 39174 90108 39238
rect 66368 39070 66374 39102
rect 24414 39038 24415 39070
rect 24349 39037 24415 39038
rect 66373 39038 66374 39070
rect 66438 39070 66444 39102
rect 71264 39102 71340 39108
rect 66438 39038 66439 39070
rect 66373 39037 66439 39038
rect 71264 39038 71270 39102
rect 71334 39038 71340 39102
rect 71813 39102 71879 39103
rect 71813 39070 71814 39102
rect 19110 38766 19111 38798
rect 19045 38765 19111 38766
rect 19448 38766 19454 38830
rect 19518 38766 19524 38830
rect 19448 38760 19524 38766
rect 66504 38830 66580 38836
rect 66504 38766 66510 38830
rect 66574 38766 66580 38830
rect 71264 38830 71340 39038
rect 71264 38798 71270 38830
rect 18904 38694 18980 38700
rect 18904 38630 18910 38694
rect 18974 38630 18980 38694
rect 17816 38422 17892 38428
rect 17816 38358 17822 38422
rect 17886 38358 17892 38422
rect 18904 38422 18980 38630
rect 66504 38558 66580 38766
rect 71269 38766 71270 38798
rect 71334 38798 71340 38830
rect 71808 39038 71814 39070
rect 71878 39070 71879 39102
rect 71878 39038 71884 39070
rect 71808 38830 71884 39038
rect 71334 38766 71335 38798
rect 71269 38765 71335 38766
rect 71808 38766 71814 38830
rect 71878 38766 71884 38830
rect 71808 38760 71884 38766
rect 66504 38526 66510 38558
rect 66509 38494 66510 38526
rect 66574 38526 66580 38558
rect 72216 38694 72292 38700
rect 72216 38630 72222 38694
rect 72286 38630 72292 38694
rect 66574 38494 66575 38526
rect 66509 38493 66575 38494
rect 18904 38390 18910 38422
rect 17816 38150 17892 38358
rect 18909 38358 18910 38390
rect 18974 38390 18980 38422
rect 72216 38422 72292 38630
rect 72216 38390 72222 38422
rect 18974 38358 18975 38390
rect 18909 38357 18975 38358
rect 72221 38358 72222 38390
rect 72286 38390 72292 38422
rect 72896 38422 72972 38428
rect 72286 38358 72287 38390
rect 72221 38357 72287 38358
rect 72896 38358 72902 38422
rect 72966 38358 72972 38422
rect 17816 38118 17822 38150
rect 17821 38086 17822 38118
rect 17886 38118 17892 38150
rect 24621 38150 24687 38151
rect 24621 38118 24622 38150
rect 17886 38086 17887 38118
rect 17821 38085 17887 38086
rect 24616 38086 24622 38118
rect 24686 38118 24687 38150
rect 66373 38150 66439 38151
rect 66373 38118 66374 38150
rect 24686 38086 24692 38118
rect 11157 38014 11223 38015
rect 11157 37982 11158 38014
rect 952 37270 1230 37334
rect 1294 37270 1300 37334
rect 952 35702 1300 37270
rect 952 35638 1230 35702
rect 1294 35638 1300 35702
rect 952 34070 1300 35638
rect 11152 37950 11158 37982
rect 11222 37982 11223 38014
rect 17816 38014 17892 38020
rect 11222 37950 11228 37982
rect 11152 35294 11228 37950
rect 17816 37950 17822 38014
rect 17886 37950 17892 38014
rect 18501 38014 18567 38015
rect 18501 37982 18502 38014
rect 17816 37742 17892 37950
rect 17816 37710 17822 37742
rect 17821 37678 17822 37710
rect 17886 37710 17892 37742
rect 18496 37950 18502 37982
rect 18566 37982 18567 38014
rect 18566 37950 18572 37982
rect 18496 37742 18572 37950
rect 24616 37878 24692 38086
rect 24616 37814 24622 37878
rect 24686 37814 24692 37878
rect 24616 37808 24692 37814
rect 66368 38086 66374 38118
rect 66438 38118 66439 38150
rect 66504 38150 66580 38156
rect 66438 38086 66444 38118
rect 66368 37878 66444 38086
rect 66368 37814 66374 37878
rect 66438 37814 66444 37878
rect 66368 37808 66444 37814
rect 66504 38086 66510 38150
rect 66574 38086 66580 38150
rect 72896 38150 72972 38358
rect 72896 38118 72902 38150
rect 17886 37678 17887 37710
rect 17821 37677 17887 37678
rect 18496 37678 18502 37742
rect 18566 37678 18572 37742
rect 66504 37742 66580 38086
rect 72901 38086 72902 38118
rect 72966 38118 72972 38150
rect 72966 38086 72967 38118
rect 72901 38085 72967 38086
rect 72085 38014 72151 38015
rect 72085 37982 72086 38014
rect 66504 37710 66510 37742
rect 18496 37672 18572 37678
rect 66509 37678 66510 37710
rect 66574 37710 66580 37742
rect 72080 37950 72086 37982
rect 72150 37982 72151 38014
rect 72901 38014 72967 38015
rect 72901 37982 72902 38014
rect 72150 37950 72156 37982
rect 72080 37742 72156 37950
rect 66574 37678 66575 37710
rect 66509 37677 66575 37678
rect 72080 37678 72086 37742
rect 72150 37678 72156 37742
rect 72080 37672 72156 37678
rect 72896 37950 72902 37982
rect 72966 37982 72967 38014
rect 72966 37950 72972 37982
rect 72896 37742 72972 37950
rect 72896 37678 72902 37742
rect 72966 37678 72972 37742
rect 72896 37672 72972 37678
rect 17952 37606 18028 37612
rect 17952 37542 17958 37606
rect 18022 37542 18028 37606
rect 19045 37606 19111 37607
rect 19045 37574 19046 37606
rect 17952 37334 18028 37542
rect 17952 37302 17958 37334
rect 17957 37270 17958 37302
rect 18022 37302 18028 37334
rect 19040 37542 19046 37574
rect 19110 37574 19111 37606
rect 19584 37606 19660 37612
rect 19110 37542 19116 37574
rect 19040 37334 19116 37542
rect 18022 37270 18023 37302
rect 17957 37269 18023 37270
rect 19040 37270 19046 37334
rect 19110 37270 19116 37334
rect 19584 37542 19590 37606
rect 19654 37542 19660 37606
rect 19584 37334 19660 37542
rect 19584 37302 19590 37334
rect 19040 37264 19116 37270
rect 19589 37270 19590 37302
rect 19654 37302 19660 37334
rect 71264 37606 71340 37612
rect 71264 37542 71270 37606
rect 71334 37542 71340 37606
rect 71677 37606 71743 37607
rect 71677 37574 71678 37606
rect 71264 37334 71340 37542
rect 71264 37302 71270 37334
rect 19654 37270 19655 37302
rect 19589 37269 19655 37270
rect 71269 37270 71270 37302
rect 71334 37302 71340 37334
rect 71672 37542 71678 37574
rect 71742 37574 71743 37606
rect 73032 37606 73108 37612
rect 71742 37542 71748 37574
rect 71672 37334 71748 37542
rect 71334 37270 71335 37302
rect 71269 37269 71335 37270
rect 71672 37270 71678 37334
rect 71742 37270 71748 37334
rect 73032 37542 73038 37606
rect 73102 37542 73108 37606
rect 73032 37334 73108 37542
rect 73032 37302 73038 37334
rect 71672 37264 71748 37270
rect 73037 37270 73038 37302
rect 73102 37302 73108 37334
rect 89760 37334 90108 39174
rect 73102 37270 73103 37302
rect 73037 37269 73103 37270
rect 89760 37270 89766 37334
rect 89830 37270 90108 37334
rect 17821 37198 17887 37199
rect 17821 37166 17822 37198
rect 17816 37134 17822 37166
rect 17886 37166 17887 37198
rect 18365 37198 18431 37199
rect 18365 37166 18366 37198
rect 17886 37134 17892 37166
rect 17816 36926 17892 37134
rect 17816 36862 17822 36926
rect 17886 36862 17892 36926
rect 17816 36856 17892 36862
rect 18360 37134 18366 37166
rect 18430 37166 18431 37198
rect 19176 37198 19252 37204
rect 18430 37134 18436 37166
rect 18360 36926 18436 37134
rect 18360 36862 18366 36926
rect 18430 36862 18436 36926
rect 19176 37134 19182 37198
rect 19246 37134 19252 37198
rect 19453 37198 19519 37199
rect 19453 37166 19454 37198
rect 19176 36926 19252 37134
rect 19176 36894 19182 36926
rect 18360 36856 18436 36862
rect 19181 36862 19182 36894
rect 19246 36894 19252 36926
rect 19448 37134 19454 37166
rect 19518 37166 19519 37198
rect 71405 37198 71471 37199
rect 71405 37166 71406 37198
rect 19518 37134 19524 37166
rect 19448 36926 19524 37134
rect 71400 37134 71406 37166
rect 71470 37166 71471 37198
rect 71677 37198 71743 37199
rect 71677 37166 71678 37198
rect 71470 37134 71476 37166
rect 19246 36862 19247 36894
rect 19181 36861 19247 36862
rect 19448 36862 19454 36926
rect 19518 36862 19524 36926
rect 24621 36926 24687 36927
rect 24621 36894 24622 36926
rect 19448 36856 19524 36862
rect 24616 36862 24622 36894
rect 24686 36894 24687 36926
rect 66373 36926 66439 36927
rect 66373 36894 66374 36926
rect 24686 36862 24692 36894
rect 17957 36790 18023 36791
rect 17957 36758 17958 36790
rect 17952 36726 17958 36758
rect 18022 36758 18023 36790
rect 18224 36790 18300 36796
rect 18022 36726 18028 36758
rect 11152 35230 11158 35294
rect 11222 35230 11228 35294
rect 11152 35224 11228 35230
rect 11288 36518 11364 36524
rect 11288 36454 11294 36518
rect 11358 36454 11364 36518
rect 952 34006 1230 34070
rect 1294 34006 1300 34070
rect 952 32302 1300 34006
rect 11016 35158 11092 35164
rect 11016 35094 11022 35158
rect 11086 35094 11092 35158
rect 11016 32438 11092 35094
rect 11288 33934 11364 36454
rect 17952 36518 18028 36726
rect 17952 36454 17958 36518
rect 18022 36454 18028 36518
rect 18224 36726 18230 36790
rect 18294 36726 18300 36790
rect 18224 36518 18300 36726
rect 18224 36486 18230 36518
rect 17952 36448 18028 36454
rect 18229 36454 18230 36486
rect 18294 36486 18300 36518
rect 18904 36790 18980 36796
rect 18904 36726 18910 36790
rect 18974 36726 18980 36790
rect 19181 36790 19247 36791
rect 19181 36758 19182 36790
rect 18904 36518 18980 36726
rect 18904 36486 18910 36518
rect 18294 36454 18295 36486
rect 18229 36453 18295 36454
rect 18909 36454 18910 36486
rect 18974 36486 18980 36518
rect 19176 36726 19182 36758
rect 19246 36758 19247 36790
rect 19589 36790 19655 36791
rect 19589 36758 19590 36790
rect 19246 36726 19252 36758
rect 19176 36518 19252 36726
rect 18974 36454 18975 36486
rect 18909 36453 18975 36454
rect 19176 36454 19182 36518
rect 19246 36454 19252 36518
rect 19176 36448 19252 36454
rect 19584 36726 19590 36758
rect 19654 36758 19655 36790
rect 19654 36726 19660 36758
rect 19584 36518 19660 36726
rect 24616 36654 24692 36862
rect 24616 36590 24622 36654
rect 24686 36590 24692 36654
rect 24616 36584 24692 36590
rect 66368 36862 66374 36894
rect 66438 36894 66439 36926
rect 71400 36926 71476 37134
rect 66438 36862 66444 36894
rect 66368 36654 66444 36862
rect 71400 36862 71406 36926
rect 71470 36862 71476 36926
rect 71400 36856 71476 36862
rect 71672 37134 71678 37166
rect 71742 37166 71743 37198
rect 72493 37198 72559 37199
rect 72493 37166 72494 37198
rect 71742 37134 71748 37166
rect 71672 36926 71748 37134
rect 71672 36862 71678 36926
rect 71742 36862 71748 36926
rect 71672 36856 71748 36862
rect 72488 37134 72494 37166
rect 72558 37166 72559 37198
rect 72901 37198 72967 37199
rect 72901 37166 72902 37198
rect 72558 37134 72564 37166
rect 72488 36926 72564 37134
rect 72488 36862 72494 36926
rect 72558 36862 72564 36926
rect 72488 36856 72564 36862
rect 72896 37134 72902 37166
rect 72966 37166 72967 37198
rect 72966 37134 72972 37166
rect 72896 36926 72972 37134
rect 72896 36862 72902 36926
rect 72966 36862 72972 36926
rect 72896 36856 72972 36862
rect 66368 36590 66374 36654
rect 66438 36590 66444 36654
rect 66368 36584 66444 36590
rect 71264 36790 71340 36796
rect 71264 36726 71270 36790
rect 71334 36726 71340 36790
rect 19584 36454 19590 36518
rect 19654 36454 19660 36518
rect 71264 36518 71340 36726
rect 71264 36486 71270 36518
rect 19584 36448 19660 36454
rect 71269 36454 71270 36486
rect 71334 36486 71340 36518
rect 71672 36790 71748 36796
rect 71672 36726 71678 36790
rect 71742 36726 71748 36790
rect 72085 36790 72151 36791
rect 72085 36758 72086 36790
rect 71672 36518 71748 36726
rect 71672 36486 71678 36518
rect 71334 36454 71335 36486
rect 71269 36453 71335 36454
rect 71677 36454 71678 36486
rect 71742 36486 71748 36518
rect 72080 36726 72086 36758
rect 72150 36758 72151 36790
rect 72352 36790 72428 36796
rect 72150 36726 72156 36758
rect 72080 36518 72156 36726
rect 71742 36454 71743 36486
rect 71677 36453 71743 36454
rect 72080 36454 72086 36518
rect 72150 36454 72156 36518
rect 72352 36726 72358 36790
rect 72422 36726 72428 36790
rect 72352 36518 72428 36726
rect 72352 36486 72358 36518
rect 72080 36448 72156 36454
rect 72357 36454 72358 36486
rect 72422 36486 72428 36518
rect 73032 36790 73108 36796
rect 73032 36726 73038 36790
rect 73102 36726 73108 36790
rect 73032 36518 73108 36726
rect 73032 36486 73038 36518
rect 72422 36454 72423 36486
rect 72357 36453 72423 36454
rect 73037 36454 73038 36486
rect 73102 36486 73108 36518
rect 73102 36454 73103 36486
rect 73037 36453 73103 36454
rect 17816 36382 17892 36388
rect 17816 36318 17822 36382
rect 17886 36318 17892 36382
rect 19045 36382 19111 36383
rect 19045 36350 19046 36382
rect 17816 36110 17892 36318
rect 17816 36078 17822 36110
rect 17821 36046 17822 36078
rect 17886 36078 17892 36110
rect 19040 36318 19046 36350
rect 19110 36350 19111 36382
rect 19448 36382 19524 36388
rect 19110 36318 19116 36350
rect 19040 36110 19116 36318
rect 17886 36046 17887 36078
rect 17821 36045 17887 36046
rect 19040 36046 19046 36110
rect 19110 36046 19116 36110
rect 19448 36318 19454 36382
rect 19518 36318 19524 36382
rect 71269 36382 71335 36383
rect 71269 36350 71270 36382
rect 19448 36110 19524 36318
rect 19448 36078 19454 36110
rect 19040 36040 19116 36046
rect 19453 36046 19454 36078
rect 19518 36078 19524 36110
rect 71264 36318 71270 36350
rect 71334 36350 71335 36382
rect 71672 36382 71748 36388
rect 71334 36318 71340 36350
rect 71264 36110 71340 36318
rect 19518 36046 19519 36078
rect 19453 36045 19519 36046
rect 71264 36046 71270 36110
rect 71334 36046 71340 36110
rect 71672 36318 71678 36382
rect 71742 36318 71748 36382
rect 71672 36110 71748 36318
rect 71672 36078 71678 36110
rect 71264 36040 71340 36046
rect 71677 36046 71678 36078
rect 71742 36078 71748 36110
rect 72488 36382 72564 36388
rect 72488 36318 72494 36382
rect 72558 36318 72564 36382
rect 72488 36110 72564 36318
rect 72488 36078 72494 36110
rect 71742 36046 71743 36078
rect 71677 36045 71743 36046
rect 72493 36046 72494 36078
rect 72558 36078 72564 36110
rect 72896 36382 72972 36388
rect 72896 36318 72902 36382
rect 72966 36318 72972 36382
rect 72896 36110 72972 36318
rect 72896 36078 72902 36110
rect 72558 36046 72559 36078
rect 72493 36045 72559 36046
rect 72901 36046 72902 36078
rect 72966 36078 72972 36110
rect 72966 36046 72967 36078
rect 72901 36045 72967 36046
rect 17821 35974 17887 35975
rect 17821 35942 17822 35974
rect 17816 35910 17822 35942
rect 17886 35942 17887 35974
rect 18909 35974 18975 35975
rect 18909 35942 18910 35974
rect 17886 35910 17892 35942
rect 17816 35702 17892 35910
rect 17816 35638 17822 35702
rect 17886 35638 17892 35702
rect 17816 35632 17892 35638
rect 18904 35910 18910 35942
rect 18974 35942 18975 35974
rect 19176 35974 19252 35980
rect 18974 35910 18980 35942
rect 18904 35702 18980 35910
rect 18904 35638 18910 35702
rect 18974 35638 18980 35702
rect 19176 35910 19182 35974
rect 19246 35910 19252 35974
rect 19453 35974 19519 35975
rect 19453 35942 19454 35974
rect 19176 35702 19252 35910
rect 19176 35670 19182 35702
rect 18904 35632 18980 35638
rect 19181 35638 19182 35670
rect 19246 35670 19252 35702
rect 19448 35910 19454 35942
rect 19518 35942 19519 35974
rect 71400 35974 71476 35980
rect 19518 35910 19524 35942
rect 19448 35702 19524 35910
rect 19246 35638 19247 35670
rect 19181 35637 19247 35638
rect 19448 35638 19454 35702
rect 19518 35638 19524 35702
rect 71400 35910 71406 35974
rect 71470 35910 71476 35974
rect 71677 35974 71743 35975
rect 71677 35942 71678 35974
rect 71400 35702 71476 35910
rect 71400 35670 71406 35702
rect 19448 35632 19524 35638
rect 71405 35638 71406 35670
rect 71470 35670 71476 35702
rect 71672 35910 71678 35942
rect 71742 35942 71743 35974
rect 72085 35974 72151 35975
rect 72085 35942 72086 35974
rect 71742 35910 71748 35942
rect 71672 35702 71748 35910
rect 71470 35638 71471 35670
rect 71405 35637 71471 35638
rect 71672 35638 71678 35702
rect 71742 35638 71748 35702
rect 71672 35632 71748 35638
rect 72080 35910 72086 35942
rect 72150 35942 72151 35974
rect 72352 35974 72428 35980
rect 72150 35910 72156 35942
rect 72080 35702 72156 35910
rect 72080 35638 72086 35702
rect 72150 35638 72156 35702
rect 72352 35910 72358 35974
rect 72422 35910 72428 35974
rect 72901 35974 72967 35975
rect 72901 35942 72902 35974
rect 72352 35702 72428 35910
rect 72352 35670 72358 35702
rect 72080 35632 72156 35638
rect 72357 35638 72358 35670
rect 72422 35670 72428 35702
rect 72896 35910 72902 35942
rect 72966 35942 72967 35974
rect 72966 35910 72972 35942
rect 72896 35702 72972 35910
rect 72422 35638 72423 35670
rect 72357 35637 72423 35638
rect 72896 35638 72902 35702
rect 72966 35638 72972 35702
rect 72896 35632 72972 35638
rect 89760 35702 90108 37270
rect 89760 35638 89766 35702
rect 89830 35638 90108 35702
rect 18501 35566 18567 35567
rect 18501 35534 18502 35566
rect 18496 35502 18502 35534
rect 18566 35534 18567 35566
rect 18909 35566 18975 35567
rect 18909 35534 18910 35566
rect 18566 35502 18572 35534
rect 18496 35294 18572 35502
rect 18496 35230 18502 35294
rect 18566 35230 18572 35294
rect 18496 35224 18572 35230
rect 18904 35502 18910 35534
rect 18974 35534 18975 35566
rect 19040 35566 19116 35572
rect 18974 35502 18980 35534
rect 18904 35294 18980 35502
rect 18904 35230 18910 35294
rect 18974 35230 18980 35294
rect 19040 35502 19046 35566
rect 19110 35502 19116 35566
rect 19040 35294 19116 35502
rect 19040 35262 19046 35294
rect 18904 35224 18980 35230
rect 19045 35230 19046 35262
rect 19110 35262 19116 35294
rect 19584 35566 19660 35572
rect 19584 35502 19590 35566
rect 19654 35502 19660 35566
rect 71269 35566 71335 35567
rect 71269 35534 71270 35566
rect 19584 35294 19660 35502
rect 19584 35262 19590 35294
rect 19110 35230 19111 35262
rect 19045 35229 19111 35230
rect 19589 35230 19590 35262
rect 19654 35262 19660 35294
rect 71264 35502 71270 35534
rect 71334 35534 71335 35566
rect 71808 35566 71884 35572
rect 71334 35502 71340 35534
rect 71264 35294 71340 35502
rect 19654 35230 19655 35262
rect 19589 35229 19655 35230
rect 71264 35230 71270 35294
rect 71334 35230 71340 35294
rect 71808 35502 71814 35566
rect 71878 35502 71884 35566
rect 71808 35294 71884 35502
rect 71808 35262 71814 35294
rect 71264 35224 71340 35230
rect 71813 35230 71814 35262
rect 71878 35262 71884 35294
rect 72216 35566 72292 35572
rect 72216 35502 72222 35566
rect 72286 35502 72292 35566
rect 72216 35294 72292 35502
rect 72216 35262 72222 35294
rect 71878 35230 71879 35262
rect 71813 35229 71879 35230
rect 72221 35230 72222 35262
rect 72286 35262 72292 35294
rect 72352 35566 72428 35572
rect 72352 35502 72358 35566
rect 72422 35502 72428 35566
rect 72352 35294 72428 35502
rect 72352 35262 72358 35294
rect 72286 35230 72287 35262
rect 72221 35229 72287 35230
rect 72357 35230 72358 35262
rect 72422 35262 72428 35294
rect 72422 35230 72423 35262
rect 72357 35229 72423 35230
rect 19045 35158 19111 35159
rect 19045 35126 19046 35158
rect 19040 35094 19046 35126
rect 19110 35126 19111 35158
rect 19448 35158 19524 35164
rect 19110 35094 19116 35126
rect 19040 34886 19116 35094
rect 19040 34822 19046 34886
rect 19110 34822 19116 34886
rect 19448 35094 19454 35158
rect 19518 35094 19524 35158
rect 71269 35158 71335 35159
rect 71269 35126 71270 35158
rect 19448 34886 19524 35094
rect 19448 34854 19454 34886
rect 19040 34816 19116 34822
rect 19453 34822 19454 34854
rect 19518 34854 19524 34886
rect 71264 35094 71270 35126
rect 71334 35126 71335 35158
rect 71813 35158 71879 35159
rect 71813 35126 71814 35158
rect 71334 35094 71340 35126
rect 71264 34886 71340 35094
rect 19518 34822 19519 34854
rect 19453 34821 19519 34822
rect 71264 34822 71270 34886
rect 71334 34822 71340 34886
rect 71264 34816 71340 34822
rect 71808 35094 71814 35126
rect 71878 35126 71879 35158
rect 71878 35094 71884 35126
rect 71808 34886 71884 35094
rect 71808 34822 71814 34886
rect 71878 34822 71884 34886
rect 71808 34816 71884 34822
rect 18637 34750 18703 34751
rect 18637 34718 18638 34750
rect 18632 34686 18638 34718
rect 18702 34718 18703 34750
rect 19040 34750 19116 34756
rect 18702 34686 18708 34718
rect 17952 34478 18028 34484
rect 17952 34414 17958 34478
rect 18022 34414 18028 34478
rect 17952 34206 18028 34414
rect 18632 34478 18708 34686
rect 18632 34414 18638 34478
rect 18702 34414 18708 34478
rect 19040 34686 19046 34750
rect 19110 34686 19116 34750
rect 19453 34750 19519 34751
rect 19453 34718 19454 34750
rect 19040 34478 19116 34686
rect 19040 34446 19046 34478
rect 18632 34408 18708 34414
rect 19045 34414 19046 34446
rect 19110 34446 19116 34478
rect 19448 34686 19454 34718
rect 19518 34718 19519 34750
rect 71264 34750 71340 34756
rect 19518 34686 19524 34718
rect 19448 34478 19524 34686
rect 71264 34686 71270 34750
rect 71334 34686 71340 34750
rect 24621 34614 24687 34615
rect 24621 34582 24622 34614
rect 19110 34414 19111 34446
rect 19045 34413 19111 34414
rect 19448 34414 19454 34478
rect 19518 34414 19524 34478
rect 19448 34408 19524 34414
rect 24616 34550 24622 34582
rect 24686 34582 24687 34614
rect 24686 34550 24692 34582
rect 24616 34342 24692 34550
rect 71264 34478 71340 34686
rect 71264 34446 71270 34478
rect 71269 34414 71270 34446
rect 71334 34446 71340 34478
rect 71672 34750 71748 34756
rect 71672 34686 71678 34750
rect 71742 34686 71748 34750
rect 71672 34478 71748 34686
rect 71672 34446 71678 34478
rect 71334 34414 71335 34446
rect 71269 34413 71335 34414
rect 71677 34414 71678 34446
rect 71742 34446 71748 34478
rect 72216 34750 72292 34756
rect 72216 34686 72222 34750
rect 72286 34686 72292 34750
rect 72216 34478 72292 34686
rect 72216 34446 72222 34478
rect 71742 34414 71743 34446
rect 71677 34413 71743 34414
rect 72221 34414 72222 34446
rect 72286 34446 72292 34478
rect 73032 34478 73108 34484
rect 72286 34414 72287 34446
rect 72221 34413 72287 34414
rect 73032 34414 73038 34478
rect 73102 34414 73108 34478
rect 24616 34278 24622 34342
rect 24686 34278 24692 34342
rect 24616 34272 24692 34278
rect 17952 34174 17958 34206
rect 17957 34142 17958 34174
rect 18022 34174 18028 34206
rect 24616 34206 24692 34212
rect 18022 34142 18023 34174
rect 17957 34141 18023 34142
rect 24616 34142 24622 34206
rect 24686 34142 24692 34206
rect 66509 34206 66575 34207
rect 66509 34174 66510 34206
rect 11288 33902 11294 33934
rect 11293 33870 11294 33902
rect 11358 33902 11364 33934
rect 17816 34070 17892 34076
rect 17816 34006 17822 34070
rect 17886 34006 17892 34070
rect 18229 34070 18295 34071
rect 18229 34038 18230 34070
rect 11358 33870 11359 33902
rect 11293 33869 11359 33870
rect 17816 33798 17892 34006
rect 17816 33766 17822 33798
rect 17821 33734 17822 33766
rect 17886 33766 17892 33798
rect 18224 34006 18230 34038
rect 18294 34038 18295 34070
rect 18632 34070 18708 34076
rect 18294 34006 18300 34038
rect 18224 33798 18300 34006
rect 17886 33734 17887 33766
rect 17821 33733 17887 33734
rect 18224 33734 18230 33798
rect 18294 33734 18300 33798
rect 18632 34006 18638 34070
rect 18702 34006 18708 34070
rect 18632 33798 18708 34006
rect 18632 33766 18638 33798
rect 18224 33728 18300 33734
rect 18637 33734 18638 33766
rect 18702 33766 18708 33798
rect 24480 33798 24556 33804
rect 18702 33734 18703 33766
rect 18637 33733 18703 33734
rect 24480 33734 24486 33798
rect 24550 33734 24556 33798
rect 24616 33798 24692 34142
rect 66504 34142 66510 34174
rect 66574 34174 66575 34206
rect 73032 34206 73108 34414
rect 73032 34174 73038 34206
rect 66574 34142 66580 34174
rect 66504 33934 66580 34142
rect 73037 34142 73038 34174
rect 73102 34174 73108 34206
rect 73102 34142 73103 34174
rect 73037 34141 73103 34142
rect 72629 34070 72695 34071
rect 72629 34038 72630 34070
rect 66504 33870 66510 33934
rect 66574 33870 66580 33934
rect 66504 33864 66580 33870
rect 72624 34006 72630 34038
rect 72694 34038 72695 34070
rect 72896 34070 72972 34076
rect 72694 34006 72700 34038
rect 24616 33766 24622 33798
rect 11157 33662 11223 33663
rect 11157 33630 11158 33662
rect 11016 32406 11022 32438
rect 11021 32374 11022 32406
rect 11086 32406 11092 32438
rect 11152 33598 11158 33630
rect 11222 33630 11223 33662
rect 17816 33662 17892 33668
rect 11222 33598 11228 33630
rect 11086 32374 11087 32406
rect 11021 32373 11087 32374
rect 952 32238 1230 32302
rect 1294 32238 1300 32302
rect 11021 32302 11087 32303
rect 11021 32270 11022 32302
rect 952 30806 1300 32238
rect 952 30742 1230 30806
rect 1294 30742 1300 30806
rect 952 28902 1300 30742
rect 11016 32238 11022 32270
rect 11086 32270 11087 32302
rect 11086 32238 11092 32270
rect 11016 29582 11092 32238
rect 11152 31078 11228 33598
rect 17816 33598 17822 33662
rect 17886 33598 17892 33662
rect 18501 33662 18567 33663
rect 18501 33630 18502 33662
rect 17816 33390 17892 33598
rect 17816 33358 17822 33390
rect 17821 33326 17822 33358
rect 17886 33358 17892 33390
rect 18496 33598 18502 33630
rect 18566 33630 18567 33662
rect 19181 33662 19247 33663
rect 19181 33630 19182 33662
rect 18566 33598 18572 33630
rect 18496 33390 18572 33598
rect 17886 33326 17887 33358
rect 17821 33325 17887 33326
rect 18496 33326 18502 33390
rect 18566 33326 18572 33390
rect 18496 33320 18572 33326
rect 19176 33598 19182 33630
rect 19246 33630 19247 33662
rect 19589 33662 19655 33663
rect 19589 33630 19590 33662
rect 19246 33598 19252 33630
rect 19176 33390 19252 33598
rect 19176 33326 19182 33390
rect 19246 33326 19252 33390
rect 19176 33320 19252 33326
rect 19584 33598 19590 33630
rect 19654 33630 19655 33662
rect 19654 33598 19660 33630
rect 19584 33390 19660 33598
rect 24480 33526 24556 33734
rect 24621 33734 24622 33766
rect 24686 33766 24692 33798
rect 66368 33798 66444 33804
rect 24686 33734 24687 33766
rect 24621 33733 24687 33734
rect 66368 33734 66374 33798
rect 66438 33734 66444 33798
rect 24480 33494 24486 33526
rect 24485 33462 24486 33494
rect 24550 33494 24556 33526
rect 66368 33526 66444 33734
rect 72624 33798 72700 34006
rect 72624 33734 72630 33798
rect 72694 33734 72700 33798
rect 72896 34006 72902 34070
rect 72966 34006 72972 34070
rect 72896 33798 72972 34006
rect 72896 33766 72902 33798
rect 72624 33728 72700 33734
rect 72901 33734 72902 33766
rect 72966 33766 72972 33798
rect 89760 34070 90108 35638
rect 89760 34006 89766 34070
rect 89830 34006 90108 34070
rect 72966 33734 72967 33766
rect 72901 33733 72967 33734
rect 71405 33662 71471 33663
rect 71405 33630 71406 33662
rect 66368 33494 66374 33526
rect 24550 33462 24551 33494
rect 24485 33461 24551 33462
rect 66373 33462 66374 33494
rect 66438 33494 66444 33526
rect 71400 33598 71406 33630
rect 71470 33630 71471 33662
rect 71813 33662 71879 33663
rect 71813 33630 71814 33662
rect 71470 33598 71476 33630
rect 66438 33462 66439 33494
rect 66373 33461 66439 33462
rect 19584 33326 19590 33390
rect 19654 33326 19660 33390
rect 19584 33320 19660 33326
rect 71400 33390 71476 33598
rect 71400 33326 71406 33390
rect 71470 33326 71476 33390
rect 71400 33320 71476 33326
rect 71808 33598 71814 33630
rect 71878 33630 71879 33662
rect 72901 33662 72967 33663
rect 72901 33630 72902 33662
rect 71878 33598 71884 33630
rect 71808 33390 71884 33598
rect 72896 33598 72902 33630
rect 72966 33630 72967 33662
rect 72966 33598 72972 33630
rect 71808 33326 71814 33390
rect 71878 33326 71884 33390
rect 71808 33320 71884 33326
rect 72352 33526 72428 33532
rect 72352 33462 72358 33526
rect 72422 33462 72428 33526
rect 17952 33254 18028 33260
rect 17952 33190 17958 33254
rect 18022 33190 18028 33254
rect 17952 32982 18028 33190
rect 17952 32950 17958 32982
rect 17957 32918 17958 32950
rect 18022 32950 18028 32982
rect 18632 33254 18708 33260
rect 18632 33190 18638 33254
rect 18702 33190 18708 33254
rect 19045 33254 19111 33255
rect 19045 33222 19046 33254
rect 18632 32982 18708 33190
rect 18632 32950 18638 32982
rect 18022 32918 18023 32950
rect 17957 32917 18023 32918
rect 18637 32918 18638 32950
rect 18702 32950 18708 32982
rect 19040 33190 19046 33222
rect 19110 33222 19111 33254
rect 19584 33254 19660 33260
rect 19110 33190 19116 33222
rect 19040 32982 19116 33190
rect 18702 32918 18703 32950
rect 18637 32917 18703 32918
rect 19040 32918 19046 32982
rect 19110 32918 19116 32982
rect 19584 33190 19590 33254
rect 19654 33190 19660 33254
rect 19584 32982 19660 33190
rect 71264 33254 71340 33260
rect 71264 33190 71270 33254
rect 71334 33190 71340 33254
rect 19584 32950 19590 32982
rect 19040 32912 19116 32918
rect 19589 32918 19590 32950
rect 19654 32950 19660 32982
rect 66368 32982 66444 32988
rect 19654 32918 19655 32950
rect 19589 32917 19655 32918
rect 66368 32918 66374 32982
rect 66438 32918 66444 32982
rect 71264 32982 71340 33190
rect 71264 32950 71270 32982
rect 17821 32846 17887 32847
rect 17821 32814 17822 32846
rect 17816 32782 17822 32814
rect 17886 32814 17887 32846
rect 18365 32846 18431 32847
rect 18365 32814 18366 32846
rect 17886 32782 17892 32814
rect 17816 32574 17892 32782
rect 17816 32510 17822 32574
rect 17886 32510 17892 32574
rect 17816 32504 17892 32510
rect 18360 32782 18366 32814
rect 18430 32814 18431 32846
rect 19176 32846 19252 32852
rect 18430 32782 18436 32814
rect 18360 32574 18436 32782
rect 18360 32510 18366 32574
rect 18430 32510 18436 32574
rect 19176 32782 19182 32846
rect 19246 32782 19252 32846
rect 19453 32846 19519 32847
rect 19453 32814 19454 32846
rect 19176 32574 19252 32782
rect 19176 32542 19182 32574
rect 18360 32504 18436 32510
rect 19181 32510 19182 32542
rect 19246 32542 19252 32574
rect 19448 32782 19454 32814
rect 19518 32814 19519 32846
rect 19518 32782 19524 32814
rect 19448 32574 19524 32782
rect 66368 32710 66444 32918
rect 71269 32918 71270 32950
rect 71334 32950 71340 32982
rect 71808 33254 71884 33260
rect 71808 33190 71814 33254
rect 71878 33190 71884 33254
rect 72352 33254 72428 33462
rect 72896 33390 72972 33598
rect 72896 33326 72902 33390
rect 72966 33326 72972 33390
rect 72896 33320 72972 33326
rect 72352 33222 72358 33254
rect 71808 32982 71884 33190
rect 72357 33190 72358 33222
rect 72422 33222 72428 33254
rect 72629 33254 72695 33255
rect 72629 33222 72630 33254
rect 72422 33190 72423 33222
rect 72357 33189 72423 33190
rect 72624 33190 72630 33222
rect 72694 33222 72695 33254
rect 73032 33254 73108 33260
rect 72694 33190 72700 33222
rect 71808 32950 71814 32982
rect 71334 32918 71335 32950
rect 71269 32917 71335 32918
rect 71813 32918 71814 32950
rect 71878 32950 71884 32982
rect 72624 32982 72700 33190
rect 71878 32918 71879 32950
rect 71813 32917 71879 32918
rect 72624 32918 72630 32982
rect 72694 32918 72700 32982
rect 73032 33190 73038 33254
rect 73102 33190 73108 33254
rect 73032 32982 73108 33190
rect 73032 32950 73038 32982
rect 72624 32912 72700 32918
rect 73037 32918 73038 32950
rect 73102 32950 73108 32982
rect 73102 32918 73103 32950
rect 73037 32917 73103 32918
rect 66368 32678 66374 32710
rect 66373 32646 66374 32678
rect 66438 32678 66444 32710
rect 71400 32846 71476 32852
rect 71400 32782 71406 32846
rect 71470 32782 71476 32846
rect 71677 32846 71743 32847
rect 71677 32814 71678 32846
rect 66438 32646 66439 32678
rect 66373 32645 66439 32646
rect 19246 32510 19247 32542
rect 19181 32509 19247 32510
rect 19448 32510 19454 32574
rect 19518 32510 19524 32574
rect 71400 32574 71476 32782
rect 71400 32542 71406 32574
rect 19448 32504 19524 32510
rect 71405 32510 71406 32542
rect 71470 32542 71476 32574
rect 71672 32782 71678 32814
rect 71742 32814 71743 32846
rect 72357 32846 72423 32847
rect 72357 32814 72358 32846
rect 71742 32782 71748 32814
rect 71672 32574 71748 32782
rect 71470 32510 71471 32542
rect 71405 32509 71471 32510
rect 71672 32510 71678 32574
rect 71742 32510 71748 32574
rect 71672 32504 71748 32510
rect 72352 32782 72358 32814
rect 72422 32814 72423 32846
rect 72901 32846 72967 32847
rect 72901 32814 72902 32846
rect 72422 32782 72428 32814
rect 72352 32574 72428 32782
rect 72352 32510 72358 32574
rect 72422 32510 72428 32574
rect 72352 32504 72428 32510
rect 72896 32782 72902 32814
rect 72966 32814 72967 32846
rect 72966 32782 72972 32814
rect 72896 32574 72972 32782
rect 72896 32510 72902 32574
rect 72966 32510 72972 32574
rect 72896 32504 72972 32510
rect 17957 32438 18023 32439
rect 17957 32406 17958 32438
rect 17952 32374 17958 32406
rect 18022 32406 18023 32438
rect 18365 32438 18431 32439
rect 18365 32406 18366 32438
rect 18022 32374 18028 32406
rect 17952 32166 18028 32374
rect 17952 32102 17958 32166
rect 18022 32102 18028 32166
rect 17952 32096 18028 32102
rect 18360 32374 18366 32406
rect 18430 32406 18431 32438
rect 18773 32438 18839 32439
rect 18773 32406 18774 32438
rect 18430 32374 18436 32406
rect 18360 32166 18436 32374
rect 18360 32102 18366 32166
rect 18430 32102 18436 32166
rect 18360 32096 18436 32102
rect 18768 32374 18774 32406
rect 18838 32406 18839 32438
rect 19181 32438 19247 32439
rect 19181 32406 19182 32438
rect 18838 32374 18844 32406
rect 18768 32166 18844 32374
rect 18768 32102 18774 32166
rect 18838 32102 18844 32166
rect 18768 32096 18844 32102
rect 19176 32374 19182 32406
rect 19246 32406 19247 32438
rect 19589 32438 19655 32439
rect 19589 32406 19590 32438
rect 19246 32374 19252 32406
rect 19176 32166 19252 32374
rect 19176 32102 19182 32166
rect 19246 32102 19252 32166
rect 19176 32096 19252 32102
rect 19584 32374 19590 32406
rect 19654 32406 19655 32438
rect 71405 32438 71471 32439
rect 71405 32406 71406 32438
rect 19654 32374 19660 32406
rect 19584 32166 19660 32374
rect 19584 32102 19590 32166
rect 19654 32102 19660 32166
rect 19584 32096 19660 32102
rect 71400 32374 71406 32406
rect 71470 32406 71471 32438
rect 71808 32438 71884 32444
rect 71470 32374 71476 32406
rect 71400 32166 71476 32374
rect 71400 32102 71406 32166
rect 71470 32102 71476 32166
rect 71808 32374 71814 32438
rect 71878 32374 71884 32438
rect 72085 32438 72151 32439
rect 72085 32406 72086 32438
rect 71808 32166 71884 32374
rect 71808 32134 71814 32166
rect 71400 32096 71476 32102
rect 71813 32102 71814 32134
rect 71878 32134 71884 32166
rect 72080 32374 72086 32406
rect 72150 32406 72151 32438
rect 72624 32438 72700 32444
rect 72150 32374 72156 32406
rect 72080 32166 72156 32374
rect 71878 32102 71879 32134
rect 71813 32101 71879 32102
rect 72080 32102 72086 32166
rect 72150 32102 72156 32166
rect 72624 32374 72630 32438
rect 72694 32374 72700 32438
rect 72624 32166 72700 32374
rect 72624 32134 72630 32166
rect 72080 32096 72156 32102
rect 72629 32102 72630 32134
rect 72694 32134 72700 32166
rect 73032 32438 73108 32444
rect 73032 32374 73038 32438
rect 73102 32374 73108 32438
rect 73032 32166 73108 32374
rect 73032 32134 73038 32166
rect 72694 32102 72695 32134
rect 72629 32101 72695 32102
rect 73037 32102 73038 32134
rect 73102 32134 73108 32166
rect 89760 32438 90108 34006
rect 89760 32374 89766 32438
rect 89830 32374 90108 32438
rect 73102 32102 73103 32134
rect 73037 32101 73103 32102
rect 17957 32030 18023 32031
rect 17957 31998 17958 32030
rect 17952 31966 17958 31998
rect 18022 31998 18023 32030
rect 18496 32030 18572 32036
rect 18022 31966 18028 31998
rect 17952 31758 18028 31966
rect 17952 31694 17958 31758
rect 18022 31694 18028 31758
rect 18496 31966 18502 32030
rect 18566 31966 18572 32030
rect 19045 32030 19111 32031
rect 19045 31998 19046 32030
rect 18496 31758 18572 31966
rect 18496 31726 18502 31758
rect 17952 31688 18028 31694
rect 18501 31694 18502 31726
rect 18566 31726 18572 31758
rect 19040 31966 19046 31998
rect 19110 31998 19111 32030
rect 19448 32030 19524 32036
rect 19110 31966 19116 31998
rect 19040 31758 19116 31966
rect 18566 31694 18567 31726
rect 18501 31693 18567 31694
rect 19040 31694 19046 31758
rect 19110 31694 19116 31758
rect 19448 31966 19454 32030
rect 19518 31966 19524 32030
rect 19448 31758 19524 31966
rect 19448 31726 19454 31758
rect 19040 31688 19116 31694
rect 19453 31694 19454 31726
rect 19518 31726 19524 31758
rect 71400 32030 71476 32036
rect 71400 31966 71406 32030
rect 71470 31966 71476 32030
rect 71677 32030 71743 32031
rect 71677 31998 71678 32030
rect 71400 31758 71476 31966
rect 71400 31726 71406 31758
rect 19518 31694 19519 31726
rect 19453 31693 19519 31694
rect 71405 31694 71406 31726
rect 71470 31726 71476 31758
rect 71672 31966 71678 31998
rect 71742 31998 71743 32030
rect 72488 32030 72564 32036
rect 71742 31966 71748 31998
rect 71672 31758 71748 31966
rect 71470 31694 71471 31726
rect 71405 31693 71471 31694
rect 71672 31694 71678 31758
rect 71742 31694 71748 31758
rect 72488 31966 72494 32030
rect 72558 31966 72564 32030
rect 73037 32030 73103 32031
rect 73037 31998 73038 32030
rect 72488 31758 72564 31966
rect 72488 31726 72494 31758
rect 71672 31688 71748 31694
rect 72493 31694 72494 31726
rect 72558 31726 72564 31758
rect 73032 31966 73038 31998
rect 73102 31998 73103 32030
rect 73102 31966 73108 31998
rect 73032 31758 73108 31966
rect 72558 31694 72559 31726
rect 72493 31693 72559 31694
rect 73032 31694 73038 31758
rect 73102 31694 73108 31758
rect 73032 31688 73108 31694
rect 18360 31622 18436 31628
rect 18360 31558 18366 31622
rect 18430 31558 18436 31622
rect 18360 31350 18436 31558
rect 18360 31318 18366 31350
rect 18365 31286 18366 31318
rect 18430 31318 18436 31350
rect 19176 31622 19252 31628
rect 19176 31558 19182 31622
rect 19246 31558 19252 31622
rect 19453 31622 19519 31623
rect 19453 31590 19454 31622
rect 19176 31350 19252 31558
rect 19176 31318 19182 31350
rect 18430 31286 18431 31318
rect 18365 31285 18431 31286
rect 19181 31286 19182 31318
rect 19246 31318 19252 31350
rect 19448 31558 19454 31590
rect 19518 31590 19519 31622
rect 71400 31622 71476 31628
rect 19518 31558 19524 31590
rect 19448 31350 19524 31558
rect 71400 31558 71406 31622
rect 71470 31558 71476 31622
rect 71677 31622 71743 31623
rect 71677 31590 71678 31622
rect 19246 31286 19247 31318
rect 19181 31285 19247 31286
rect 19448 31286 19454 31350
rect 19518 31286 19524 31350
rect 19448 31280 19524 31286
rect 24480 31486 24556 31492
rect 24480 31422 24486 31486
rect 24550 31422 24556 31486
rect 19045 31214 19111 31215
rect 19045 31182 19046 31214
rect 11152 31014 11158 31078
rect 11222 31014 11228 31078
rect 11152 31008 11228 31014
rect 19040 31150 19046 31182
rect 19110 31182 19111 31214
rect 19453 31214 19519 31215
rect 19453 31182 19454 31214
rect 19110 31150 19116 31182
rect 11016 29518 11022 29582
rect 11086 29518 11092 29582
rect 11016 29512 11092 29518
rect 11152 30942 11228 30948
rect 11152 30878 11158 30942
rect 11222 30878 11228 30942
rect 952 28838 1230 28902
rect 1294 28838 1300 28902
rect 952 27270 1300 28838
rect 11152 28222 11228 30878
rect 19040 30942 19116 31150
rect 19040 30878 19046 30942
rect 19110 30878 19116 30942
rect 19040 30872 19116 30878
rect 19448 31150 19454 31182
rect 19518 31182 19519 31214
rect 24480 31214 24556 31422
rect 71400 31350 71476 31558
rect 71400 31318 71406 31350
rect 71405 31286 71406 31318
rect 71470 31318 71476 31350
rect 71672 31558 71678 31590
rect 71742 31590 71743 31622
rect 72085 31622 72151 31623
rect 72085 31590 72086 31622
rect 71742 31558 71748 31590
rect 71672 31350 71748 31558
rect 71470 31286 71471 31318
rect 71405 31285 71471 31286
rect 71672 31286 71678 31350
rect 71742 31286 71748 31350
rect 71672 31280 71748 31286
rect 72080 31558 72086 31590
rect 72150 31590 72151 31622
rect 72150 31558 72156 31590
rect 72080 31350 72156 31558
rect 72080 31286 72086 31350
rect 72150 31286 72156 31350
rect 72080 31280 72156 31286
rect 24480 31182 24486 31214
rect 19518 31150 19524 31182
rect 19448 30942 19524 31150
rect 24485 31150 24486 31182
rect 24550 31182 24556 31214
rect 71269 31214 71335 31215
rect 71269 31182 71270 31214
rect 24550 31150 24551 31182
rect 24485 31149 24551 31150
rect 71264 31150 71270 31182
rect 71334 31182 71335 31214
rect 71808 31214 71884 31220
rect 71334 31150 71340 31182
rect 19448 30878 19454 30942
rect 19518 30878 19524 30942
rect 19448 30872 19524 30878
rect 71264 30942 71340 31150
rect 71264 30878 71270 30942
rect 71334 30878 71340 30942
rect 71808 31150 71814 31214
rect 71878 31150 71884 31214
rect 71808 30942 71884 31150
rect 71808 30910 71814 30942
rect 71264 30872 71340 30878
rect 71813 30878 71814 30910
rect 71878 30910 71884 30942
rect 71878 30878 71879 30910
rect 71813 30877 71879 30878
rect 18496 30806 18572 30812
rect 18496 30742 18502 30806
rect 18566 30742 18572 30806
rect 17821 30534 17887 30535
rect 17821 30502 17822 30534
rect 17816 30470 17822 30502
rect 17886 30502 17887 30534
rect 18496 30534 18572 30742
rect 18496 30502 18502 30534
rect 17886 30470 17892 30502
rect 17816 30262 17892 30470
rect 18501 30470 18502 30502
rect 18566 30502 18572 30534
rect 19176 30806 19252 30812
rect 19176 30742 19182 30806
rect 19246 30742 19252 30806
rect 19589 30806 19655 30807
rect 19589 30774 19590 30806
rect 19176 30534 19252 30742
rect 19176 30502 19182 30534
rect 18566 30470 18567 30502
rect 18501 30469 18567 30470
rect 19181 30470 19182 30502
rect 19246 30502 19252 30534
rect 19584 30742 19590 30774
rect 19654 30774 19655 30806
rect 71400 30806 71476 30812
rect 19654 30742 19660 30774
rect 19584 30534 19660 30742
rect 71400 30742 71406 30806
rect 71470 30742 71476 30806
rect 71813 30806 71879 30807
rect 71813 30774 71814 30806
rect 24621 30670 24687 30671
rect 24621 30638 24622 30670
rect 19246 30470 19247 30502
rect 19181 30469 19247 30470
rect 19584 30470 19590 30534
rect 19654 30470 19660 30534
rect 19584 30464 19660 30470
rect 24616 30606 24622 30638
rect 24686 30638 24687 30670
rect 24686 30606 24692 30638
rect 24616 30398 24692 30606
rect 71400 30534 71476 30742
rect 71400 30502 71406 30534
rect 71405 30470 71406 30502
rect 71470 30502 71476 30534
rect 71808 30742 71814 30774
rect 71878 30774 71879 30806
rect 72080 30806 72156 30812
rect 71878 30742 71884 30774
rect 71808 30534 71884 30742
rect 71470 30470 71471 30502
rect 71405 30469 71471 30470
rect 71808 30470 71814 30534
rect 71878 30470 71884 30534
rect 72080 30742 72086 30806
rect 72150 30742 72156 30806
rect 72080 30534 72156 30742
rect 89760 30670 90108 32374
rect 89760 30606 89766 30670
rect 89830 30606 90108 30670
rect 72080 30502 72086 30534
rect 71808 30464 71884 30470
rect 72085 30470 72086 30502
rect 72150 30502 72156 30534
rect 72896 30534 72972 30540
rect 72150 30470 72151 30502
rect 72085 30469 72151 30470
rect 72896 30470 72902 30534
rect 72966 30470 72972 30534
rect 24616 30334 24622 30398
rect 24686 30334 24692 30398
rect 24616 30328 24692 30334
rect 17816 30198 17822 30262
rect 17886 30198 17892 30262
rect 17816 30192 17892 30198
rect 24480 30262 24556 30268
rect 24480 30198 24486 30262
rect 24550 30198 24556 30262
rect 66373 30262 66439 30263
rect 66373 30230 66374 30262
rect 17821 30126 17887 30127
rect 17821 30094 17822 30126
rect 17816 30062 17822 30094
rect 17886 30094 17887 30126
rect 18632 30126 18708 30132
rect 17886 30062 17892 30094
rect 17816 29854 17892 30062
rect 17816 29790 17822 29854
rect 17886 29790 17892 29854
rect 18632 30062 18638 30126
rect 18702 30062 18708 30126
rect 18632 29854 18708 30062
rect 24480 29990 24556 30198
rect 24480 29958 24486 29990
rect 24485 29926 24486 29958
rect 24550 29958 24556 29990
rect 66368 30198 66374 30230
rect 66438 30230 66439 30262
rect 72896 30262 72972 30470
rect 72896 30230 72902 30262
rect 66438 30198 66444 30230
rect 66368 29990 66444 30198
rect 72901 30198 72902 30230
rect 72966 30230 72972 30262
rect 72966 30198 72967 30230
rect 72901 30197 72967 30198
rect 72221 30126 72287 30127
rect 72221 30094 72222 30126
rect 24550 29926 24551 29958
rect 24485 29925 24551 29926
rect 66368 29926 66374 29990
rect 66438 29926 66444 29990
rect 66368 29920 66444 29926
rect 72216 30062 72222 30094
rect 72286 30094 72287 30126
rect 72629 30126 72695 30127
rect 72629 30094 72630 30126
rect 72286 30062 72292 30094
rect 18632 29822 18638 29854
rect 17816 29784 17892 29790
rect 18637 29790 18638 29822
rect 18702 29822 18708 29854
rect 66509 29854 66575 29855
rect 66509 29822 66510 29854
rect 18702 29790 18703 29822
rect 18637 29789 18703 29790
rect 66504 29790 66510 29822
rect 66574 29822 66575 29854
rect 72216 29854 72292 30062
rect 66574 29790 66580 29822
rect 17816 29718 17892 29724
rect 17816 29654 17822 29718
rect 17886 29654 17892 29718
rect 14829 29446 14895 29447
rect 14829 29414 14830 29446
rect 11152 28190 11158 28222
rect 11157 28158 11158 28190
rect 11222 28190 11228 28222
rect 14824 29382 14830 29414
rect 14894 29414 14895 29446
rect 17816 29446 17892 29654
rect 66504 29582 66580 29790
rect 72216 29790 72222 29854
rect 72286 29790 72292 29854
rect 72216 29784 72292 29790
rect 72624 30062 72630 30094
rect 72694 30094 72695 30126
rect 73037 30126 73103 30127
rect 73037 30094 73038 30126
rect 72694 30062 72700 30094
rect 72624 29854 72700 30062
rect 72624 29790 72630 29854
rect 72694 29790 72700 29854
rect 72624 29784 72700 29790
rect 73032 30062 73038 30094
rect 73102 30094 73103 30126
rect 73102 30062 73108 30094
rect 73032 29854 73108 30062
rect 73032 29790 73038 29854
rect 73102 29790 73108 29854
rect 73032 29784 73108 29790
rect 73037 29718 73103 29719
rect 73037 29686 73038 29718
rect 66504 29518 66510 29582
rect 66574 29518 66580 29582
rect 66504 29512 66580 29518
rect 73032 29654 73038 29686
rect 73102 29686 73103 29718
rect 73102 29654 73108 29686
rect 17816 29414 17822 29446
rect 14894 29382 14900 29414
rect 11222 28158 11223 28190
rect 11157 28157 11223 28158
rect 12925 28086 12991 28087
rect 12925 28054 12926 28086
rect 952 27206 1230 27270
rect 1294 27206 1300 27270
rect 952 25638 1300 27206
rect 12920 28022 12926 28054
rect 12990 28054 12991 28086
rect 12990 28022 12996 28054
rect 2460 25732 2526 25733
rect 2460 25668 2461 25732
rect 2525 25668 2526 25732
rect 2460 25667 2526 25668
rect 952 25574 1230 25638
rect 1294 25574 1300 25638
rect 2181 25638 2247 25639
rect 2181 25606 2182 25638
rect 952 23870 1300 25574
rect 2176 25574 2182 25606
rect 2246 25606 2247 25638
rect 2246 25574 2252 25606
rect 2176 25094 2252 25574
rect 2176 25030 2182 25094
rect 2246 25030 2252 25094
rect 2176 25024 2252 25030
rect 952 23806 1230 23870
rect 1294 23806 1300 23870
rect 952 22238 1300 23806
rect 952 22174 1230 22238
rect 1294 22174 1300 22238
rect 952 20470 1300 22174
rect 952 20406 1230 20470
rect 1294 20406 1300 20470
rect 952 18838 1300 20406
rect 952 18774 1230 18838
rect 1294 18774 1300 18838
rect 952 17206 1300 18774
rect 2463 18326 2523 25667
rect 12920 25502 12996 28022
rect 14824 27814 14900 29382
rect 17821 29382 17822 29414
rect 17886 29414 17892 29446
rect 73032 29446 73108 29654
rect 17886 29382 17887 29414
rect 17821 29381 17887 29382
rect 73032 29382 73038 29446
rect 73102 29382 73108 29446
rect 73032 29376 73108 29382
rect 17821 29310 17887 29311
rect 17821 29278 17822 29310
rect 17816 29246 17822 29278
rect 17886 29278 17887 29310
rect 18768 29310 18844 29316
rect 17886 29246 17892 29278
rect 17816 29038 17892 29246
rect 17816 28974 17822 29038
rect 17886 28974 17892 29038
rect 18768 29246 18774 29310
rect 18838 29246 18844 29310
rect 18768 29038 18844 29246
rect 18768 29006 18774 29038
rect 17816 28968 17892 28974
rect 18773 28974 18774 29006
rect 18838 29006 18844 29038
rect 19040 29310 19116 29316
rect 19040 29246 19046 29310
rect 19110 29246 19116 29310
rect 19453 29310 19519 29311
rect 19453 29278 19454 29310
rect 19040 29038 19116 29246
rect 19040 29006 19046 29038
rect 18838 28974 18839 29006
rect 18773 28973 18839 28974
rect 19045 28974 19046 29006
rect 19110 29006 19116 29038
rect 19448 29246 19454 29278
rect 19518 29278 19519 29310
rect 71405 29310 71471 29311
rect 71405 29278 71406 29310
rect 19518 29246 19524 29278
rect 19448 29038 19524 29246
rect 71400 29246 71406 29278
rect 71470 29278 71471 29310
rect 71813 29310 71879 29311
rect 71813 29278 71814 29310
rect 71470 29246 71476 29278
rect 19110 28974 19111 29006
rect 19045 28973 19111 28974
rect 19448 28974 19454 29038
rect 19518 28974 19524 29038
rect 19448 28968 19524 28974
rect 66504 29038 66580 29044
rect 66504 28974 66510 29038
rect 66574 28974 66580 29038
rect 17821 28902 17887 28903
rect 17821 28870 17822 28902
rect 17816 28838 17822 28870
rect 17886 28870 17887 28902
rect 18224 28902 18300 28908
rect 17886 28838 17892 28870
rect 17816 28630 17892 28838
rect 17816 28566 17822 28630
rect 17886 28566 17892 28630
rect 18224 28838 18230 28902
rect 18294 28838 18300 28902
rect 18224 28630 18300 28838
rect 18224 28598 18230 28630
rect 17816 28560 17892 28566
rect 18229 28566 18230 28598
rect 18294 28598 18300 28630
rect 18496 28902 18572 28908
rect 18496 28838 18502 28902
rect 18566 28838 18572 28902
rect 19045 28902 19111 28903
rect 19045 28870 19046 28902
rect 18496 28630 18572 28838
rect 18496 28598 18502 28630
rect 18294 28566 18295 28598
rect 18229 28565 18295 28566
rect 18501 28566 18502 28598
rect 18566 28598 18572 28630
rect 19040 28838 19046 28870
rect 19110 28870 19111 28902
rect 19584 28902 19660 28908
rect 19110 28838 19116 28870
rect 19040 28630 19116 28838
rect 18566 28566 18567 28598
rect 18501 28565 18567 28566
rect 19040 28566 19046 28630
rect 19110 28566 19116 28630
rect 19584 28838 19590 28902
rect 19654 28838 19660 28902
rect 19584 28630 19660 28838
rect 66504 28766 66580 28974
rect 71400 29038 71476 29246
rect 71400 28974 71406 29038
rect 71470 28974 71476 29038
rect 71400 28968 71476 28974
rect 71808 29246 71814 29278
rect 71878 29278 71879 29310
rect 73032 29310 73108 29316
rect 71878 29246 71884 29278
rect 71808 29038 71884 29246
rect 71808 28974 71814 29038
rect 71878 28974 71884 29038
rect 73032 29246 73038 29310
rect 73102 29246 73108 29310
rect 73032 29038 73108 29246
rect 73032 29006 73038 29038
rect 71808 28968 71884 28974
rect 73037 28974 73038 29006
rect 73102 29006 73108 29038
rect 89760 29038 90108 30606
rect 73102 28974 73103 29006
rect 73037 28973 73103 28974
rect 89760 28974 89766 29038
rect 89830 28974 90108 29038
rect 66504 28734 66510 28766
rect 66509 28702 66510 28734
rect 66574 28734 66580 28766
rect 71264 28902 71340 28908
rect 71264 28838 71270 28902
rect 71334 28838 71340 28902
rect 66574 28702 66575 28734
rect 66509 28701 66575 28702
rect 19584 28598 19590 28630
rect 19040 28560 19116 28566
rect 19589 28566 19590 28598
rect 19654 28598 19660 28630
rect 71264 28630 71340 28838
rect 71264 28598 71270 28630
rect 19654 28566 19655 28598
rect 19589 28565 19655 28566
rect 71269 28566 71270 28598
rect 71334 28598 71340 28630
rect 71808 28902 71884 28908
rect 71808 28838 71814 28902
rect 71878 28838 71884 28902
rect 71808 28630 71884 28838
rect 71808 28598 71814 28630
rect 71334 28566 71335 28598
rect 71269 28565 71335 28566
rect 71813 28566 71814 28598
rect 71878 28598 71884 28630
rect 72488 28902 72564 28908
rect 72488 28838 72494 28902
rect 72558 28838 72564 28902
rect 72488 28630 72564 28838
rect 72488 28598 72494 28630
rect 71878 28566 71879 28598
rect 71813 28565 71879 28566
rect 72493 28566 72494 28598
rect 72558 28598 72564 28630
rect 73032 28902 73108 28908
rect 73032 28838 73038 28902
rect 73102 28838 73108 28902
rect 73032 28630 73108 28838
rect 73032 28598 73038 28630
rect 72558 28566 72559 28598
rect 72493 28565 72559 28566
rect 73037 28566 73038 28598
rect 73102 28598 73108 28630
rect 73102 28566 73103 28598
rect 73037 28565 73103 28566
rect 17821 28494 17887 28495
rect 17821 28462 17822 28494
rect 17816 28430 17822 28462
rect 17886 28462 17887 28494
rect 18365 28494 18431 28495
rect 18365 28462 18366 28494
rect 17886 28430 17892 28462
rect 17816 28222 17892 28430
rect 17816 28158 17822 28222
rect 17886 28158 17892 28222
rect 17816 28152 17892 28158
rect 18360 28430 18366 28462
rect 18430 28462 18431 28494
rect 19176 28494 19252 28500
rect 18430 28430 18436 28462
rect 18360 28222 18436 28430
rect 18360 28158 18366 28222
rect 18430 28158 18436 28222
rect 19176 28430 19182 28494
rect 19246 28430 19252 28494
rect 19176 28222 19252 28430
rect 19176 28190 19182 28222
rect 18360 28152 18436 28158
rect 19181 28158 19182 28190
rect 19246 28190 19252 28222
rect 19584 28494 19660 28500
rect 19584 28430 19590 28494
rect 19654 28430 19660 28494
rect 71405 28494 71471 28495
rect 71405 28462 71406 28494
rect 19584 28222 19660 28430
rect 19584 28190 19590 28222
rect 19246 28158 19247 28190
rect 19181 28157 19247 28158
rect 19589 28158 19590 28190
rect 19654 28190 19660 28222
rect 71400 28430 71406 28462
rect 71470 28462 71471 28494
rect 71677 28494 71743 28495
rect 71677 28462 71678 28494
rect 71470 28430 71476 28462
rect 71400 28222 71476 28430
rect 19654 28158 19655 28190
rect 19589 28157 19655 28158
rect 71400 28158 71406 28222
rect 71470 28158 71476 28222
rect 71400 28152 71476 28158
rect 71672 28430 71678 28462
rect 71742 28462 71743 28494
rect 72085 28494 72151 28495
rect 72085 28462 72086 28494
rect 71742 28430 71748 28462
rect 71672 28222 71748 28430
rect 71672 28158 71678 28222
rect 71742 28158 71748 28222
rect 71672 28152 71748 28158
rect 72080 28430 72086 28462
rect 72150 28462 72151 28494
rect 72488 28494 72564 28500
rect 72150 28430 72156 28462
rect 72080 28222 72156 28430
rect 72080 28158 72086 28222
rect 72150 28158 72156 28222
rect 72488 28430 72494 28494
rect 72558 28430 72564 28494
rect 72901 28494 72967 28495
rect 72901 28462 72902 28494
rect 72488 28222 72564 28430
rect 72488 28190 72494 28222
rect 72080 28152 72156 28158
rect 72493 28158 72494 28190
rect 72558 28190 72564 28222
rect 72896 28430 72902 28462
rect 72966 28462 72967 28494
rect 72966 28430 72972 28462
rect 72896 28222 72972 28430
rect 72558 28158 72559 28190
rect 72493 28157 72559 28158
rect 72896 28158 72902 28222
rect 72966 28158 72972 28222
rect 72896 28152 72972 28158
rect 14824 27750 14830 27814
rect 14894 27750 14900 27814
rect 17816 28086 17892 28092
rect 17816 28022 17822 28086
rect 17886 28022 17892 28086
rect 17816 27814 17892 28022
rect 17816 27782 17822 27814
rect 14824 27744 14900 27750
rect 17821 27750 17822 27782
rect 17886 27782 17892 27814
rect 18224 28086 18300 28092
rect 18224 28022 18230 28086
rect 18294 28022 18300 28086
rect 18773 28086 18839 28087
rect 18773 28054 18774 28086
rect 18224 27814 18300 28022
rect 18224 27782 18230 27814
rect 17886 27750 17887 27782
rect 17821 27749 17887 27750
rect 18229 27750 18230 27782
rect 18294 27782 18300 27814
rect 18768 28022 18774 28054
rect 18838 28054 18839 28086
rect 19040 28086 19116 28092
rect 18838 28022 18844 28054
rect 18768 27814 18844 28022
rect 18294 27750 18295 27782
rect 18229 27749 18295 27750
rect 18768 27750 18774 27814
rect 18838 27750 18844 27814
rect 19040 28022 19046 28086
rect 19110 28022 19116 28086
rect 19589 28086 19655 28087
rect 19589 28054 19590 28086
rect 19040 27814 19116 28022
rect 19040 27782 19046 27814
rect 18768 27744 18844 27750
rect 19045 27750 19046 27782
rect 19110 27782 19116 27814
rect 19584 28022 19590 28054
rect 19654 28054 19655 28086
rect 71264 28086 71340 28092
rect 19654 28022 19660 28054
rect 19584 27814 19660 28022
rect 19110 27750 19111 27782
rect 19045 27749 19111 27750
rect 19584 27750 19590 27814
rect 19654 27750 19660 27814
rect 71264 28022 71270 28086
rect 71334 28022 71340 28086
rect 71264 27814 71340 28022
rect 71264 27782 71270 27814
rect 19584 27744 19660 27750
rect 71269 27750 71270 27782
rect 71334 27782 71340 27814
rect 71672 28086 71748 28092
rect 71672 28022 71678 28086
rect 71742 28022 71748 28086
rect 71672 27814 71748 28022
rect 71672 27782 71678 27814
rect 71334 27750 71335 27782
rect 71269 27749 71335 27750
rect 71677 27750 71678 27782
rect 71742 27782 71748 27814
rect 72216 28086 72292 28092
rect 72216 28022 72222 28086
rect 72286 28022 72292 28086
rect 72901 28086 72967 28087
rect 72901 28054 72902 28086
rect 72216 27814 72292 28022
rect 72216 27782 72222 27814
rect 71742 27750 71743 27782
rect 71677 27749 71743 27750
rect 72221 27750 72222 27782
rect 72286 27782 72292 27814
rect 72896 28022 72902 28054
rect 72966 28054 72967 28086
rect 72966 28022 72972 28054
rect 72896 27814 72972 28022
rect 72286 27750 72287 27782
rect 72221 27749 72287 27750
rect 72896 27750 72902 27814
rect 72966 27750 72972 27814
rect 72896 27744 72972 27750
rect 14557 27678 14623 27679
rect 14557 27646 14558 27678
rect 14552 27614 14558 27646
rect 14622 27646 14623 27678
rect 15373 27678 15439 27679
rect 15373 27646 15374 27678
rect 14622 27614 14628 27646
rect 14552 26998 14628 27614
rect 14552 26934 14558 26998
rect 14622 26934 14628 26998
rect 14552 26928 14628 26934
rect 15368 27614 15374 27646
rect 15438 27646 15439 27678
rect 15776 27678 15852 27684
rect 15438 27614 15444 27646
rect 15368 26998 15444 27614
rect 15368 26934 15374 26998
rect 15438 26934 15444 26998
rect 15776 27614 15782 27678
rect 15846 27614 15852 27678
rect 15776 26998 15852 27614
rect 18496 27678 18572 27684
rect 18496 27614 18502 27678
rect 18566 27614 18572 27678
rect 18496 27406 18572 27614
rect 18496 27374 18502 27406
rect 18501 27342 18502 27374
rect 18566 27374 18572 27406
rect 18768 27678 18844 27684
rect 18768 27614 18774 27678
rect 18838 27614 18844 27678
rect 19045 27678 19111 27679
rect 19045 27646 19046 27678
rect 18768 27406 18844 27614
rect 18768 27374 18774 27406
rect 18566 27342 18567 27374
rect 18501 27341 18567 27342
rect 18773 27342 18774 27374
rect 18838 27374 18844 27406
rect 19040 27614 19046 27646
rect 19110 27646 19111 27678
rect 19453 27678 19519 27679
rect 19453 27646 19454 27678
rect 19110 27614 19116 27646
rect 19040 27406 19116 27614
rect 18838 27342 18839 27374
rect 18773 27341 18839 27342
rect 19040 27342 19046 27406
rect 19110 27342 19116 27406
rect 19040 27336 19116 27342
rect 19448 27614 19454 27646
rect 19518 27646 19519 27678
rect 71269 27678 71335 27679
rect 71269 27646 71270 27678
rect 19518 27614 19524 27646
rect 19448 27406 19524 27614
rect 19448 27342 19454 27406
rect 19518 27342 19524 27406
rect 19448 27336 19524 27342
rect 71264 27614 71270 27646
rect 71334 27646 71335 27678
rect 71677 27678 71743 27679
rect 71677 27646 71678 27678
rect 71334 27614 71340 27646
rect 71264 27406 71340 27614
rect 71264 27342 71270 27406
rect 71334 27342 71340 27406
rect 71264 27336 71340 27342
rect 71672 27614 71678 27646
rect 71742 27646 71743 27678
rect 72629 27678 72695 27679
rect 72629 27646 72630 27678
rect 71742 27614 71748 27646
rect 71672 27406 71748 27614
rect 71672 27342 71678 27406
rect 71742 27342 71748 27406
rect 71672 27336 71748 27342
rect 72624 27614 72630 27646
rect 72694 27646 72695 27678
rect 74805 27678 74871 27679
rect 74805 27646 74806 27678
rect 72694 27614 72700 27646
rect 72624 27406 72700 27614
rect 72624 27342 72630 27406
rect 72694 27342 72700 27406
rect 72624 27336 72700 27342
rect 74800 27614 74806 27646
rect 74870 27646 74871 27678
rect 75213 27678 75279 27679
rect 75213 27646 75214 27678
rect 74870 27614 74876 27646
rect 17821 27270 17887 27271
rect 17821 27238 17822 27270
rect 15776 26966 15782 26998
rect 15368 26928 15444 26934
rect 15781 26934 15782 26966
rect 15846 26966 15852 26998
rect 17816 27206 17822 27238
rect 17886 27238 17887 27270
rect 18632 27270 18708 27276
rect 17886 27206 17892 27238
rect 17816 26998 17892 27206
rect 15846 26934 15847 26966
rect 15781 26933 15847 26934
rect 17816 26934 17822 26998
rect 17886 26934 17892 26998
rect 18632 27206 18638 27270
rect 18702 27206 18708 27270
rect 19181 27270 19247 27271
rect 19181 27238 19182 27270
rect 18632 26998 18708 27206
rect 18632 26966 18638 26998
rect 17816 26928 17892 26934
rect 18637 26934 18638 26966
rect 18702 26966 18708 26998
rect 19176 27206 19182 27238
rect 19246 27238 19247 27270
rect 19584 27270 19660 27276
rect 19246 27206 19252 27238
rect 19176 26998 19252 27206
rect 18702 26934 18703 26966
rect 18637 26933 18703 26934
rect 19176 26934 19182 26998
rect 19246 26934 19252 26998
rect 19584 27206 19590 27270
rect 19654 27206 19660 27270
rect 19584 26998 19660 27206
rect 19584 26966 19590 26998
rect 19176 26928 19252 26934
rect 19589 26934 19590 26966
rect 19654 26966 19660 26998
rect 71400 27270 71476 27276
rect 71400 27206 71406 27270
rect 71470 27206 71476 27270
rect 71677 27270 71743 27271
rect 71677 27238 71678 27270
rect 71400 26998 71476 27206
rect 71400 26966 71406 26998
rect 19654 26934 19655 26966
rect 19589 26933 19655 26934
rect 71405 26934 71406 26966
rect 71470 26966 71476 26998
rect 71672 27206 71678 27238
rect 71742 27238 71743 27270
rect 72488 27270 72564 27276
rect 71742 27206 71748 27238
rect 71672 26998 71748 27206
rect 71470 26934 71471 26966
rect 71405 26933 71471 26934
rect 71672 26934 71678 26998
rect 71742 26934 71748 26998
rect 72488 27206 72494 27270
rect 72558 27206 72564 27270
rect 72488 26998 72564 27206
rect 72488 26966 72494 26998
rect 71672 26928 71748 26934
rect 72493 26934 72494 26966
rect 72558 26966 72564 26998
rect 72896 27270 72972 27276
rect 72896 27206 72902 27270
rect 72966 27206 72972 27270
rect 72896 26998 72972 27206
rect 72896 26966 72902 26998
rect 72558 26934 72559 26966
rect 72493 26933 72559 26934
rect 72901 26934 72902 26966
rect 72966 26966 72972 26998
rect 74800 26998 74876 27614
rect 72966 26934 72967 26966
rect 72901 26933 72967 26934
rect 74800 26934 74806 26998
rect 74870 26934 74876 26998
rect 74800 26928 74876 26934
rect 75208 27614 75214 27646
rect 75278 27646 75279 27678
rect 76437 27678 76503 27679
rect 76437 27646 76438 27678
rect 75278 27614 75284 27646
rect 75208 26998 75284 27614
rect 75208 26934 75214 26998
rect 75278 26934 75284 26998
rect 75208 26928 75284 26934
rect 76432 27614 76438 27646
rect 76502 27646 76503 27678
rect 76502 27614 76508 27646
rect 76432 26998 76508 27614
rect 76432 26934 76438 26998
rect 76502 26934 76508 26998
rect 76432 26928 76508 26934
rect 89760 27406 90108 28974
rect 89760 27342 89766 27406
rect 89830 27342 90108 27406
rect 14416 26862 14492 26868
rect 14416 26798 14422 26862
rect 14486 26798 14492 26862
rect 14416 26318 14492 26798
rect 14416 26286 14422 26318
rect 14421 26254 14422 26286
rect 14486 26286 14492 26318
rect 15096 26862 15172 26868
rect 15096 26798 15102 26862
rect 15166 26798 15172 26862
rect 15096 26318 15172 26798
rect 15096 26286 15102 26318
rect 14486 26254 14487 26286
rect 14421 26253 14487 26254
rect 15101 26254 15102 26286
rect 15166 26286 15172 26318
rect 15640 26862 15716 26868
rect 15640 26798 15646 26862
rect 15710 26798 15716 26862
rect 15166 26254 15167 26286
rect 15101 26253 15167 26254
rect 15640 26182 15716 26798
rect 16184 26862 16260 26868
rect 16184 26798 16190 26862
rect 16254 26798 16260 26862
rect 18501 26862 18567 26863
rect 18501 26830 18502 26862
rect 15640 26150 15646 26182
rect 15645 26118 15646 26150
rect 15710 26150 15716 26182
rect 15912 26318 15988 26324
rect 15912 26254 15918 26318
rect 15982 26254 15988 26318
rect 15710 26118 15711 26150
rect 15645 26117 15711 26118
rect 14421 26046 14487 26047
rect 14421 26014 14422 26046
rect 12920 25438 12926 25502
rect 12990 25438 12996 25502
rect 12920 25432 12996 25438
rect 14416 25982 14422 26014
rect 14486 26014 14487 26046
rect 14824 26046 14900 26052
rect 14486 25982 14492 26014
rect 14416 25502 14492 25982
rect 14824 25982 14830 26046
rect 14894 25982 14900 26046
rect 15101 26046 15167 26047
rect 15101 26014 15102 26046
rect 14824 25638 14900 25982
rect 14824 25606 14830 25638
rect 14829 25574 14830 25606
rect 14894 25606 14900 25638
rect 15096 25982 15102 26014
rect 15166 26014 15167 26046
rect 15781 26046 15847 26047
rect 15781 26014 15782 26046
rect 15166 25982 15172 26014
rect 14894 25574 14895 25606
rect 14829 25573 14895 25574
rect 14416 25438 14422 25502
rect 14486 25438 14492 25502
rect 14416 25432 14492 25438
rect 15096 25502 15172 25982
rect 15096 25438 15102 25502
rect 15166 25438 15172 25502
rect 15096 25432 15172 25438
rect 15776 25982 15782 26014
rect 15846 26014 15847 26046
rect 15846 25982 15852 26014
rect 15776 25502 15852 25982
rect 15776 25438 15782 25502
rect 15846 25438 15852 25502
rect 15912 25502 15988 26254
rect 16184 26182 16260 26798
rect 18496 26798 18502 26830
rect 18566 26830 18567 26862
rect 18909 26862 18975 26863
rect 18909 26830 18910 26862
rect 18566 26798 18572 26830
rect 17957 26590 18023 26591
rect 17957 26558 17958 26590
rect 17952 26526 17958 26558
rect 18022 26558 18023 26590
rect 18496 26590 18572 26798
rect 18022 26526 18028 26558
rect 17952 26318 18028 26526
rect 18496 26526 18502 26590
rect 18566 26526 18572 26590
rect 18496 26520 18572 26526
rect 18904 26798 18910 26830
rect 18974 26830 18975 26862
rect 19045 26862 19111 26863
rect 19045 26830 19046 26862
rect 18974 26798 18980 26830
rect 18904 26590 18980 26798
rect 18904 26526 18910 26590
rect 18974 26526 18980 26590
rect 18904 26520 18980 26526
rect 19040 26798 19046 26830
rect 19110 26830 19111 26862
rect 19453 26862 19519 26863
rect 19453 26830 19454 26862
rect 19110 26798 19116 26830
rect 19040 26590 19116 26798
rect 19040 26526 19046 26590
rect 19110 26526 19116 26590
rect 19040 26520 19116 26526
rect 19448 26798 19454 26830
rect 19518 26830 19519 26862
rect 71269 26862 71335 26863
rect 71269 26830 71270 26862
rect 19518 26798 19524 26830
rect 19448 26590 19524 26798
rect 19448 26526 19454 26590
rect 19518 26526 19524 26590
rect 19448 26520 19524 26526
rect 71264 26798 71270 26830
rect 71334 26830 71335 26862
rect 71808 26862 71884 26868
rect 71334 26798 71340 26830
rect 71264 26590 71340 26798
rect 71264 26526 71270 26590
rect 71334 26526 71340 26590
rect 71808 26798 71814 26862
rect 71878 26798 71884 26862
rect 72357 26862 72423 26863
rect 72357 26830 72358 26862
rect 71808 26590 71884 26798
rect 71808 26558 71814 26590
rect 71264 26520 71340 26526
rect 71813 26526 71814 26558
rect 71878 26558 71884 26590
rect 72352 26798 72358 26830
rect 72422 26830 72423 26862
rect 75213 26862 75279 26863
rect 75213 26830 75214 26862
rect 72422 26798 72428 26830
rect 72352 26590 72428 26798
rect 75208 26798 75214 26830
rect 75278 26830 75279 26862
rect 76024 26862 76100 26868
rect 75278 26798 75284 26830
rect 71878 26526 71879 26558
rect 71813 26525 71879 26526
rect 72352 26526 72358 26590
rect 72422 26526 72428 26590
rect 73037 26590 73103 26591
rect 73037 26558 73038 26590
rect 72352 26520 72428 26526
rect 73032 26526 73038 26558
rect 73102 26558 73103 26590
rect 73102 26526 73108 26558
rect 17952 26254 17958 26318
rect 18022 26254 18028 26318
rect 17952 26248 18028 26254
rect 19176 26454 19252 26460
rect 19176 26390 19182 26454
rect 19246 26390 19252 26454
rect 16184 26150 16190 26182
rect 16189 26118 16190 26150
rect 16254 26150 16260 26182
rect 19176 26182 19252 26390
rect 19176 26150 19182 26182
rect 16254 26118 16255 26150
rect 16189 26117 16255 26118
rect 19181 26118 19182 26150
rect 19246 26150 19252 26182
rect 19448 26454 19524 26460
rect 19448 26390 19454 26454
rect 19518 26390 19524 26454
rect 71269 26454 71335 26455
rect 71269 26422 71270 26454
rect 19448 26182 19524 26390
rect 19448 26150 19454 26182
rect 19246 26118 19247 26150
rect 19181 26117 19247 26118
rect 19453 26118 19454 26150
rect 19518 26150 19524 26182
rect 71264 26390 71270 26422
rect 71334 26422 71335 26454
rect 71672 26454 71748 26460
rect 71334 26390 71340 26422
rect 71264 26182 71340 26390
rect 19518 26118 19519 26150
rect 19453 26117 19519 26118
rect 71264 26118 71270 26182
rect 71334 26118 71340 26182
rect 71672 26390 71678 26454
rect 71742 26390 71748 26454
rect 71672 26182 71748 26390
rect 73032 26318 73108 26526
rect 74669 26454 74735 26455
rect 74669 26422 74670 26454
rect 73032 26254 73038 26318
rect 73102 26254 73108 26318
rect 73032 26248 73108 26254
rect 74664 26390 74670 26422
rect 74734 26422 74735 26454
rect 74734 26390 74740 26422
rect 71672 26150 71678 26182
rect 71264 26112 71340 26118
rect 71677 26118 71678 26150
rect 71742 26150 71748 26182
rect 74664 26182 74740 26390
rect 71742 26118 71743 26150
rect 71677 26117 71743 26118
rect 74664 26118 74670 26182
rect 74734 26118 74740 26182
rect 74664 26112 74740 26118
rect 75208 26182 75284 26798
rect 76024 26798 76030 26862
rect 76094 26798 76100 26862
rect 76024 26318 76100 26798
rect 76024 26286 76030 26318
rect 76029 26254 76030 26286
rect 76094 26286 76100 26318
rect 76296 26862 76372 26868
rect 76296 26798 76302 26862
rect 76366 26798 76372 26862
rect 76296 26318 76372 26798
rect 76296 26286 76302 26318
rect 76094 26254 76095 26286
rect 76029 26253 76095 26254
rect 76301 26254 76302 26286
rect 76366 26286 76372 26318
rect 76366 26254 76367 26286
rect 76301 26253 76367 26254
rect 75208 26118 75214 26182
rect 75278 26118 75284 26182
rect 75208 26112 75284 26118
rect 15912 25470 15918 25502
rect 15776 25432 15852 25438
rect 15917 25438 15918 25470
rect 15982 25470 15988 25502
rect 16048 26046 16124 26052
rect 16048 25982 16054 26046
rect 16118 25982 16124 26046
rect 17685 26046 17751 26047
rect 17685 26014 17686 26046
rect 16048 25502 16124 25982
rect 17680 25982 17686 26014
rect 17750 26014 17751 26046
rect 18637 26046 18703 26047
rect 18637 26014 18638 26046
rect 17750 25982 17756 26014
rect 17680 25638 17756 25982
rect 18632 25982 18638 26014
rect 18702 26014 18703 26046
rect 72216 26046 72292 26052
rect 18702 25982 18708 26014
rect 17680 25574 17686 25638
rect 17750 25574 17756 25638
rect 17680 25568 17756 25574
rect 17952 25774 18028 25780
rect 17952 25710 17958 25774
rect 18022 25710 18028 25774
rect 16048 25470 16054 25502
rect 15982 25438 15983 25470
rect 15917 25437 15983 25438
rect 16053 25438 16054 25470
rect 16118 25470 16124 25502
rect 17952 25502 18028 25710
rect 18632 25774 18708 25982
rect 72216 25982 72222 26046
rect 72286 25982 72292 26046
rect 74669 26046 74735 26047
rect 74669 26014 74670 26046
rect 24621 25910 24687 25911
rect 24621 25878 24622 25910
rect 18632 25710 18638 25774
rect 18702 25710 18708 25774
rect 18632 25704 18708 25710
rect 24616 25846 24622 25878
rect 24686 25878 24687 25910
rect 66373 25910 66439 25911
rect 66373 25878 66374 25910
rect 24686 25846 24692 25878
rect 24616 25638 24692 25846
rect 24616 25574 24622 25638
rect 24686 25574 24692 25638
rect 24616 25568 24692 25574
rect 66368 25846 66374 25878
rect 66438 25878 66439 25910
rect 66438 25846 66444 25878
rect 66368 25638 66444 25846
rect 72216 25774 72292 25982
rect 74664 25982 74670 26014
rect 74734 26014 74735 26046
rect 75077 26046 75143 26047
rect 75077 26014 75078 26046
rect 74734 25982 74740 26014
rect 72216 25742 72222 25774
rect 72221 25710 72222 25742
rect 72286 25742 72292 25774
rect 73037 25774 73103 25775
rect 73037 25742 73038 25774
rect 72286 25710 72287 25742
rect 72221 25709 72287 25710
rect 73032 25710 73038 25742
rect 73102 25742 73103 25774
rect 73102 25710 73108 25742
rect 66368 25574 66374 25638
rect 66438 25574 66444 25638
rect 66368 25568 66444 25574
rect 17952 25470 17958 25502
rect 16118 25438 16119 25470
rect 16053 25437 16119 25438
rect 17957 25438 17958 25470
rect 18022 25470 18028 25502
rect 73032 25502 73108 25710
rect 18022 25438 18023 25470
rect 17957 25437 18023 25438
rect 73032 25438 73038 25502
rect 73102 25438 73108 25502
rect 73032 25432 73108 25438
rect 74664 25502 74740 25982
rect 74664 25438 74670 25502
rect 74734 25438 74740 25502
rect 74664 25432 74740 25438
rect 75072 25982 75078 26014
rect 75142 26014 75143 26046
rect 75757 26046 75823 26047
rect 75757 26014 75758 26046
rect 75142 25982 75148 26014
rect 75072 25502 75148 25982
rect 75072 25438 75078 25502
rect 75142 25438 75148 25502
rect 75072 25432 75148 25438
rect 75752 25982 75758 26014
rect 75822 26014 75823 26046
rect 76296 26046 76372 26052
rect 75822 25982 75828 26014
rect 75752 25502 75828 25982
rect 76296 25982 76302 26046
rect 76366 25982 76372 26046
rect 76437 26046 76503 26047
rect 76437 26014 76438 26046
rect 76296 25638 76372 25982
rect 76296 25606 76302 25638
rect 76301 25574 76302 25606
rect 76366 25606 76372 25638
rect 76432 25982 76438 26014
rect 76502 26014 76503 26046
rect 76502 25982 76508 26014
rect 76366 25574 76367 25606
rect 76301 25573 76367 25574
rect 75752 25438 75758 25502
rect 75822 25438 75828 25502
rect 75752 25432 75828 25438
rect 76432 25502 76508 25982
rect 77389 25910 77455 25911
rect 77389 25878 77390 25910
rect 76432 25438 76438 25502
rect 76502 25438 76508 25502
rect 76432 25432 76508 25438
rect 77384 25846 77390 25878
rect 77454 25878 77455 25910
rect 77454 25846 77460 25878
rect 77384 25502 77460 25846
rect 77384 25438 77390 25502
rect 77454 25438 77460 25502
rect 77384 25432 77460 25438
rect 89760 25638 90108 27342
rect 89760 25574 89766 25638
rect 89830 25574 90108 25638
rect 14693 25366 14759 25367
rect 14693 25334 14694 25366
rect 14688 25302 14694 25334
rect 14758 25334 14759 25366
rect 17816 25366 17892 25372
rect 14758 25302 14764 25334
rect 14688 23870 14764 25302
rect 17816 25302 17822 25366
rect 17886 25302 17892 25366
rect 18229 25366 18295 25367
rect 18229 25334 18230 25366
rect 15237 25230 15303 25231
rect 15237 25198 15238 25230
rect 14688 23806 14694 23870
rect 14758 23806 14764 23870
rect 14688 23800 14764 23806
rect 15232 25166 15238 25198
rect 15302 25198 15303 25230
rect 15302 25166 15308 25198
rect 15232 23870 15308 25166
rect 17816 25094 17892 25302
rect 17816 25062 17822 25094
rect 17821 25030 17822 25062
rect 17886 25062 17892 25094
rect 18224 25302 18230 25334
rect 18294 25334 18295 25366
rect 18496 25366 18572 25372
rect 18294 25302 18300 25334
rect 18224 25094 18300 25302
rect 17886 25030 17887 25062
rect 17821 25029 17887 25030
rect 18224 25030 18230 25094
rect 18294 25030 18300 25094
rect 18496 25302 18502 25366
rect 18566 25302 18572 25366
rect 19045 25366 19111 25367
rect 19045 25334 19046 25366
rect 18496 25094 18572 25302
rect 18496 25062 18502 25094
rect 18224 25024 18300 25030
rect 18501 25030 18502 25062
rect 18566 25062 18572 25094
rect 19040 25302 19046 25334
rect 19110 25334 19111 25366
rect 19589 25366 19655 25367
rect 19589 25334 19590 25366
rect 19110 25302 19116 25334
rect 19040 25094 19116 25302
rect 18566 25030 18567 25062
rect 18501 25029 18567 25030
rect 19040 25030 19046 25094
rect 19110 25030 19116 25094
rect 19040 25024 19116 25030
rect 19584 25302 19590 25334
rect 19654 25334 19655 25366
rect 71400 25366 71476 25372
rect 19654 25302 19660 25334
rect 19584 25094 19660 25302
rect 71400 25302 71406 25366
rect 71470 25302 71476 25366
rect 19584 25030 19590 25094
rect 19654 25030 19660 25094
rect 24621 25094 24687 25095
rect 24621 25062 24622 25094
rect 19584 25024 19660 25030
rect 24616 25030 24622 25062
rect 24686 25062 24687 25094
rect 66368 25094 66444 25100
rect 24686 25030 24692 25062
rect 17816 24958 17892 24964
rect 17816 24894 17822 24958
rect 17886 24894 17892 24958
rect 17816 24686 17892 24894
rect 17816 24654 17822 24686
rect 17821 24622 17822 24654
rect 17886 24654 17892 24686
rect 18768 24958 18844 24964
rect 18768 24894 18774 24958
rect 18838 24894 18844 24958
rect 19181 24958 19247 24959
rect 19181 24926 19182 24958
rect 18768 24686 18844 24894
rect 18768 24654 18774 24686
rect 17886 24622 17887 24654
rect 17821 24621 17887 24622
rect 18773 24622 18774 24654
rect 18838 24654 18844 24686
rect 19176 24894 19182 24926
rect 19246 24926 19247 24958
rect 19448 24958 19524 24964
rect 19246 24894 19252 24926
rect 19176 24686 19252 24894
rect 18838 24622 18839 24654
rect 18773 24621 18839 24622
rect 19176 24622 19182 24686
rect 19246 24622 19252 24686
rect 19448 24894 19454 24958
rect 19518 24894 19524 24958
rect 19448 24686 19524 24894
rect 24616 24822 24692 25030
rect 24616 24758 24622 24822
rect 24686 24758 24692 24822
rect 66368 25030 66374 25094
rect 66438 25030 66444 25094
rect 71400 25094 71476 25302
rect 71400 25062 71406 25094
rect 66368 24822 66444 25030
rect 71405 25030 71406 25062
rect 71470 25062 71476 25094
rect 71672 25366 71748 25372
rect 71672 25302 71678 25366
rect 71742 25302 71748 25366
rect 72221 25366 72287 25367
rect 72221 25334 72222 25366
rect 71672 25094 71748 25302
rect 71672 25062 71678 25094
rect 71470 25030 71471 25062
rect 71405 25029 71471 25030
rect 71677 25030 71678 25062
rect 71742 25062 71748 25094
rect 72216 25302 72222 25334
rect 72286 25334 72287 25366
rect 72896 25366 72972 25372
rect 72286 25302 72292 25334
rect 72216 25094 72292 25302
rect 71742 25030 71743 25062
rect 71677 25029 71743 25030
rect 72216 25030 72222 25094
rect 72286 25030 72292 25094
rect 72896 25302 72902 25366
rect 72966 25302 72972 25366
rect 72896 25094 72972 25302
rect 72896 25062 72902 25094
rect 72216 25024 72292 25030
rect 72901 25030 72902 25062
rect 72966 25062 72972 25094
rect 74664 25366 74740 25372
rect 74664 25302 74670 25366
rect 74734 25302 74740 25366
rect 72966 25030 72967 25062
rect 72901 25029 72967 25030
rect 71405 24958 71471 24959
rect 71405 24926 71406 24958
rect 66368 24790 66374 24822
rect 24616 24752 24692 24758
rect 66373 24758 66374 24790
rect 66438 24790 66444 24822
rect 71400 24894 71406 24926
rect 71470 24926 71471 24958
rect 71672 24958 71748 24964
rect 71470 24894 71476 24926
rect 66438 24758 66439 24790
rect 66373 24757 66439 24758
rect 19448 24654 19454 24686
rect 19176 24616 19252 24622
rect 19453 24622 19454 24654
rect 19518 24654 19524 24686
rect 71400 24686 71476 24894
rect 19518 24622 19519 24654
rect 19453 24621 19519 24622
rect 71400 24622 71406 24686
rect 71470 24622 71476 24686
rect 71672 24894 71678 24958
rect 71742 24894 71748 24958
rect 71672 24686 71748 24894
rect 71672 24654 71678 24686
rect 71400 24616 71476 24622
rect 71677 24622 71678 24654
rect 71742 24654 71748 24686
rect 72216 24958 72292 24964
rect 72216 24894 72222 24958
rect 72286 24894 72292 24958
rect 72216 24686 72292 24894
rect 72216 24654 72222 24686
rect 71742 24622 71743 24654
rect 71677 24621 71743 24622
rect 72221 24622 72222 24654
rect 72286 24654 72292 24686
rect 73032 24958 73108 24964
rect 73032 24894 73038 24958
rect 73102 24894 73108 24958
rect 73032 24686 73108 24894
rect 73032 24654 73038 24686
rect 72286 24622 72287 24654
rect 72221 24621 72287 24622
rect 73037 24622 73038 24654
rect 73102 24654 73108 24686
rect 73102 24622 73103 24654
rect 73037 24621 73103 24622
rect 17952 24550 18028 24556
rect 17952 24486 17958 24550
rect 18022 24486 18028 24550
rect 17952 24278 18028 24486
rect 17952 24246 17958 24278
rect 17957 24214 17958 24246
rect 18022 24246 18028 24278
rect 18224 24550 18300 24556
rect 18224 24486 18230 24550
rect 18294 24486 18300 24550
rect 18637 24550 18703 24551
rect 18637 24518 18638 24550
rect 18224 24278 18300 24486
rect 18224 24246 18230 24278
rect 18022 24214 18023 24246
rect 17957 24213 18023 24214
rect 18229 24214 18230 24246
rect 18294 24246 18300 24278
rect 18632 24486 18638 24518
rect 18702 24518 18703 24550
rect 19040 24550 19116 24556
rect 18702 24486 18708 24518
rect 18632 24278 18708 24486
rect 18294 24214 18295 24246
rect 18229 24213 18295 24214
rect 18632 24214 18638 24278
rect 18702 24214 18708 24278
rect 19040 24486 19046 24550
rect 19110 24486 19116 24550
rect 19040 24278 19116 24486
rect 19040 24246 19046 24278
rect 18632 24208 18708 24214
rect 19045 24214 19046 24246
rect 19110 24246 19116 24278
rect 19584 24550 19660 24556
rect 19584 24486 19590 24550
rect 19654 24486 19660 24550
rect 71269 24550 71335 24551
rect 71269 24518 71270 24550
rect 19584 24278 19660 24486
rect 19584 24246 19590 24278
rect 19110 24214 19111 24246
rect 19045 24213 19111 24214
rect 19589 24214 19590 24246
rect 19654 24246 19660 24278
rect 71264 24486 71270 24518
rect 71334 24518 71335 24550
rect 71677 24550 71743 24551
rect 71677 24518 71678 24550
rect 71334 24486 71340 24518
rect 71264 24278 71340 24486
rect 19654 24214 19655 24246
rect 19589 24213 19655 24214
rect 71264 24214 71270 24278
rect 71334 24214 71340 24278
rect 71264 24208 71340 24214
rect 71672 24486 71678 24518
rect 71742 24518 71743 24550
rect 72629 24550 72695 24551
rect 72629 24518 72630 24550
rect 71742 24486 71748 24518
rect 71672 24278 71748 24486
rect 71672 24214 71678 24278
rect 71742 24214 71748 24278
rect 71672 24208 71748 24214
rect 72624 24486 72630 24518
rect 72694 24518 72695 24550
rect 73037 24550 73103 24551
rect 73037 24518 73038 24550
rect 72694 24486 72700 24518
rect 72624 24278 72700 24486
rect 72624 24214 72630 24278
rect 72694 24214 72700 24278
rect 72624 24208 72700 24214
rect 73032 24486 73038 24518
rect 73102 24518 73103 24550
rect 73102 24486 73108 24518
rect 73032 24278 73108 24486
rect 73032 24214 73038 24278
rect 73102 24214 73108 24278
rect 73032 24208 73108 24214
rect 17821 24142 17887 24143
rect 17821 24110 17822 24142
rect 15232 23806 15238 23870
rect 15302 23806 15308 23870
rect 15232 23800 15308 23806
rect 17816 24078 17822 24110
rect 17886 24110 17887 24142
rect 18365 24142 18431 24143
rect 18365 24110 18366 24142
rect 17886 24078 17892 24110
rect 17816 23870 17892 24078
rect 17816 23806 17822 23870
rect 17886 23806 17892 23870
rect 17816 23800 17892 23806
rect 18360 24078 18366 24110
rect 18430 24110 18431 24142
rect 18501 24142 18567 24143
rect 18501 24110 18502 24142
rect 18430 24078 18436 24110
rect 18360 23870 18436 24078
rect 18360 23806 18366 23870
rect 18430 23806 18436 23870
rect 18360 23800 18436 23806
rect 18496 24078 18502 24110
rect 18566 24110 18567 24142
rect 19181 24142 19247 24143
rect 19181 24110 19182 24142
rect 18566 24078 18572 24110
rect 18496 23870 18572 24078
rect 18496 23806 18502 23870
rect 18566 23806 18572 23870
rect 18496 23800 18572 23806
rect 19176 24078 19182 24110
rect 19246 24110 19247 24142
rect 19453 24142 19519 24143
rect 19453 24110 19454 24142
rect 19246 24078 19252 24110
rect 19176 23870 19252 24078
rect 19176 23806 19182 23870
rect 19246 23806 19252 23870
rect 19176 23800 19252 23806
rect 19448 24078 19454 24110
rect 19518 24110 19519 24142
rect 71400 24142 71476 24148
rect 19518 24078 19524 24110
rect 19448 23870 19524 24078
rect 19448 23806 19454 23870
rect 19518 23806 19524 23870
rect 71400 24078 71406 24142
rect 71470 24078 71476 24142
rect 71677 24142 71743 24143
rect 71677 24110 71678 24142
rect 71400 23870 71476 24078
rect 71400 23838 71406 23870
rect 19448 23800 19524 23806
rect 71405 23806 71406 23838
rect 71470 23838 71476 23870
rect 71672 24078 71678 24110
rect 71742 24110 71743 24142
rect 72085 24142 72151 24143
rect 72085 24110 72086 24142
rect 71742 24078 71748 24110
rect 71672 23870 71748 24078
rect 71470 23806 71471 23838
rect 71405 23805 71471 23806
rect 71672 23806 71678 23870
rect 71742 23806 71748 23870
rect 71672 23800 71748 23806
rect 72080 24078 72086 24110
rect 72150 24110 72151 24142
rect 72488 24142 72564 24148
rect 72150 24078 72156 24110
rect 72080 23870 72156 24078
rect 72080 23806 72086 23870
rect 72150 23806 72156 23870
rect 72488 24078 72494 24142
rect 72558 24078 72564 24142
rect 72901 24142 72967 24143
rect 72901 24110 72902 24142
rect 72488 23870 72564 24078
rect 72488 23838 72494 23870
rect 72080 23800 72156 23806
rect 72493 23806 72494 23838
rect 72558 23838 72564 23870
rect 72896 24078 72902 24110
rect 72966 24110 72967 24142
rect 72966 24078 72972 24110
rect 72896 23870 72972 24078
rect 72558 23806 72559 23838
rect 72493 23805 72559 23806
rect 72896 23806 72902 23870
rect 72966 23806 72972 23870
rect 74664 23870 74740 25302
rect 76296 25366 76372 25372
rect 76296 25302 76302 25366
rect 76366 25302 76372 25366
rect 75077 24142 75143 24143
rect 75077 24110 75078 24142
rect 74664 23838 74670 23870
rect 72896 23800 72972 23806
rect 74669 23806 74670 23838
rect 74734 23838 74740 23870
rect 75072 24078 75078 24110
rect 75142 24110 75143 24142
rect 75142 24078 75148 24110
rect 75072 23870 75148 24078
rect 74734 23806 74735 23838
rect 74669 23805 74735 23806
rect 75072 23806 75078 23870
rect 75142 23806 75148 23870
rect 76296 23870 76372 25302
rect 76296 23838 76302 23870
rect 75072 23800 75148 23806
rect 76301 23806 76302 23838
rect 76366 23838 76372 23870
rect 89760 23870 90108 25574
rect 76366 23806 76367 23838
rect 76301 23805 76367 23806
rect 89760 23806 89766 23870
rect 89830 23806 90108 23870
rect 15237 23734 15303 23735
rect 15237 23702 15238 23734
rect 15232 23670 15238 23702
rect 15302 23702 15303 23734
rect 15781 23734 15847 23735
rect 15781 23702 15782 23734
rect 15302 23670 15308 23702
rect 3672 23462 3748 23468
rect 3672 23398 3678 23462
rect 3742 23398 3748 23462
rect 3672 20878 3748 23398
rect 15232 23054 15308 23670
rect 15232 22990 15238 23054
rect 15302 22990 15308 23054
rect 15232 22984 15308 22990
rect 15776 23670 15782 23702
rect 15846 23702 15847 23734
rect 16189 23734 16255 23735
rect 16189 23702 16190 23734
rect 15846 23670 15852 23702
rect 15776 23054 15852 23670
rect 15776 22990 15782 23054
rect 15846 22990 15852 23054
rect 15776 22984 15852 22990
rect 16184 23670 16190 23702
rect 16254 23702 16255 23734
rect 17816 23734 17892 23740
rect 16254 23670 16260 23702
rect 16184 23054 16260 23670
rect 17816 23670 17822 23734
rect 17886 23670 17892 23734
rect 17816 23462 17892 23670
rect 17816 23430 17822 23462
rect 17821 23398 17822 23430
rect 17886 23430 17892 23462
rect 18224 23734 18300 23740
rect 18224 23670 18230 23734
rect 18294 23670 18300 23734
rect 19181 23734 19247 23735
rect 19181 23702 19182 23734
rect 18224 23462 18300 23670
rect 18224 23430 18230 23462
rect 17886 23398 17887 23430
rect 17821 23397 17887 23398
rect 18229 23398 18230 23430
rect 18294 23430 18300 23462
rect 19176 23670 19182 23702
rect 19246 23702 19247 23734
rect 19448 23734 19524 23740
rect 19246 23670 19252 23702
rect 19176 23462 19252 23670
rect 18294 23398 18295 23430
rect 18229 23397 18295 23398
rect 19176 23398 19182 23462
rect 19246 23398 19252 23462
rect 19448 23670 19454 23734
rect 19518 23670 19524 23734
rect 19448 23462 19524 23670
rect 19448 23430 19454 23462
rect 19176 23392 19252 23398
rect 19453 23398 19454 23430
rect 19518 23430 19524 23462
rect 71264 23734 71340 23740
rect 71264 23670 71270 23734
rect 71334 23670 71340 23734
rect 71264 23462 71340 23670
rect 71264 23430 71270 23462
rect 19518 23398 19519 23430
rect 19453 23397 19519 23398
rect 71269 23398 71270 23430
rect 71334 23430 71340 23462
rect 71672 23734 71748 23740
rect 71672 23670 71678 23734
rect 71742 23670 71748 23734
rect 72085 23734 72151 23735
rect 72085 23702 72086 23734
rect 71672 23462 71748 23670
rect 71672 23430 71678 23462
rect 71334 23398 71335 23430
rect 71269 23397 71335 23398
rect 71677 23398 71678 23430
rect 71742 23430 71748 23462
rect 72080 23670 72086 23702
rect 72150 23702 72151 23734
rect 73032 23734 73108 23740
rect 72150 23670 72156 23702
rect 72080 23462 72156 23670
rect 71742 23398 71743 23430
rect 71677 23397 71743 23398
rect 72080 23398 72086 23462
rect 72150 23398 72156 23462
rect 73032 23670 73038 23734
rect 73102 23670 73108 23734
rect 73032 23462 73108 23670
rect 73032 23430 73038 23462
rect 72080 23392 72156 23398
rect 73037 23398 73038 23430
rect 73102 23430 73108 23462
rect 74664 23734 74740 23740
rect 74664 23670 74670 23734
rect 74734 23670 74740 23734
rect 73102 23398 73103 23430
rect 73037 23397 73103 23398
rect 17821 23326 17887 23327
rect 17821 23294 17822 23326
rect 16184 22990 16190 23054
rect 16254 22990 16260 23054
rect 16184 22984 16260 22990
rect 17816 23262 17822 23294
rect 17886 23294 17887 23326
rect 18496 23326 18572 23332
rect 17886 23262 17892 23294
rect 17816 23054 17892 23262
rect 17816 22990 17822 23054
rect 17886 22990 17892 23054
rect 18496 23262 18502 23326
rect 18566 23262 18572 23326
rect 18496 23054 18572 23262
rect 18496 23022 18502 23054
rect 17816 22984 17892 22990
rect 18501 22990 18502 23022
rect 18566 23022 18572 23054
rect 19176 23326 19252 23332
rect 19176 23262 19182 23326
rect 19246 23262 19252 23326
rect 19589 23326 19655 23327
rect 19589 23294 19590 23326
rect 19176 23054 19252 23262
rect 19176 23022 19182 23054
rect 18566 22990 18567 23022
rect 18501 22989 18567 22990
rect 19181 22990 19182 23022
rect 19246 23022 19252 23054
rect 19584 23262 19590 23294
rect 19654 23294 19655 23326
rect 71269 23326 71335 23327
rect 71269 23294 71270 23326
rect 19654 23262 19660 23294
rect 19584 23054 19660 23262
rect 19246 22990 19247 23022
rect 19181 22989 19247 22990
rect 19584 22990 19590 23054
rect 19654 22990 19660 23054
rect 19584 22984 19660 22990
rect 71264 23262 71270 23294
rect 71334 23294 71335 23326
rect 71677 23326 71743 23327
rect 71677 23294 71678 23326
rect 71334 23262 71340 23294
rect 71264 23054 71340 23262
rect 71264 22990 71270 23054
rect 71334 22990 71340 23054
rect 71264 22984 71340 22990
rect 71672 23262 71678 23294
rect 71742 23294 71743 23326
rect 72080 23326 72156 23332
rect 71742 23262 71748 23294
rect 71672 23054 71748 23262
rect 71672 22990 71678 23054
rect 71742 22990 71748 23054
rect 72080 23262 72086 23326
rect 72150 23262 72156 23326
rect 72080 23054 72156 23262
rect 72080 23022 72086 23054
rect 71672 22984 71748 22990
rect 72085 22990 72086 23022
rect 72150 23022 72156 23054
rect 72896 23326 72972 23332
rect 72896 23262 72902 23326
rect 72966 23262 72972 23326
rect 72896 23054 72972 23262
rect 72896 23022 72902 23054
rect 72150 22990 72151 23022
rect 72085 22989 72151 22990
rect 72901 22990 72902 23022
rect 72966 23022 72972 23054
rect 74664 23054 74740 23670
rect 74664 23022 74670 23054
rect 72966 22990 72967 23022
rect 72901 22989 72967 22990
rect 74669 22990 74670 23022
rect 74734 23022 74740 23054
rect 75480 23734 75556 23740
rect 75480 23670 75486 23734
rect 75550 23670 75556 23734
rect 75480 23054 75556 23670
rect 75480 23022 75486 23054
rect 74734 22990 74735 23022
rect 74669 22989 74735 22990
rect 75485 22990 75486 23022
rect 75550 23022 75556 23054
rect 76024 23734 76100 23740
rect 76024 23670 76030 23734
rect 76094 23670 76100 23734
rect 76024 23054 76100 23670
rect 76024 23022 76030 23054
rect 75550 22990 75551 23022
rect 75485 22989 75551 22990
rect 76029 22990 76030 23022
rect 76094 23022 76100 23054
rect 76094 22990 76095 23022
rect 76029 22989 76095 22990
rect 15237 22918 15303 22919
rect 15237 22886 15238 22918
rect 15232 22854 15238 22886
rect 15302 22886 15303 22918
rect 15640 22918 15716 22924
rect 15302 22854 15308 22886
rect 15096 22646 15172 22652
rect 15096 22582 15102 22646
rect 15166 22582 15172 22646
rect 15096 21558 15172 22582
rect 15096 21526 15102 21558
rect 15101 21494 15102 21526
rect 15166 21526 15172 21558
rect 15232 21558 15308 22854
rect 15640 22854 15646 22918
rect 15710 22854 15716 22918
rect 19181 22918 19247 22919
rect 19181 22886 19182 22918
rect 15640 22646 15716 22854
rect 19176 22854 19182 22886
rect 19246 22886 19247 22918
rect 19584 22918 19660 22924
rect 19246 22854 19252 22886
rect 15640 22614 15646 22646
rect 15645 22582 15646 22614
rect 15710 22614 15716 22646
rect 17957 22646 18023 22647
rect 17957 22614 17958 22646
rect 15710 22582 15711 22614
rect 15645 22581 15711 22582
rect 17952 22582 17958 22614
rect 18022 22614 18023 22646
rect 19176 22646 19252 22854
rect 18022 22582 18028 22614
rect 17952 22374 18028 22582
rect 19176 22582 19182 22646
rect 19246 22582 19252 22646
rect 19584 22854 19590 22918
rect 19654 22854 19660 22918
rect 19584 22646 19660 22854
rect 19584 22614 19590 22646
rect 19176 22576 19252 22582
rect 19589 22582 19590 22614
rect 19654 22614 19660 22646
rect 71400 22918 71476 22924
rect 71400 22854 71406 22918
rect 71470 22854 71476 22918
rect 71400 22646 71476 22854
rect 71400 22614 71406 22646
rect 19654 22582 19655 22614
rect 19589 22581 19655 22582
rect 71405 22582 71406 22614
rect 71470 22614 71476 22646
rect 71808 22918 71884 22924
rect 71808 22854 71814 22918
rect 71878 22854 71884 22918
rect 72085 22918 72151 22919
rect 72085 22886 72086 22918
rect 71808 22646 71884 22854
rect 71808 22614 71814 22646
rect 71470 22582 71471 22614
rect 71405 22581 71471 22582
rect 71813 22582 71814 22614
rect 71878 22614 71884 22646
rect 72080 22854 72086 22886
rect 72150 22886 72151 22918
rect 72488 22918 72564 22924
rect 72150 22854 72156 22886
rect 72080 22646 72156 22854
rect 71878 22582 71879 22614
rect 71813 22581 71879 22582
rect 72080 22582 72086 22646
rect 72150 22582 72156 22646
rect 72488 22854 72494 22918
rect 72558 22854 72564 22918
rect 72488 22646 72564 22854
rect 75072 22918 75148 22924
rect 75072 22854 75078 22918
rect 75142 22854 75148 22918
rect 75485 22918 75551 22919
rect 75485 22886 75486 22918
rect 72488 22614 72494 22646
rect 72080 22576 72156 22582
rect 72493 22582 72494 22614
rect 72558 22614 72564 22646
rect 72901 22646 72967 22647
rect 72901 22614 72902 22646
rect 72558 22582 72559 22614
rect 72493 22581 72559 22582
rect 72896 22582 72902 22614
rect 72966 22614 72967 22646
rect 72966 22582 72972 22614
rect 19045 22510 19111 22511
rect 19045 22478 19046 22510
rect 17952 22310 17958 22374
rect 18022 22310 18028 22374
rect 17952 22304 18028 22310
rect 19040 22446 19046 22478
rect 19110 22478 19111 22510
rect 19453 22510 19519 22511
rect 19453 22478 19454 22510
rect 19110 22446 19116 22478
rect 19040 22238 19116 22446
rect 19040 22174 19046 22238
rect 19110 22174 19116 22238
rect 19040 22168 19116 22174
rect 19448 22446 19454 22478
rect 19518 22478 19519 22510
rect 71269 22510 71335 22511
rect 71269 22478 71270 22510
rect 19518 22446 19524 22478
rect 19448 22238 19524 22446
rect 19448 22174 19454 22238
rect 19518 22174 19524 22238
rect 19448 22168 19524 22174
rect 71264 22446 71270 22478
rect 71334 22478 71335 22510
rect 71677 22510 71743 22511
rect 71677 22478 71678 22510
rect 71334 22446 71340 22478
rect 71264 22238 71340 22446
rect 71264 22174 71270 22238
rect 71334 22174 71340 22238
rect 71264 22168 71340 22174
rect 71672 22446 71678 22478
rect 71742 22478 71743 22510
rect 71742 22446 71748 22478
rect 71672 22238 71748 22446
rect 72896 22374 72972 22582
rect 72896 22310 72902 22374
rect 72966 22310 72972 22374
rect 72896 22304 72972 22310
rect 71672 22174 71678 22238
rect 71742 22174 71748 22238
rect 71672 22168 71748 22174
rect 18360 22102 18436 22108
rect 18360 22038 18366 22102
rect 18430 22038 18436 22102
rect 17821 21830 17887 21831
rect 17821 21798 17822 21830
rect 15166 21494 15167 21526
rect 15101 21493 15167 21494
rect 15232 21494 15238 21558
rect 15302 21494 15308 21558
rect 15232 21488 15308 21494
rect 17816 21766 17822 21798
rect 17886 21798 17887 21830
rect 18360 21830 18436 22038
rect 18360 21798 18366 21830
rect 17886 21766 17892 21798
rect 17816 21558 17892 21766
rect 18365 21766 18366 21798
rect 18430 21798 18436 21830
rect 18768 22102 18844 22108
rect 18768 22038 18774 22102
rect 18838 22038 18844 22102
rect 18768 21830 18844 22038
rect 72080 22102 72156 22108
rect 72080 22038 72086 22102
rect 72150 22038 72156 22102
rect 18768 21798 18774 21830
rect 18430 21766 18431 21798
rect 18365 21765 18431 21766
rect 18773 21766 18774 21798
rect 18838 21798 18844 21830
rect 24344 21966 24420 21972
rect 24344 21902 24350 21966
rect 24414 21902 24420 21966
rect 66373 21966 66439 21967
rect 66373 21934 66374 21966
rect 18838 21766 18839 21798
rect 18773 21765 18839 21766
rect 24344 21694 24420 21902
rect 66368 21902 66374 21934
rect 66438 21934 66439 21966
rect 66438 21902 66444 21934
rect 24344 21662 24350 21694
rect 24349 21630 24350 21662
rect 24414 21662 24420 21694
rect 24480 21694 24556 21700
rect 24414 21630 24415 21662
rect 24349 21629 24415 21630
rect 24480 21630 24486 21694
rect 24550 21630 24556 21694
rect 17816 21494 17822 21558
rect 17886 21494 17892 21558
rect 17816 21488 17892 21494
rect 17952 21422 18028 21428
rect 17952 21358 17958 21422
rect 18022 21358 18028 21422
rect 18909 21422 18975 21423
rect 18909 21390 18910 21422
rect 15781 21286 15847 21287
rect 15781 21254 15782 21286
rect 3672 20846 3678 20878
rect 3677 20814 3678 20846
rect 3742 20846 3748 20878
rect 15776 21222 15782 21254
rect 15846 21254 15847 21286
rect 16189 21286 16255 21287
rect 16189 21254 16190 21286
rect 15846 21222 15852 21254
rect 3742 20814 3743 20846
rect 3677 20813 3743 20814
rect 15776 20742 15852 21222
rect 15776 20678 15782 20742
rect 15846 20678 15852 20742
rect 15776 20672 15852 20678
rect 16184 21222 16190 21254
rect 16254 21254 16255 21286
rect 16254 21222 16260 21254
rect 16184 20742 16260 21222
rect 17952 21150 18028 21358
rect 17952 21118 17958 21150
rect 17957 21086 17958 21118
rect 18022 21118 18028 21150
rect 18904 21358 18910 21390
rect 18974 21390 18975 21422
rect 18974 21358 18980 21390
rect 18904 21150 18980 21358
rect 24480 21286 24556 21630
rect 66368 21694 66444 21902
rect 72080 21830 72156 22038
rect 72080 21798 72086 21830
rect 72085 21766 72086 21798
rect 72150 21798 72156 21830
rect 72896 21830 72972 21836
rect 72150 21766 72151 21798
rect 72085 21765 72151 21766
rect 72896 21766 72902 21830
rect 72966 21766 72972 21830
rect 66368 21630 66374 21694
rect 66438 21630 66444 21694
rect 66368 21624 66444 21630
rect 24621 21558 24687 21559
rect 24621 21526 24622 21558
rect 24480 21254 24486 21286
rect 24485 21222 24486 21254
rect 24550 21254 24556 21286
rect 24616 21494 24622 21526
rect 24686 21526 24687 21558
rect 66504 21558 66580 21564
rect 24686 21494 24692 21526
rect 24616 21286 24692 21494
rect 24550 21222 24551 21254
rect 24485 21221 24551 21222
rect 24616 21222 24622 21286
rect 24686 21222 24692 21286
rect 66504 21494 66510 21558
rect 66574 21494 66580 21558
rect 72896 21558 72972 21766
rect 72896 21526 72902 21558
rect 66504 21286 66580 21494
rect 72901 21494 72902 21526
rect 72966 21526 72972 21558
rect 75072 21558 75148 22854
rect 75072 21526 75078 21558
rect 72966 21494 72967 21526
rect 72901 21493 72967 21494
rect 75077 21494 75078 21526
rect 75142 21526 75148 21558
rect 75480 22854 75486 22886
rect 75550 22886 75551 22918
rect 75550 22854 75556 22886
rect 75480 21558 75556 22854
rect 75142 21494 75143 21526
rect 75077 21493 75143 21494
rect 75480 21494 75486 21558
rect 75550 21494 75556 21558
rect 75480 21488 75556 21494
rect 89760 22238 90108 23806
rect 89760 22174 89766 22238
rect 89830 22174 90108 22238
rect 72221 21422 72287 21423
rect 72221 21390 72222 21422
rect 66504 21254 66510 21286
rect 24616 21216 24692 21222
rect 66509 21222 66510 21254
rect 66574 21254 66580 21286
rect 72216 21358 72222 21390
rect 72286 21390 72287 21422
rect 73037 21422 73103 21423
rect 73037 21390 73038 21422
rect 72286 21358 72292 21390
rect 66574 21222 66575 21254
rect 66509 21221 66575 21222
rect 18022 21086 18023 21118
rect 17957 21085 18023 21086
rect 18904 21086 18910 21150
rect 18974 21086 18980 21150
rect 66509 21150 66575 21151
rect 66509 21118 66510 21150
rect 18904 21080 18980 21086
rect 66504 21086 66510 21118
rect 66574 21118 66575 21150
rect 72216 21150 72292 21358
rect 66574 21086 66580 21118
rect 17957 21014 18023 21015
rect 17957 20982 17958 21014
rect 16184 20678 16190 20742
rect 16254 20678 16260 20742
rect 16184 20672 16260 20678
rect 17952 20950 17958 20982
rect 18022 20982 18023 21014
rect 19045 21014 19111 21015
rect 19045 20982 19046 21014
rect 18022 20950 18028 20982
rect 17952 20742 18028 20950
rect 19040 20950 19046 20982
rect 19110 20982 19111 21014
rect 19589 21014 19655 21015
rect 19589 20982 19590 21014
rect 19110 20950 19116 20982
rect 17952 20678 17958 20742
rect 18022 20678 18028 20742
rect 17952 20672 18028 20678
rect 18496 20878 18572 20884
rect 18496 20814 18502 20878
rect 18566 20814 18572 20878
rect 3949 20606 4015 20607
rect 3949 20574 3950 20606
rect 3944 20542 3950 20574
rect 4014 20574 4015 20606
rect 13600 20606 13676 20612
rect 4014 20542 4020 20574
rect 3128 19246 3204 19252
rect 3128 19182 3134 19246
rect 3198 19182 3204 19246
rect 3128 18974 3204 19182
rect 3128 18942 3134 18974
rect 3133 18910 3134 18942
rect 3198 18942 3204 18974
rect 3198 18910 3199 18942
rect 3133 18909 3199 18910
rect 2460 18325 2526 18326
rect 2460 18261 2461 18325
rect 2525 18261 2526 18325
rect 2460 18260 2526 18261
rect 3944 18022 4020 20542
rect 13600 20542 13606 20606
rect 13670 20542 13676 20606
rect 13600 19382 13676 20542
rect 13600 19350 13606 19382
rect 13605 19318 13606 19350
rect 13670 19350 13676 19382
rect 14008 20606 14084 20612
rect 14008 20542 14014 20606
rect 14078 20542 14084 20606
rect 18496 20606 18572 20814
rect 19040 20742 19116 20950
rect 19040 20678 19046 20742
rect 19110 20678 19116 20742
rect 19040 20672 19116 20678
rect 19584 20950 19590 20982
rect 19654 20982 19655 21014
rect 19654 20950 19660 20982
rect 19584 20742 19660 20950
rect 66504 20878 66580 21086
rect 72216 21086 72222 21150
rect 72286 21086 72292 21150
rect 72216 21080 72292 21086
rect 73032 21358 73038 21390
rect 73102 21390 73103 21422
rect 75485 21422 75551 21423
rect 75485 21390 75486 21422
rect 73102 21358 73108 21390
rect 73032 21150 73108 21358
rect 75480 21358 75486 21390
rect 75550 21390 75551 21422
rect 75893 21422 75959 21423
rect 75893 21390 75894 21422
rect 75550 21358 75556 21390
rect 74805 21286 74871 21287
rect 74805 21254 74806 21286
rect 73032 21086 73038 21150
rect 73102 21086 73108 21150
rect 73032 21080 73108 21086
rect 74800 21222 74806 21254
rect 74870 21254 74871 21286
rect 75072 21286 75148 21292
rect 74870 21222 74876 21254
rect 66504 20814 66510 20878
rect 66574 20814 66580 20878
rect 66504 20808 66580 20814
rect 71400 21014 71476 21020
rect 71400 20950 71406 21014
rect 71470 20950 71476 21014
rect 71813 21014 71879 21015
rect 71813 20982 71814 21014
rect 19584 20678 19590 20742
rect 19654 20678 19660 20742
rect 71400 20742 71476 20950
rect 71400 20710 71406 20742
rect 19584 20672 19660 20678
rect 71405 20678 71406 20710
rect 71470 20710 71476 20742
rect 71808 20950 71814 20982
rect 71878 20982 71879 21014
rect 73037 21014 73103 21015
rect 73037 20982 73038 21014
rect 71878 20950 71884 20982
rect 71808 20742 71884 20950
rect 71470 20678 71471 20710
rect 71405 20677 71471 20678
rect 71808 20678 71814 20742
rect 71878 20678 71884 20742
rect 71808 20672 71884 20678
rect 73032 20950 73038 20982
rect 73102 20982 73103 21014
rect 73102 20950 73108 20982
rect 73032 20742 73108 20950
rect 73032 20678 73038 20742
rect 73102 20678 73108 20742
rect 73032 20672 73108 20678
rect 74800 20742 74876 21222
rect 74800 20678 74806 20742
rect 74870 20678 74876 20742
rect 75072 21222 75078 21286
rect 75142 21222 75148 21286
rect 75072 20742 75148 21222
rect 75072 20710 75078 20742
rect 74800 20672 74876 20678
rect 75077 20678 75078 20710
rect 75142 20710 75148 20742
rect 75480 20742 75556 21358
rect 75142 20678 75143 20710
rect 75077 20677 75143 20678
rect 75480 20678 75486 20742
rect 75550 20678 75556 20742
rect 75480 20672 75556 20678
rect 75888 21358 75894 21390
rect 75958 21390 75959 21422
rect 75958 21358 75964 21390
rect 75888 20742 75964 21358
rect 75888 20678 75894 20742
rect 75958 20678 75964 20742
rect 75888 20672 75964 20678
rect 18496 20574 18502 20606
rect 13670 19318 13671 19350
rect 13605 19317 13671 19318
rect 3944 17958 3950 18022
rect 4014 17958 4020 18022
rect 3944 17952 4020 17958
rect 11560 19246 11636 19252
rect 11560 19182 11566 19246
rect 11630 19182 11636 19246
rect 952 17142 1230 17206
rect 1294 17142 1300 17206
rect 2453 17206 2519 17207
rect 2453 17174 2454 17206
rect 952 15710 1300 17142
rect 2448 17142 2454 17174
rect 2518 17174 2519 17206
rect 2518 17142 2524 17174
rect 2448 16526 2524 17142
rect 2448 16462 2454 16526
rect 2518 16462 2524 16526
rect 11560 16526 11636 19182
rect 14008 18022 14084 20542
rect 18501 20542 18502 20574
rect 18566 20574 18572 20606
rect 19040 20606 19116 20612
rect 18566 20542 18567 20574
rect 18501 20541 18567 20542
rect 19040 20542 19046 20606
rect 19110 20542 19116 20606
rect 19453 20606 19519 20607
rect 19453 20574 19454 20606
rect 14008 17990 14014 18022
rect 14013 17958 14014 17990
rect 14078 17990 14084 18022
rect 14078 17958 14079 17990
rect 14013 17957 14079 17958
rect 11701 17886 11767 17887
rect 11701 17854 11702 17886
rect 11560 16494 11566 16526
rect 2448 16456 2524 16462
rect 11565 16462 11566 16494
rect 11630 16494 11636 16526
rect 11696 17822 11702 17854
rect 11766 17854 11767 17886
rect 11766 17822 11772 17854
rect 11630 16462 11631 16494
rect 11565 16461 11631 16462
rect 11429 16390 11495 16391
rect 11429 16358 11430 16390
rect 952 15646 1230 15710
rect 1294 15646 1300 15710
rect 952 13806 1300 15646
rect 952 13742 1230 13806
rect 1294 13742 1300 13806
rect 952 12310 1300 13742
rect 11424 16326 11430 16358
rect 11494 16358 11495 16390
rect 11494 16326 11500 16358
rect 11424 13806 11500 16326
rect 11696 15166 11772 17822
rect 19040 17750 19116 20542
rect 19448 20542 19454 20574
rect 19518 20574 19519 20606
rect 77117 20606 77183 20607
rect 77117 20574 77118 20606
rect 19518 20542 19524 20574
rect 19448 20198 19524 20542
rect 77112 20542 77118 20574
rect 77182 20574 77183 20606
rect 79837 20606 79903 20607
rect 79837 20574 79838 20606
rect 77182 20542 77188 20574
rect 19448 20134 19454 20198
rect 19518 20134 19524 20198
rect 19448 20128 19524 20134
rect 66368 20198 66444 20204
rect 66368 20134 66374 20198
rect 66438 20134 66444 20198
rect 19040 17718 19046 17750
rect 19045 17686 19046 17718
rect 19110 17718 19116 17750
rect 19176 19926 19252 19932
rect 19176 19862 19182 19926
rect 19246 19862 19252 19926
rect 19110 17686 19111 17718
rect 19045 17685 19111 17686
rect 16592 17614 16668 17620
rect 16592 17550 16598 17614
rect 16662 17550 16668 17614
rect 11696 15102 11702 15166
rect 11766 15102 11772 15166
rect 11696 15096 11772 15102
rect 16456 16254 16532 16260
rect 16456 16190 16462 16254
rect 16526 16190 16532 16254
rect 11424 13742 11430 13806
rect 11494 13742 11500 13806
rect 11424 13736 11500 13742
rect 11560 15030 11636 15036
rect 11560 14966 11566 15030
rect 11630 14966 11636 15030
rect 952 12246 1230 12310
rect 1294 12246 1300 12310
rect 11560 12310 11636 14966
rect 11701 13534 11767 13535
rect 11701 13502 11702 13534
rect 11560 12278 11566 12310
rect 952 10542 1300 12246
rect 11565 12246 11566 12278
rect 11630 12278 11636 12310
rect 11696 13470 11702 13502
rect 11766 13502 11767 13534
rect 16456 13534 16532 16190
rect 16592 14894 16668 17550
rect 19176 16390 19252 19862
rect 25301 19654 25367 19655
rect 25301 19622 25302 19654
rect 25296 19590 25302 19622
rect 25366 19622 25367 19654
rect 26525 19654 26591 19655
rect 26525 19622 26526 19654
rect 25366 19590 25372 19622
rect 25296 19110 25372 19590
rect 25296 19046 25302 19110
rect 25366 19046 25372 19110
rect 25296 19040 25372 19046
rect 26520 19590 26526 19622
rect 26590 19622 26591 19654
rect 28152 19654 28228 19660
rect 26590 19590 26596 19622
rect 26520 19110 26596 19590
rect 26520 19046 26526 19110
rect 26590 19046 26596 19110
rect 28152 19590 28158 19654
rect 28222 19590 28228 19654
rect 28152 19110 28228 19590
rect 28152 19078 28158 19110
rect 26520 19040 26596 19046
rect 28157 19046 28158 19078
rect 28222 19078 28228 19110
rect 29512 19654 29588 19660
rect 29512 19590 29518 19654
rect 29582 19590 29588 19654
rect 29653 19654 29719 19655
rect 29653 19622 29654 19654
rect 29512 19110 29588 19590
rect 29512 19078 29518 19110
rect 28222 19046 28223 19078
rect 28157 19045 28223 19046
rect 29517 19046 29518 19078
rect 29582 19078 29588 19110
rect 29648 19590 29654 19622
rect 29718 19622 29719 19654
rect 30328 19654 30404 19660
rect 29718 19590 29724 19622
rect 29648 19110 29724 19590
rect 29582 19046 29583 19078
rect 29517 19045 29583 19046
rect 29648 19046 29654 19110
rect 29718 19046 29724 19110
rect 30328 19590 30334 19654
rect 30398 19590 30404 19654
rect 31557 19654 31623 19655
rect 31557 19622 31558 19654
rect 30328 19110 30404 19590
rect 30328 19078 30334 19110
rect 29648 19040 29724 19046
rect 30333 19046 30334 19078
rect 30398 19078 30404 19110
rect 31552 19590 31558 19622
rect 31622 19622 31623 19654
rect 31960 19654 32036 19660
rect 31622 19590 31628 19622
rect 31552 19110 31628 19590
rect 30398 19046 30399 19078
rect 30333 19045 30399 19046
rect 31552 19046 31558 19110
rect 31622 19046 31628 19110
rect 31960 19590 31966 19654
rect 32030 19590 32036 19654
rect 32645 19654 32711 19655
rect 32645 19622 32646 19654
rect 31960 19110 32036 19590
rect 31960 19078 31966 19110
rect 31552 19040 31628 19046
rect 31965 19046 31966 19078
rect 32030 19078 32036 19110
rect 32640 19590 32646 19622
rect 32710 19622 32711 19654
rect 33184 19654 33260 19660
rect 32710 19590 32716 19622
rect 32640 19110 32716 19590
rect 32030 19046 32031 19078
rect 31965 19045 32031 19046
rect 32640 19046 32646 19110
rect 32710 19046 32716 19110
rect 33184 19590 33190 19654
rect 33254 19590 33260 19654
rect 33184 19110 33260 19590
rect 33184 19078 33190 19110
rect 32640 19040 32716 19046
rect 33189 19046 33190 19078
rect 33254 19078 33260 19110
rect 34544 19654 34620 19660
rect 34544 19590 34550 19654
rect 34614 19590 34620 19654
rect 35229 19654 35295 19655
rect 35229 19622 35230 19654
rect 34544 19110 34620 19590
rect 34544 19078 34550 19110
rect 33254 19046 33255 19078
rect 33189 19045 33255 19046
rect 34549 19046 34550 19078
rect 34614 19078 34620 19110
rect 35224 19590 35230 19622
rect 35294 19622 35295 19654
rect 35768 19654 35844 19660
rect 35294 19590 35300 19622
rect 35224 19110 35300 19590
rect 34614 19046 34615 19078
rect 34549 19045 34615 19046
rect 35224 19046 35230 19110
rect 35294 19046 35300 19110
rect 35768 19590 35774 19654
rect 35838 19590 35844 19654
rect 36453 19654 36519 19655
rect 36453 19622 36454 19654
rect 35768 19110 35844 19590
rect 35768 19078 35774 19110
rect 35224 19040 35300 19046
rect 35773 19046 35774 19078
rect 35838 19078 35844 19110
rect 36448 19590 36454 19622
rect 36518 19622 36519 19654
rect 38357 19654 38423 19655
rect 38357 19622 38358 19654
rect 36518 19590 36524 19622
rect 36448 19110 36524 19590
rect 35838 19046 35839 19078
rect 35773 19045 35839 19046
rect 36448 19046 36454 19110
rect 36518 19046 36524 19110
rect 36448 19040 36524 19046
rect 38352 19590 38358 19622
rect 38422 19622 38423 19654
rect 40800 19654 40876 19660
rect 38422 19590 38428 19622
rect 38352 19110 38428 19590
rect 38352 19046 38358 19110
rect 38422 19046 38428 19110
rect 40800 19590 40806 19654
rect 40870 19590 40876 19654
rect 41485 19654 41551 19655
rect 41485 19622 41486 19654
rect 40800 19110 40876 19590
rect 40800 19078 40806 19110
rect 38352 19040 38428 19046
rect 40805 19046 40806 19078
rect 40870 19078 40876 19110
rect 41480 19590 41486 19622
rect 41550 19622 41551 19654
rect 42709 19654 42775 19655
rect 42709 19622 42710 19654
rect 41550 19590 41556 19622
rect 41480 19110 41556 19590
rect 40870 19046 40871 19078
rect 40805 19045 40871 19046
rect 41480 19046 41486 19110
rect 41550 19046 41556 19110
rect 41480 19040 41556 19046
rect 42704 19590 42710 19622
rect 42774 19622 42775 19654
rect 43933 19654 43999 19655
rect 43933 19622 43934 19654
rect 42774 19590 42780 19622
rect 42704 19110 42780 19590
rect 42704 19046 42710 19110
rect 42774 19046 42780 19110
rect 42704 19040 42780 19046
rect 43928 19590 43934 19622
rect 43998 19622 43999 19654
rect 44472 19654 44548 19660
rect 43998 19590 44004 19622
rect 43928 19110 44004 19590
rect 43928 19046 43934 19110
rect 43998 19046 44004 19110
rect 44472 19590 44478 19654
rect 44542 19590 44548 19654
rect 45565 19654 45631 19655
rect 45565 19622 45566 19654
rect 44472 19110 44548 19590
rect 44472 19078 44478 19110
rect 43928 19040 44004 19046
rect 44477 19046 44478 19078
rect 44542 19078 44548 19110
rect 45560 19590 45566 19622
rect 45630 19622 45631 19654
rect 46920 19654 46996 19660
rect 45630 19590 45636 19622
rect 45560 19110 45636 19590
rect 44542 19046 44543 19078
rect 44477 19045 44543 19046
rect 45560 19046 45566 19110
rect 45630 19046 45636 19110
rect 46920 19590 46926 19654
rect 46990 19590 46996 19654
rect 46920 19110 46996 19590
rect 46920 19078 46926 19110
rect 45560 19040 45636 19046
rect 46925 19046 46926 19078
rect 46990 19078 46996 19110
rect 47872 19654 47948 19660
rect 47872 19590 47878 19654
rect 47942 19590 47948 19654
rect 47872 19110 47948 19590
rect 47872 19078 47878 19110
rect 46990 19046 46991 19078
rect 46925 19045 46991 19046
rect 47877 19046 47878 19078
rect 47942 19078 47948 19110
rect 49368 19654 49444 19660
rect 49368 19590 49374 19654
rect 49438 19590 49444 19654
rect 50189 19654 50255 19655
rect 50189 19622 50190 19654
rect 49368 19110 49444 19590
rect 49368 19078 49374 19110
rect 47942 19046 47943 19078
rect 47877 19045 47943 19046
rect 49373 19046 49374 19078
rect 49438 19078 49444 19110
rect 50184 19590 50190 19622
rect 50254 19622 50255 19654
rect 50728 19654 50804 19660
rect 50254 19590 50260 19622
rect 50184 19110 50260 19590
rect 49438 19046 49439 19078
rect 49373 19045 49439 19046
rect 50184 19046 50190 19110
rect 50254 19046 50260 19110
rect 50728 19590 50734 19654
rect 50798 19590 50804 19654
rect 50728 19110 50804 19590
rect 50728 19078 50734 19110
rect 50184 19040 50260 19046
rect 50733 19046 50734 19078
rect 50798 19078 50804 19110
rect 51952 19654 52028 19660
rect 51952 19590 51958 19654
rect 52022 19590 52028 19654
rect 51952 19110 52028 19590
rect 51952 19078 51958 19110
rect 50798 19046 50799 19078
rect 50733 19045 50799 19046
rect 51957 19046 51958 19078
rect 52022 19078 52028 19110
rect 53176 19654 53252 19660
rect 53176 19590 53182 19654
rect 53246 19590 53252 19654
rect 53176 19110 53252 19590
rect 53176 19078 53182 19110
rect 52022 19046 52023 19078
rect 51957 19045 52023 19046
rect 53181 19046 53182 19078
rect 53246 19078 53252 19110
rect 54128 19654 54204 19660
rect 54128 19590 54134 19654
rect 54198 19590 54204 19654
rect 54128 19110 54204 19590
rect 54128 19078 54134 19110
rect 53246 19046 53247 19078
rect 53181 19045 53247 19046
rect 54133 19046 54134 19078
rect 54198 19078 54204 19110
rect 55760 19654 55836 19660
rect 55760 19590 55766 19654
rect 55830 19590 55836 19654
rect 55760 19110 55836 19590
rect 55760 19078 55766 19110
rect 54198 19046 54199 19078
rect 54133 19045 54199 19046
rect 55765 19046 55766 19078
rect 55830 19078 55836 19110
rect 56984 19654 57060 19660
rect 56984 19590 56990 19654
rect 57054 19590 57060 19654
rect 56984 19110 57060 19590
rect 56984 19078 56990 19110
rect 55830 19046 55831 19078
rect 55765 19045 55831 19046
rect 56989 19046 56990 19078
rect 57054 19078 57060 19110
rect 58208 19654 58284 19660
rect 58208 19590 58214 19654
rect 58278 19590 58284 19654
rect 58893 19654 58959 19655
rect 58893 19622 58894 19654
rect 58208 19110 58284 19590
rect 58208 19078 58214 19110
rect 57054 19046 57055 19078
rect 56989 19045 57055 19046
rect 58213 19046 58214 19078
rect 58278 19078 58284 19110
rect 58888 19590 58894 19622
rect 58958 19622 58959 19654
rect 59432 19654 59508 19660
rect 58958 19590 58964 19622
rect 58888 19110 58964 19590
rect 58278 19046 58279 19078
rect 58213 19045 58279 19046
rect 58888 19046 58894 19110
rect 58958 19046 58964 19110
rect 59432 19590 59438 19654
rect 59502 19590 59508 19654
rect 60117 19654 60183 19655
rect 60117 19622 60118 19654
rect 59432 19110 59508 19590
rect 59432 19078 59438 19110
rect 58888 19040 58964 19046
rect 59437 19046 59438 19078
rect 59502 19078 59508 19110
rect 60112 19590 60118 19622
rect 60182 19622 60183 19654
rect 60656 19654 60732 19660
rect 60182 19590 60188 19622
rect 60112 19110 60188 19590
rect 59502 19046 59503 19078
rect 59437 19045 59503 19046
rect 60112 19046 60118 19110
rect 60182 19046 60188 19110
rect 60656 19590 60662 19654
rect 60726 19590 60732 19654
rect 60656 19110 60732 19590
rect 60656 19078 60662 19110
rect 60112 19040 60188 19046
rect 60661 19046 60662 19078
rect 60726 19078 60732 19110
rect 61880 19654 61956 19660
rect 61880 19590 61886 19654
rect 61950 19590 61956 19654
rect 61880 19110 61956 19590
rect 61880 19078 61886 19110
rect 60726 19046 60727 19078
rect 60661 19045 60727 19046
rect 61885 19046 61886 19078
rect 61950 19078 61956 19110
rect 62832 19654 62908 19660
rect 62832 19590 62838 19654
rect 62902 19590 62908 19654
rect 63925 19654 63991 19655
rect 63925 19622 63926 19654
rect 62832 19110 62908 19590
rect 62832 19078 62838 19110
rect 61950 19046 61951 19078
rect 61885 19045 61951 19046
rect 62837 19046 62838 19078
rect 62902 19078 62908 19110
rect 63920 19590 63926 19622
rect 63990 19622 63991 19654
rect 65688 19654 65764 19660
rect 63990 19590 63996 19622
rect 63920 19110 63996 19590
rect 62902 19046 62903 19078
rect 62837 19045 62903 19046
rect 63920 19046 63926 19110
rect 63990 19046 63996 19110
rect 65688 19590 65694 19654
rect 65758 19590 65764 19654
rect 65688 19110 65764 19590
rect 65688 19078 65694 19110
rect 63920 19040 63996 19046
rect 65693 19046 65694 19078
rect 65758 19078 65764 19110
rect 65758 19046 65759 19078
rect 65693 19045 65759 19046
rect 26792 18974 26868 18980
rect 26792 18910 26798 18974
rect 26862 18910 26868 18974
rect 30741 18974 30807 18975
rect 30741 18942 30742 18974
rect 19176 16358 19182 16390
rect 19181 16326 19182 16358
rect 19246 16358 19252 16390
rect 25976 17478 26052 17484
rect 25976 17414 25982 17478
rect 26046 17414 26052 17478
rect 19246 16326 19247 16358
rect 19181 16325 19247 16326
rect 25976 15030 26052 17414
rect 25976 14998 25982 15030
rect 25981 14966 25982 14998
rect 26046 14998 26052 15030
rect 26112 15030 26188 15036
rect 26046 14966 26047 14998
rect 25981 14965 26047 14966
rect 26112 14966 26118 15030
rect 26182 14966 26188 15030
rect 16592 14862 16598 14894
rect 16597 14830 16598 14862
rect 16662 14862 16668 14894
rect 16662 14830 16663 14862
rect 16597 14829 16663 14830
rect 16456 13502 16462 13534
rect 11766 13470 11772 13502
rect 11630 12246 11631 12278
rect 11565 12245 11631 12246
rect 952 10478 1230 10542
rect 1294 10478 1300 10542
rect 952 8910 1300 10478
rect 11560 12174 11636 12180
rect 11560 12110 11566 12174
rect 11630 12110 11636 12174
rect 11560 9454 11636 12110
rect 11696 10950 11772 13470
rect 16461 13470 16462 13502
rect 16526 13502 16532 13534
rect 16592 14758 16668 14764
rect 16592 14694 16598 14758
rect 16662 14694 16668 14758
rect 16526 13470 16527 13502
rect 16461 13469 16527 13470
rect 16592 12174 16668 14694
rect 25981 14214 26047 14215
rect 25981 14182 25982 14214
rect 25976 14150 25982 14182
rect 26046 14182 26047 14214
rect 26046 14150 26052 14182
rect 25976 13534 26052 14150
rect 25976 13470 25982 13534
rect 26046 13470 26052 13534
rect 25976 13464 26052 13470
rect 16592 12142 16598 12174
rect 16597 12110 16598 12142
rect 16662 12142 16668 12174
rect 17952 13398 18028 13404
rect 17952 13334 17958 13398
rect 18022 13334 18028 13398
rect 16662 12110 16663 12142
rect 16597 12109 16663 12110
rect 16597 11902 16663 11903
rect 16597 11870 16598 11902
rect 11696 10886 11702 10950
rect 11766 10886 11772 10950
rect 11696 10880 11772 10886
rect 16592 11838 16598 11870
rect 16662 11870 16663 11902
rect 16662 11838 16668 11870
rect 11560 9422 11566 9454
rect 11565 9390 11566 9422
rect 11630 9422 11636 9454
rect 11696 10814 11772 10820
rect 11696 10750 11702 10814
rect 11766 10750 11772 10814
rect 11630 9390 11631 9422
rect 11565 9389 11631 9390
rect 952 8846 1230 8910
rect 1294 8846 1300 8910
rect 2448 9318 2524 9324
rect 2448 9254 2454 9318
rect 2518 9254 2524 9318
rect 2448 8910 2524 9254
rect 2448 8878 2454 8910
rect 952 7142 1300 8846
rect 2453 8846 2454 8878
rect 2518 8878 2524 8910
rect 2518 8846 2519 8878
rect 2453 8845 2519 8846
rect 2861 8638 2927 8639
rect 2861 8606 2862 8638
rect 2856 8574 2862 8606
rect 2926 8606 2927 8638
rect 2926 8574 2932 8606
rect 2856 8366 2932 8574
rect 2856 8302 2862 8366
rect 2926 8302 2932 8366
rect 2856 8296 2932 8302
rect 11696 8094 11772 10750
rect 16461 10542 16527 10543
rect 16461 10510 16462 10542
rect 11696 8062 11702 8094
rect 11701 8030 11702 8062
rect 11766 8062 11772 8094
rect 16456 10478 16462 10510
rect 16526 10510 16527 10542
rect 16526 10478 16532 10510
rect 11766 8030 11767 8062
rect 11701 8029 11767 8030
rect 16456 7822 16532 10478
rect 16592 9318 16668 11838
rect 17952 10678 18028 13334
rect 25976 13398 26052 13404
rect 25976 13334 25982 13398
rect 26046 13334 26052 13398
rect 25301 12990 25367 12991
rect 25301 12958 25302 12990
rect 25296 12926 25302 12958
rect 25366 12958 25367 12990
rect 25366 12926 25372 12958
rect 17952 10646 17958 10678
rect 17957 10614 17958 10646
rect 18022 10646 18028 10678
rect 25160 11222 25236 11228
rect 25160 11158 25166 11222
rect 25230 11158 25236 11222
rect 18022 10614 18023 10646
rect 17957 10613 18023 10614
rect 25160 9454 25236 11158
rect 25160 9422 25166 9454
rect 25165 9390 25166 9422
rect 25230 9422 25236 9454
rect 25230 9390 25231 9422
rect 25165 9389 25231 9390
rect 16592 9254 16598 9318
rect 16662 9254 16668 9318
rect 16592 9248 16668 9254
rect 16456 7758 16462 7822
rect 16526 7758 16532 7822
rect 16456 7752 16532 7758
rect 16592 9182 16668 9188
rect 16592 9118 16598 9182
rect 16662 9118 16668 9182
rect 952 7078 1230 7142
rect 1294 7078 1300 7142
rect 952 5374 1300 7078
rect 952 5310 1230 5374
rect 1294 5310 1300 5374
rect 952 3742 1300 5310
rect 16456 7686 16532 7692
rect 16456 7622 16462 7686
rect 16526 7622 16532 7686
rect 16456 4014 16532 7622
rect 16592 6462 16668 9118
rect 16592 6430 16598 6462
rect 16597 6398 16598 6430
rect 16662 6430 16668 6462
rect 16662 6398 16663 6430
rect 16597 6397 16663 6398
rect 16456 3982 16462 4014
rect 16461 3950 16462 3982
rect 16526 3982 16532 4014
rect 16526 3950 16527 3982
rect 16461 3949 16527 3950
rect 952 3678 1230 3742
rect 1294 3678 1300 3742
rect 25165 3742 25231 3743
rect 25165 3710 25166 3742
rect 952 1294 1300 3678
rect 25160 3678 25166 3710
rect 25230 3710 25231 3742
rect 25230 3678 25236 3710
rect 12925 2926 12991 2927
rect 12925 2894 12926 2926
rect 12920 2862 12926 2894
rect 12990 2894 12991 2926
rect 14285 2926 14351 2927
rect 14285 2894 14286 2926
rect 12990 2862 12996 2894
rect 1909 2110 1975 2111
rect 1909 2078 1910 2110
rect 1904 2046 1910 2078
rect 1974 2078 1975 2110
rect 1974 2046 1980 2078
rect 1904 1838 1980 2046
rect 1904 1774 1910 1838
rect 1974 1774 1980 1838
rect 1904 1768 1980 1774
rect 1909 1702 1975 1703
rect 1909 1670 1910 1702
rect 952 1230 958 1294
rect 1022 1230 1094 1294
rect 1158 1230 1230 1294
rect 1294 1230 1300 1294
rect 952 1158 1300 1230
rect 1904 1638 1910 1670
rect 1974 1670 1975 1702
rect 3677 1702 3743 1703
rect 3677 1670 3678 1702
rect 1974 1638 1980 1670
rect 1904 1294 1980 1638
rect 1904 1230 1910 1294
rect 1974 1230 1980 1294
rect 1904 1224 1980 1230
rect 3672 1638 3678 1670
rect 3742 1670 3743 1702
rect 5309 1702 5375 1703
rect 5309 1670 5310 1702
rect 3742 1638 3748 1670
rect 3672 1294 3748 1638
rect 3672 1230 3678 1294
rect 3742 1230 3748 1294
rect 3672 1224 3748 1230
rect 5304 1638 5310 1670
rect 5374 1670 5375 1702
rect 7077 1702 7143 1703
rect 7077 1670 7078 1702
rect 5374 1638 5380 1670
rect 5304 1294 5380 1638
rect 5304 1230 5310 1294
rect 5374 1230 5380 1294
rect 5304 1224 5380 1230
rect 7072 1638 7078 1670
rect 7142 1670 7143 1702
rect 8845 1702 8911 1703
rect 8845 1670 8846 1702
rect 7142 1638 7148 1670
rect 7072 1294 7148 1638
rect 7072 1230 7078 1294
rect 7142 1230 7148 1294
rect 7072 1224 7148 1230
rect 8840 1638 8846 1670
rect 8910 1670 8911 1702
rect 10341 1702 10407 1703
rect 10341 1670 10342 1702
rect 8910 1638 8916 1670
rect 8840 1294 8916 1638
rect 8840 1230 8846 1294
rect 8910 1230 8916 1294
rect 8840 1224 8916 1230
rect 10336 1638 10342 1670
rect 10406 1670 10407 1702
rect 12109 1702 12175 1703
rect 12109 1670 12110 1702
rect 10406 1638 10412 1670
rect 10336 1294 10412 1638
rect 10336 1230 10342 1294
rect 10406 1230 10412 1294
rect 10336 1224 10412 1230
rect 12104 1638 12110 1670
rect 12174 1670 12175 1702
rect 12174 1638 12180 1670
rect 12104 1294 12180 1638
rect 12104 1230 12110 1294
rect 12174 1230 12180 1294
rect 12104 1224 12180 1230
rect 952 1094 958 1158
rect 1022 1094 1094 1158
rect 1158 1094 1230 1158
rect 1294 1094 1300 1158
rect 952 1022 1300 1094
rect 952 958 958 1022
rect 1022 958 1094 1022
rect 1158 958 1230 1022
rect 1294 958 1300 1022
rect 952 952 1300 958
rect 272 550 278 614
rect 342 550 414 614
rect 478 550 550 614
rect 614 550 620 614
rect 272 478 620 550
rect 272 414 278 478
rect 342 414 414 478
rect 478 414 550 478
rect 614 414 620 478
rect 272 342 620 414
rect 272 278 278 342
rect 342 278 414 342
rect 478 278 550 342
rect 614 278 620 342
rect 272 272 620 278
rect 12920 0 12996 2862
rect 14280 2862 14286 2894
rect 14350 2894 14351 2926
rect 15373 2926 15439 2927
rect 15373 2894 15374 2926
rect 14350 2862 14356 2894
rect 13333 2382 13399 2383
rect 13333 2350 13334 2382
rect 13328 2318 13334 2350
rect 13398 2350 13399 2382
rect 13398 2318 13404 2350
rect 13328 614 13404 2318
rect 13877 1702 13943 1703
rect 13877 1670 13878 1702
rect 13872 1638 13878 1670
rect 13942 1670 13943 1702
rect 13942 1638 13948 1670
rect 13872 1294 13948 1638
rect 13872 1230 13878 1294
rect 13942 1230 13948 1294
rect 13872 1224 13948 1230
rect 13328 550 13334 614
rect 13398 550 13404 614
rect 13328 544 13404 550
rect 14280 0 14356 2862
rect 15368 2862 15374 2894
rect 15438 2894 15439 2926
rect 16461 2926 16527 2927
rect 16461 2894 16462 2926
rect 15438 2862 15444 2894
rect 15368 0 15444 2862
rect 16456 2862 16462 2894
rect 16526 2894 16527 2926
rect 17685 2926 17751 2927
rect 17685 2894 17686 2926
rect 16526 2862 16532 2894
rect 15509 1702 15575 1703
rect 15509 1670 15510 1702
rect 15504 1638 15510 1670
rect 15574 1670 15575 1702
rect 15574 1638 15580 1670
rect 15504 1294 15580 1638
rect 15504 1230 15510 1294
rect 15574 1230 15580 1294
rect 15504 1224 15580 1230
rect 16456 0 16532 2862
rect 17680 2862 17686 2894
rect 17750 2894 17751 2926
rect 18909 2926 18975 2927
rect 18909 2894 18910 2926
rect 17750 2862 17756 2894
rect 17141 1702 17207 1703
rect 17141 1670 17142 1702
rect 17136 1638 17142 1670
rect 17206 1670 17207 1702
rect 17206 1638 17212 1670
rect 17136 1294 17212 1638
rect 17136 1230 17142 1294
rect 17206 1230 17212 1294
rect 17136 1224 17212 1230
rect 17680 0 17756 2862
rect 18904 2862 18910 2894
rect 18974 2894 18975 2926
rect 19997 2926 20063 2927
rect 19997 2894 19998 2926
rect 18974 2862 18980 2894
rect 18773 1702 18839 1703
rect 18773 1670 18774 1702
rect 18768 1638 18774 1670
rect 18838 1670 18839 1702
rect 18838 1638 18844 1670
rect 18768 1294 18844 1638
rect 18768 1230 18774 1294
rect 18838 1230 18844 1294
rect 18768 1224 18844 1230
rect 18904 0 18980 2862
rect 19992 2862 19998 2894
rect 20062 2894 20063 2926
rect 21085 2926 21151 2927
rect 21085 2894 21086 2926
rect 20062 2862 20068 2894
rect 19992 0 20068 2862
rect 21080 2862 21086 2894
rect 21150 2894 21151 2926
rect 22309 2926 22375 2927
rect 22309 2894 22310 2926
rect 21150 2862 21156 2894
rect 20405 1702 20471 1703
rect 20405 1670 20406 1702
rect 20400 1638 20406 1670
rect 20470 1670 20471 1702
rect 20470 1638 20476 1670
rect 20400 1294 20476 1638
rect 20400 1230 20406 1294
rect 20470 1230 20476 1294
rect 20400 1224 20476 1230
rect 21080 0 21156 2862
rect 22304 2862 22310 2894
rect 22374 2894 22375 2926
rect 23397 2926 23463 2927
rect 23397 2894 23398 2926
rect 22374 2862 22380 2894
rect 22173 1702 22239 1703
rect 22173 1670 22174 1702
rect 22168 1638 22174 1670
rect 22238 1670 22239 1702
rect 22238 1638 22244 1670
rect 22168 1294 22244 1638
rect 22168 1230 22174 1294
rect 22238 1230 22244 1294
rect 22168 1224 22244 1230
rect 22304 0 22380 2862
rect 23392 2862 23398 2894
rect 23462 2894 23463 2926
rect 24757 2926 24823 2927
rect 24757 2894 24758 2926
rect 23462 2862 23468 2894
rect 23392 0 23468 2862
rect 24752 2862 24758 2894
rect 24822 2894 24823 2926
rect 24822 2862 24828 2894
rect 23805 1702 23871 1703
rect 23805 1670 23806 1702
rect 23800 1638 23806 1670
rect 23870 1670 23871 1702
rect 23870 1638 23876 1670
rect 23800 1294 23876 1638
rect 23800 1230 23806 1294
rect 23870 1230 23876 1294
rect 23800 1224 23876 1230
rect 24752 0 24828 2862
rect 25160 1838 25236 3678
rect 25160 1774 25166 1838
rect 25230 1774 25236 1838
rect 25160 1768 25236 1774
rect 25296 0 25372 12926
rect 25840 12854 25916 12860
rect 25840 12790 25846 12854
rect 25910 12790 25916 12854
rect 25840 12446 25916 12790
rect 25840 12414 25846 12446
rect 25845 12382 25846 12414
rect 25910 12414 25916 12446
rect 25910 12382 25911 12414
rect 25845 12381 25911 12382
rect 25845 12310 25911 12311
rect 25845 12278 25846 12310
rect 25840 12246 25846 12278
rect 25910 12278 25911 12310
rect 25910 12246 25916 12278
rect 25709 11766 25775 11767
rect 25709 11734 25710 11766
rect 25704 11702 25710 11734
rect 25774 11734 25775 11766
rect 25774 11702 25780 11734
rect 25568 10950 25644 10956
rect 25568 10886 25574 10950
rect 25638 10886 25644 10950
rect 25568 10542 25644 10886
rect 25704 10950 25780 11702
rect 25840 11630 25916 12246
rect 25976 11902 26052 13334
rect 26112 13262 26188 14966
rect 26792 14350 26868 18910
rect 26792 14318 26798 14350
rect 26797 14286 26798 14318
rect 26862 14318 26868 14350
rect 30736 18910 30742 18942
rect 30806 18942 30807 18974
rect 36448 18974 36524 18980
rect 30806 18910 30812 18942
rect 30736 14350 30812 18910
rect 36448 18910 36454 18974
rect 36518 18910 36524 18974
rect 31144 17478 31220 17484
rect 31144 17414 31150 17478
rect 31214 17414 31220 17478
rect 26862 14286 26863 14318
rect 26797 14285 26863 14286
rect 30736 14286 30742 14350
rect 30806 14286 30812 14350
rect 30736 14280 30812 14286
rect 31008 15030 31084 15036
rect 31008 14966 31014 15030
rect 31078 14966 31084 15030
rect 31144 15030 31220 17414
rect 36176 17478 36252 17484
rect 36176 17414 36182 17478
rect 36246 17414 36252 17478
rect 31144 14998 31150 15030
rect 30741 14214 30807 14215
rect 30741 14182 30742 14214
rect 30736 14150 30742 14182
rect 30806 14182 30807 14214
rect 30806 14150 30812 14182
rect 30736 13534 30812 14150
rect 30736 13470 30742 13534
rect 30806 13470 30812 13534
rect 30736 13464 30812 13470
rect 26112 13230 26118 13262
rect 26117 13198 26118 13230
rect 26182 13230 26188 13262
rect 30872 13398 30948 13404
rect 30872 13334 30878 13398
rect 30942 13334 30948 13398
rect 26182 13198 26183 13230
rect 26117 13197 26183 13198
rect 30469 12990 30535 12991
rect 30469 12958 30470 12990
rect 25976 11870 25982 11902
rect 25981 11838 25982 11870
rect 26046 11870 26052 11902
rect 30464 12926 30470 12958
rect 30534 12958 30535 12990
rect 30534 12926 30540 12958
rect 26046 11838 26047 11870
rect 25981 11837 26047 11838
rect 25840 11566 25846 11630
rect 25910 11566 25916 11630
rect 25840 11560 25916 11566
rect 25704 10886 25710 10950
rect 25774 10886 25780 10950
rect 25704 10880 25780 10886
rect 25568 10510 25574 10542
rect 25573 10478 25574 10510
rect 25638 10510 25644 10542
rect 25638 10478 25639 10510
rect 25573 10477 25639 10478
rect 25709 2926 25775 2927
rect 25709 2894 25710 2926
rect 25704 2862 25710 2894
rect 25774 2894 25775 2926
rect 25774 2862 25780 2894
rect 25573 1702 25639 1703
rect 25573 1670 25574 1702
rect 25568 1638 25574 1670
rect 25638 1670 25639 1702
rect 25638 1638 25644 1670
rect 25568 1294 25644 1638
rect 25568 1230 25574 1294
rect 25638 1230 25644 1294
rect 25568 1224 25644 1230
rect 25704 0 25780 2862
rect 27341 1702 27407 1703
rect 27341 1670 27342 1702
rect 27336 1638 27342 1670
rect 27406 1670 27407 1702
rect 28837 1702 28903 1703
rect 28837 1670 28838 1702
rect 27406 1638 27412 1670
rect 27336 1294 27412 1638
rect 27336 1230 27342 1294
rect 27406 1230 27412 1294
rect 27336 1224 27412 1230
rect 28832 1638 28838 1670
rect 28902 1670 28903 1702
rect 28902 1638 28908 1670
rect 28832 1294 28908 1638
rect 28832 1230 28838 1294
rect 28902 1230 28908 1294
rect 28832 1224 28908 1230
rect 30464 0 30540 12926
rect 30741 12310 30807 12311
rect 30741 12278 30742 12310
rect 30736 12246 30742 12278
rect 30806 12278 30807 12310
rect 30806 12246 30812 12278
rect 30736 11630 30812 12246
rect 30872 11902 30948 13334
rect 31008 13262 31084 14966
rect 31149 14966 31150 14998
rect 31214 14998 31220 15030
rect 36040 15030 36116 15036
rect 31214 14966 31215 14998
rect 31149 14965 31215 14966
rect 36040 14966 36046 15030
rect 36110 14966 36116 15030
rect 36176 15030 36252 17414
rect 36176 14998 36182 15030
rect 35773 14214 35839 14215
rect 35773 14182 35774 14214
rect 35768 14150 35774 14182
rect 35838 14182 35839 14214
rect 35838 14150 35844 14182
rect 35768 13534 35844 14150
rect 35768 13470 35774 13534
rect 35838 13470 35844 13534
rect 35768 13464 35844 13470
rect 31008 13230 31014 13262
rect 31013 13198 31014 13230
rect 31078 13230 31084 13262
rect 35904 13398 35980 13404
rect 35904 13334 35910 13398
rect 35974 13334 35980 13398
rect 31078 13198 31079 13230
rect 31013 13197 31079 13198
rect 31008 12990 31084 12996
rect 31008 12926 31014 12990
rect 31078 12926 31084 12990
rect 35501 12990 35567 12991
rect 35501 12958 35502 12990
rect 31008 12446 31084 12926
rect 31008 12414 31014 12446
rect 31013 12382 31014 12414
rect 31078 12414 31084 12446
rect 35496 12926 35502 12958
rect 35566 12958 35567 12990
rect 35566 12926 35572 12958
rect 31078 12382 31079 12414
rect 31013 12381 31079 12382
rect 30872 11870 30878 11902
rect 30877 11838 30878 11870
rect 30942 11870 30948 11902
rect 30942 11838 30943 11870
rect 30877 11837 30943 11838
rect 30877 11766 30943 11767
rect 30877 11734 30878 11766
rect 30736 11566 30742 11630
rect 30806 11566 30812 11630
rect 30736 11560 30812 11566
rect 30872 11702 30878 11734
rect 30942 11734 30943 11766
rect 30942 11702 30948 11734
rect 30872 10950 30948 11702
rect 30872 10886 30878 10950
rect 30942 10886 30948 10950
rect 30872 10880 30948 10886
rect 30741 1702 30807 1703
rect 30741 1670 30742 1702
rect 30736 1638 30742 1670
rect 30806 1670 30807 1702
rect 32373 1702 32439 1703
rect 32373 1670 32374 1702
rect 30806 1638 30812 1670
rect 30736 1294 30812 1638
rect 30736 1230 30742 1294
rect 30806 1230 30812 1294
rect 30736 1224 30812 1230
rect 32368 1638 32374 1670
rect 32438 1670 32439 1702
rect 33869 1702 33935 1703
rect 33869 1670 33870 1702
rect 32438 1638 32444 1670
rect 32368 1294 32444 1638
rect 32368 1230 32374 1294
rect 32438 1230 32444 1294
rect 32368 1224 32444 1230
rect 33864 1638 33870 1670
rect 33934 1670 33935 1702
rect 33934 1638 33940 1670
rect 33864 1294 33940 1638
rect 33864 1230 33870 1294
rect 33934 1230 33940 1294
rect 33864 1224 33940 1230
rect 35496 0 35572 12926
rect 35768 12854 35844 12860
rect 35768 12790 35774 12854
rect 35838 12790 35844 12854
rect 35768 12446 35844 12790
rect 35768 12414 35774 12446
rect 35773 12382 35774 12414
rect 35838 12414 35844 12446
rect 35838 12382 35839 12414
rect 35773 12381 35839 12382
rect 35637 12310 35703 12311
rect 35637 12278 35638 12310
rect 35632 12246 35638 12278
rect 35702 12278 35703 12310
rect 35702 12246 35708 12278
rect 35632 11630 35708 12246
rect 35904 11902 35980 13334
rect 36040 13262 36116 14966
rect 36181 14966 36182 14998
rect 36246 14998 36252 15030
rect 36246 14966 36247 14998
rect 36181 14965 36247 14966
rect 36448 14350 36524 18910
rect 41480 18974 41556 18980
rect 41480 18910 41486 18974
rect 41550 18910 41556 18974
rect 45701 18974 45767 18975
rect 45701 18942 45702 18974
rect 40936 17478 41012 17484
rect 40936 17414 40942 17478
rect 41006 17414 41012 17478
rect 40936 15030 41012 17414
rect 40936 14998 40942 15030
rect 40941 14966 40942 14998
rect 41006 14998 41012 15030
rect 41072 15030 41148 15036
rect 41006 14966 41007 14998
rect 40941 14965 41007 14966
rect 41072 14966 41078 15030
rect 41142 14966 41148 15030
rect 36448 14318 36454 14350
rect 36453 14286 36454 14318
rect 36518 14318 36524 14350
rect 36518 14286 36519 14318
rect 36453 14285 36519 14286
rect 40941 14214 41007 14215
rect 40941 14182 40942 14214
rect 40936 14150 40942 14182
rect 41006 14182 41007 14214
rect 41006 14150 41012 14182
rect 40936 13534 41012 14150
rect 40936 13470 40942 13534
rect 41006 13470 41012 13534
rect 40936 13464 41012 13470
rect 36040 13230 36046 13262
rect 36045 13198 36046 13230
rect 36110 13230 36116 13262
rect 40936 13398 41012 13404
rect 40936 13334 40942 13398
rect 41006 13334 41012 13398
rect 36110 13198 36111 13230
rect 36045 13197 36111 13198
rect 40533 12990 40599 12991
rect 40533 12958 40534 12990
rect 35904 11870 35910 11902
rect 35909 11838 35910 11870
rect 35974 11870 35980 11902
rect 40528 12926 40534 12958
rect 40598 12958 40599 12990
rect 40598 12926 40604 12958
rect 35974 11838 35975 11870
rect 35909 11837 35975 11838
rect 35773 11766 35839 11767
rect 35773 11734 35774 11766
rect 35632 11566 35638 11630
rect 35702 11566 35708 11630
rect 35632 11560 35708 11566
rect 35768 11702 35774 11734
rect 35838 11734 35839 11766
rect 35838 11702 35844 11734
rect 35768 10950 35844 11702
rect 35768 10886 35774 10950
rect 35838 10886 35844 10950
rect 35768 10880 35844 10886
rect 35637 1702 35703 1703
rect 35637 1670 35638 1702
rect 35632 1638 35638 1670
rect 35702 1670 35703 1702
rect 37405 1702 37471 1703
rect 37405 1670 37406 1702
rect 35702 1638 35708 1670
rect 35632 1294 35708 1638
rect 35632 1230 35638 1294
rect 35702 1230 35708 1294
rect 35632 1224 35708 1230
rect 37400 1638 37406 1670
rect 37470 1670 37471 1702
rect 38901 1702 38967 1703
rect 38901 1670 38902 1702
rect 37470 1638 37476 1670
rect 37400 1294 37476 1638
rect 37400 1230 37406 1294
rect 37470 1230 37476 1294
rect 37400 1224 37476 1230
rect 38896 1638 38902 1670
rect 38966 1670 38967 1702
rect 38966 1638 38972 1670
rect 38896 1294 38972 1638
rect 38896 1230 38902 1294
rect 38966 1230 38972 1294
rect 38896 1224 38972 1230
rect 40528 0 40604 12926
rect 40800 12854 40876 12860
rect 40800 12790 40806 12854
rect 40870 12790 40876 12854
rect 40800 12446 40876 12790
rect 40800 12414 40806 12446
rect 40805 12382 40806 12414
rect 40870 12414 40876 12446
rect 40870 12382 40871 12414
rect 40805 12381 40871 12382
rect 40936 11902 41012 13334
rect 41072 13262 41148 14966
rect 41480 14350 41556 18910
rect 41480 14318 41486 14350
rect 41485 14286 41486 14318
rect 41550 14318 41556 14350
rect 45696 18910 45702 18942
rect 45766 18942 45767 18974
rect 51408 18974 51484 18980
rect 45766 18910 45772 18942
rect 45696 14350 45772 18910
rect 51408 18910 51414 18974
rect 51478 18910 51484 18974
rect 55765 18974 55831 18975
rect 55765 18942 55766 18974
rect 45968 17478 46044 17484
rect 45968 17414 45974 17478
rect 46038 17414 46044 17478
rect 41550 14286 41551 14318
rect 41485 14285 41551 14286
rect 45696 14286 45702 14350
rect 45766 14286 45772 14350
rect 45696 14280 45772 14286
rect 45832 15030 45908 15036
rect 45832 14966 45838 15030
rect 45902 14966 45908 15030
rect 45968 15030 46044 17414
rect 51136 17478 51212 17484
rect 51136 17414 51142 17478
rect 51206 17414 51212 17478
rect 45968 14998 45974 15030
rect 41072 13230 41078 13262
rect 41077 13198 41078 13230
rect 41142 13230 41148 13262
rect 45696 13398 45772 13404
rect 45696 13334 45702 13398
rect 45766 13334 45772 13398
rect 41142 13198 41143 13230
rect 41077 13197 41143 13198
rect 45565 12990 45631 12991
rect 45565 12958 45566 12990
rect 45560 12926 45566 12958
rect 45630 12958 45631 12990
rect 45630 12926 45636 12958
rect 41077 12310 41143 12311
rect 41077 12278 41078 12310
rect 40936 11870 40942 11902
rect 40941 11838 40942 11870
rect 41006 11870 41012 11902
rect 41072 12246 41078 12278
rect 41142 12278 41143 12310
rect 41142 12246 41148 12278
rect 41006 11838 41007 11870
rect 40941 11837 41007 11838
rect 40805 11766 40871 11767
rect 40805 11734 40806 11766
rect 40800 11702 40806 11734
rect 40870 11734 40871 11766
rect 40870 11702 40876 11734
rect 40800 10950 40876 11702
rect 41072 11630 41148 12246
rect 41072 11566 41078 11630
rect 41142 11566 41148 11630
rect 41072 11560 41148 11566
rect 40800 10886 40806 10950
rect 40870 10886 40876 10950
rect 40800 10880 40876 10886
rect 40805 1702 40871 1703
rect 40805 1670 40806 1702
rect 40800 1638 40806 1670
rect 40870 1670 40871 1702
rect 42301 1702 42367 1703
rect 42301 1670 42302 1702
rect 40870 1638 40876 1670
rect 40800 1294 40876 1638
rect 40800 1230 40806 1294
rect 40870 1230 40876 1294
rect 40800 1224 40876 1230
rect 42296 1638 42302 1670
rect 42366 1670 42367 1702
rect 43933 1702 43999 1703
rect 43933 1670 43934 1702
rect 42366 1638 42372 1670
rect 42296 1294 42372 1638
rect 42296 1230 42302 1294
rect 42366 1230 42372 1294
rect 42296 1224 42372 1230
rect 43928 1638 43934 1670
rect 43998 1670 43999 1702
rect 43998 1638 44004 1670
rect 43928 1294 44004 1638
rect 43928 1230 43934 1294
rect 43998 1230 44004 1294
rect 43928 1224 44004 1230
rect 45560 0 45636 12926
rect 45696 11902 45772 13334
rect 45832 13262 45908 14966
rect 45973 14966 45974 14998
rect 46038 14998 46044 15030
rect 51000 15030 51076 15036
rect 46038 14966 46039 14998
rect 45973 14965 46039 14966
rect 51000 14966 51006 15030
rect 51070 14966 51076 15030
rect 51136 15030 51212 17414
rect 51136 14998 51142 15030
rect 45973 14214 46039 14215
rect 45973 14182 45974 14214
rect 45968 14150 45974 14182
rect 46038 14182 46039 14214
rect 50733 14214 50799 14215
rect 50733 14182 50734 14214
rect 46038 14150 46044 14182
rect 45968 13534 46044 14150
rect 45968 13470 45974 13534
rect 46038 13470 46044 13534
rect 45968 13464 46044 13470
rect 50728 14150 50734 14182
rect 50798 14182 50799 14214
rect 50798 14150 50804 14182
rect 50728 13534 50804 14150
rect 50728 13470 50734 13534
rect 50798 13470 50804 13534
rect 50728 13464 50804 13470
rect 45832 13230 45838 13262
rect 45837 13198 45838 13230
rect 45902 13230 45908 13262
rect 50864 13398 50940 13404
rect 50864 13334 50870 13398
rect 50934 13334 50940 13398
rect 45902 13198 45903 13230
rect 45837 13197 45903 13198
rect 45832 12990 45908 12996
rect 45832 12926 45838 12990
rect 45902 12926 45908 12990
rect 50461 12990 50527 12991
rect 50461 12958 50462 12990
rect 45832 12446 45908 12926
rect 45832 12414 45838 12446
rect 45837 12382 45838 12414
rect 45902 12414 45908 12446
rect 50456 12926 50462 12958
rect 50526 12958 50527 12990
rect 50526 12926 50532 12958
rect 45902 12382 45903 12414
rect 45837 12381 45903 12382
rect 45837 12310 45903 12311
rect 45837 12278 45838 12310
rect 45696 11870 45702 11902
rect 45701 11838 45702 11870
rect 45766 11870 45772 11902
rect 45832 12246 45838 12278
rect 45902 12278 45903 12310
rect 45902 12246 45908 12278
rect 45766 11838 45767 11870
rect 45701 11837 45767 11838
rect 45701 11766 45767 11767
rect 45701 11734 45702 11766
rect 45696 11702 45702 11734
rect 45766 11734 45767 11766
rect 45766 11702 45772 11734
rect 45696 10950 45772 11702
rect 45832 11630 45908 12246
rect 45832 11566 45838 11630
rect 45902 11566 45908 11630
rect 45832 11560 45908 11566
rect 45696 10886 45702 10950
rect 45766 10886 45772 10950
rect 45696 10880 45772 10886
rect 45837 1702 45903 1703
rect 45837 1670 45838 1702
rect 45832 1638 45838 1670
rect 45902 1670 45903 1702
rect 47333 1702 47399 1703
rect 47333 1670 47334 1702
rect 45902 1638 45908 1670
rect 45832 1294 45908 1638
rect 45832 1230 45838 1294
rect 45902 1230 45908 1294
rect 45832 1224 45908 1230
rect 47328 1638 47334 1670
rect 47398 1670 47399 1702
rect 49101 1702 49167 1703
rect 49101 1670 49102 1702
rect 47398 1638 47404 1670
rect 47328 1294 47404 1638
rect 47328 1230 47334 1294
rect 47398 1230 47404 1294
rect 47328 1224 47404 1230
rect 49096 1638 49102 1670
rect 49166 1670 49167 1702
rect 49166 1638 49172 1670
rect 49096 1294 49172 1638
rect 49096 1230 49102 1294
rect 49166 1230 49172 1294
rect 49096 1224 49172 1230
rect 50456 0 50532 12926
rect 50728 12854 50804 12860
rect 50728 12790 50734 12854
rect 50798 12790 50804 12854
rect 50728 12446 50804 12790
rect 50728 12414 50734 12446
rect 50733 12382 50734 12414
rect 50798 12414 50804 12446
rect 50798 12382 50799 12414
rect 50733 12381 50799 12382
rect 50864 11902 50940 13334
rect 51000 13262 51076 14966
rect 51141 14966 51142 14998
rect 51206 14998 51212 15030
rect 51206 14966 51207 14998
rect 51141 14965 51207 14966
rect 51408 14350 51484 18910
rect 51408 14318 51414 14350
rect 51413 14286 51414 14318
rect 51478 14318 51484 14350
rect 55760 18910 55766 18942
rect 55830 18942 55831 18974
rect 61472 18974 61548 18980
rect 55830 18910 55836 18942
rect 55760 14350 55836 18910
rect 61472 18910 61478 18974
rect 61542 18910 61548 18974
rect 56168 17478 56244 17484
rect 56168 17414 56174 17478
rect 56238 17414 56244 17478
rect 51478 14286 51479 14318
rect 51413 14285 51479 14286
rect 55760 14286 55766 14350
rect 55830 14286 55836 14350
rect 55760 14280 55836 14286
rect 56032 15030 56108 15036
rect 56032 14966 56038 15030
rect 56102 14966 56108 15030
rect 56168 15030 56244 17414
rect 56168 14998 56174 15030
rect 55765 14214 55831 14215
rect 55765 14182 55766 14214
rect 55760 14150 55766 14182
rect 55830 14182 55831 14214
rect 55830 14150 55836 14182
rect 55760 13534 55836 14150
rect 55760 13470 55766 13534
rect 55830 13470 55836 13534
rect 55760 13464 55836 13470
rect 51000 13230 51006 13262
rect 51005 13198 51006 13230
rect 51070 13230 51076 13262
rect 55896 13398 55972 13404
rect 55896 13334 55902 13398
rect 55966 13334 55972 13398
rect 51070 13198 51071 13230
rect 51005 13197 51071 13198
rect 55493 12990 55559 12991
rect 55493 12958 55494 12990
rect 55488 12926 55494 12958
rect 55558 12958 55559 12990
rect 55558 12926 55564 12958
rect 51005 12310 51071 12311
rect 51005 12278 51006 12310
rect 50864 11870 50870 11902
rect 50869 11838 50870 11870
rect 50934 11870 50940 11902
rect 51000 12246 51006 12278
rect 51070 12278 51071 12310
rect 51070 12246 51076 12278
rect 50934 11838 50935 11870
rect 50869 11837 50935 11838
rect 50733 11766 50799 11767
rect 50733 11734 50734 11766
rect 50728 11702 50734 11734
rect 50798 11734 50799 11766
rect 50798 11702 50804 11734
rect 50728 10950 50804 11702
rect 51000 11630 51076 12246
rect 51000 11566 51006 11630
rect 51070 11566 51076 11630
rect 51000 11560 51076 11566
rect 50728 10886 50734 10950
rect 50798 10886 50804 10950
rect 50728 10880 50804 10886
rect 50869 1702 50935 1703
rect 50869 1670 50870 1702
rect 50864 1638 50870 1670
rect 50934 1670 50935 1702
rect 52365 1702 52431 1703
rect 52365 1670 52366 1702
rect 50934 1638 50940 1670
rect 50864 1294 50940 1638
rect 50864 1230 50870 1294
rect 50934 1230 50940 1294
rect 50864 1224 50940 1230
rect 52360 1638 52366 1670
rect 52430 1670 52431 1702
rect 54133 1702 54199 1703
rect 54133 1670 54134 1702
rect 52430 1638 52436 1670
rect 52360 1294 52436 1638
rect 52360 1230 52366 1294
rect 52430 1230 52436 1294
rect 52360 1224 52436 1230
rect 54128 1638 54134 1670
rect 54198 1670 54199 1702
rect 54198 1638 54204 1670
rect 54128 1294 54204 1638
rect 54128 1230 54134 1294
rect 54198 1230 54204 1294
rect 54128 1224 54204 1230
rect 55488 0 55564 12926
rect 55760 12854 55836 12860
rect 55760 12790 55766 12854
rect 55830 12790 55836 12854
rect 55760 12446 55836 12790
rect 55760 12414 55766 12446
rect 55765 12382 55766 12414
rect 55830 12414 55836 12446
rect 55830 12382 55831 12414
rect 55765 12381 55831 12382
rect 55896 11902 55972 13334
rect 56032 13262 56108 14966
rect 56173 14966 56174 14998
rect 56238 14998 56244 15030
rect 60928 17478 61004 17484
rect 60928 17414 60934 17478
rect 60998 17414 61004 17478
rect 60928 15030 61004 17414
rect 60928 14998 60934 15030
rect 56238 14966 56239 14998
rect 56173 14965 56239 14966
rect 60933 14966 60934 14998
rect 60998 14998 61004 15030
rect 61064 15030 61140 15036
rect 60998 14966 60999 14998
rect 60933 14965 60999 14966
rect 61064 14966 61070 15030
rect 61134 14966 61140 15030
rect 60797 14214 60863 14215
rect 60797 14182 60798 14214
rect 60792 14150 60798 14182
rect 60862 14182 60863 14214
rect 60862 14150 60868 14182
rect 60792 13534 60868 14150
rect 60792 13470 60798 13534
rect 60862 13470 60868 13534
rect 60792 13464 60868 13470
rect 56032 13230 56038 13262
rect 56037 13198 56038 13230
rect 56102 13230 56108 13262
rect 60928 13398 61004 13404
rect 60928 13334 60934 13398
rect 60998 13334 61004 13398
rect 56102 13198 56103 13230
rect 56037 13197 56103 13198
rect 60525 12990 60591 12991
rect 60525 12958 60526 12990
rect 60520 12926 60526 12958
rect 60590 12958 60591 12990
rect 60590 12926 60596 12958
rect 56037 12310 56103 12311
rect 56037 12278 56038 12310
rect 55896 11870 55902 11902
rect 55901 11838 55902 11870
rect 55966 11870 55972 11902
rect 56032 12246 56038 12278
rect 56102 12278 56103 12310
rect 56102 12246 56108 12278
rect 55966 11838 55967 11870
rect 55901 11837 55967 11838
rect 55765 11766 55831 11767
rect 55765 11734 55766 11766
rect 55760 11702 55766 11734
rect 55830 11734 55831 11766
rect 55830 11702 55836 11734
rect 55760 10950 55836 11702
rect 56032 11630 56108 12246
rect 56032 11566 56038 11630
rect 56102 11566 56108 11630
rect 56032 11560 56108 11566
rect 55760 10886 55766 10950
rect 55830 10886 55836 10950
rect 55760 10880 55836 10886
rect 55901 1702 55967 1703
rect 55901 1670 55902 1702
rect 55896 1638 55902 1670
rect 55966 1670 55967 1702
rect 57397 1702 57463 1703
rect 57397 1670 57398 1702
rect 55966 1638 55972 1670
rect 55896 1294 55972 1638
rect 55896 1230 55902 1294
rect 55966 1230 55972 1294
rect 55896 1224 55972 1230
rect 57392 1638 57398 1670
rect 57462 1670 57463 1702
rect 59301 1702 59367 1703
rect 59301 1670 59302 1702
rect 57462 1638 57468 1670
rect 57392 1294 57468 1638
rect 57392 1230 57398 1294
rect 57462 1230 57468 1294
rect 57392 1224 57468 1230
rect 59296 1638 59302 1670
rect 59366 1670 59367 1702
rect 59366 1638 59372 1670
rect 59296 1294 59372 1638
rect 59296 1230 59302 1294
rect 59366 1230 59372 1294
rect 59296 1224 59372 1230
rect 60520 0 60596 12926
rect 60792 12854 60868 12860
rect 60792 12790 60798 12854
rect 60862 12790 60868 12854
rect 60792 12446 60868 12790
rect 60792 12414 60798 12446
rect 60797 12382 60798 12414
rect 60862 12414 60868 12446
rect 60862 12382 60863 12414
rect 60797 12381 60863 12382
rect 60661 12310 60727 12311
rect 60661 12278 60662 12310
rect 60656 12246 60662 12278
rect 60726 12278 60727 12310
rect 60726 12246 60732 12278
rect 60656 11630 60732 12246
rect 60928 11902 61004 13334
rect 61064 13262 61140 14966
rect 61472 14350 61548 18910
rect 66368 17614 66444 20134
rect 77112 18974 77188 20542
rect 79832 20542 79838 20574
rect 79902 20574 79903 20606
rect 89760 20606 90108 22174
rect 79902 20542 79908 20574
rect 79832 20334 79908 20542
rect 79832 20270 79838 20334
rect 79902 20270 79908 20334
rect 79832 20264 79908 20270
rect 89760 20542 89766 20606
rect 89830 20542 90108 20606
rect 79973 20198 80039 20199
rect 79973 20166 79974 20198
rect 77112 18910 77118 18974
rect 77182 18910 77188 18974
rect 77112 18904 77188 18910
rect 79968 20134 79974 20166
rect 80038 20166 80039 20198
rect 80038 20134 80044 20166
rect 79837 18702 79903 18703
rect 79837 18670 79838 18702
rect 66368 17582 66374 17614
rect 66373 17550 66374 17582
rect 66438 17582 66444 17614
rect 79832 18638 79838 18670
rect 79902 18670 79903 18702
rect 79902 18638 79908 18670
rect 66438 17550 66439 17582
rect 66373 17549 66439 17550
rect 79832 16118 79908 18638
rect 79968 17478 80044 20134
rect 79968 17414 79974 17478
rect 80038 17414 80044 17478
rect 79968 17408 80044 17414
rect 89760 18838 90108 20542
rect 89760 18774 89766 18838
rect 89830 18774 90108 18838
rect 79832 16054 79838 16118
rect 79902 16054 79908 16118
rect 79832 16048 79908 16054
rect 79968 17342 80044 17348
rect 79968 17278 79974 17342
rect 80038 17278 80044 17342
rect 61472 14318 61478 14350
rect 61477 14286 61478 14318
rect 61542 14318 61548 14350
rect 79832 15982 79908 15988
rect 79832 15918 79838 15982
rect 79902 15918 79908 15982
rect 61542 14286 61543 14318
rect 61477 14285 61543 14286
rect 61064 13230 61070 13262
rect 61069 13198 61070 13230
rect 61134 13230 61140 13262
rect 79832 13262 79908 15918
rect 79968 14622 80044 17278
rect 79968 14590 79974 14622
rect 79973 14558 79974 14590
rect 80038 14590 80044 14622
rect 89760 17206 90108 18774
rect 89760 17142 89766 17206
rect 89830 17142 90108 17206
rect 89760 15574 90108 17142
rect 89760 15510 89766 15574
rect 89830 15510 90108 15574
rect 80038 14558 80039 14590
rect 79973 14557 80039 14558
rect 79832 13230 79838 13262
rect 61134 13198 61135 13230
rect 61069 13197 61135 13198
rect 79837 13198 79838 13230
rect 79902 13230 79908 13262
rect 79968 14486 80044 14492
rect 79968 14422 79974 14486
rect 80038 14422 80044 14486
rect 79902 13198 79903 13230
rect 79837 13197 79903 13198
rect 79837 13126 79903 13127
rect 79837 13094 79838 13126
rect 60928 11870 60934 11902
rect 60933 11838 60934 11870
rect 60998 11870 61004 11902
rect 79832 13062 79838 13094
rect 79902 13094 79903 13126
rect 79902 13062 79908 13094
rect 60998 11838 60999 11870
rect 60933 11837 60999 11838
rect 60797 11766 60863 11767
rect 60797 11734 60798 11766
rect 60656 11566 60662 11630
rect 60726 11566 60732 11630
rect 60656 11560 60732 11566
rect 60792 11702 60798 11734
rect 60862 11734 60863 11766
rect 60862 11702 60868 11734
rect 60792 10950 60868 11702
rect 65421 11494 65487 11495
rect 65421 11462 65422 11494
rect 65416 11430 65422 11462
rect 65486 11462 65487 11494
rect 65486 11430 65492 11462
rect 60792 10886 60798 10950
rect 60862 10886 60868 10950
rect 65285 10950 65351 10951
rect 65285 10918 65286 10950
rect 60792 10880 60868 10886
rect 65280 10886 65286 10918
rect 65350 10918 65351 10950
rect 65350 10886 65356 10918
rect 65280 10542 65356 10886
rect 65280 10478 65286 10542
rect 65350 10478 65356 10542
rect 65280 10472 65356 10478
rect 65416 9454 65492 11430
rect 79832 10406 79908 13062
rect 79968 11902 80044 14422
rect 79968 11870 79974 11902
rect 79973 11838 79974 11870
rect 80038 11870 80044 11902
rect 89760 13942 90108 15510
rect 89760 13878 89766 13942
rect 89830 13878 90108 13942
rect 89760 12310 90108 13878
rect 89760 12246 89766 12310
rect 89830 12246 90108 12310
rect 80038 11838 80039 11870
rect 79973 11837 80039 11838
rect 79832 10342 79838 10406
rect 79902 10342 79908 10406
rect 79832 10336 79908 10342
rect 89760 10406 90108 12246
rect 89760 10342 89766 10406
rect 89830 10342 90108 10406
rect 65416 9390 65422 9454
rect 65486 9390 65492 9454
rect 65416 9384 65492 9390
rect 89760 8774 90108 10342
rect 89760 8710 89766 8774
rect 89830 8710 90108 8774
rect 89760 7278 90108 8710
rect 89760 7214 89766 7278
rect 89830 7214 90108 7278
rect 89760 5374 90108 7214
rect 89760 5310 89766 5374
rect 89830 5310 90108 5374
rect 89760 3742 90108 5310
rect 89760 3678 89766 3742
rect 89830 3678 90108 3742
rect 89760 2110 90108 3678
rect 89760 2046 89766 2110
rect 89830 2046 90108 2110
rect 60797 1702 60863 1703
rect 60797 1670 60798 1702
rect 60792 1638 60798 1670
rect 60862 1670 60863 1702
rect 62429 1702 62495 1703
rect 62429 1670 62430 1702
rect 60862 1638 60868 1670
rect 60792 1294 60868 1638
rect 60792 1230 60798 1294
rect 60862 1230 60868 1294
rect 60792 1224 60868 1230
rect 62424 1638 62430 1670
rect 62494 1670 62495 1702
rect 64333 1702 64399 1703
rect 64333 1670 64334 1702
rect 62494 1638 62500 1670
rect 62424 1294 62500 1638
rect 62424 1230 62430 1294
rect 62494 1230 62500 1294
rect 62424 1224 62500 1230
rect 64328 1638 64334 1670
rect 64398 1670 64399 1702
rect 65829 1702 65895 1703
rect 65829 1670 65830 1702
rect 64398 1638 64404 1670
rect 64328 1294 64404 1638
rect 64328 1230 64334 1294
rect 64398 1230 64404 1294
rect 64328 1224 64404 1230
rect 65824 1638 65830 1670
rect 65894 1670 65895 1702
rect 67597 1702 67663 1703
rect 67597 1670 67598 1702
rect 65894 1638 65900 1670
rect 65824 1294 65900 1638
rect 65824 1230 65830 1294
rect 65894 1230 65900 1294
rect 65824 1224 65900 1230
rect 67592 1638 67598 1670
rect 67662 1670 67663 1702
rect 69365 1702 69431 1703
rect 69365 1670 69366 1702
rect 67662 1638 67668 1670
rect 67592 1294 67668 1638
rect 67592 1230 67598 1294
rect 67662 1230 67668 1294
rect 67592 1224 67668 1230
rect 69360 1638 69366 1670
rect 69430 1670 69431 1702
rect 70861 1702 70927 1703
rect 70861 1670 70862 1702
rect 69430 1638 69436 1670
rect 69360 1294 69436 1638
rect 69360 1230 69366 1294
rect 69430 1230 69436 1294
rect 69360 1224 69436 1230
rect 70856 1638 70862 1670
rect 70926 1670 70927 1702
rect 72629 1702 72695 1703
rect 72629 1670 72630 1702
rect 70926 1638 70932 1670
rect 70856 1294 70932 1638
rect 70856 1230 70862 1294
rect 70926 1230 70932 1294
rect 70856 1224 70932 1230
rect 72624 1638 72630 1670
rect 72694 1670 72695 1702
rect 74397 1702 74463 1703
rect 74397 1670 74398 1702
rect 72694 1638 72700 1670
rect 72624 1294 72700 1638
rect 72624 1230 72630 1294
rect 72694 1230 72700 1294
rect 72624 1224 72700 1230
rect 74392 1638 74398 1670
rect 74462 1670 74463 1702
rect 75893 1702 75959 1703
rect 75893 1670 75894 1702
rect 74462 1638 74468 1670
rect 74392 1294 74468 1638
rect 74392 1230 74398 1294
rect 74462 1230 74468 1294
rect 74392 1224 74468 1230
rect 75888 1638 75894 1670
rect 75958 1670 75959 1702
rect 77661 1702 77727 1703
rect 77661 1670 77662 1702
rect 75958 1638 75964 1670
rect 75888 1294 75964 1638
rect 75888 1230 75894 1294
rect 75958 1230 75964 1294
rect 75888 1224 75964 1230
rect 77656 1638 77662 1670
rect 77726 1670 77727 1702
rect 79293 1702 79359 1703
rect 79293 1670 79294 1702
rect 77726 1638 77732 1670
rect 77656 1294 77732 1638
rect 77656 1230 77662 1294
rect 77726 1230 77732 1294
rect 77656 1224 77732 1230
rect 79288 1638 79294 1670
rect 79358 1670 79359 1702
rect 80925 1702 80991 1703
rect 80925 1670 80926 1702
rect 79358 1638 79364 1670
rect 79288 1294 79364 1638
rect 79288 1230 79294 1294
rect 79358 1230 79364 1294
rect 79288 1224 79364 1230
rect 80920 1638 80926 1670
rect 80990 1670 80991 1702
rect 82829 1702 82895 1703
rect 82829 1670 82830 1702
rect 80990 1638 80996 1670
rect 80920 1294 80996 1638
rect 80920 1230 80926 1294
rect 80990 1230 80996 1294
rect 80920 1224 80996 1230
rect 82824 1638 82830 1670
rect 82894 1670 82895 1702
rect 84325 1702 84391 1703
rect 84325 1670 84326 1702
rect 82894 1638 82900 1670
rect 82824 1294 82900 1638
rect 82824 1230 82830 1294
rect 82894 1230 82900 1294
rect 82824 1224 82900 1230
rect 84320 1638 84326 1670
rect 84390 1670 84391 1702
rect 86093 1702 86159 1703
rect 86093 1670 86094 1702
rect 84390 1638 84396 1670
rect 84320 1294 84396 1638
rect 84320 1230 84326 1294
rect 84390 1230 84396 1294
rect 84320 1224 84396 1230
rect 86088 1638 86094 1670
rect 86158 1670 86159 1702
rect 87589 1702 87655 1703
rect 87589 1670 87590 1702
rect 86158 1638 86164 1670
rect 86088 1294 86164 1638
rect 86088 1230 86094 1294
rect 86158 1230 86164 1294
rect 86088 1224 86164 1230
rect 87584 1638 87590 1670
rect 87654 1670 87655 1702
rect 87654 1638 87660 1670
rect 87584 1294 87660 1638
rect 87584 1230 87590 1294
rect 87654 1230 87660 1294
rect 87584 1224 87660 1230
rect 89760 1294 90108 2046
rect 89760 1230 89766 1294
rect 89830 1230 89902 1294
rect 89966 1230 90038 1294
rect 90102 1230 90108 1294
rect 89760 1158 90108 1230
rect 89760 1094 89766 1158
rect 89830 1094 89902 1158
rect 89966 1094 90038 1158
rect 90102 1094 90108 1158
rect 89760 1022 90108 1094
rect 89760 958 89766 1022
rect 89830 958 89902 1022
rect 89966 958 90038 1022
rect 90102 958 90108 1022
rect 89760 952 90108 958
rect 90440 80174 90788 88678
rect 90440 80110 90446 80174
rect 90510 80110 90788 80174
rect 90440 73238 90788 80110
rect 90440 73174 90446 73238
rect 90510 73174 90788 73238
rect 90440 70246 90788 73174
rect 90440 70182 90446 70246
rect 90510 70182 90788 70246
rect 90440 64534 90788 70182
rect 90440 64470 90446 64534
rect 90510 64470 90788 64534
rect 90440 614 90788 64470
rect 90440 550 90446 614
rect 90510 550 90582 614
rect 90646 550 90718 614
rect 90782 550 90788 614
rect 90440 478 90788 550
rect 90440 414 90446 478
rect 90510 414 90582 478
rect 90646 414 90718 478
rect 90782 414 90788 478
rect 90440 342 90788 414
rect 90440 278 90446 342
rect 90510 278 90582 342
rect 90646 278 90718 342
rect 90782 278 90788 342
rect 90440 272 90788 278
use sky130_sram_1kbyte_1rw1r_8x1024_8_bank  sky130_sram_1kbyte_1rw1r_8x1024_8_bank_0
timestamp 1704896540
transform 1 0 11870 0 1 6294
box 0 0 67334 78433
use sky130_sram_1kbyte_1rw1r_8x1024_8_col_addr_dff  sky130_sram_1kbyte_1rw1r_8x1024_8_col_addr_dff_0
timestamp 1704896540
transform 1 0 12870 0 1 2440
box -36 -49 3540 1467
use sky130_sram_1kbyte_1rw1r_8x1024_8_col_addr_dff  sky130_sram_1kbyte_1rw1r_8x1024_8_col_addr_dff_1
timestamp 1704896540
transform -1 0 77036 0 -1 86824
box -36 -49 3540 1467
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_0
timestamp 1704896540
transform 1 0 89211 0 1 5427
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_1
timestamp 1704896540
transform 1 0 89211 0 1 3747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_2
timestamp 1704896540
transform 1 0 89211 0 1 2067
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_3
timestamp 1704896540
transform 1 0 87729 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_4
timestamp 1704896540
transform 1 0 86049 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_5
timestamp 1704896540
transform 1 0 84369 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_6
timestamp 1704896540
transform 1 0 82689 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_7
timestamp 1704896540
transform 1 0 81009 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_8
timestamp 1704896540
transform 1 0 80337 0 1 11128
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_9
timestamp 1704896540
transform 1 0 89211 0 1 8787
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_10
timestamp 1704896540
transform 1 0 89211 0 1 7107
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_11
timestamp 1704896540
transform 1 0 89211 0 1 10467
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_12
timestamp 1704896540
transform 1 0 72609 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_13
timestamp 1704896540
transform 1 0 70929 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_14
timestamp 1704896540
transform 1 0 78574 0 1 11057
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_15
timestamp 1704896540
transform 1 0 79392 0 1 11057
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_16
timestamp 1704896540
transform 1 0 69249 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_17
timestamp 1704896540
transform 1 0 79329 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_18
timestamp 1704896540
transform 1 0 77649 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_19
timestamp 1704896540
transform 1 0 75969 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_20
timestamp 1704896540
transform 1 0 74289 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_21
timestamp 1704896540
transform 1 0 78974 0 1 17983
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_22
timestamp 1704896540
transform 1 0 79392 0 1 17983
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_23
timestamp 1704896540
transform 1 0 79054 0 1 19541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_24
timestamp 1704896540
transform 1 0 79392 0 1 19541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_25
timestamp 1704896540
transform 1 0 78654 0 1 12327
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_26
timestamp 1704896540
transform 1 0 79392 0 1 12327
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_27
timestamp 1704896540
transform 1 0 78734 0 1 13885
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_28
timestamp 1704896540
transform 1 0 79392 0 1 13885
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_29
timestamp 1704896540
transform 1 0 78814 0 1 15155
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_30
timestamp 1704896540
transform 1 0 79392 0 1 15155
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_31
timestamp 1704896540
transform 1 0 78894 0 1 16713
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_32
timestamp 1704896540
transform 1 0 79392 0 1 16713
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_33
timestamp 1704896540
transform 1 0 89211 0 1 13827
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_34
timestamp 1704896540
transform 1 0 89211 0 1 12147
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_35
timestamp 1704896540
transform 1 0 89211 0 1 15507
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_36
timestamp 1704896540
transform 1 0 80337 0 1 16784
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_37
timestamp 1704896540
transform 1 0 80337 0 1 12256
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_38
timestamp 1704896540
transform 1 0 80337 0 1 13956
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_39
timestamp 1704896540
transform 1 0 80337 0 1 15084
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_40
timestamp 1704896540
transform 1 0 80337 0 1 17912
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_41
timestamp 1704896540
transform 1 0 80337 0 1 19612
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_42
timestamp 1704896540
transform 1 0 89211 0 1 22227
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_43
timestamp 1704896540
transform 1 0 89211 0 1 20547
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_44
timestamp 1704896540
transform 1 0 89211 0 1 18867
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_45
timestamp 1704896540
transform 1 0 89211 0 1 17187
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_46
timestamp 1704896540
transform 1 0 67569 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_47
timestamp 1704896540
transform 1 0 65889 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_48
timestamp 1704896540
transform 1 0 64209 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_49
timestamp 1704896540
transform 1 0 60849 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_50
timestamp 1704896540
transform 1 0 62529 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_51
timestamp 1704896540
transform 1 0 59169 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_52
timestamp 1704896540
transform 1 0 57489 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_53
timestamp 1704896540
transform 1 0 50769 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_54
timestamp 1704896540
transform 1 0 54129 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_55
timestamp 1704896540
transform 1 0 47409 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_56
timestamp 1704896540
transform 1 0 55809 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_57
timestamp 1704896540
transform 1 0 49089 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_58
timestamp 1704896540
transform 1 0 45729 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_59
timestamp 1704896540
transform 1 0 52449 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_60
timestamp 1704896540
transform 1 0 55573 0 1 13067
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_61
timestamp 1704896540
transform 1 0 50581 0 1 13067
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_62
timestamp 1704896540
transform 1 0 45589 0 1 13067
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_63
timestamp 1704896540
transform 1 0 60565 0 1 13067
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_64
timestamp 1704896540
transform 1 0 89211 0 1 27267
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_65
timestamp 1704896540
transform 1 0 89211 0 1 23907
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_66
timestamp 1704896540
transform 1 0 89211 0 1 25587
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_67
timestamp 1704896540
transform 1 0 89211 0 1 28947
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_68
timestamp 1704896540
transform 1 0 89211 0 1 32307
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_69
timestamp 1704896540
transform 1 0 89211 0 1 30627
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_70
timestamp 1704896540
transform 1 0 89211 0 1 37347
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_71
timestamp 1704896540
transform 1 0 89211 0 1 35667
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_72
timestamp 1704896540
transform 1 0 89211 0 1 33987
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_73
timestamp 1704896540
transform 1 0 89211 0 1 44067
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_74
timestamp 1704896540
transform 1 0 89211 0 1 42387
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_75
timestamp 1704896540
transform 1 0 89211 0 1 40707
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_76
timestamp 1704896540
transform 1 0 89211 0 1 39027
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_77
timestamp 1704896540
transform 1 0 39009 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_78
timestamp 1704896540
transform 1 0 44049 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_79
timestamp 1704896540
transform 1 0 40689 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_80
timestamp 1704896540
transform 1 0 35649 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_81
timestamp 1704896540
transform 1 0 42369 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_82
timestamp 1704896540
transform 1 0 37329 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_83
timestamp 1704896540
transform 1 0 33969 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_84
timestamp 1704896540
transform 1 0 28929 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_85
timestamp 1704896540
transform 1 0 32289 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_86
timestamp 1704896540
transform 1 0 30609 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_87
timestamp 1704896540
transform 1 0 23889 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_88
timestamp 1704896540
transform 1 0 25855 0 1 2967
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_89
timestamp 1704896540
transform 1 0 24687 0 1 2967
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_90
timestamp 1704896540
transform 1 0 23519 0 1 2967
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_91
timestamp 1704896540
transform 1 0 27249 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_92
timestamp 1704896540
transform 1 0 25569 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_93
timestamp 1704896540
transform 1 0 30613 0 1 13067
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_94
timestamp 1704896540
transform 1 0 25621 0 1 13067
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_95
timestamp 1704896540
transform 1 0 23762 0 1 14313
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_96
timestamp 1704896540
transform 1 0 23638 0 1 12915
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_97
timestamp 1704896540
transform 1 0 23514 0 1 15707
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_98
timestamp 1704896540
transform 1 0 40597 0 1 13067
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_99
timestamp 1704896540
transform 1 0 35605 0 1 13067
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_100
timestamp 1704896540
transform 1 0 18849 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_101
timestamp 1704896540
transform 1 0 20529 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_102
timestamp 1704896540
transform 1 0 22209 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_103
timestamp 1704896540
transform 1 0 22351 0 1 2967
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_104
timestamp 1704896540
transform 1 0 21183 0 1 2967
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_105
timestamp 1704896540
transform 1 0 20015 0 1 2967
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_106
timestamp 1704896540
transform 1 0 18847 0 1 2967
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_107
timestamp 1704896540
transform 1 0 17679 0 1 2967
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_108
timestamp 1704896540
transform 1 0 16511 0 1 2967
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_109
timestamp 1704896540
transform 1 0 13809 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_110
timestamp 1704896540
transform 1 0 15343 0 1 2967
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_111
timestamp 1704896540
transform 1 0 14175 0 1 2967
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_112
timestamp 1704896540
transform 1 0 13007 0 1 2967
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_113
timestamp 1704896540
transform 1 0 17169 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_114
timestamp 1704896540
transform 1 0 12129 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_115
timestamp 1704896540
transform 1 0 15489 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_116
timestamp 1704896540
transform 1 0 7089 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_117
timestamp 1704896540
transform 1 0 10449 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_118
timestamp 1704896540
transform 1 0 8769 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_119
timestamp 1704896540
transform 1 0 1713 0 1 2067
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_120
timestamp 1704896540
transform 1 0 1713 0 1 5427
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_121
timestamp 1704896540
transform 1 0 5409 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_122
timestamp 1704896540
transform 1 0 3729 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_123
timestamp 1704896540
transform 1 0 1713 0 1 3747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_124
timestamp 1704896540
transform 1 0 2049 0 1 1731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_125
timestamp 1704896540
transform 1 0 1713 0 1 10467
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_126
timestamp 1704896540
transform 1 0 1713 0 1 8787
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_127
timestamp 1704896540
transform 1 0 2673 0 1 10214
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_128
timestamp 1704896540
transform 1 0 2673 0 1 8514
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_129
timestamp 1704896540
transform 1 0 1713 0 1 7107
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_130
timestamp 1704896540
transform 1 0 5894 0 1 8619
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_131
timestamp 1704896540
transform 1 0 1713 0 1 13827
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_132
timestamp 1704896540
transform 1 0 1713 0 1 15507
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_133
timestamp 1704896540
transform 1 0 1713 0 1 12147
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_134
timestamp 1704896540
transform 1 0 1713 0 1 22227
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_135
timestamp 1704896540
transform 1 0 1713 0 1 20547
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_136
timestamp 1704896540
transform 1 0 1713 0 1 18867
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_137
timestamp 1704896540
transform 1 0 1713 0 1 17187
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_138
timestamp 1704896540
transform 1 0 11669 0 1 12915
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_139
timestamp 1704896540
transform 1 0 19811 0 1 18555
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_140
timestamp 1704896540
transform 1 0 11669 0 1 18555
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_141
timestamp 1704896540
transform 1 0 11669 0 1 15727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_142
timestamp 1704896540
transform 1 0 11669 0 1 14313
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_143
timestamp 1704896540
transform 1 0 11616 0 1 33097
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_144
timestamp 1704896540
transform 1 0 12030 0 1 31539
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_145
timestamp 1704896540
transform 1 0 11950 0 1 30269
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_146
timestamp 1704896540
transform 1 0 11616 0 1 30269
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_147
timestamp 1704896540
transform 1 0 11870 0 1 28711
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_148
timestamp 1704896540
transform 1 0 11616 0 1 28711
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_149
timestamp 1704896540
transform 1 0 12110 0 1 33097
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_150
timestamp 1704896540
transform 1 0 11616 0 1 31539
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_151
timestamp 1704896540
transform 1 0 1713 0 1 23907
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_152
timestamp 1704896540
transform 1 0 1713 0 1 27267
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_153
timestamp 1704896540
transform 1 0 2460 0 1 25663
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_154
timestamp 1704896540
transform 1 0 1713 0 1 25587
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_155
timestamp 1704896540
transform 1 0 1713 0 1 28947
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_156
timestamp 1704896540
transform 1 0 1713 0 1 30627
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_157
timestamp 1704896540
transform 1 0 1713 0 1 32307
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_158
timestamp 1704896540
transform 1 0 10671 0 1 33168
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_159
timestamp 1704896540
transform 1 0 10671 0 1 31468
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_160
timestamp 1704896540
transform 1 0 10671 0 1 30340
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_161
timestamp 1704896540
transform 1 0 10671 0 1 28640
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_162
timestamp 1704896540
transform 1 0 10671 0 1 34296
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_163
timestamp 1704896540
transform 1 0 10671 0 1 37124
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_164
timestamp 1704896540
transform 1 0 10671 0 1 35996
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_165
timestamp 1704896540
transform 1 0 1713 0 1 33987
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_166
timestamp 1704896540
transform 1 0 1713 0 1 37347
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_167
timestamp 1704896540
transform 1 0 1713 0 1 35667
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_168
timestamp 1704896540
transform 1 0 1713 0 1 44067
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_169
timestamp 1704896540
transform 1 0 1713 0 1 42387
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_170
timestamp 1704896540
transform 1 0 1713 0 1 40707
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_171
timestamp 1704896540
transform 1 0 1713 0 1 39027
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_172
timestamp 1704896540
transform 1 0 11616 0 1 35925
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_173
timestamp 1704896540
transform 1 0 12190 0 1 34367
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_174
timestamp 1704896540
transform 1 0 11616 0 1 34367
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_175
timestamp 1704896540
transform 1 0 12350 0 1 37195
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_176
timestamp 1704896540
transform 1 0 11616 0 1 37195
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_177
timestamp 1704896540
transform 1 0 12270 0 1 35925
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_178
timestamp 1704896540
transform 1 0 1713 0 1 47427
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_179
timestamp 1704896540
transform 1 0 1713 0 1 45747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_180
timestamp 1704896540
transform 1 0 1713 0 1 49107
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_181
timestamp 1704896540
transform 1 0 1713 0 1 52467
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_182
timestamp 1704896540
transform 1 0 1713 0 1 50787
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_183
timestamp 1704896540
transform 1 0 1713 0 1 54147
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_184
timestamp 1704896540
transform 1 0 1713 0 1 57507
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_185
timestamp 1704896540
transform 1 0 1713 0 1 55827
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_186
timestamp 1704896540
transform 1 0 1713 0 1 60867
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_187
timestamp 1704896540
transform 1 0 1713 0 1 59187
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_188
timestamp 1704896540
transform 1 0 1713 0 1 64227
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_189
timestamp 1704896540
transform 1 0 1713 0 1 62547
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_190
timestamp 1704896540
transform 1 0 1713 0 1 65907
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_191
timestamp 1704896540
transform 1 0 1713 0 1 70947
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_192
timestamp 1704896540
transform 1 0 1713 0 1 69267
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_193
timestamp 1704896540
transform 1 0 1713 0 1 67587
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_194
timestamp 1704896540
transform 1 0 1713 0 1 75987
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_195
timestamp 1704896540
transform 1 0 1713 0 1 74307
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_196
timestamp 1704896540
transform 1 0 1713 0 1 72627
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_197
timestamp 1704896540
transform 1 0 1713 0 1 77667
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_198
timestamp 1704896540
transform 1 0 1713 0 1 81027
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_199
timestamp 1704896540
transform 1 0 1713 0 1 79347
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_200
timestamp 1704896540
transform 1 0 1713 0 1 82707
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_201
timestamp 1704896540
transform 1 0 1713 0 1 86067
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_202
timestamp 1704896540
transform 1 0 1713 0 1 84387
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_203
timestamp 1704896540
transform 1 0 5409 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_204
timestamp 1704896540
transform 1 0 3729 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_205
timestamp 1704896540
transform 1 0 2049 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_206
timestamp 1704896540
transform 1 0 10449 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_207
timestamp 1704896540
transform 1 0 8769 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_208
timestamp 1704896540
transform 1 0 7089 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_209
timestamp 1704896540
transform 1 0 22209 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_210
timestamp 1704896540
transform 1 0 20529 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_211
timestamp 1704896540
transform 1 0 18849 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_212
timestamp 1704896540
transform 1 0 17169 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_213
timestamp 1704896540
transform 1 0 15489 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_214
timestamp 1704896540
transform 1 0 13809 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_215
timestamp 1704896540
transform 1 0 12129 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_216
timestamp 1704896540
transform 1 0 40597 0 1 77845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_217
timestamp 1704896540
transform 1 0 35605 0 1 77845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_218
timestamp 1704896540
transform 1 0 25621 0 1 77845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_219
timestamp 1704896540
transform 1 0 30613 0 1 77845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_220
timestamp 1704896540
transform 1 0 28929 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_221
timestamp 1704896540
transform 1 0 27249 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_222
timestamp 1704896540
transform 1 0 25569 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_223
timestamp 1704896540
transform 1 0 23889 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_224
timestamp 1704896540
transform 1 0 33969 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_225
timestamp 1704896540
transform 1 0 32289 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_226
timestamp 1704896540
transform 1 0 30609 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_227
timestamp 1704896540
transform 1 0 42369 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_228
timestamp 1704896540
transform 1 0 40689 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_229
timestamp 1704896540
transform 1 0 39009 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_230
timestamp 1704896540
transform 1 0 37329 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_231
timestamp 1704896540
transform 1 0 35649 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_232
timestamp 1704896540
transform 1 0 44049 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_233
timestamp 1704896540
transform 1 0 89211 0 1 45747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_234
timestamp 1704896540
transform 1 0 89211 0 1 49107
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_235
timestamp 1704896540
transform 1 0 89211 0 1 47427
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_236
timestamp 1704896540
transform 1 0 89211 0 1 54147
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_237
timestamp 1704896540
transform 1 0 89211 0 1 50787
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_238
timestamp 1704896540
transform 1 0 89211 0 1 52467
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_239
timestamp 1704896540
transform 1 0 89211 0 1 55827
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_240
timestamp 1704896540
transform 1 0 89211 0 1 60867
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_241
timestamp 1704896540
transform 1 0 89211 0 1 59187
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_242
timestamp 1704896540
transform 1 0 89211 0 1 57507
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_243
timestamp 1704896540
transform 1 0 88464 0 1 62421
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_244
timestamp 1704896540
transform 1 0 89211 0 1 65907
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_245
timestamp 1704896540
transform 1 0 89211 0 1 64227
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_246
timestamp 1704896540
transform 1 0 89211 0 1 62547
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_247
timestamp 1704896540
transform 1 0 60565 0 1 77845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_248
timestamp 1704896540
transform 1 0 67128 0 1 75189
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_249
timestamp 1704896540
transform 1 0 67252 0 1 73771
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_250
timestamp 1704896540
transform 1 0 45589 0 1 77845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_251
timestamp 1704896540
transform 1 0 55573 0 1 77845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_252
timestamp 1704896540
transform 1 0 50581 0 1 77845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_253
timestamp 1704896540
transform 1 0 54129 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_254
timestamp 1704896540
transform 1 0 52449 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_255
timestamp 1704896540
transform 1 0 50769 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_256
timestamp 1704896540
transform 1 0 49089 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_257
timestamp 1704896540
transform 1 0 47409 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_258
timestamp 1704896540
transform 1 0 45729 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_259
timestamp 1704896540
transform 1 0 55809 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_260
timestamp 1704896540
transform 1 0 67569 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_261
timestamp 1704896540
transform 1 0 65889 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_262
timestamp 1704896540
transform 1 0 64209 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_263
timestamp 1704896540
transform 1 0 62529 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_264
timestamp 1704896540
transform 1 0 60849 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_265
timestamp 1704896540
transform 1 0 59169 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_266
timestamp 1704896540
transform 1 0 57489 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_267
timestamp 1704896540
transform 1 0 89211 0 1 69267
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_268
timestamp 1704896540
transform 1 0 89211 0 1 67587
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_269
timestamp 1704896540
transform 1 0 89211 0 1 70947
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_270
timestamp 1704896540
transform 1 0 89211 0 1 77667
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_271
timestamp 1704896540
transform 1 0 89211 0 1 75987
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_272
timestamp 1704896540
transform 1 0 89211 0 1 74307
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_273
timestamp 1704896540
transform 1 0 89211 0 1 72627
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_274
timestamp 1704896540
transform 1 0 79339 0 1 73771
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_275
timestamp 1704896540
transform 1 0 71113 0 1 72357
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_276
timestamp 1704896540
transform 1 0 79339 0 1 72357
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_277
timestamp 1704896540
transform 1 0 79339 0 1 75169
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_278
timestamp 1704896540
transform 1 0 70929 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_279
timestamp 1704896540
transform 1 0 69249 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_280
timestamp 1704896540
transform 1 0 72609 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_281
timestamp 1704896540
transform 1 0 74497 0 1 86223
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_282
timestamp 1704896540
transform 1 0 75665 0 1 86223
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_283
timestamp 1704896540
transform 1 0 76833 0 1 86223
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_284
timestamp 1704896540
transform 1 0 79329 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_285
timestamp 1704896540
transform 1 0 77649 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_286
timestamp 1704896540
transform 1 0 75969 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_287
timestamp 1704896540
transform 1 0 74289 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_288
timestamp 1704896540
transform 1 0 89211 0 1 79347
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_289
timestamp 1704896540
transform 1 0 88251 0 1 79570
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_290
timestamp 1704896540
transform 1 0 89211 0 1 82707
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_291
timestamp 1704896540
transform 1 0 89211 0 1 81027
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_292
timestamp 1704896540
transform 1 0 81009 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_293
timestamp 1704896540
transform 1 0 84369 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_294
timestamp 1704896540
transform 1 0 82689 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_295
timestamp 1704896540
transform 1 0 89211 0 1 86067
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_296
timestamp 1704896540
transform 1 0 89211 0 1 84387
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_297
timestamp 1704896540
transform 1 0 87729 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_298
timestamp 1704896540
transform 1 0 86049 0 1 87459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_299
timestamp 1704896540
transform 1 0 85114 0 1 79465
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_0
timestamp 1704896540
transform 1 0 89219 0 1 5423
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_1
timestamp 1704896540
transform 1 0 89219 0 1 5087
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_2
timestamp 1704896540
transform 1 0 89219 0 1 4751
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_3
timestamp 1704896540
transform 1 0 89219 0 1 4415
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_4
timestamp 1704896540
transform 1 0 89219 0 1 4079
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_5
timestamp 1704896540
transform 1 0 89219 0 1 3743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_6
timestamp 1704896540
transform 1 0 89219 0 1 3407
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_7
timestamp 1704896540
transform 1 0 89219 0 1 3071
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_8
timestamp 1704896540
transform 1 0 89219 0 1 2735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_9
timestamp 1704896540
transform 1 0 88745 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_10
timestamp 1704896540
transform 1 0 89219 0 1 2399
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_11
timestamp 1704896540
transform 1 0 88409 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_12
timestamp 1704896540
transform 1 0 89219 0 1 2063
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_13
timestamp 1704896540
transform 1 0 88073 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_14
timestamp 1704896540
transform 1 0 87737 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_15
timestamp 1704896540
transform 1 0 87401 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_16
timestamp 1704896540
transform 1 0 87065 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_17
timestamp 1704896540
transform 1 0 86729 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_18
timestamp 1704896540
transform 1 0 86393 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_19
timestamp 1704896540
transform 1 0 86057 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_20
timestamp 1704896540
transform 1 0 85721 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_21
timestamp 1704896540
transform 1 0 85385 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_22
timestamp 1704896540
transform 1 0 84713 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_23
timestamp 1704896540
transform 1 0 84377 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_24
timestamp 1704896540
transform 1 0 84041 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_25
timestamp 1704896540
transform 1 0 83705 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_26
timestamp 1704896540
transform 1 0 83369 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_27
timestamp 1704896540
transform 1 0 83033 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_28
timestamp 1704896540
transform 1 0 82697 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_29
timestamp 1704896540
transform 1 0 82361 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_30
timestamp 1704896540
transform 1 0 82025 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_31
timestamp 1704896540
transform 1 0 81689 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_32
timestamp 1704896540
transform 1 0 81353 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_33
timestamp 1704896540
transform 1 0 81017 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_34
timestamp 1704896540
transform 1 0 80681 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_35
timestamp 1704896540
transform 1 0 80345 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_36
timestamp 1704896540
transform 1 0 80009 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_37
timestamp 1704896540
transform 1 0 79673 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_38
timestamp 1704896540
transform 1 0 89219 0 1 9791
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_39
timestamp 1704896540
transform 1 0 89219 0 1 9455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_40
timestamp 1704896540
transform 1 0 89219 0 1 9119
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_41
timestamp 1704896540
transform 1 0 89219 0 1 8783
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_42
timestamp 1704896540
transform 1 0 89219 0 1 8447
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_43
timestamp 1704896540
transform 1 0 89219 0 1 8111
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_44
timestamp 1704896540
transform 1 0 89219 0 1 7775
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_45
timestamp 1704896540
transform 1 0 89219 0 1 7439
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_46
timestamp 1704896540
transform 1 0 89219 0 1 7103
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_47
timestamp 1704896540
transform 1 0 89219 0 1 6767
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_48
timestamp 1704896540
transform 1 0 89219 0 1 6431
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_49
timestamp 1704896540
transform 1 0 89219 0 1 6095
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_50
timestamp 1704896540
transform 1 0 89219 0 1 10127
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_51
timestamp 1704896540
transform 1 0 89219 0 1 11135
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_52
timestamp 1704896540
transform 1 0 89219 0 1 10799
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_53
timestamp 1704896540
transform 1 0 89219 0 1 10463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_54
timestamp 1704896540
transform 1 0 85049 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_55
timestamp 1704896540
transform 1 0 89219 0 1 5759
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_56
timestamp 1704896540
transform 1 0 74297 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_57
timestamp 1704896540
transform 1 0 73961 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_58
timestamp 1704896540
transform 1 0 73625 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_59
timestamp 1704896540
transform 1 0 73289 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_60
timestamp 1704896540
transform 1 0 72953 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_61
timestamp 1704896540
transform 1 0 72617 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_62
timestamp 1704896540
transform 1 0 72281 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_63
timestamp 1704896540
transform 1 0 71945 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_64
timestamp 1704896540
transform 1 0 71609 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_65
timestamp 1704896540
transform 1 0 71273 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_66
timestamp 1704896540
transform 1 0 70937 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_67
timestamp 1704896540
transform 1 0 68921 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_68
timestamp 1704896540
transform 1 0 68585 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_69
timestamp 1704896540
transform 1 0 68249 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_70
timestamp 1704896540
transform 1 0 70601 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_71
timestamp 1704896540
transform 1 0 70265 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_72
timestamp 1704896540
transform 1 0 69929 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_73
timestamp 1704896540
transform 1 0 69593 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_74
timestamp 1704896540
transform 1 0 79337 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_75
timestamp 1704896540
transform 1 0 79001 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_76
timestamp 1704896540
transform 1 0 78665 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_77
timestamp 1704896540
transform 1 0 78329 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_78
timestamp 1704896540
transform 1 0 77993 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_79
timestamp 1704896540
transform 1 0 77657 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_80
timestamp 1704896540
transform 1 0 77321 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_81
timestamp 1704896540
transform 1 0 76985 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_82
timestamp 1704896540
transform 1 0 76649 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_83
timestamp 1704896540
transform 1 0 76313 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_84
timestamp 1704896540
transform 1 0 75977 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_85
timestamp 1704896540
transform 1 0 75641 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_86
timestamp 1704896540
transform 1 0 75305 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_87
timestamp 1704896540
transform 1 0 74969 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_88
timestamp 1704896540
transform 1 0 69257 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_89
timestamp 1704896540
transform 1 0 74633 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_90
timestamp 1704896540
transform 1 0 89219 0 1 14159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_91
timestamp 1704896540
transform 1 0 89219 0 1 13823
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_92
timestamp 1704896540
transform 1 0 89219 0 1 13487
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_93
timestamp 1704896540
transform 1 0 89219 0 1 11471
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_94
timestamp 1704896540
transform 1 0 89219 0 1 13151
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_95
timestamp 1704896540
transform 1 0 89219 0 1 12815
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_96
timestamp 1704896540
transform 1 0 89219 0 1 12479
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_97
timestamp 1704896540
transform 1 0 89219 0 1 12143
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_98
timestamp 1704896540
transform 1 0 89219 0 1 11807
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_99
timestamp 1704896540
transform 1 0 89219 0 1 16511
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_100
timestamp 1704896540
transform 1 0 89219 0 1 16175
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_101
timestamp 1704896540
transform 1 0 89219 0 1 15839
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_102
timestamp 1704896540
transform 1 0 89219 0 1 15503
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_103
timestamp 1704896540
transform 1 0 89219 0 1 15167
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_104
timestamp 1704896540
transform 1 0 89219 0 1 14831
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_105
timestamp 1704896540
transform 1 0 89219 0 1 14495
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_106
timestamp 1704896540
transform 1 0 89219 0 1 22223
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_107
timestamp 1704896540
transform 1 0 89219 0 1 21887
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_108
timestamp 1704896540
transform 1 0 89219 0 1 21551
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_109
timestamp 1704896540
transform 1 0 89219 0 1 21215
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_110
timestamp 1704896540
transform 1 0 89219 0 1 20879
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_111
timestamp 1704896540
transform 1 0 89219 0 1 20543
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_112
timestamp 1704896540
transform 1 0 89219 0 1 20207
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_113
timestamp 1704896540
transform 1 0 89219 0 1 19871
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_114
timestamp 1704896540
transform 1 0 89219 0 1 19535
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_115
timestamp 1704896540
transform 1 0 89219 0 1 19199
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_116
timestamp 1704896540
transform 1 0 89219 0 1 18863
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_117
timestamp 1704896540
transform 1 0 89219 0 1 18527
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_118
timestamp 1704896540
transform 1 0 89219 0 1 18191
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_119
timestamp 1704896540
transform 1 0 89219 0 1 17855
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_120
timestamp 1704896540
transform 1 0 89219 0 1 17519
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_121
timestamp 1704896540
transform 1 0 89219 0 1 17183
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_122
timestamp 1704896540
transform 1 0 89219 0 1 16847
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_123
timestamp 1704896540
transform 1 0 67577 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_124
timestamp 1704896540
transform 1 0 67241 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_125
timestamp 1704896540
transform 1 0 66905 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_126
timestamp 1704896540
transform 1 0 57161 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_127
timestamp 1704896540
transform 1 0 66569 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_128
timestamp 1704896540
transform 1 0 66233 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_129
timestamp 1704896540
transform 1 0 65897 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_130
timestamp 1704896540
transform 1 0 65561 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_131
timestamp 1704896540
transform 1 0 65225 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_132
timestamp 1704896540
transform 1 0 64889 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_133
timestamp 1704896540
transform 1 0 64553 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_134
timestamp 1704896540
transform 1 0 64217 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_135
timestamp 1704896540
transform 1 0 60521 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_136
timestamp 1704896540
transform 1 0 63881 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_137
timestamp 1704896540
transform 1 0 63545 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_138
timestamp 1704896540
transform 1 0 58841 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_139
timestamp 1704896540
transform 1 0 60185 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_140
timestamp 1704896540
transform 1 0 59849 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_141
timestamp 1704896540
transform 1 0 57833 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_142
timestamp 1704896540
transform 1 0 57497 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_143
timestamp 1704896540
transform 1 0 61193 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_144
timestamp 1704896540
transform 1 0 58505 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_145
timestamp 1704896540
transform 1 0 59513 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_146
timestamp 1704896540
transform 1 0 63209 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_147
timestamp 1704896540
transform 1 0 62873 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_148
timestamp 1704896540
transform 1 0 62537 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_149
timestamp 1704896540
transform 1 0 62201 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_150
timestamp 1704896540
transform 1 0 61865 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_151
timestamp 1704896540
transform 1 0 61529 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_152
timestamp 1704896540
transform 1 0 60857 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_153
timestamp 1704896540
transform 1 0 67913 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_154
timestamp 1704896540
transform 1 0 59177 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_155
timestamp 1704896540
transform 1 0 58169 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_156
timestamp 1704896540
transform 1 0 48425 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_157
timestamp 1704896540
transform 1 0 46409 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_158
timestamp 1704896540
transform 1 0 55145 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_159
timestamp 1704896540
transform 1 0 51113 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_160
timestamp 1704896540
transform 1 0 46745 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_161
timestamp 1704896540
transform 1 0 50777 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_162
timestamp 1704896540
transform 1 0 48089 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_163
timestamp 1704896540
transform 1 0 54809 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_164
timestamp 1704896540
transform 1 0 54473 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_165
timestamp 1704896540
transform 1 0 56489 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_166
timestamp 1704896540
transform 1 0 47753 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_167
timestamp 1704896540
transform 1 0 54137 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_168
timestamp 1704896540
transform 1 0 56153 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_169
timestamp 1704896540
transform 1 0 48761 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_170
timestamp 1704896540
transform 1 0 49433 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_171
timestamp 1704896540
transform 1 0 53129 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_172
timestamp 1704896540
transform 1 0 50441 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_173
timestamp 1704896540
transform 1 0 50105 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_174
timestamp 1704896540
transform 1 0 49097 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_175
timestamp 1704896540
transform 1 0 49769 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_176
timestamp 1704896540
transform 1 0 52457 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_177
timestamp 1704896540
transform 1 0 53801 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_178
timestamp 1704896540
transform 1 0 51785 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_179
timestamp 1704896540
transform 1 0 52121 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_180
timestamp 1704896540
transform 1 0 51449 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_181
timestamp 1704896540
transform 1 0 46073 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_182
timestamp 1704896540
transform 1 0 45737 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_183
timestamp 1704896540
transform 1 0 53465 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_184
timestamp 1704896540
transform 1 0 52793 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_185
timestamp 1704896540
transform 1 0 47417 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_186
timestamp 1704896540
transform 1 0 55817 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_187
timestamp 1704896540
transform 1 0 47081 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_188
timestamp 1704896540
transform 1 0 55481 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_189
timestamp 1704896540
transform 1 0 56825 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_190
timestamp 1704896540
transform 1 0 89219 0 1 25583
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_191
timestamp 1704896540
transform 1 0 89219 0 1 25247
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_192
timestamp 1704896540
transform 1 0 89219 0 1 24911
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_193
timestamp 1704896540
transform 1 0 89219 0 1 24575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_194
timestamp 1704896540
transform 1 0 89219 0 1 22895
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_195
timestamp 1704896540
transform 1 0 89219 0 1 22559
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_196
timestamp 1704896540
transform 1 0 89219 0 1 24239
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_197
timestamp 1704896540
transform 1 0 89219 0 1 27599
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_198
timestamp 1704896540
transform 1 0 89219 0 1 27263
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_199
timestamp 1704896540
transform 1 0 89219 0 1 26927
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_200
timestamp 1704896540
transform 1 0 89219 0 1 26591
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_201
timestamp 1704896540
transform 1 0 89219 0 1 26255
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_202
timestamp 1704896540
transform 1 0 89219 0 1 23903
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_203
timestamp 1704896540
transform 1 0 89219 0 1 23567
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_204
timestamp 1704896540
transform 1 0 89219 0 1 25919
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_205
timestamp 1704896540
transform 1 0 89219 0 1 23231
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_206
timestamp 1704896540
transform 1 0 89219 0 1 30287
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_207
timestamp 1704896540
transform 1 0 89219 0 1 29951
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_208
timestamp 1704896540
transform 1 0 89219 0 1 29615
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_209
timestamp 1704896540
transform 1 0 89219 0 1 29279
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_210
timestamp 1704896540
transform 1 0 89219 0 1 28943
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_211
timestamp 1704896540
transform 1 0 89219 0 1 28607
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_212
timestamp 1704896540
transform 1 0 89219 0 1 28271
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_213
timestamp 1704896540
transform 1 0 89219 0 1 30623
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_214
timestamp 1704896540
transform 1 0 89219 0 1 33311
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_215
timestamp 1704896540
transform 1 0 89219 0 1 32975
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_216
timestamp 1704896540
transform 1 0 89219 0 1 32639
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_217
timestamp 1704896540
transform 1 0 89219 0 1 32303
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_218
timestamp 1704896540
transform 1 0 89219 0 1 31967
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_219
timestamp 1704896540
transform 1 0 89219 0 1 31631
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_220
timestamp 1704896540
transform 1 0 89219 0 1 31295
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_221
timestamp 1704896540
transform 1 0 89219 0 1 30959
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_222
timestamp 1704896540
transform 1 0 89219 0 1 27935
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_223
timestamp 1704896540
transform 1 0 89219 0 1 38687
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_224
timestamp 1704896540
transform 1 0 89219 0 1 38351
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_225
timestamp 1704896540
transform 1 0 89219 0 1 38015
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_226
timestamp 1704896540
transform 1 0 89219 0 1 37679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_227
timestamp 1704896540
transform 1 0 89219 0 1 37343
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_228
timestamp 1704896540
transform 1 0 89219 0 1 37007
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_229
timestamp 1704896540
transform 1 0 89219 0 1 36671
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_230
timestamp 1704896540
transform 1 0 89219 0 1 36335
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_231
timestamp 1704896540
transform 1 0 89219 0 1 35999
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_232
timestamp 1704896540
transform 1 0 89219 0 1 35663
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_233
timestamp 1704896540
transform 1 0 89219 0 1 35327
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_234
timestamp 1704896540
transform 1 0 89219 0 1 34991
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_235
timestamp 1704896540
transform 1 0 89219 0 1 34655
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_236
timestamp 1704896540
transform 1 0 89219 0 1 34319
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_237
timestamp 1704896540
transform 1 0 89219 0 1 33983
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_238
timestamp 1704896540
transform 1 0 89219 0 1 33647
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_239
timestamp 1704896540
transform 1 0 89219 0 1 44399
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_240
timestamp 1704896540
transform 1 0 89219 0 1 44063
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_241
timestamp 1704896540
transform 1 0 89219 0 1 43727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_242
timestamp 1704896540
transform 1 0 89219 0 1 43391
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_243
timestamp 1704896540
transform 1 0 89219 0 1 43055
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_244
timestamp 1704896540
transform 1 0 89219 0 1 42719
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_245
timestamp 1704896540
transform 1 0 89219 0 1 42383
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_246
timestamp 1704896540
transform 1 0 89219 0 1 42047
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_247
timestamp 1704896540
transform 1 0 89219 0 1 41711
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_248
timestamp 1704896540
transform 1 0 89219 0 1 41375
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_249
timestamp 1704896540
transform 1 0 89219 0 1 41039
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_250
timestamp 1704896540
transform 1 0 89219 0 1 40703
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_251
timestamp 1704896540
transform 1 0 89219 0 1 40367
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_252
timestamp 1704896540
transform 1 0 89219 0 1 40031
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_253
timestamp 1704896540
transform 1 0 89219 0 1 39695
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_254
timestamp 1704896540
transform 1 0 89219 0 1 39359
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_255
timestamp 1704896540
transform 1 0 89219 0 1 39023
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_256
timestamp 1704896540
transform 1 0 45065 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_257
timestamp 1704896540
transform 1 0 40697 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_258
timestamp 1704896540
transform 1 0 44729 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_259
timestamp 1704896540
transform 1 0 37337 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_260
timestamp 1704896540
transform 1 0 37001 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_261
timestamp 1704896540
transform 1 0 40361 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_262
timestamp 1704896540
transform 1 0 39017 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_263
timestamp 1704896540
transform 1 0 41033 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_264
timestamp 1704896540
transform 1 0 44393 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_265
timestamp 1704896540
transform 1 0 44057 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_266
timestamp 1704896540
transform 1 0 38681 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_267
timestamp 1704896540
transform 1 0 36665 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_268
timestamp 1704896540
transform 1 0 41705 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_269
timestamp 1704896540
transform 1 0 38345 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_270
timestamp 1704896540
transform 1 0 36329 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_271
timestamp 1704896540
transform 1 0 35993 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_272
timestamp 1704896540
transform 1 0 39353 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_273
timestamp 1704896540
transform 1 0 42041 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_274
timestamp 1704896540
transform 1 0 43721 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_275
timestamp 1704896540
transform 1 0 41369 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_276
timestamp 1704896540
transform 1 0 35657 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_277
timestamp 1704896540
transform 1 0 45401 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_278
timestamp 1704896540
transform 1 0 40025 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_279
timestamp 1704896540
transform 1 0 43385 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_280
timestamp 1704896540
transform 1 0 39689 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_281
timestamp 1704896540
transform 1 0 35321 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_282
timestamp 1704896540
transform 1 0 43049 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_283
timestamp 1704896540
transform 1 0 34985 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_284
timestamp 1704896540
transform 1 0 42713 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_285
timestamp 1704896540
transform 1 0 38009 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_286
timestamp 1704896540
transform 1 0 34649 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_287
timestamp 1704896540
transform 1 0 37673 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_288
timestamp 1704896540
transform 1 0 34313 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_289
timestamp 1704896540
transform 1 0 42377 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_290
timestamp 1704896540
transform 1 0 29945 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_291
timestamp 1704896540
transform 1 0 33977 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_292
timestamp 1704896540
transform 1 0 29609 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_293
timestamp 1704896540
transform 1 0 28937 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_294
timestamp 1704896540
transform 1 0 32297 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_295
timestamp 1704896540
transform 1 0 31961 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_296
timestamp 1704896540
transform 1 0 31625 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_297
timestamp 1704896540
transform 1 0 31289 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_298
timestamp 1704896540
transform 1 0 32633 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_299
timestamp 1704896540
transform 1 0 30953 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_300
timestamp 1704896540
transform 1 0 33641 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_301
timestamp 1704896540
transform 1 0 33305 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_302
timestamp 1704896540
transform 1 0 32969 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_303
timestamp 1704896540
transform 1 0 29273 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_304
timestamp 1704896540
transform 1 0 30617 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_305
timestamp 1704896540
transform 1 0 30281 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_306
timestamp 1704896540
transform 1 0 23225 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_307
timestamp 1704896540
transform 1 0 24569 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_308
timestamp 1704896540
transform 1 0 24233 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_309
timestamp 1704896540
transform 1 0 25577 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_310
timestamp 1704896540
transform 1 0 23561 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_311
timestamp 1704896540
transform 1 0 25241 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_312
timestamp 1704896540
transform 1 0 23897 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_313
timestamp 1704896540
transform 1 0 28265 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_314
timestamp 1704896540
transform 1 0 27929 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_315
timestamp 1704896540
transform 1 0 27593 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_316
timestamp 1704896540
transform 1 0 27257 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_317
timestamp 1704896540
transform 1 0 26921 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_318
timestamp 1704896540
transform 1 0 26585 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_319
timestamp 1704896540
transform 1 0 26249 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_320
timestamp 1704896540
transform 1 0 25913 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_321
timestamp 1704896540
transform 1 0 24905 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_322
timestamp 1704896540
transform 1 0 28601 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_323
timestamp 1704896540
transform 1 0 21881 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_324
timestamp 1704896540
transform 1 0 21545 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_325
timestamp 1704896540
transform 1 0 18857 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_326
timestamp 1704896540
transform 1 0 18521 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_327
timestamp 1704896540
transform 1 0 18185 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_328
timestamp 1704896540
transform 1 0 19865 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_329
timestamp 1704896540
transform 1 0 20873 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_330
timestamp 1704896540
transform 1 0 19193 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_331
timestamp 1704896540
transform 1 0 21209 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_332
timestamp 1704896540
transform 1 0 22217 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_333
timestamp 1704896540
transform 1 0 17849 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_334
timestamp 1704896540
transform 1 0 19529 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_335
timestamp 1704896540
transform 1 0 20537 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_336
timestamp 1704896540
transform 1 0 22553 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_337
timestamp 1704896540
transform 1 0 17513 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_338
timestamp 1704896540
transform 1 0 20201 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_339
timestamp 1704896540
transform 1 0 12137 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_340
timestamp 1704896540
transform 1 0 11801 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_341
timestamp 1704896540
transform 1 0 14825 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_342
timestamp 1704896540
transform 1 0 13481 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_343
timestamp 1704896540
transform 1 0 14489 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_344
timestamp 1704896540
transform 1 0 15497 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_345
timestamp 1704896540
transform 1 0 13145 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_346
timestamp 1704896540
transform 1 0 12809 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_347
timestamp 1704896540
transform 1 0 12473 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_348
timestamp 1704896540
transform 1 0 14153 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_349
timestamp 1704896540
transform 1 0 16841 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_350
timestamp 1704896540
transform 1 0 13817 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_351
timestamp 1704896540
transform 1 0 16505 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_352
timestamp 1704896540
transform 1 0 15161 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_353
timestamp 1704896540
transform 1 0 16169 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_354
timestamp 1704896540
transform 1 0 15833 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_355
timestamp 1704896540
transform 1 0 17177 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_356
timestamp 1704896540
transform 1 0 8105 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_357
timestamp 1704896540
transform 1 0 7769 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_358
timestamp 1704896540
transform 1 0 11465 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_359
timestamp 1704896540
transform 1 0 7433 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_360
timestamp 1704896540
transform 1 0 11129 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_361
timestamp 1704896540
transform 1 0 10793 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_362
timestamp 1704896540
transform 1 0 10457 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_363
timestamp 1704896540
transform 1 0 10121 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_364
timestamp 1704896540
transform 1 0 9785 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_365
timestamp 1704896540
transform 1 0 7097 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_366
timestamp 1704896540
transform 1 0 9449 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_367
timestamp 1704896540
transform 1 0 9113 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_368
timestamp 1704896540
transform 1 0 6089 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_369
timestamp 1704896540
transform 1 0 6761 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_370
timestamp 1704896540
transform 1 0 6425 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_371
timestamp 1704896540
transform 1 0 8777 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_372
timestamp 1704896540
transform 1 0 8441 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_373
timestamp 1704896540
transform 1 0 1721 0 1 2399
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_374
timestamp 1704896540
transform 1 0 1721 0 1 2063
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_375
timestamp 1704896540
transform 1 0 1721 0 1 5423
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_376
timestamp 1704896540
transform 1 0 1721 0 1 5087
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_377
timestamp 1704896540
transform 1 0 1721 0 1 4751
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_378
timestamp 1704896540
transform 1 0 1721 0 1 4415
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_379
timestamp 1704896540
transform 1 0 5753 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_380
timestamp 1704896540
transform 1 0 5417 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_381
timestamp 1704896540
transform 1 0 5081 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_382
timestamp 1704896540
transform 1 0 4745 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_383
timestamp 1704896540
transform 1 0 4409 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_384
timestamp 1704896540
transform 1 0 4073 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_385
timestamp 1704896540
transform 1 0 3737 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_386
timestamp 1704896540
transform 1 0 1721 0 1 4079
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_387
timestamp 1704896540
transform 1 0 3401 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_388
timestamp 1704896540
transform 1 0 3065 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_389
timestamp 1704896540
transform 1 0 2729 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_390
timestamp 1704896540
transform 1 0 2393 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_391
timestamp 1704896540
transform 1 0 1721 0 1 3743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_392
timestamp 1704896540
transform 1 0 1721 0 1 3407
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_393
timestamp 1704896540
transform 1 0 2057 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_394
timestamp 1704896540
transform 1 0 1721 0 1 3071
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_395
timestamp 1704896540
transform 1 0 1721 0 1 2735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_396
timestamp 1704896540
transform 1 0 1721 0 1 11135
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_397
timestamp 1704896540
transform 1 0 1721 0 1 10799
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_398
timestamp 1704896540
transform 1 0 1721 0 1 10463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_399
timestamp 1704896540
transform 1 0 1721 0 1 10127
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_400
timestamp 1704896540
transform 1 0 1721 0 1 9791
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_401
timestamp 1704896540
transform 1 0 1721 0 1 9455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_402
timestamp 1704896540
transform 1 0 1721 0 1 9119
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_403
timestamp 1704896540
transform 1 0 1721 0 1 8783
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_404
timestamp 1704896540
transform 1 0 1721 0 1 8447
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_405
timestamp 1704896540
transform 1 0 1721 0 1 8111
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_406
timestamp 1704896540
transform 1 0 1721 0 1 6095
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_407
timestamp 1704896540
transform 1 0 1721 0 1 7775
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_408
timestamp 1704896540
transform 1 0 1721 0 1 7439
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_409
timestamp 1704896540
transform 1 0 1721 0 1 7103
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_410
timestamp 1704896540
transform 1 0 1721 0 1 6767
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_411
timestamp 1704896540
transform 1 0 1721 0 1 6431
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_412
timestamp 1704896540
transform 1 0 1721 0 1 5759
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_413
timestamp 1704896540
transform 1 0 1721 0 1 14831
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_414
timestamp 1704896540
transform 1 0 1721 0 1 12143
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_415
timestamp 1704896540
transform 1 0 1721 0 1 11471
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_416
timestamp 1704896540
transform 1 0 1721 0 1 14495
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_417
timestamp 1704896540
transform 1 0 1721 0 1 14159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_418
timestamp 1704896540
transform 1 0 1721 0 1 13487
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_419
timestamp 1704896540
transform 1 0 1721 0 1 13151
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_420
timestamp 1704896540
transform 1 0 1721 0 1 12815
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_421
timestamp 1704896540
transform 1 0 1721 0 1 12479
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_422
timestamp 1704896540
transform 1 0 1721 0 1 16511
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_423
timestamp 1704896540
transform 1 0 1721 0 1 16175
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_424
timestamp 1704896540
transform 1 0 1721 0 1 15839
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_425
timestamp 1704896540
transform 1 0 1721 0 1 13823
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_426
timestamp 1704896540
transform 1 0 1721 0 1 15167
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_427
timestamp 1704896540
transform 1 0 1721 0 1 11807
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_428
timestamp 1704896540
transform 1 0 1721 0 1 15503
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_429
timestamp 1704896540
transform 1 0 1721 0 1 22223
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_430
timestamp 1704896540
transform 1 0 1721 0 1 21887
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_431
timestamp 1704896540
transform 1 0 1721 0 1 21551
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_432
timestamp 1704896540
transform 1 0 1721 0 1 21215
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_433
timestamp 1704896540
transform 1 0 1721 0 1 20879
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_434
timestamp 1704896540
transform 1 0 1721 0 1 20543
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_435
timestamp 1704896540
transform 1 0 1721 0 1 20207
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_436
timestamp 1704896540
transform 1 0 1721 0 1 19871
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_437
timestamp 1704896540
transform 1 0 1721 0 1 19535
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_438
timestamp 1704896540
transform 1 0 1721 0 1 19199
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_439
timestamp 1704896540
transform 1 0 1721 0 1 18863
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_440
timestamp 1704896540
transform 1 0 1721 0 1 18527
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_441
timestamp 1704896540
transform 1 0 1721 0 1 18191
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_442
timestamp 1704896540
transform 1 0 1721 0 1 17855
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_443
timestamp 1704896540
transform 1 0 1721 0 1 17519
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_444
timestamp 1704896540
transform 1 0 1721 0 1 17183
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_445
timestamp 1704896540
transform 1 0 1721 0 1 16847
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_446
timestamp 1704896540
transform 1 0 1721 0 1 25247
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_447
timestamp 1704896540
transform 1 0 1721 0 1 24911
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_448
timestamp 1704896540
transform 1 0 1721 0 1 24575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_449
timestamp 1704896540
transform 1 0 1721 0 1 22559
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_450
timestamp 1704896540
transform 1 0 1721 0 1 24239
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_451
timestamp 1704896540
transform 1 0 1721 0 1 23903
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_452
timestamp 1704896540
transform 1 0 1721 0 1 23567
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_453
timestamp 1704896540
transform 1 0 1721 0 1 23231
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_454
timestamp 1704896540
transform 1 0 1721 0 1 27599
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_455
timestamp 1704896540
transform 1 0 1721 0 1 27263
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_456
timestamp 1704896540
transform 1 0 1721 0 1 26927
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_457
timestamp 1704896540
transform 1 0 1721 0 1 26591
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_458
timestamp 1704896540
transform 1 0 1721 0 1 26255
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_459
timestamp 1704896540
transform 1 0 1721 0 1 25919
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_460
timestamp 1704896540
transform 1 0 1721 0 1 25583
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_461
timestamp 1704896540
transform 1 0 1721 0 1 22895
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_462
timestamp 1704896540
transform 1 0 1721 0 1 30287
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_463
timestamp 1704896540
transform 1 0 1721 0 1 29951
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_464
timestamp 1704896540
transform 1 0 1721 0 1 29615
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_465
timestamp 1704896540
transform 1 0 1721 0 1 29279
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_466
timestamp 1704896540
transform 1 0 1721 0 1 31631
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_467
timestamp 1704896540
transform 1 0 1721 0 1 28943
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_468
timestamp 1704896540
transform 1 0 1721 0 1 28607
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_469
timestamp 1704896540
transform 1 0 1721 0 1 28271
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_470
timestamp 1704896540
transform 1 0 1721 0 1 31295
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_471
timestamp 1704896540
transform 1 0 1721 0 1 30959
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_472
timestamp 1704896540
transform 1 0 1721 0 1 30623
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_473
timestamp 1704896540
transform 1 0 1721 0 1 33311
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_474
timestamp 1704896540
transform 1 0 1721 0 1 32975
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_475
timestamp 1704896540
transform 1 0 1721 0 1 32639
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_476
timestamp 1704896540
transform 1 0 1721 0 1 32303
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_477
timestamp 1704896540
transform 1 0 1721 0 1 31967
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_478
timestamp 1704896540
transform 1 0 1721 0 1 27935
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_479
timestamp 1704896540
transform 1 0 1721 0 1 34655
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_480
timestamp 1704896540
transform 1 0 1721 0 1 34319
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_481
timestamp 1704896540
transform 1 0 1721 0 1 38687
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_482
timestamp 1704896540
transform 1 0 1721 0 1 38351
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_483
timestamp 1704896540
transform 1 0 1721 0 1 38015
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_484
timestamp 1704896540
transform 1 0 1721 0 1 37679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_485
timestamp 1704896540
transform 1 0 1721 0 1 37343
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_486
timestamp 1704896540
transform 1 0 1721 0 1 37007
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_487
timestamp 1704896540
transform 1 0 1721 0 1 36671
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_488
timestamp 1704896540
transform 1 0 1721 0 1 36335
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_489
timestamp 1704896540
transform 1 0 1721 0 1 35999
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_490
timestamp 1704896540
transform 1 0 1721 0 1 35663
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_491
timestamp 1704896540
transform 1 0 1721 0 1 33983
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_492
timestamp 1704896540
transform 1 0 1721 0 1 35327
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_493
timestamp 1704896540
transform 1 0 1721 0 1 34991
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_494
timestamp 1704896540
transform 1 0 1721 0 1 33647
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_495
timestamp 1704896540
transform 1 0 1721 0 1 39695
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_496
timestamp 1704896540
transform 1 0 1721 0 1 39359
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_497
timestamp 1704896540
transform 1 0 1721 0 1 40031
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_498
timestamp 1704896540
transform 1 0 1721 0 1 44399
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_499
timestamp 1704896540
transform 1 0 1721 0 1 44063
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_500
timestamp 1704896540
transform 1 0 1721 0 1 43727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_501
timestamp 1704896540
transform 1 0 1721 0 1 43391
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_502
timestamp 1704896540
transform 1 0 1721 0 1 43055
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_503
timestamp 1704896540
transform 1 0 1721 0 1 42719
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_504
timestamp 1704896540
transform 1 0 1721 0 1 42383
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_505
timestamp 1704896540
transform 1 0 1721 0 1 42047
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_506
timestamp 1704896540
transform 1 0 1721 0 1 41711
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_507
timestamp 1704896540
transform 1 0 1721 0 1 41375
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_508
timestamp 1704896540
transform 1 0 1721 0 1 41039
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_509
timestamp 1704896540
transform 1 0 1721 0 1 40703
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_510
timestamp 1704896540
transform 1 0 1721 0 1 40367
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_511
timestamp 1704896540
transform 1 0 1721 0 1 39023
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_512
timestamp 1704896540
transform 1 0 22889 0 1 1727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_513
timestamp 1704896540
transform 1 0 1721 0 1 47759
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_514
timestamp 1704896540
transform 1 0 1721 0 1 47423
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_515
timestamp 1704896540
transform 1 0 1721 0 1 47087
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_516
timestamp 1704896540
transform 1 0 1721 0 1 46751
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_517
timestamp 1704896540
transform 1 0 1721 0 1 46415
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_518
timestamp 1704896540
transform 1 0 1721 0 1 46079
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_519
timestamp 1704896540
transform 1 0 1721 0 1 45743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_520
timestamp 1704896540
transform 1 0 1721 0 1 45407
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_521
timestamp 1704896540
transform 1 0 1721 0 1 45071
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_522
timestamp 1704896540
transform 1 0 1721 0 1 44735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_523
timestamp 1704896540
transform 1 0 1721 0 1 49775
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_524
timestamp 1704896540
transform 1 0 1721 0 1 49439
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_525
timestamp 1704896540
transform 1 0 1721 0 1 49103
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_526
timestamp 1704896540
transform 1 0 1721 0 1 48767
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_527
timestamp 1704896540
transform 1 0 1721 0 1 48431
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_528
timestamp 1704896540
transform 1 0 1721 0 1 48095
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_529
timestamp 1704896540
transform 1 0 1721 0 1 53471
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_530
timestamp 1704896540
transform 1 0 1721 0 1 53135
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_531
timestamp 1704896540
transform 1 0 1721 0 1 52799
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_532
timestamp 1704896540
transform 1 0 1721 0 1 52463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_533
timestamp 1704896540
transform 1 0 1721 0 1 52127
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_534
timestamp 1704896540
transform 1 0 1721 0 1 51791
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_535
timestamp 1704896540
transform 1 0 1721 0 1 51455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_536
timestamp 1704896540
transform 1 0 1721 0 1 51119
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_537
timestamp 1704896540
transform 1 0 1721 0 1 50783
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_538
timestamp 1704896540
transform 1 0 1721 0 1 50447
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_539
timestamp 1704896540
transform 1 0 1721 0 1 54815
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_540
timestamp 1704896540
transform 1 0 1721 0 1 55487
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_541
timestamp 1704896540
transform 1 0 1721 0 1 54143
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_542
timestamp 1704896540
transform 1 0 1721 0 1 53807
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_543
timestamp 1704896540
transform 1 0 1721 0 1 55151
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_544
timestamp 1704896540
transform 1 0 1721 0 1 54479
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_545
timestamp 1704896540
transform 1 0 1721 0 1 50111
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_546
timestamp 1704896540
transform 1 0 1721 0 1 55823
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_547
timestamp 1704896540
transform 1 0 1721 0 1 57839
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_548
timestamp 1704896540
transform 1 0 1721 0 1 56495
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_549
timestamp 1704896540
transform 1 0 1721 0 1 57503
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_550
timestamp 1704896540
transform 1 0 1721 0 1 57167
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_551
timestamp 1704896540
transform 1 0 1721 0 1 56159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_552
timestamp 1704896540
transform 1 0 1721 0 1 58847
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_553
timestamp 1704896540
transform 1 0 1721 0 1 58511
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_554
timestamp 1704896540
transform 1 0 1721 0 1 58175
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_555
timestamp 1704896540
transform 1 0 1721 0 1 60863
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_556
timestamp 1704896540
transform 1 0 1721 0 1 60527
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_557
timestamp 1704896540
transform 1 0 1721 0 1 60191
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_558
timestamp 1704896540
transform 1 0 1721 0 1 59855
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_559
timestamp 1704896540
transform 1 0 1721 0 1 56831
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_560
timestamp 1704896540
transform 1 0 1721 0 1 59519
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_561
timestamp 1704896540
transform 1 0 1721 0 1 59183
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_562
timestamp 1704896540
transform 1 0 1721 0 1 65231
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_563
timestamp 1704896540
transform 1 0 1721 0 1 64895
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_564
timestamp 1704896540
transform 1 0 1721 0 1 64559
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_565
timestamp 1704896540
transform 1 0 1721 0 1 64223
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_566
timestamp 1704896540
transform 1 0 1721 0 1 63887
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_567
timestamp 1704896540
transform 1 0 1721 0 1 63551
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_568
timestamp 1704896540
transform 1 0 1721 0 1 63215
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_569
timestamp 1704896540
transform 1 0 1721 0 1 62879
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_570
timestamp 1704896540
transform 1 0 1721 0 1 62543
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_571
timestamp 1704896540
transform 1 0 1721 0 1 62207
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_572
timestamp 1704896540
transform 1 0 1721 0 1 61871
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_573
timestamp 1704896540
transform 1 0 1721 0 1 61535
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_574
timestamp 1704896540
transform 1 0 1721 0 1 66575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_575
timestamp 1704896540
transform 1 0 1721 0 1 66239
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_576
timestamp 1704896540
transform 1 0 1721 0 1 65903
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_577
timestamp 1704896540
transform 1 0 1721 0 1 65567
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_578
timestamp 1704896540
transform 1 0 1721 0 1 61199
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_579
timestamp 1704896540
transform 1 0 1721 0 1 71615
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_580
timestamp 1704896540
transform 1 0 1721 0 1 71279
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_581
timestamp 1704896540
transform 1 0 1721 0 1 70943
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_582
timestamp 1704896540
transform 1 0 1721 0 1 70607
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_583
timestamp 1704896540
transform 1 0 1721 0 1 70271
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_584
timestamp 1704896540
transform 1 0 1721 0 1 69935
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_585
timestamp 1704896540
transform 1 0 1721 0 1 69599
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_586
timestamp 1704896540
transform 1 0 1721 0 1 69263
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_587
timestamp 1704896540
transform 1 0 1721 0 1 68927
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_588
timestamp 1704896540
transform 1 0 1721 0 1 68591
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_589
timestamp 1704896540
transform 1 0 1721 0 1 68255
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_590
timestamp 1704896540
transform 1 0 1721 0 1 67919
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_591
timestamp 1704896540
transform 1 0 1721 0 1 67583
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_592
timestamp 1704896540
transform 1 0 1721 0 1 67247
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_593
timestamp 1704896540
transform 1 0 1721 0 1 66911
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_594
timestamp 1704896540
transform 1 0 1721 0 1 71951
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_595
timestamp 1704896540
transform 1 0 1721 0 1 77663
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_596
timestamp 1704896540
transform 1 0 1721 0 1 77327
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_597
timestamp 1704896540
transform 1 0 1721 0 1 76991
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_598
timestamp 1704896540
transform 1 0 1721 0 1 76655
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_599
timestamp 1704896540
transform 1 0 1721 0 1 76319
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_600
timestamp 1704896540
transform 1 0 1721 0 1 75983
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_601
timestamp 1704896540
transform 1 0 1721 0 1 75647
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_602
timestamp 1704896540
transform 1 0 1721 0 1 75311
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_603
timestamp 1704896540
transform 1 0 1721 0 1 74975
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_604
timestamp 1704896540
transform 1 0 1721 0 1 74639
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_605
timestamp 1704896540
transform 1 0 1721 0 1 74303
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_606
timestamp 1704896540
transform 1 0 1721 0 1 73967
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_607
timestamp 1704896540
transform 1 0 1721 0 1 73631
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_608
timestamp 1704896540
transform 1 0 1721 0 1 73295
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_609
timestamp 1704896540
transform 1 0 1721 0 1 72959
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_610
timestamp 1704896540
transform 1 0 1721 0 1 72623
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_611
timestamp 1704896540
transform 1 0 1721 0 1 72287
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_612
timestamp 1704896540
transform 1 0 1721 0 1 82367
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_613
timestamp 1704896540
transform 1 0 1721 0 1 82031
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_614
timestamp 1704896540
transform 1 0 1721 0 1 81695
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_615
timestamp 1704896540
transform 1 0 1721 0 1 79007
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_616
timestamp 1704896540
transform 1 0 1721 0 1 78671
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_617
timestamp 1704896540
transform 1 0 1721 0 1 78335
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_618
timestamp 1704896540
transform 1 0 1721 0 1 77999
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_619
timestamp 1704896540
transform 1 0 1721 0 1 81359
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_620
timestamp 1704896540
transform 1 0 1721 0 1 81023
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_621
timestamp 1704896540
transform 1 0 1721 0 1 80687
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_622
timestamp 1704896540
transform 1 0 1721 0 1 80351
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_623
timestamp 1704896540
transform 1 0 1721 0 1 80015
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_624
timestamp 1704896540
transform 1 0 1721 0 1 79679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_625
timestamp 1704896540
transform 1 0 1721 0 1 79343
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_626
timestamp 1704896540
transform 1 0 1721 0 1 83039
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_627
timestamp 1704896540
transform 1 0 1721 0 1 82703
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_628
timestamp 1704896540
transform 1 0 1721 0 1 87071
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_629
timestamp 1704896540
transform 1 0 1721 0 1 86735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_630
timestamp 1704896540
transform 1 0 1721 0 1 86399
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_631
timestamp 1704896540
transform 1 0 1721 0 1 86063
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_632
timestamp 1704896540
transform 1 0 1721 0 1 85727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_633
timestamp 1704896540
transform 1 0 1721 0 1 85391
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_634
timestamp 1704896540
transform 1 0 1721 0 1 85055
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_635
timestamp 1704896540
transform 1 0 1721 0 1 84719
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_636
timestamp 1704896540
transform 1 0 1721 0 1 84383
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_637
timestamp 1704896540
transform 1 0 1721 0 1 84047
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_638
timestamp 1704896540
transform 1 0 1721 0 1 83711
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_639
timestamp 1704896540
transform 1 0 5753 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_640
timestamp 1704896540
transform 1 0 5417 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_641
timestamp 1704896540
transform 1 0 5081 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_642
timestamp 1704896540
transform 1 0 4745 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_643
timestamp 1704896540
transform 1 0 4409 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_644
timestamp 1704896540
transform 1 0 4073 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_645
timestamp 1704896540
transform 1 0 3737 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_646
timestamp 1704896540
transform 1 0 3401 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_647
timestamp 1704896540
transform 1 0 3065 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_648
timestamp 1704896540
transform 1 0 2729 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_649
timestamp 1704896540
transform 1 0 2393 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_650
timestamp 1704896540
transform 1 0 2057 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_651
timestamp 1704896540
transform 1 0 6089 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_652
timestamp 1704896540
transform 1 0 11465 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_653
timestamp 1704896540
transform 1 0 11129 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_654
timestamp 1704896540
transform 1 0 10793 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_655
timestamp 1704896540
transform 1 0 10457 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_656
timestamp 1704896540
transform 1 0 10121 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_657
timestamp 1704896540
transform 1 0 9785 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_658
timestamp 1704896540
transform 1 0 9449 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_659
timestamp 1704896540
transform 1 0 9113 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_660
timestamp 1704896540
transform 1 0 8777 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_661
timestamp 1704896540
transform 1 0 8441 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_662
timestamp 1704896540
transform 1 0 8105 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_663
timestamp 1704896540
transform 1 0 7769 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_664
timestamp 1704896540
transform 1 0 7433 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_665
timestamp 1704896540
transform 1 0 7097 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_666
timestamp 1704896540
transform 1 0 6761 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_667
timestamp 1704896540
transform 1 0 6425 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_668
timestamp 1704896540
transform 1 0 1721 0 1 83375
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_669
timestamp 1704896540
transform 1 0 22553 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_670
timestamp 1704896540
transform 1 0 22217 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_671
timestamp 1704896540
transform 1 0 21881 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_672
timestamp 1704896540
transform 1 0 21545 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_673
timestamp 1704896540
transform 1 0 21209 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_674
timestamp 1704896540
transform 1 0 20873 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_675
timestamp 1704896540
transform 1 0 20537 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_676
timestamp 1704896540
transform 1 0 20201 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_677
timestamp 1704896540
transform 1 0 19865 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_678
timestamp 1704896540
transform 1 0 19529 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_679
timestamp 1704896540
transform 1 0 19193 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_680
timestamp 1704896540
transform 1 0 18857 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_681
timestamp 1704896540
transform 1 0 18521 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_682
timestamp 1704896540
transform 1 0 18185 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_683
timestamp 1704896540
transform 1 0 17849 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_684
timestamp 1704896540
transform 1 0 17513 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_685
timestamp 1704896540
transform 1 0 17177 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_686
timestamp 1704896540
transform 1 0 16841 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_687
timestamp 1704896540
transform 1 0 16505 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_688
timestamp 1704896540
transform 1 0 16169 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_689
timestamp 1704896540
transform 1 0 15833 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_690
timestamp 1704896540
transform 1 0 15497 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_691
timestamp 1704896540
transform 1 0 15161 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_692
timestamp 1704896540
transform 1 0 14825 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_693
timestamp 1704896540
transform 1 0 14489 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_694
timestamp 1704896540
transform 1 0 14153 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_695
timestamp 1704896540
transform 1 0 13817 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_696
timestamp 1704896540
transform 1 0 13481 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_697
timestamp 1704896540
transform 1 0 13145 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_698
timestamp 1704896540
transform 1 0 12809 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_699
timestamp 1704896540
transform 1 0 12473 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_700
timestamp 1704896540
transform 1 0 12137 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_701
timestamp 1704896540
transform 1 0 11801 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_702
timestamp 1704896540
transform 1 0 30617 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_703
timestamp 1704896540
transform 1 0 30281 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_704
timestamp 1704896540
transform 1 0 29945 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_705
timestamp 1704896540
transform 1 0 29609 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_706
timestamp 1704896540
transform 1 0 29273 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_707
timestamp 1704896540
transform 1 0 28937 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_708
timestamp 1704896540
transform 1 0 28601 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_709
timestamp 1704896540
transform 1 0 28265 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_710
timestamp 1704896540
transform 1 0 27929 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_711
timestamp 1704896540
transform 1 0 27593 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_712
timestamp 1704896540
transform 1 0 27257 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_713
timestamp 1704896540
transform 1 0 26921 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_714
timestamp 1704896540
transform 1 0 26585 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_715
timestamp 1704896540
transform 1 0 26249 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_716
timestamp 1704896540
transform 1 0 25913 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_717
timestamp 1704896540
transform 1 0 25577 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_718
timestamp 1704896540
transform 1 0 25241 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_719
timestamp 1704896540
transform 1 0 24905 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_720
timestamp 1704896540
transform 1 0 24569 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_721
timestamp 1704896540
transform 1 0 24233 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_722
timestamp 1704896540
transform 1 0 23897 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_723
timestamp 1704896540
transform 1 0 23561 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_724
timestamp 1704896540
transform 1 0 23225 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_725
timestamp 1704896540
transform 1 0 33977 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_726
timestamp 1704896540
transform 1 0 33641 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_727
timestamp 1704896540
transform 1 0 33305 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_728
timestamp 1704896540
transform 1 0 32969 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_729
timestamp 1704896540
transform 1 0 32633 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_730
timestamp 1704896540
transform 1 0 32297 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_731
timestamp 1704896540
transform 1 0 31961 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_732
timestamp 1704896540
transform 1 0 31625 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_733
timestamp 1704896540
transform 1 0 31289 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_734
timestamp 1704896540
transform 1 0 30953 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_735
timestamp 1704896540
transform 1 0 44057 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_736
timestamp 1704896540
transform 1 0 43721 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_737
timestamp 1704896540
transform 1 0 43385 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_738
timestamp 1704896540
transform 1 0 43049 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_739
timestamp 1704896540
transform 1 0 42713 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_740
timestamp 1704896540
transform 1 0 42377 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_741
timestamp 1704896540
transform 1 0 42041 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_742
timestamp 1704896540
transform 1 0 41705 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_743
timestamp 1704896540
transform 1 0 41369 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_744
timestamp 1704896540
transform 1 0 41033 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_745
timestamp 1704896540
transform 1 0 40697 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_746
timestamp 1704896540
transform 1 0 40361 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_747
timestamp 1704896540
transform 1 0 40025 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_748
timestamp 1704896540
transform 1 0 39689 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_749
timestamp 1704896540
transform 1 0 39353 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_750
timestamp 1704896540
transform 1 0 39017 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_751
timestamp 1704896540
transform 1 0 38681 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_752
timestamp 1704896540
transform 1 0 38345 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_753
timestamp 1704896540
transform 1 0 38009 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_754
timestamp 1704896540
transform 1 0 37673 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_755
timestamp 1704896540
transform 1 0 37337 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_756
timestamp 1704896540
transform 1 0 37001 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_757
timestamp 1704896540
transform 1 0 36665 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_758
timestamp 1704896540
transform 1 0 36329 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_759
timestamp 1704896540
transform 1 0 35993 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_760
timestamp 1704896540
transform 1 0 35657 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_761
timestamp 1704896540
transform 1 0 35321 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_762
timestamp 1704896540
transform 1 0 34985 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_763
timestamp 1704896540
transform 1 0 34649 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_764
timestamp 1704896540
transform 1 0 34313 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_765
timestamp 1704896540
transform 1 0 45401 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_766
timestamp 1704896540
transform 1 0 45065 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_767
timestamp 1704896540
transform 1 0 44729 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_768
timestamp 1704896540
transform 1 0 44393 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_769
timestamp 1704896540
transform 1 0 22889 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_770
timestamp 1704896540
transform 1 0 89219 0 1 47423
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_771
timestamp 1704896540
transform 1 0 89219 0 1 47087
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_772
timestamp 1704896540
transform 1 0 89219 0 1 46751
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_773
timestamp 1704896540
transform 1 0 89219 0 1 46415
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_774
timestamp 1704896540
transform 1 0 89219 0 1 48431
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_775
timestamp 1704896540
transform 1 0 89219 0 1 49775
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_776
timestamp 1704896540
transform 1 0 89219 0 1 49439
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_777
timestamp 1704896540
transform 1 0 89219 0 1 46079
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_778
timestamp 1704896540
transform 1 0 89219 0 1 49103
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_779
timestamp 1704896540
transform 1 0 89219 0 1 48095
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_780
timestamp 1704896540
transform 1 0 89219 0 1 45743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_781
timestamp 1704896540
transform 1 0 89219 0 1 47759
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_782
timestamp 1704896540
transform 1 0 89219 0 1 45407
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_783
timestamp 1704896540
transform 1 0 89219 0 1 48767
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_784
timestamp 1704896540
transform 1 0 89219 0 1 45071
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_785
timestamp 1704896540
transform 1 0 89219 0 1 44735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_786
timestamp 1704896540
transform 1 0 89219 0 1 55487
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_787
timestamp 1704896540
transform 1 0 89219 0 1 55151
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_788
timestamp 1704896540
transform 1 0 89219 0 1 54815
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_789
timestamp 1704896540
transform 1 0 89219 0 1 54479
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_790
timestamp 1704896540
transform 1 0 89219 0 1 54143
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_791
timestamp 1704896540
transform 1 0 89219 0 1 53807
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_792
timestamp 1704896540
transform 1 0 89219 0 1 53471
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_793
timestamp 1704896540
transform 1 0 89219 0 1 50783
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_794
timestamp 1704896540
transform 1 0 89219 0 1 52127
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_795
timestamp 1704896540
transform 1 0 89219 0 1 51791
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_796
timestamp 1704896540
transform 1 0 89219 0 1 50447
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_797
timestamp 1704896540
transform 1 0 89219 0 1 51455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_798
timestamp 1704896540
transform 1 0 89219 0 1 51119
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_799
timestamp 1704896540
transform 1 0 89219 0 1 53135
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_800
timestamp 1704896540
transform 1 0 89219 0 1 52799
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_801
timestamp 1704896540
transform 1 0 89219 0 1 52463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_802
timestamp 1704896540
transform 1 0 89219 0 1 50111
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_803
timestamp 1704896540
transform 1 0 89219 0 1 56159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_804
timestamp 1704896540
transform 1 0 89219 0 1 57503
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_805
timestamp 1704896540
transform 1 0 89219 0 1 55823
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_806
timestamp 1704896540
transform 1 0 89219 0 1 57167
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_807
timestamp 1704896540
transform 1 0 89219 0 1 56831
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_808
timestamp 1704896540
transform 1 0 89219 0 1 56495
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_809
timestamp 1704896540
transform 1 0 89219 0 1 60863
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_810
timestamp 1704896540
transform 1 0 89219 0 1 60527
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_811
timestamp 1704896540
transform 1 0 89219 0 1 60191
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_812
timestamp 1704896540
transform 1 0 89219 0 1 59855
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_813
timestamp 1704896540
transform 1 0 89219 0 1 59519
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_814
timestamp 1704896540
transform 1 0 89219 0 1 59183
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_815
timestamp 1704896540
transform 1 0 89219 0 1 58847
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_816
timestamp 1704896540
transform 1 0 89219 0 1 58511
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_817
timestamp 1704896540
transform 1 0 89219 0 1 58175
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_818
timestamp 1704896540
transform 1 0 89219 0 1 57839
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_819
timestamp 1704896540
transform 1 0 89219 0 1 66575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_820
timestamp 1704896540
transform 1 0 89219 0 1 66239
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_821
timestamp 1704896540
transform 1 0 89219 0 1 65903
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_822
timestamp 1704896540
transform 1 0 89219 0 1 65567
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_823
timestamp 1704896540
transform 1 0 89219 0 1 65231
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_824
timestamp 1704896540
transform 1 0 89219 0 1 64895
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_825
timestamp 1704896540
transform 1 0 89219 0 1 64559
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_826
timestamp 1704896540
transform 1 0 89219 0 1 64223
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_827
timestamp 1704896540
transform 1 0 89219 0 1 63887
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_828
timestamp 1704896540
transform 1 0 89219 0 1 63551
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_829
timestamp 1704896540
transform 1 0 89219 0 1 63215
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_830
timestamp 1704896540
transform 1 0 89219 0 1 62879
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_831
timestamp 1704896540
transform 1 0 89219 0 1 62543
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_832
timestamp 1704896540
transform 1 0 89219 0 1 62207
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_833
timestamp 1704896540
transform 1 0 89219 0 1 61871
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_834
timestamp 1704896540
transform 1 0 89219 0 1 61535
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_835
timestamp 1704896540
transform 1 0 89219 0 1 61199
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_836
timestamp 1704896540
transform 1 0 45737 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_837
timestamp 1704896540
transform 1 0 55481 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_838
timestamp 1704896540
transform 1 0 55145 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_839
timestamp 1704896540
transform 1 0 54809 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_840
timestamp 1704896540
transform 1 0 54473 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_841
timestamp 1704896540
transform 1 0 54137 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_842
timestamp 1704896540
transform 1 0 53801 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_843
timestamp 1704896540
transform 1 0 53465 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_844
timestamp 1704896540
transform 1 0 53129 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_845
timestamp 1704896540
transform 1 0 52793 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_846
timestamp 1704896540
transform 1 0 52457 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_847
timestamp 1704896540
transform 1 0 52121 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_848
timestamp 1704896540
transform 1 0 51785 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_849
timestamp 1704896540
transform 1 0 51449 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_850
timestamp 1704896540
transform 1 0 51113 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_851
timestamp 1704896540
transform 1 0 50777 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_852
timestamp 1704896540
transform 1 0 50441 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_853
timestamp 1704896540
transform 1 0 50105 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_854
timestamp 1704896540
transform 1 0 49769 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_855
timestamp 1704896540
transform 1 0 49433 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_856
timestamp 1704896540
transform 1 0 49097 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_857
timestamp 1704896540
transform 1 0 48761 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_858
timestamp 1704896540
transform 1 0 47753 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_859
timestamp 1704896540
transform 1 0 47417 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_860
timestamp 1704896540
transform 1 0 47081 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_861
timestamp 1704896540
transform 1 0 46745 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_862
timestamp 1704896540
transform 1 0 46409 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_863
timestamp 1704896540
transform 1 0 46073 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_864
timestamp 1704896540
transform 1 0 48425 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_865
timestamp 1704896540
transform 1 0 48089 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_866
timestamp 1704896540
transform 1 0 56489 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_867
timestamp 1704896540
transform 1 0 56153 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_868
timestamp 1704896540
transform 1 0 55817 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_869
timestamp 1704896540
transform 1 0 67913 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_870
timestamp 1704896540
transform 1 0 67577 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_871
timestamp 1704896540
transform 1 0 67241 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_872
timestamp 1704896540
transform 1 0 66905 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_873
timestamp 1704896540
transform 1 0 66569 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_874
timestamp 1704896540
transform 1 0 66233 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_875
timestamp 1704896540
transform 1 0 65897 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_876
timestamp 1704896540
transform 1 0 65561 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_877
timestamp 1704896540
transform 1 0 65225 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_878
timestamp 1704896540
transform 1 0 64889 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_879
timestamp 1704896540
transform 1 0 64553 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_880
timestamp 1704896540
transform 1 0 64217 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_881
timestamp 1704896540
transform 1 0 63881 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_882
timestamp 1704896540
transform 1 0 63545 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_883
timestamp 1704896540
transform 1 0 63209 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_884
timestamp 1704896540
transform 1 0 62873 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_885
timestamp 1704896540
transform 1 0 62537 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_886
timestamp 1704896540
transform 1 0 62201 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_887
timestamp 1704896540
transform 1 0 61865 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_888
timestamp 1704896540
transform 1 0 61529 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_889
timestamp 1704896540
transform 1 0 61193 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_890
timestamp 1704896540
transform 1 0 60857 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_891
timestamp 1704896540
transform 1 0 60521 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_892
timestamp 1704896540
transform 1 0 60185 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_893
timestamp 1704896540
transform 1 0 59849 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_894
timestamp 1704896540
transform 1 0 59513 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_895
timestamp 1704896540
transform 1 0 59177 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_896
timestamp 1704896540
transform 1 0 58841 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_897
timestamp 1704896540
transform 1 0 58505 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_898
timestamp 1704896540
transform 1 0 58169 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_899
timestamp 1704896540
transform 1 0 57833 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_900
timestamp 1704896540
transform 1 0 57497 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_901
timestamp 1704896540
transform 1 0 57161 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_902
timestamp 1704896540
transform 1 0 56825 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_903
timestamp 1704896540
transform 1 0 89219 0 1 70943
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_904
timestamp 1704896540
transform 1 0 89219 0 1 70607
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_905
timestamp 1704896540
transform 1 0 89219 0 1 70271
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_906
timestamp 1704896540
transform 1 0 89219 0 1 69935
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_907
timestamp 1704896540
transform 1 0 89219 0 1 69599
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_908
timestamp 1704896540
transform 1 0 89219 0 1 69263
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_909
timestamp 1704896540
transform 1 0 89219 0 1 68927
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_910
timestamp 1704896540
transform 1 0 89219 0 1 68591
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_911
timestamp 1704896540
transform 1 0 89219 0 1 68255
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_912
timestamp 1704896540
transform 1 0 89219 0 1 67919
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_913
timestamp 1704896540
transform 1 0 89219 0 1 67583
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_914
timestamp 1704896540
transform 1 0 89219 0 1 67247
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_915
timestamp 1704896540
transform 1 0 89219 0 1 66911
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_916
timestamp 1704896540
transform 1 0 89219 0 1 71951
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_917
timestamp 1704896540
transform 1 0 89219 0 1 71615
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_918
timestamp 1704896540
transform 1 0 89219 0 1 71279
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_919
timestamp 1704896540
transform 1 0 89219 0 1 77663
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_920
timestamp 1704896540
transform 1 0 89219 0 1 77327
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_921
timestamp 1704896540
transform 1 0 89219 0 1 76991
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_922
timestamp 1704896540
transform 1 0 89219 0 1 76655
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_923
timestamp 1704896540
transform 1 0 89219 0 1 76319
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_924
timestamp 1704896540
transform 1 0 89219 0 1 75983
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_925
timestamp 1704896540
transform 1 0 89219 0 1 75647
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_926
timestamp 1704896540
transform 1 0 89219 0 1 75311
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_927
timestamp 1704896540
transform 1 0 89219 0 1 74975
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_928
timestamp 1704896540
transform 1 0 89219 0 1 74639
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_929
timestamp 1704896540
transform 1 0 89219 0 1 74303
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_930
timestamp 1704896540
transform 1 0 89219 0 1 73967
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_931
timestamp 1704896540
transform 1 0 89219 0 1 73631
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_932
timestamp 1704896540
transform 1 0 89219 0 1 73295
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_933
timestamp 1704896540
transform 1 0 89219 0 1 72959
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_934
timestamp 1704896540
transform 1 0 89219 0 1 72623
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_935
timestamp 1704896540
transform 1 0 89219 0 1 72287
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_936
timestamp 1704896540
transform 1 0 71609 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_937
timestamp 1704896540
transform 1 0 68585 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_938
timestamp 1704896540
transform 1 0 68249 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_939
timestamp 1704896540
transform 1 0 72617 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_940
timestamp 1704896540
transform 1 0 71273 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_941
timestamp 1704896540
transform 1 0 70937 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_942
timestamp 1704896540
transform 1 0 70601 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_943
timestamp 1704896540
transform 1 0 70265 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_944
timestamp 1704896540
transform 1 0 69929 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_945
timestamp 1704896540
transform 1 0 69593 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_946
timestamp 1704896540
transform 1 0 69257 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_947
timestamp 1704896540
transform 1 0 68921 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_948
timestamp 1704896540
transform 1 0 72281 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_949
timestamp 1704896540
transform 1 0 71945 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_950
timestamp 1704896540
transform 1 0 73625 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_951
timestamp 1704896540
transform 1 0 73289 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_952
timestamp 1704896540
transform 1 0 72953 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_953
timestamp 1704896540
transform 1 0 73961 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_954
timestamp 1704896540
transform 1 0 79337 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_955
timestamp 1704896540
transform 1 0 79001 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_956
timestamp 1704896540
transform 1 0 78665 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_957
timestamp 1704896540
transform 1 0 78329 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_958
timestamp 1704896540
transform 1 0 77993 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_959
timestamp 1704896540
transform 1 0 77657 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_960
timestamp 1704896540
transform 1 0 77321 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_961
timestamp 1704896540
transform 1 0 76985 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_962
timestamp 1704896540
transform 1 0 76649 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_963
timestamp 1704896540
transform 1 0 76313 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_964
timestamp 1704896540
transform 1 0 75977 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_965
timestamp 1704896540
transform 1 0 75641 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_966
timestamp 1704896540
transform 1 0 75305 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_967
timestamp 1704896540
transform 1 0 74969 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_968
timestamp 1704896540
transform 1 0 74633 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_969
timestamp 1704896540
transform 1 0 74297 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_970
timestamp 1704896540
transform 1 0 89219 0 1 79679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_971
timestamp 1704896540
transform 1 0 89219 0 1 79343
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_972
timestamp 1704896540
transform 1 0 89219 0 1 79007
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_973
timestamp 1704896540
transform 1 0 89219 0 1 78671
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_974
timestamp 1704896540
transform 1 0 89219 0 1 78335
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_975
timestamp 1704896540
transform 1 0 89219 0 1 77999
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_976
timestamp 1704896540
transform 1 0 89219 0 1 83039
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_977
timestamp 1704896540
transform 1 0 89219 0 1 82703
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_978
timestamp 1704896540
transform 1 0 89219 0 1 82367
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_979
timestamp 1704896540
transform 1 0 89219 0 1 82031
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_980
timestamp 1704896540
transform 1 0 89219 0 1 81695
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_981
timestamp 1704896540
transform 1 0 89219 0 1 81359
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_982
timestamp 1704896540
transform 1 0 89219 0 1 81023
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_983
timestamp 1704896540
transform 1 0 89219 0 1 80687
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_984
timestamp 1704896540
transform 1 0 89219 0 1 80351
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_985
timestamp 1704896540
transform 1 0 89219 0 1 80015
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_986
timestamp 1704896540
transform 1 0 79673 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_987
timestamp 1704896540
transform 1 0 82025 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_988
timestamp 1704896540
transform 1 0 81689 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_989
timestamp 1704896540
transform 1 0 81353 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_990
timestamp 1704896540
transform 1 0 81017 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_991
timestamp 1704896540
transform 1 0 80681 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_992
timestamp 1704896540
transform 1 0 80345 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_993
timestamp 1704896540
transform 1 0 80009 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_994
timestamp 1704896540
transform 1 0 84713 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_995
timestamp 1704896540
transform 1 0 84377 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_996
timestamp 1704896540
transform 1 0 84041 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_997
timestamp 1704896540
transform 1 0 83705 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_998
timestamp 1704896540
transform 1 0 83369 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_999
timestamp 1704896540
transform 1 0 83033 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_1000
timestamp 1704896540
transform 1 0 82697 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_1001
timestamp 1704896540
transform 1 0 82361 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_1002
timestamp 1704896540
transform 1 0 89219 0 1 87071
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_1003
timestamp 1704896540
transform 1 0 89219 0 1 86735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_1004
timestamp 1704896540
transform 1 0 89219 0 1 86399
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_1005
timestamp 1704896540
transform 1 0 89219 0 1 86063
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_1006
timestamp 1704896540
transform 1 0 89219 0 1 85727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_1007
timestamp 1704896540
transform 1 0 89219 0 1 85391
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_1008
timestamp 1704896540
transform 1 0 89219 0 1 85055
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_1009
timestamp 1704896540
transform 1 0 89219 0 1 84719
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_1010
timestamp 1704896540
transform 1 0 89219 0 1 84383
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_1011
timestamp 1704896540
transform 1 0 89219 0 1 84047
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_1012
timestamp 1704896540
transform 1 0 89219 0 1 83711
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_1013
timestamp 1704896540
transform 1 0 85385 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_1014
timestamp 1704896540
transform 1 0 88745 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_1015
timestamp 1704896540
transform 1 0 88409 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_1016
timestamp 1704896540
transform 1 0 88073 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_1017
timestamp 1704896540
transform 1 0 87737 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_1018
timestamp 1704896540
transform 1 0 87401 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_1019
timestamp 1704896540
transform 1 0 87065 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_1020
timestamp 1704896540
transform 1 0 86729 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_1021
timestamp 1704896540
transform 1 0 86393 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_1022
timestamp 1704896540
transform 1 0 86057 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_1023
timestamp 1704896540
transform 1 0 85721 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_1024
timestamp 1704896540
transform 1 0 89219 0 1 83375
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_13_1025
timestamp 1704896540
transform 1 0 85049 0 1 87455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_0
timestamp 1704896540
transform 1 0 89215 0 1 5431
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_1
timestamp 1704896540
transform 1 0 89215 0 1 5095
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_2
timestamp 1704896540
transform 1 0 89215 0 1 4759
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_3
timestamp 1704896540
transform 1 0 89215 0 1 4423
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_4
timestamp 1704896540
transform 1 0 89215 0 1 4087
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_5
timestamp 1704896540
transform 1 0 89215 0 1 3751
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_6
timestamp 1704896540
transform 1 0 89215 0 1 3415
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_7
timestamp 1704896540
transform 1 0 89215 0 1 3079
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_8
timestamp 1704896540
transform 1 0 89215 0 1 2743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_9
timestamp 1704896540
transform 1 0 88741 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_10
timestamp 1704896540
transform 1 0 89215 0 1 2407
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_11
timestamp 1704896540
transform 1 0 88405 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_12
timestamp 1704896540
transform 1 0 89215 0 1 2071
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_13
timestamp 1704896540
transform 1 0 88069 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_14
timestamp 1704896540
transform 1 0 87733 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_15
timestamp 1704896540
transform 1 0 87397 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_16
timestamp 1704896540
transform 1 0 87061 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_17
timestamp 1704896540
transform 1 0 86725 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_18
timestamp 1704896540
transform 1 0 86389 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_19
timestamp 1704896540
transform 1 0 86053 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_20
timestamp 1704896540
transform 1 0 85717 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_21
timestamp 1704896540
transform 1 0 85381 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_22
timestamp 1704896540
transform 1 0 84709 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_23
timestamp 1704896540
transform 1 0 84373 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_24
timestamp 1704896540
transform 1 0 84037 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_25
timestamp 1704896540
transform 1 0 83701 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_26
timestamp 1704896540
transform 1 0 83365 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_27
timestamp 1704896540
transform 1 0 83029 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_28
timestamp 1704896540
transform 1 0 82693 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_29
timestamp 1704896540
transform 1 0 82357 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_30
timestamp 1704896540
transform 1 0 82021 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_31
timestamp 1704896540
transform 1 0 81685 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_32
timestamp 1704896540
transform 1 0 81349 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_33
timestamp 1704896540
transform 1 0 81013 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_34
timestamp 1704896540
transform 1 0 80677 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_35
timestamp 1704896540
transform 1 0 80341 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_36
timestamp 1704896540
transform 1 0 80005 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_37
timestamp 1704896540
transform 1 0 79669 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_38
timestamp 1704896540
transform 1 0 85045 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_39
timestamp 1704896540
transform 1 0 89215 0 1 9463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_40
timestamp 1704896540
transform 1 0 89215 0 1 9127
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_41
timestamp 1704896540
transform 1 0 89215 0 1 8791
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_42
timestamp 1704896540
transform 1 0 89215 0 1 8455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_43
timestamp 1704896540
transform 1 0 89215 0 1 8119
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_44
timestamp 1704896540
transform 1 0 89215 0 1 7783
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_45
timestamp 1704896540
transform 1 0 89215 0 1 7447
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_46
timestamp 1704896540
transform 1 0 89215 0 1 7111
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_47
timestamp 1704896540
transform 1 0 89215 0 1 6775
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_48
timestamp 1704896540
transform 1 0 89215 0 1 6439
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_49
timestamp 1704896540
transform 1 0 89215 0 1 6103
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_50
timestamp 1704896540
transform 1 0 89215 0 1 10135
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_51
timestamp 1704896540
transform 1 0 89215 0 1 11143
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_52
timestamp 1704896540
transform 1 0 89215 0 1 10807
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_53
timestamp 1704896540
transform 1 0 89215 0 1 9799
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_54
timestamp 1704896540
transform 1 0 89215 0 1 10471
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_55
timestamp 1704896540
transform 1 0 89215 0 1 5767
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_56
timestamp 1704896540
transform 1 0 73957 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_57
timestamp 1704896540
transform 1 0 73621 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_58
timestamp 1704896540
transform 1 0 73285 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_59
timestamp 1704896540
transform 1 0 72949 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_60
timestamp 1704896540
transform 1 0 72613 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_61
timestamp 1704896540
transform 1 0 72277 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_62
timestamp 1704896540
transform 1 0 71941 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_63
timestamp 1704896540
transform 1 0 68917 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_64
timestamp 1704896540
transform 1 0 71605 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_65
timestamp 1704896540
transform 1 0 71269 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_66
timestamp 1704896540
transform 1 0 70933 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_67
timestamp 1704896540
transform 1 0 68245 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_68
timestamp 1704896540
transform 1 0 70597 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_69
timestamp 1704896540
transform 1 0 70261 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_70
timestamp 1704896540
transform 1 0 69925 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_71
timestamp 1704896540
transform 1 0 68581 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_72
timestamp 1704896540
transform 1 0 69253 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_73
timestamp 1704896540
transform 1 0 69589 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_74
timestamp 1704896540
transform 1 0 79333 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_75
timestamp 1704896540
transform 1 0 78997 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_76
timestamp 1704896540
transform 1 0 78661 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_77
timestamp 1704896540
transform 1 0 78325 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_78
timestamp 1704896540
transform 1 0 77989 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_79
timestamp 1704896540
transform 1 0 77653 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_80
timestamp 1704896540
transform 1 0 77317 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_81
timestamp 1704896540
transform 1 0 76981 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_82
timestamp 1704896540
transform 1 0 76645 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_83
timestamp 1704896540
transform 1 0 76309 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_84
timestamp 1704896540
transform 1 0 75973 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_85
timestamp 1704896540
transform 1 0 75637 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_86
timestamp 1704896540
transform 1 0 75301 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_87
timestamp 1704896540
transform 1 0 74965 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_88
timestamp 1704896540
transform 1 0 74629 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_89
timestamp 1704896540
transform 1 0 74293 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_90
timestamp 1704896540
transform 1 0 89215 0 1 13831
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_91
timestamp 1704896540
transform 1 0 89215 0 1 13495
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_92
timestamp 1704896540
transform 1 0 89215 0 1 13159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_93
timestamp 1704896540
transform 1 0 89215 0 1 12823
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_94
timestamp 1704896540
transform 1 0 89215 0 1 12487
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_95
timestamp 1704896540
transform 1 0 89215 0 1 12151
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_96
timestamp 1704896540
transform 1 0 89215 0 1 11815
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_97
timestamp 1704896540
transform 1 0 89215 0 1 11479
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_98
timestamp 1704896540
transform 1 0 89215 0 1 16519
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_99
timestamp 1704896540
transform 1 0 89215 0 1 16183
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_100
timestamp 1704896540
transform 1 0 89215 0 1 15847
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_101
timestamp 1704896540
transform 1 0 89215 0 1 15511
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_102
timestamp 1704896540
transform 1 0 89215 0 1 15175
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_103
timestamp 1704896540
transform 1 0 89215 0 1 14839
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_104
timestamp 1704896540
transform 1 0 89215 0 1 14503
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_105
timestamp 1704896540
transform 1 0 89215 0 1 14167
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_106
timestamp 1704896540
transform 1 0 89215 0 1 22231
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_107
timestamp 1704896540
transform 1 0 89215 0 1 21895
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_108
timestamp 1704896540
transform 1 0 89215 0 1 21559
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_109
timestamp 1704896540
transform 1 0 89215 0 1 21223
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_110
timestamp 1704896540
transform 1 0 89215 0 1 20887
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_111
timestamp 1704896540
transform 1 0 89215 0 1 20551
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_112
timestamp 1704896540
transform 1 0 89215 0 1 20215
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_113
timestamp 1704896540
transform 1 0 89215 0 1 19879
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_114
timestamp 1704896540
transform 1 0 89215 0 1 19543
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_115
timestamp 1704896540
transform 1 0 89215 0 1 19207
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_116
timestamp 1704896540
transform 1 0 89215 0 1 18871
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_117
timestamp 1704896540
transform 1 0 89215 0 1 18535
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_118
timestamp 1704896540
transform 1 0 89215 0 1 18199
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_119
timestamp 1704896540
transform 1 0 89215 0 1 17863
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_120
timestamp 1704896540
transform 1 0 89215 0 1 17527
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_121
timestamp 1704896540
transform 1 0 89215 0 1 17191
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_122
timestamp 1704896540
transform 1 0 89215 0 1 16855
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_123
timestamp 1704896540
transform 1 0 67573 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_124
timestamp 1704896540
transform 1 0 67237 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_125
timestamp 1704896540
transform 1 0 66901 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_126
timestamp 1704896540
transform 1 0 66565 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_127
timestamp 1704896540
transform 1 0 66229 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_128
timestamp 1704896540
transform 1 0 65893 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_129
timestamp 1704896540
transform 1 0 65557 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_130
timestamp 1704896540
transform 1 0 65221 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_131
timestamp 1704896540
transform 1 0 64885 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_132
timestamp 1704896540
transform 1 0 64549 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_133
timestamp 1704896540
transform 1 0 64213 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_134
timestamp 1704896540
transform 1 0 63877 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_135
timestamp 1704896540
transform 1 0 57829 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_136
timestamp 1704896540
transform 1 0 60181 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_137
timestamp 1704896540
transform 1 0 63541 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_138
timestamp 1704896540
transform 1 0 63205 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_139
timestamp 1704896540
transform 1 0 58837 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_140
timestamp 1704896540
transform 1 0 59845 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_141
timestamp 1704896540
transform 1 0 58501 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_142
timestamp 1704896540
transform 1 0 59509 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_143
timestamp 1704896540
transform 1 0 62869 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_144
timestamp 1704896540
transform 1 0 62533 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_145
timestamp 1704896540
transform 1 0 62197 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_146
timestamp 1704896540
transform 1 0 61861 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_147
timestamp 1704896540
transform 1 0 61525 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_148
timestamp 1704896540
transform 1 0 61189 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_149
timestamp 1704896540
transform 1 0 60853 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_150
timestamp 1704896540
transform 1 0 57157 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_151
timestamp 1704896540
transform 1 0 58165 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_152
timestamp 1704896540
transform 1 0 57493 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_153
timestamp 1704896540
transform 1 0 60517 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_154
timestamp 1704896540
transform 1 0 59173 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_155
timestamp 1704896540
transform 1 0 67909 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_156
timestamp 1704896540
transform 1 0 46405 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_157
timestamp 1704896540
transform 1 0 48421 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_158
timestamp 1704896540
transform 1 0 46069 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_159
timestamp 1704896540
transform 1 0 49093 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_160
timestamp 1704896540
transform 1 0 54805 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_161
timestamp 1704896540
transform 1 0 48085 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_162
timestamp 1704896540
transform 1 0 54469 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_163
timestamp 1704896540
transform 1 0 47749 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_164
timestamp 1704896540
transform 1 0 56485 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_165
timestamp 1704896540
transform 1 0 56149 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_166
timestamp 1704896540
transform 1 0 54133 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_167
timestamp 1704896540
transform 1 0 53797 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_168
timestamp 1704896540
transform 1 0 50437 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_169
timestamp 1704896540
transform 1 0 52453 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_170
timestamp 1704896540
transform 1 0 50101 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_171
timestamp 1704896540
transform 1 0 49765 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_172
timestamp 1704896540
transform 1 0 51109 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_173
timestamp 1704896540
transform 1 0 52117 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_174
timestamp 1704896540
transform 1 0 51445 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_175
timestamp 1704896540
transform 1 0 48757 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_176
timestamp 1704896540
transform 1 0 53461 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_177
timestamp 1704896540
transform 1 0 45733 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_178
timestamp 1704896540
transform 1 0 51781 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_179
timestamp 1704896540
transform 1 0 52789 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_180
timestamp 1704896540
transform 1 0 53125 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_181
timestamp 1704896540
transform 1 0 47413 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_182
timestamp 1704896540
transform 1 0 55813 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_183
timestamp 1704896540
transform 1 0 50773 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_184
timestamp 1704896540
transform 1 0 47077 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_185
timestamp 1704896540
transform 1 0 55477 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_186
timestamp 1704896540
transform 1 0 46741 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_187
timestamp 1704896540
transform 1 0 55141 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_188
timestamp 1704896540
transform 1 0 49429 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_189
timestamp 1704896540
transform 1 0 56821 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_190
timestamp 1704896540
transform 1 0 89215 0 1 25591
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_191
timestamp 1704896540
transform 1 0 89215 0 1 25255
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_192
timestamp 1704896540
transform 1 0 89215 0 1 24919
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_193
timestamp 1704896540
transform 1 0 89215 0 1 24583
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_194
timestamp 1704896540
transform 1 0 89215 0 1 24247
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_195
timestamp 1704896540
transform 1 0 89215 0 1 22903
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_196
timestamp 1704896540
transform 1 0 89215 0 1 22567
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_197
timestamp 1704896540
transform 1 0 89215 0 1 27607
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_198
timestamp 1704896540
transform 1 0 89215 0 1 27271
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_199
timestamp 1704896540
transform 1 0 89215 0 1 26935
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_200
timestamp 1704896540
transform 1 0 89215 0 1 26599
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_201
timestamp 1704896540
transform 1 0 89215 0 1 26263
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_202
timestamp 1704896540
transform 1 0 89215 0 1 23911
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_203
timestamp 1704896540
transform 1 0 89215 0 1 23575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_204
timestamp 1704896540
transform 1 0 89215 0 1 23239
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_205
timestamp 1704896540
transform 1 0 89215 0 1 25927
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_206
timestamp 1704896540
transform 1 0 89215 0 1 29959
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_207
timestamp 1704896540
transform 1 0 89215 0 1 29623
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_208
timestamp 1704896540
transform 1 0 89215 0 1 29287
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_209
timestamp 1704896540
transform 1 0 89215 0 1 28951
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_210
timestamp 1704896540
transform 1 0 89215 0 1 28615
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_211
timestamp 1704896540
transform 1 0 89215 0 1 28279
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_212
timestamp 1704896540
transform 1 0 89215 0 1 30295
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_213
timestamp 1704896540
transform 1 0 89215 0 1 33319
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_214
timestamp 1704896540
transform 1 0 89215 0 1 32983
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_215
timestamp 1704896540
transform 1 0 89215 0 1 32647
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_216
timestamp 1704896540
transform 1 0 89215 0 1 32311
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_217
timestamp 1704896540
transform 1 0 89215 0 1 31975
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_218
timestamp 1704896540
transform 1 0 89215 0 1 31639
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_219
timestamp 1704896540
transform 1 0 89215 0 1 31303
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_220
timestamp 1704896540
transform 1 0 89215 0 1 30967
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_221
timestamp 1704896540
transform 1 0 89215 0 1 30631
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_222
timestamp 1704896540
transform 1 0 89215 0 1 27943
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_223
timestamp 1704896540
transform 1 0 89215 0 1 38695
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_224
timestamp 1704896540
transform 1 0 89215 0 1 38359
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_225
timestamp 1704896540
transform 1 0 89215 0 1 38023
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_226
timestamp 1704896540
transform 1 0 89215 0 1 37687
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_227
timestamp 1704896540
transform 1 0 89215 0 1 37351
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_228
timestamp 1704896540
transform 1 0 89215 0 1 37015
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_229
timestamp 1704896540
transform 1 0 89215 0 1 36679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_230
timestamp 1704896540
transform 1 0 89215 0 1 36343
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_231
timestamp 1704896540
transform 1 0 89215 0 1 36007
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_232
timestamp 1704896540
transform 1 0 89215 0 1 35671
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_233
timestamp 1704896540
transform 1 0 89215 0 1 35335
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_234
timestamp 1704896540
transform 1 0 89215 0 1 34999
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_235
timestamp 1704896540
transform 1 0 89215 0 1 34663
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_236
timestamp 1704896540
transform 1 0 89215 0 1 34327
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_237
timestamp 1704896540
transform 1 0 89215 0 1 33991
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_238
timestamp 1704896540
transform 1 0 89215 0 1 33655
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_239
timestamp 1704896540
transform 1 0 89215 0 1 39031
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_240
timestamp 1704896540
transform 1 0 89215 0 1 44407
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_241
timestamp 1704896540
transform 1 0 89215 0 1 44071
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_242
timestamp 1704896540
transform 1 0 89215 0 1 43735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_243
timestamp 1704896540
transform 1 0 89215 0 1 43399
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_244
timestamp 1704896540
transform 1 0 89215 0 1 43063
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_245
timestamp 1704896540
transform 1 0 89215 0 1 42727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_246
timestamp 1704896540
transform 1 0 89215 0 1 42391
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_247
timestamp 1704896540
transform 1 0 89215 0 1 42055
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_248
timestamp 1704896540
transform 1 0 89215 0 1 41719
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_249
timestamp 1704896540
transform 1 0 89215 0 1 41383
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_250
timestamp 1704896540
transform 1 0 89215 0 1 41047
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_251
timestamp 1704896540
transform 1 0 89215 0 1 40711
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_252
timestamp 1704896540
transform 1 0 89215 0 1 40375
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_253
timestamp 1704896540
transform 1 0 89215 0 1 40039
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_254
timestamp 1704896540
transform 1 0 89215 0 1 39703
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_255
timestamp 1704896540
transform 1 0 89215 0 1 39367
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_256
timestamp 1704896540
transform 1 0 37333 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_257
timestamp 1704896540
transform 1 0 40357 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_258
timestamp 1704896540
transform 1 0 36997 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_259
timestamp 1704896540
transform 1 0 44389 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_260
timestamp 1704896540
transform 1 0 40021 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_261
timestamp 1704896540
transform 1 0 40693 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_262
timestamp 1704896540
transform 1 0 39013 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_263
timestamp 1704896540
transform 1 0 36661 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_264
timestamp 1704896540
transform 1 0 38677 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_265
timestamp 1704896540
transform 1 0 44053 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_266
timestamp 1704896540
transform 1 0 43717 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_267
timestamp 1704896540
transform 1 0 44725 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_268
timestamp 1704896540
transform 1 0 45061 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_269
timestamp 1704896540
transform 1 0 36325 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_270
timestamp 1704896540
transform 1 0 38341 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_271
timestamp 1704896540
transform 1 0 41365 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_272
timestamp 1704896540
transform 1 0 38005 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_273
timestamp 1704896540
transform 1 0 35989 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_274
timestamp 1704896540
transform 1 0 41701 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_275
timestamp 1704896540
transform 1 0 35653 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_276
timestamp 1704896540
transform 1 0 41029 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_277
timestamp 1704896540
transform 1 0 45397 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_278
timestamp 1704896540
transform 1 0 35317 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_279
timestamp 1704896540
transform 1 0 39685 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_280
timestamp 1704896540
transform 1 0 43381 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_281
timestamp 1704896540
transform 1 0 43045 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_282
timestamp 1704896540
transform 1 0 34981 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_283
timestamp 1704896540
transform 1 0 39349 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_284
timestamp 1704896540
transform 1 0 42709 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_285
timestamp 1704896540
transform 1 0 42373 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_286
timestamp 1704896540
transform 1 0 34645 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_287
timestamp 1704896540
transform 1 0 37669 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_288
timestamp 1704896540
transform 1 0 34309 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_289
timestamp 1704896540
transform 1 0 42037 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_290
timestamp 1704896540
transform 1 0 33973 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_291
timestamp 1704896540
transform 1 0 28933 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_292
timestamp 1704896540
transform 1 0 32629 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_293
timestamp 1704896540
transform 1 0 29605 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_294
timestamp 1704896540
transform 1 0 32293 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_295
timestamp 1704896540
transform 1 0 31957 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_296
timestamp 1704896540
transform 1 0 32965 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_297
timestamp 1704896540
transform 1 0 31621 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_298
timestamp 1704896540
transform 1 0 33637 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_299
timestamp 1704896540
transform 1 0 28597 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_300
timestamp 1704896540
transform 1 0 31285 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_301
timestamp 1704896540
transform 1 0 30949 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_302
timestamp 1704896540
transform 1 0 33301 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_303
timestamp 1704896540
transform 1 0 30613 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_304
timestamp 1704896540
transform 1 0 29269 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_305
timestamp 1704896540
transform 1 0 30277 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_306
timestamp 1704896540
transform 1 0 29941 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_307
timestamp 1704896540
transform 1 0 24229 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_308
timestamp 1704896540
transform 1 0 25573 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_309
timestamp 1704896540
transform 1 0 25237 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_310
timestamp 1704896540
transform 1 0 23893 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_311
timestamp 1704896540
transform 1 0 23221 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_312
timestamp 1704896540
transform 1 0 23557 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_313
timestamp 1704896540
transform 1 0 24901 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_314
timestamp 1704896540
transform 1 0 28261 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_315
timestamp 1704896540
transform 1 0 27925 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_316
timestamp 1704896540
transform 1 0 27589 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_317
timestamp 1704896540
transform 1 0 27253 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_318
timestamp 1704896540
transform 1 0 26917 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_319
timestamp 1704896540
transform 1 0 26581 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_320
timestamp 1704896540
transform 1 0 26245 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_321
timestamp 1704896540
transform 1 0 25909 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_322
timestamp 1704896540
transform 1 0 24565 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_323
timestamp 1704896540
transform 1 0 21541 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_324
timestamp 1704896540
transform 1 0 21205 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_325
timestamp 1704896540
transform 1 0 20869 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_326
timestamp 1704896540
transform 1 0 18517 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_327
timestamp 1704896540
transform 1 0 18181 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_328
timestamp 1704896540
transform 1 0 17845 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_329
timestamp 1704896540
transform 1 0 19525 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_330
timestamp 1704896540
transform 1 0 18853 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_331
timestamp 1704896540
transform 1 0 19189 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_332
timestamp 1704896540
transform 1 0 21877 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_333
timestamp 1704896540
transform 1 0 17509 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_334
timestamp 1704896540
transform 1 0 20533 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_335
timestamp 1704896540
transform 1 0 22549 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_336
timestamp 1704896540
transform 1 0 20197 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_337
timestamp 1704896540
transform 1 0 19861 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_338
timestamp 1704896540
transform 1 0 22213 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_339
timestamp 1704896540
transform 1 0 12133 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_340
timestamp 1704896540
transform 1 0 11797 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_341
timestamp 1704896540
transform 1 0 14485 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_342
timestamp 1704896540
transform 1 0 13813 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_343
timestamp 1704896540
transform 1 0 13141 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_344
timestamp 1704896540
transform 1 0 14149 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_345
timestamp 1704896540
transform 1 0 15493 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_346
timestamp 1704896540
transform 1 0 12805 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_347
timestamp 1704896540
transform 1 0 12469 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_348
timestamp 1704896540
transform 1 0 17173 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_349
timestamp 1704896540
transform 1 0 16837 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_350
timestamp 1704896540
transform 1 0 16501 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_351
timestamp 1704896540
transform 1 0 13477 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_352
timestamp 1704896540
transform 1 0 15157 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_353
timestamp 1704896540
transform 1 0 16165 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_354
timestamp 1704896540
transform 1 0 15829 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_355
timestamp 1704896540
transform 1 0 14821 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_356
timestamp 1704896540
transform 1 0 11461 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_357
timestamp 1704896540
transform 1 0 8101 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_358
timestamp 1704896540
transform 1 0 7765 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_359
timestamp 1704896540
transform 1 0 11125 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_360
timestamp 1704896540
transform 1 0 7429 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_361
timestamp 1704896540
transform 1 0 10789 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_362
timestamp 1704896540
transform 1 0 10453 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_363
timestamp 1704896540
transform 1 0 10117 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_364
timestamp 1704896540
transform 1 0 9781 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_365
timestamp 1704896540
transform 1 0 7093 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_366
timestamp 1704896540
transform 1 0 9445 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_367
timestamp 1704896540
transform 1 0 9109 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_368
timestamp 1704896540
transform 1 0 6085 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_369
timestamp 1704896540
transform 1 0 6757 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_370
timestamp 1704896540
transform 1 0 6421 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_371
timestamp 1704896540
transform 1 0 8773 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_372
timestamp 1704896540
transform 1 0 8437 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_373
timestamp 1704896540
transform 1 0 1717 0 1 2071
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_374
timestamp 1704896540
transform 1 0 1717 0 1 5431
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_375
timestamp 1704896540
transform 1 0 1717 0 1 5095
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_376
timestamp 1704896540
transform 1 0 1717 0 1 4759
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_377
timestamp 1704896540
transform 1 0 1717 0 1 4423
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_378
timestamp 1704896540
transform 1 0 5749 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_379
timestamp 1704896540
transform 1 0 5413 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_380
timestamp 1704896540
transform 1 0 5077 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_381
timestamp 1704896540
transform 1 0 4741 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_382
timestamp 1704896540
transform 1 0 1717 0 1 4087
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_383
timestamp 1704896540
transform 1 0 4405 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_384
timestamp 1704896540
transform 1 0 4069 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_385
timestamp 1704896540
transform 1 0 3733 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_386
timestamp 1704896540
transform 1 0 1717 0 1 3751
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_387
timestamp 1704896540
transform 1 0 3397 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_388
timestamp 1704896540
transform 1 0 3061 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_389
timestamp 1704896540
transform 1 0 2725 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_390
timestamp 1704896540
transform 1 0 2389 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_391
timestamp 1704896540
transform 1 0 1717 0 1 3415
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_392
timestamp 1704896540
transform 1 0 2053 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_393
timestamp 1704896540
transform 1 0 1717 0 1 3079
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_394
timestamp 1704896540
transform 1 0 1717 0 1 2743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_395
timestamp 1704896540
transform 1 0 1717 0 1 2407
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_396
timestamp 1704896540
transform 1 0 1717 0 1 6103
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_397
timestamp 1704896540
transform 1 0 1717 0 1 11143
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_398
timestamp 1704896540
transform 1 0 1717 0 1 10807
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_399
timestamp 1704896540
transform 1 0 1717 0 1 10471
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_400
timestamp 1704896540
transform 1 0 1717 0 1 10135
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_401
timestamp 1704896540
transform 1 0 1717 0 1 9799
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_402
timestamp 1704896540
transform 1 0 1717 0 1 9463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_403
timestamp 1704896540
transform 1 0 1717 0 1 9127
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_404
timestamp 1704896540
transform 1 0 1717 0 1 8791
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_405
timestamp 1704896540
transform 1 0 1717 0 1 8455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_406
timestamp 1704896540
transform 1 0 1717 0 1 8119
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_407
timestamp 1704896540
transform 1 0 1717 0 1 7783
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_408
timestamp 1704896540
transform 1 0 1717 0 1 7447
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_409
timestamp 1704896540
transform 1 0 1717 0 1 7111
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_410
timestamp 1704896540
transform 1 0 1717 0 1 6775
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_411
timestamp 1704896540
transform 1 0 1717 0 1 6439
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_412
timestamp 1704896540
transform 1 0 1717 0 1 5767
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_413
timestamp 1704896540
transform 1 0 1717 0 1 14839
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_414
timestamp 1704896540
transform 1 0 1717 0 1 14503
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_415
timestamp 1704896540
transform 1 0 1717 0 1 12151
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_416
timestamp 1704896540
transform 1 0 1717 0 1 14167
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_417
timestamp 1704896540
transform 1 0 1717 0 1 13159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_418
timestamp 1704896540
transform 1 0 1717 0 1 12823
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_419
timestamp 1704896540
transform 1 0 1717 0 1 12487
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_420
timestamp 1704896540
transform 1 0 1717 0 1 13831
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_421
timestamp 1704896540
transform 1 0 1717 0 1 16183
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_422
timestamp 1704896540
transform 1 0 1717 0 1 15847
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_423
timestamp 1704896540
transform 1 0 1717 0 1 15175
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_424
timestamp 1704896540
transform 1 0 1717 0 1 11479
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_425
timestamp 1704896540
transform 1 0 1717 0 1 15511
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_426
timestamp 1704896540
transform 1 0 1717 0 1 11815
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_427
timestamp 1704896540
transform 1 0 1717 0 1 13495
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_428
timestamp 1704896540
transform 1 0 1717 0 1 16519
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_429
timestamp 1704896540
transform 1 0 1717 0 1 22231
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_430
timestamp 1704896540
transform 1 0 1717 0 1 21895
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_431
timestamp 1704896540
transform 1 0 1717 0 1 21559
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_432
timestamp 1704896540
transform 1 0 1717 0 1 21223
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_433
timestamp 1704896540
transform 1 0 1717 0 1 20887
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_434
timestamp 1704896540
transform 1 0 1717 0 1 20551
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_435
timestamp 1704896540
transform 1 0 1717 0 1 20215
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_436
timestamp 1704896540
transform 1 0 1717 0 1 19879
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_437
timestamp 1704896540
transform 1 0 1717 0 1 19543
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_438
timestamp 1704896540
transform 1 0 1717 0 1 19207
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_439
timestamp 1704896540
transform 1 0 1717 0 1 18871
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_440
timestamp 1704896540
transform 1 0 1717 0 1 18535
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_441
timestamp 1704896540
transform 1 0 1717 0 1 18199
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_442
timestamp 1704896540
transform 1 0 1717 0 1 17863
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_443
timestamp 1704896540
transform 1 0 1717 0 1 17527
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_444
timestamp 1704896540
transform 1 0 1717 0 1 17191
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_445
timestamp 1704896540
transform 1 0 1717 0 1 16855
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_446
timestamp 1704896540
transform 1 0 1717 0 1 25255
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_447
timestamp 1704896540
transform 1 0 1717 0 1 24919
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_448
timestamp 1704896540
transform 1 0 1717 0 1 24583
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_449
timestamp 1704896540
transform 1 0 1717 0 1 24247
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_450
timestamp 1704896540
transform 1 0 1717 0 1 23911
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_451
timestamp 1704896540
transform 1 0 1717 0 1 23575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_452
timestamp 1704896540
transform 1 0 1717 0 1 23239
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_453
timestamp 1704896540
transform 1 0 1717 0 1 27607
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_454
timestamp 1704896540
transform 1 0 1717 0 1 22903
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_455
timestamp 1704896540
transform 1 0 1717 0 1 27271
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_456
timestamp 1704896540
transform 1 0 1717 0 1 26935
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_457
timestamp 1704896540
transform 1 0 1717 0 1 26599
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_458
timestamp 1704896540
transform 1 0 1717 0 1 26263
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_459
timestamp 1704896540
transform 1 0 1717 0 1 25927
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_460
timestamp 1704896540
transform 1 0 1717 0 1 25591
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_461
timestamp 1704896540
transform 1 0 1717 0 1 22567
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_462
timestamp 1704896540
transform 1 0 1717 0 1 30295
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_463
timestamp 1704896540
transform 1 0 1717 0 1 29959
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_464
timestamp 1704896540
transform 1 0 1717 0 1 29623
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_465
timestamp 1704896540
transform 1 0 1717 0 1 29287
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_466
timestamp 1704896540
transform 1 0 1717 0 1 31639
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_467
timestamp 1704896540
transform 1 0 1717 0 1 28951
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_468
timestamp 1704896540
transform 1 0 1717 0 1 28615
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_469
timestamp 1704896540
transform 1 0 1717 0 1 28279
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_470
timestamp 1704896540
transform 1 0 1717 0 1 31303
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_471
timestamp 1704896540
transform 1 0 1717 0 1 30967
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_472
timestamp 1704896540
transform 1 0 1717 0 1 30631
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_473
timestamp 1704896540
transform 1 0 1717 0 1 33319
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_474
timestamp 1704896540
transform 1 0 1717 0 1 32983
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_475
timestamp 1704896540
transform 1 0 1717 0 1 32647
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_476
timestamp 1704896540
transform 1 0 1717 0 1 32311
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_477
timestamp 1704896540
transform 1 0 1717 0 1 31975
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_478
timestamp 1704896540
transform 1 0 1717 0 1 27943
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_479
timestamp 1704896540
transform 1 0 1717 0 1 34327
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_480
timestamp 1704896540
transform 1 0 1717 0 1 39031
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_481
timestamp 1704896540
transform 1 0 1717 0 1 33991
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_482
timestamp 1704896540
transform 1 0 1717 0 1 38695
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_483
timestamp 1704896540
transform 1 0 1717 0 1 38359
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_484
timestamp 1704896540
transform 1 0 1717 0 1 38023
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_485
timestamp 1704896540
transform 1 0 1717 0 1 37687
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_486
timestamp 1704896540
transform 1 0 1717 0 1 37351
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_487
timestamp 1704896540
transform 1 0 1717 0 1 37015
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_488
timestamp 1704896540
transform 1 0 1717 0 1 36679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_489
timestamp 1704896540
transform 1 0 1717 0 1 36343
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_490
timestamp 1704896540
transform 1 0 1717 0 1 36007
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_491
timestamp 1704896540
transform 1 0 1717 0 1 35671
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_492
timestamp 1704896540
transform 1 0 1717 0 1 35335
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_493
timestamp 1704896540
transform 1 0 1717 0 1 33655
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_494
timestamp 1704896540
transform 1 0 1717 0 1 34999
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_495
timestamp 1704896540
transform 1 0 1717 0 1 34663
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_496
timestamp 1704896540
transform 1 0 1717 0 1 39703
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_497
timestamp 1704896540
transform 1 0 1717 0 1 39367
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_498
timestamp 1704896540
transform 1 0 1717 0 1 40039
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_499
timestamp 1704896540
transform 1 0 1717 0 1 44407
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_500
timestamp 1704896540
transform 1 0 1717 0 1 44071
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_501
timestamp 1704896540
transform 1 0 1717 0 1 43735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_502
timestamp 1704896540
transform 1 0 1717 0 1 43399
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_503
timestamp 1704896540
transform 1 0 1717 0 1 43063
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_504
timestamp 1704896540
transform 1 0 1717 0 1 42727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_505
timestamp 1704896540
transform 1 0 1717 0 1 42391
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_506
timestamp 1704896540
transform 1 0 1717 0 1 42055
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_507
timestamp 1704896540
transform 1 0 1717 0 1 41719
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_508
timestamp 1704896540
transform 1 0 1717 0 1 41383
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_509
timestamp 1704896540
transform 1 0 1717 0 1 41047
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_510
timestamp 1704896540
transform 1 0 1717 0 1 40711
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_511
timestamp 1704896540
transform 1 0 1717 0 1 40375
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_512
timestamp 1704896540
transform 1 0 22885 0 1 1735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_513
timestamp 1704896540
transform 1 0 1717 0 1 47431
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_514
timestamp 1704896540
transform 1 0 1717 0 1 47095
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_515
timestamp 1704896540
transform 1 0 1717 0 1 46759
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_516
timestamp 1704896540
transform 1 0 1717 0 1 46423
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_517
timestamp 1704896540
transform 1 0 1717 0 1 46087
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_518
timestamp 1704896540
transform 1 0 1717 0 1 45751
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_519
timestamp 1704896540
transform 1 0 1717 0 1 45415
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_520
timestamp 1704896540
transform 1 0 1717 0 1 45079
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_521
timestamp 1704896540
transform 1 0 1717 0 1 44743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_522
timestamp 1704896540
transform 1 0 1717 0 1 50119
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_523
timestamp 1704896540
transform 1 0 1717 0 1 49783
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_524
timestamp 1704896540
transform 1 0 1717 0 1 49447
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_525
timestamp 1704896540
transform 1 0 1717 0 1 49111
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_526
timestamp 1704896540
transform 1 0 1717 0 1 48775
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_527
timestamp 1704896540
transform 1 0 1717 0 1 48439
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_528
timestamp 1704896540
transform 1 0 1717 0 1 48103
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_529
timestamp 1704896540
transform 1 0 1717 0 1 47767
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_530
timestamp 1704896540
transform 1 0 1717 0 1 53479
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_531
timestamp 1704896540
transform 1 0 1717 0 1 53143
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_532
timestamp 1704896540
transform 1 0 1717 0 1 52807
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_533
timestamp 1704896540
transform 1 0 1717 0 1 52471
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_534
timestamp 1704896540
transform 1 0 1717 0 1 52135
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_535
timestamp 1704896540
transform 1 0 1717 0 1 51799
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_536
timestamp 1704896540
transform 1 0 1717 0 1 51463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_537
timestamp 1704896540
transform 1 0 1717 0 1 51127
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_538
timestamp 1704896540
transform 1 0 1717 0 1 50791
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_539
timestamp 1704896540
transform 1 0 1717 0 1 50455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_540
timestamp 1704896540
transform 1 0 1717 0 1 54823
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_541
timestamp 1704896540
transform 1 0 1717 0 1 54151
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_542
timestamp 1704896540
transform 1 0 1717 0 1 55159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_543
timestamp 1704896540
transform 1 0 1717 0 1 54487
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_544
timestamp 1704896540
transform 1 0 1717 0 1 55495
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_545
timestamp 1704896540
transform 1 0 1717 0 1 53815
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_546
timestamp 1704896540
transform 1 0 1717 0 1 57847
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_547
timestamp 1704896540
transform 1 0 1717 0 1 56167
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_548
timestamp 1704896540
transform 1 0 1717 0 1 57511
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_549
timestamp 1704896540
transform 1 0 1717 0 1 57175
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_550
timestamp 1704896540
transform 1 0 1717 0 1 56839
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_551
timestamp 1704896540
transform 1 0 1717 0 1 61207
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_552
timestamp 1704896540
transform 1 0 1717 0 1 58855
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_553
timestamp 1704896540
transform 1 0 1717 0 1 58519
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_554
timestamp 1704896540
transform 1 0 1717 0 1 58183
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_555
timestamp 1704896540
transform 1 0 1717 0 1 60871
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_556
timestamp 1704896540
transform 1 0 1717 0 1 60535
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_557
timestamp 1704896540
transform 1 0 1717 0 1 60199
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_558
timestamp 1704896540
transform 1 0 1717 0 1 55831
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_559
timestamp 1704896540
transform 1 0 1717 0 1 59863
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_560
timestamp 1704896540
transform 1 0 1717 0 1 56503
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_561
timestamp 1704896540
transform 1 0 1717 0 1 59527
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_562
timestamp 1704896540
transform 1 0 1717 0 1 59191
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_563
timestamp 1704896540
transform 1 0 1717 0 1 65239
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_564
timestamp 1704896540
transform 1 0 1717 0 1 64903
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_565
timestamp 1704896540
transform 1 0 1717 0 1 64567
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_566
timestamp 1704896540
transform 1 0 1717 0 1 64231
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_567
timestamp 1704896540
transform 1 0 1717 0 1 63895
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_568
timestamp 1704896540
transform 1 0 1717 0 1 63559
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_569
timestamp 1704896540
transform 1 0 1717 0 1 63223
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_570
timestamp 1704896540
transform 1 0 1717 0 1 62887
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_571
timestamp 1704896540
transform 1 0 1717 0 1 62551
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_572
timestamp 1704896540
transform 1 0 1717 0 1 62215
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_573
timestamp 1704896540
transform 1 0 1717 0 1 61879
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_574
timestamp 1704896540
transform 1 0 1717 0 1 61543
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_575
timestamp 1704896540
transform 1 0 1717 0 1 66583
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_576
timestamp 1704896540
transform 1 0 1717 0 1 66247
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_577
timestamp 1704896540
transform 1 0 1717 0 1 65911
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_578
timestamp 1704896540
transform 1 0 1717 0 1 65575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_579
timestamp 1704896540
transform 1 0 1717 0 1 71623
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_580
timestamp 1704896540
transform 1 0 1717 0 1 71287
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_581
timestamp 1704896540
transform 1 0 1717 0 1 70951
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_582
timestamp 1704896540
transform 1 0 1717 0 1 70615
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_583
timestamp 1704896540
transform 1 0 1717 0 1 70279
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_584
timestamp 1704896540
transform 1 0 1717 0 1 69943
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_585
timestamp 1704896540
transform 1 0 1717 0 1 69607
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_586
timestamp 1704896540
transform 1 0 1717 0 1 69271
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_587
timestamp 1704896540
transform 1 0 1717 0 1 68935
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_588
timestamp 1704896540
transform 1 0 1717 0 1 68599
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_589
timestamp 1704896540
transform 1 0 1717 0 1 68263
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_590
timestamp 1704896540
transform 1 0 1717 0 1 67927
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_591
timestamp 1704896540
transform 1 0 1717 0 1 67591
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_592
timestamp 1704896540
transform 1 0 1717 0 1 67255
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_593
timestamp 1704896540
transform 1 0 1717 0 1 66919
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_594
timestamp 1704896540
transform 1 0 1717 0 1 72295
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_595
timestamp 1704896540
transform 1 0 1717 0 1 71959
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_596
timestamp 1704896540
transform 1 0 1717 0 1 77335
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_597
timestamp 1704896540
transform 1 0 1717 0 1 76999
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_598
timestamp 1704896540
transform 1 0 1717 0 1 76663
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_599
timestamp 1704896540
transform 1 0 1717 0 1 76327
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_600
timestamp 1704896540
transform 1 0 1717 0 1 75991
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_601
timestamp 1704896540
transform 1 0 1717 0 1 75655
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_602
timestamp 1704896540
transform 1 0 1717 0 1 75319
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_603
timestamp 1704896540
transform 1 0 1717 0 1 74983
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_604
timestamp 1704896540
transform 1 0 1717 0 1 74647
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_605
timestamp 1704896540
transform 1 0 1717 0 1 74311
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_606
timestamp 1704896540
transform 1 0 1717 0 1 73975
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_607
timestamp 1704896540
transform 1 0 1717 0 1 73639
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_608
timestamp 1704896540
transform 1 0 1717 0 1 73303
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_609
timestamp 1704896540
transform 1 0 1717 0 1 72967
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_610
timestamp 1704896540
transform 1 0 1717 0 1 72631
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_611
timestamp 1704896540
transform 1 0 1717 0 1 77671
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_612
timestamp 1704896540
transform 1 0 1717 0 1 82375
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_613
timestamp 1704896540
transform 1 0 1717 0 1 82039
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_614
timestamp 1704896540
transform 1 0 1717 0 1 81703
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_615
timestamp 1704896540
transform 1 0 1717 0 1 79015
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_616
timestamp 1704896540
transform 1 0 1717 0 1 78679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_617
timestamp 1704896540
transform 1 0 1717 0 1 78343
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_618
timestamp 1704896540
transform 1 0 1717 0 1 78007
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_619
timestamp 1704896540
transform 1 0 1717 0 1 81367
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_620
timestamp 1704896540
transform 1 0 1717 0 1 81031
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_621
timestamp 1704896540
transform 1 0 1717 0 1 80695
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_622
timestamp 1704896540
transform 1 0 1717 0 1 80359
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_623
timestamp 1704896540
transform 1 0 1717 0 1 80023
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_624
timestamp 1704896540
transform 1 0 1717 0 1 79687
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_625
timestamp 1704896540
transform 1 0 1717 0 1 79351
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_626
timestamp 1704896540
transform 1 0 1717 0 1 83383
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_627
timestamp 1704896540
transform 1 0 1717 0 1 83047
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_628
timestamp 1704896540
transform 1 0 1717 0 1 82711
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_629
timestamp 1704896540
transform 1 0 1717 0 1 87079
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_630
timestamp 1704896540
transform 1 0 1717 0 1 86743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_631
timestamp 1704896540
transform 1 0 1717 0 1 86407
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_632
timestamp 1704896540
transform 1 0 1717 0 1 86071
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_633
timestamp 1704896540
transform 1 0 1717 0 1 85735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_634
timestamp 1704896540
transform 1 0 1717 0 1 85399
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_635
timestamp 1704896540
transform 1 0 1717 0 1 85063
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_636
timestamp 1704896540
transform 1 0 1717 0 1 84727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_637
timestamp 1704896540
transform 1 0 1717 0 1 84391
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_638
timestamp 1704896540
transform 1 0 1717 0 1 84055
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_639
timestamp 1704896540
transform 1 0 1717 0 1 83719
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_640
timestamp 1704896540
transform 1 0 5749 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_641
timestamp 1704896540
transform 1 0 5413 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_642
timestamp 1704896540
transform 1 0 5077 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_643
timestamp 1704896540
transform 1 0 4741 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_644
timestamp 1704896540
transform 1 0 4405 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_645
timestamp 1704896540
transform 1 0 4069 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_646
timestamp 1704896540
transform 1 0 3733 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_647
timestamp 1704896540
transform 1 0 3397 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_648
timestamp 1704896540
transform 1 0 3061 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_649
timestamp 1704896540
transform 1 0 2725 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_650
timestamp 1704896540
transform 1 0 2389 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_651
timestamp 1704896540
transform 1 0 2053 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_652
timestamp 1704896540
transform 1 0 11461 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_653
timestamp 1704896540
transform 1 0 11125 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_654
timestamp 1704896540
transform 1 0 10789 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_655
timestamp 1704896540
transform 1 0 10453 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_656
timestamp 1704896540
transform 1 0 10117 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_657
timestamp 1704896540
transform 1 0 9781 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_658
timestamp 1704896540
transform 1 0 9445 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_659
timestamp 1704896540
transform 1 0 9109 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_660
timestamp 1704896540
transform 1 0 8773 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_661
timestamp 1704896540
transform 1 0 8437 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_662
timestamp 1704896540
transform 1 0 8101 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_663
timestamp 1704896540
transform 1 0 7765 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_664
timestamp 1704896540
transform 1 0 7429 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_665
timestamp 1704896540
transform 1 0 7093 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_666
timestamp 1704896540
transform 1 0 6757 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_667
timestamp 1704896540
transform 1 0 6421 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_668
timestamp 1704896540
transform 1 0 6085 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_669
timestamp 1704896540
transform 1 0 22549 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_670
timestamp 1704896540
transform 1 0 22213 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_671
timestamp 1704896540
transform 1 0 21877 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_672
timestamp 1704896540
transform 1 0 21541 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_673
timestamp 1704896540
transform 1 0 21205 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_674
timestamp 1704896540
transform 1 0 20869 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_675
timestamp 1704896540
transform 1 0 20533 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_676
timestamp 1704896540
transform 1 0 20197 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_677
timestamp 1704896540
transform 1 0 19861 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_678
timestamp 1704896540
transform 1 0 19525 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_679
timestamp 1704896540
transform 1 0 19189 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_680
timestamp 1704896540
transform 1 0 18853 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_681
timestamp 1704896540
transform 1 0 18517 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_682
timestamp 1704896540
transform 1 0 18181 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_683
timestamp 1704896540
transform 1 0 17845 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_684
timestamp 1704896540
transform 1 0 17509 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_685
timestamp 1704896540
transform 1 0 17173 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_686
timestamp 1704896540
transform 1 0 16837 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_687
timestamp 1704896540
transform 1 0 16501 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_688
timestamp 1704896540
transform 1 0 16165 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_689
timestamp 1704896540
transform 1 0 15829 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_690
timestamp 1704896540
transform 1 0 15493 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_691
timestamp 1704896540
transform 1 0 15157 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_692
timestamp 1704896540
transform 1 0 14821 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_693
timestamp 1704896540
transform 1 0 14485 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_694
timestamp 1704896540
transform 1 0 14149 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_695
timestamp 1704896540
transform 1 0 13813 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_696
timestamp 1704896540
transform 1 0 13477 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_697
timestamp 1704896540
transform 1 0 13141 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_698
timestamp 1704896540
transform 1 0 12805 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_699
timestamp 1704896540
transform 1 0 12469 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_700
timestamp 1704896540
transform 1 0 12133 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_701
timestamp 1704896540
transform 1 0 11797 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_702
timestamp 1704896540
transform 1 0 30613 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_703
timestamp 1704896540
transform 1 0 30277 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_704
timestamp 1704896540
transform 1 0 29941 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_705
timestamp 1704896540
transform 1 0 29605 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_706
timestamp 1704896540
transform 1 0 29269 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_707
timestamp 1704896540
transform 1 0 28933 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_708
timestamp 1704896540
transform 1 0 28597 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_709
timestamp 1704896540
transform 1 0 28261 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_710
timestamp 1704896540
transform 1 0 27925 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_711
timestamp 1704896540
transform 1 0 27589 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_712
timestamp 1704896540
transform 1 0 27253 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_713
timestamp 1704896540
transform 1 0 26917 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_714
timestamp 1704896540
transform 1 0 26581 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_715
timestamp 1704896540
transform 1 0 26245 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_716
timestamp 1704896540
transform 1 0 25909 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_717
timestamp 1704896540
transform 1 0 25573 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_718
timestamp 1704896540
transform 1 0 25237 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_719
timestamp 1704896540
transform 1 0 24901 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_720
timestamp 1704896540
transform 1 0 24565 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_721
timestamp 1704896540
transform 1 0 24229 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_722
timestamp 1704896540
transform 1 0 23893 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_723
timestamp 1704896540
transform 1 0 23557 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_724
timestamp 1704896540
transform 1 0 23221 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_725
timestamp 1704896540
transform 1 0 33973 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_726
timestamp 1704896540
transform 1 0 33637 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_727
timestamp 1704896540
transform 1 0 33301 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_728
timestamp 1704896540
transform 1 0 32965 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_729
timestamp 1704896540
transform 1 0 32629 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_730
timestamp 1704896540
transform 1 0 32293 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_731
timestamp 1704896540
transform 1 0 31957 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_732
timestamp 1704896540
transform 1 0 31621 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_733
timestamp 1704896540
transform 1 0 31285 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_734
timestamp 1704896540
transform 1 0 30949 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_735
timestamp 1704896540
transform 1 0 44053 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_736
timestamp 1704896540
transform 1 0 43717 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_737
timestamp 1704896540
transform 1 0 43381 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_738
timestamp 1704896540
transform 1 0 43045 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_739
timestamp 1704896540
transform 1 0 42709 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_740
timestamp 1704896540
transform 1 0 42373 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_741
timestamp 1704896540
transform 1 0 42037 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_742
timestamp 1704896540
transform 1 0 41701 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_743
timestamp 1704896540
transform 1 0 41365 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_744
timestamp 1704896540
transform 1 0 41029 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_745
timestamp 1704896540
transform 1 0 40693 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_746
timestamp 1704896540
transform 1 0 40357 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_747
timestamp 1704896540
transform 1 0 40021 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_748
timestamp 1704896540
transform 1 0 39685 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_749
timestamp 1704896540
transform 1 0 39349 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_750
timestamp 1704896540
transform 1 0 39013 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_751
timestamp 1704896540
transform 1 0 38677 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_752
timestamp 1704896540
transform 1 0 38341 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_753
timestamp 1704896540
transform 1 0 38005 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_754
timestamp 1704896540
transform 1 0 37669 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_755
timestamp 1704896540
transform 1 0 37333 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_756
timestamp 1704896540
transform 1 0 36997 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_757
timestamp 1704896540
transform 1 0 36661 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_758
timestamp 1704896540
transform 1 0 36325 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_759
timestamp 1704896540
transform 1 0 35989 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_760
timestamp 1704896540
transform 1 0 35653 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_761
timestamp 1704896540
transform 1 0 35317 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_762
timestamp 1704896540
transform 1 0 34981 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_763
timestamp 1704896540
transform 1 0 34645 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_764
timestamp 1704896540
transform 1 0 34309 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_765
timestamp 1704896540
transform 1 0 45397 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_766
timestamp 1704896540
transform 1 0 45061 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_767
timestamp 1704896540
transform 1 0 44725 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_768
timestamp 1704896540
transform 1 0 44389 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_769
timestamp 1704896540
transform 1 0 22885 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_770
timestamp 1704896540
transform 1 0 89215 0 1 47095
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_771
timestamp 1704896540
transform 1 0 89215 0 1 46759
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_772
timestamp 1704896540
transform 1 0 89215 0 1 46423
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_773
timestamp 1704896540
transform 1 0 89215 0 1 48439
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_774
timestamp 1704896540
transform 1 0 89215 0 1 50119
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_775
timestamp 1704896540
transform 1 0 89215 0 1 48103
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_776
timestamp 1704896540
transform 1 0 89215 0 1 49783
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_777
timestamp 1704896540
transform 1 0 89215 0 1 49447
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_778
timestamp 1704896540
transform 1 0 89215 0 1 46087
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_779
timestamp 1704896540
transform 1 0 89215 0 1 49111
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_780
timestamp 1704896540
transform 1 0 89215 0 1 45751
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_781
timestamp 1704896540
transform 1 0 89215 0 1 45415
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_782
timestamp 1704896540
transform 1 0 89215 0 1 48775
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_783
timestamp 1704896540
transform 1 0 89215 0 1 47767
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_784
timestamp 1704896540
transform 1 0 89215 0 1 47431
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_785
timestamp 1704896540
transform 1 0 89215 0 1 45079
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_786
timestamp 1704896540
transform 1 0 89215 0 1 44743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_787
timestamp 1704896540
transform 1 0 89215 0 1 55495
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_788
timestamp 1704896540
transform 1 0 89215 0 1 55159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_789
timestamp 1704896540
transform 1 0 89215 0 1 54823
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_790
timestamp 1704896540
transform 1 0 89215 0 1 54487
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_791
timestamp 1704896540
transform 1 0 89215 0 1 54151
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_792
timestamp 1704896540
transform 1 0 89215 0 1 52135
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_793
timestamp 1704896540
transform 1 0 89215 0 1 53815
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_794
timestamp 1704896540
transform 1 0 89215 0 1 53479
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_795
timestamp 1704896540
transform 1 0 89215 0 1 51799
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_796
timestamp 1704896540
transform 1 0 89215 0 1 50455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_797
timestamp 1704896540
transform 1 0 89215 0 1 51463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_798
timestamp 1704896540
transform 1 0 89215 0 1 51127
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_799
timestamp 1704896540
transform 1 0 89215 0 1 53143
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_800
timestamp 1704896540
transform 1 0 89215 0 1 52807
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_801
timestamp 1704896540
transform 1 0 89215 0 1 52471
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_802
timestamp 1704896540
transform 1 0 89215 0 1 50791
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_803
timestamp 1704896540
transform 1 0 89215 0 1 57511
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_804
timestamp 1704896540
transform 1 0 89215 0 1 55831
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_805
timestamp 1704896540
transform 1 0 89215 0 1 57175
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_806
timestamp 1704896540
transform 1 0 89215 0 1 56839
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_807
timestamp 1704896540
transform 1 0 89215 0 1 56503
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_808
timestamp 1704896540
transform 1 0 89215 0 1 61207
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_809
timestamp 1704896540
transform 1 0 89215 0 1 56167
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_810
timestamp 1704896540
transform 1 0 89215 0 1 60871
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_811
timestamp 1704896540
transform 1 0 89215 0 1 60535
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_812
timestamp 1704896540
transform 1 0 89215 0 1 60199
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_813
timestamp 1704896540
transform 1 0 89215 0 1 59863
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_814
timestamp 1704896540
transform 1 0 89215 0 1 59527
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_815
timestamp 1704896540
transform 1 0 89215 0 1 59191
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_816
timestamp 1704896540
transform 1 0 89215 0 1 58855
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_817
timestamp 1704896540
transform 1 0 89215 0 1 58519
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_818
timestamp 1704896540
transform 1 0 89215 0 1 58183
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_819
timestamp 1704896540
transform 1 0 89215 0 1 57847
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_820
timestamp 1704896540
transform 1 0 89215 0 1 66583
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_821
timestamp 1704896540
transform 1 0 89215 0 1 66247
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_822
timestamp 1704896540
transform 1 0 89215 0 1 65911
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_823
timestamp 1704896540
transform 1 0 89215 0 1 65575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_824
timestamp 1704896540
transform 1 0 89215 0 1 65239
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_825
timestamp 1704896540
transform 1 0 89215 0 1 64903
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_826
timestamp 1704896540
transform 1 0 89215 0 1 64567
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_827
timestamp 1704896540
transform 1 0 89215 0 1 64231
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_828
timestamp 1704896540
transform 1 0 89215 0 1 63895
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_829
timestamp 1704896540
transform 1 0 89215 0 1 63559
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_830
timestamp 1704896540
transform 1 0 89215 0 1 63223
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_831
timestamp 1704896540
transform 1 0 89215 0 1 62887
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_832
timestamp 1704896540
transform 1 0 89215 0 1 62551
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_833
timestamp 1704896540
transform 1 0 89215 0 1 62215
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_834
timestamp 1704896540
transform 1 0 89215 0 1 61879
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_835
timestamp 1704896540
transform 1 0 89215 0 1 61543
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_836
timestamp 1704896540
transform 1 0 45733 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_837
timestamp 1704896540
transform 1 0 55477 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_838
timestamp 1704896540
transform 1 0 55141 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_839
timestamp 1704896540
transform 1 0 54805 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_840
timestamp 1704896540
transform 1 0 54469 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_841
timestamp 1704896540
transform 1 0 54133 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_842
timestamp 1704896540
transform 1 0 53797 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_843
timestamp 1704896540
transform 1 0 53461 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_844
timestamp 1704896540
transform 1 0 53125 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_845
timestamp 1704896540
transform 1 0 52789 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_846
timestamp 1704896540
transform 1 0 52453 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_847
timestamp 1704896540
transform 1 0 52117 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_848
timestamp 1704896540
transform 1 0 51781 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_849
timestamp 1704896540
transform 1 0 51445 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_850
timestamp 1704896540
transform 1 0 51109 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_851
timestamp 1704896540
transform 1 0 50773 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_852
timestamp 1704896540
transform 1 0 50437 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_853
timestamp 1704896540
transform 1 0 50101 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_854
timestamp 1704896540
transform 1 0 49765 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_855
timestamp 1704896540
transform 1 0 49429 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_856
timestamp 1704896540
transform 1 0 49093 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_857
timestamp 1704896540
transform 1 0 48757 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_858
timestamp 1704896540
transform 1 0 48421 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_859
timestamp 1704896540
transform 1 0 47413 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_860
timestamp 1704896540
transform 1 0 47077 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_861
timestamp 1704896540
transform 1 0 46741 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_862
timestamp 1704896540
transform 1 0 46405 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_863
timestamp 1704896540
transform 1 0 46069 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_864
timestamp 1704896540
transform 1 0 48085 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_865
timestamp 1704896540
transform 1 0 47749 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_866
timestamp 1704896540
transform 1 0 56485 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_867
timestamp 1704896540
transform 1 0 56149 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_868
timestamp 1704896540
transform 1 0 55813 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_869
timestamp 1704896540
transform 1 0 67909 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_870
timestamp 1704896540
transform 1 0 67573 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_871
timestamp 1704896540
transform 1 0 67237 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_872
timestamp 1704896540
transform 1 0 66901 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_873
timestamp 1704896540
transform 1 0 66565 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_874
timestamp 1704896540
transform 1 0 66229 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_875
timestamp 1704896540
transform 1 0 65893 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_876
timestamp 1704896540
transform 1 0 65557 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_877
timestamp 1704896540
transform 1 0 65221 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_878
timestamp 1704896540
transform 1 0 64885 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_879
timestamp 1704896540
transform 1 0 64549 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_880
timestamp 1704896540
transform 1 0 64213 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_881
timestamp 1704896540
transform 1 0 63877 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_882
timestamp 1704896540
transform 1 0 63541 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_883
timestamp 1704896540
transform 1 0 63205 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_884
timestamp 1704896540
transform 1 0 62869 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_885
timestamp 1704896540
transform 1 0 62533 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_886
timestamp 1704896540
transform 1 0 62197 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_887
timestamp 1704896540
transform 1 0 61861 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_888
timestamp 1704896540
transform 1 0 61525 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_889
timestamp 1704896540
transform 1 0 61189 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_890
timestamp 1704896540
transform 1 0 60853 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_891
timestamp 1704896540
transform 1 0 60517 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_892
timestamp 1704896540
transform 1 0 60181 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_893
timestamp 1704896540
transform 1 0 59845 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_894
timestamp 1704896540
transform 1 0 59509 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_895
timestamp 1704896540
transform 1 0 59173 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_896
timestamp 1704896540
transform 1 0 58837 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_897
timestamp 1704896540
transform 1 0 58501 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_898
timestamp 1704896540
transform 1 0 58165 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_899
timestamp 1704896540
transform 1 0 57829 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_900
timestamp 1704896540
transform 1 0 57493 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_901
timestamp 1704896540
transform 1 0 57157 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_902
timestamp 1704896540
transform 1 0 56821 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_903
timestamp 1704896540
transform 1 0 89215 0 1 70951
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_904
timestamp 1704896540
transform 1 0 89215 0 1 70615
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_905
timestamp 1704896540
transform 1 0 89215 0 1 70279
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_906
timestamp 1704896540
transform 1 0 89215 0 1 69943
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_907
timestamp 1704896540
transform 1 0 89215 0 1 69607
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_908
timestamp 1704896540
transform 1 0 89215 0 1 69271
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_909
timestamp 1704896540
transform 1 0 89215 0 1 68935
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_910
timestamp 1704896540
transform 1 0 89215 0 1 68599
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_911
timestamp 1704896540
transform 1 0 89215 0 1 68263
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_912
timestamp 1704896540
transform 1 0 89215 0 1 67927
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_913
timestamp 1704896540
transform 1 0 89215 0 1 67591
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_914
timestamp 1704896540
transform 1 0 89215 0 1 67255
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_915
timestamp 1704896540
transform 1 0 89215 0 1 66919
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_916
timestamp 1704896540
transform 1 0 89215 0 1 71959
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_917
timestamp 1704896540
transform 1 0 89215 0 1 71623
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_918
timestamp 1704896540
transform 1 0 89215 0 1 71287
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_919
timestamp 1704896540
transform 1 0 89215 0 1 72295
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_920
timestamp 1704896540
transform 1 0 89215 0 1 77671
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_921
timestamp 1704896540
transform 1 0 89215 0 1 77335
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_922
timestamp 1704896540
transform 1 0 89215 0 1 76999
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_923
timestamp 1704896540
transform 1 0 89215 0 1 76663
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_924
timestamp 1704896540
transform 1 0 89215 0 1 76327
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_925
timestamp 1704896540
transform 1 0 89215 0 1 75991
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_926
timestamp 1704896540
transform 1 0 89215 0 1 75655
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_927
timestamp 1704896540
transform 1 0 89215 0 1 75319
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_928
timestamp 1704896540
transform 1 0 89215 0 1 74983
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_929
timestamp 1704896540
transform 1 0 89215 0 1 74647
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_930
timestamp 1704896540
transform 1 0 89215 0 1 74311
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_931
timestamp 1704896540
transform 1 0 89215 0 1 73975
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_932
timestamp 1704896540
transform 1 0 89215 0 1 73639
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_933
timestamp 1704896540
transform 1 0 89215 0 1 73303
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_934
timestamp 1704896540
transform 1 0 89215 0 1 72967
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_935
timestamp 1704896540
transform 1 0 89215 0 1 72631
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_936
timestamp 1704896540
transform 1 0 71605 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_937
timestamp 1704896540
transform 1 0 71269 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_938
timestamp 1704896540
transform 1 0 68245 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_939
timestamp 1704896540
transform 1 0 72613 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_940
timestamp 1704896540
transform 1 0 72277 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_941
timestamp 1704896540
transform 1 0 70933 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_942
timestamp 1704896540
transform 1 0 70597 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_943
timestamp 1704896540
transform 1 0 70261 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_944
timestamp 1704896540
transform 1 0 69925 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_945
timestamp 1704896540
transform 1 0 69589 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_946
timestamp 1704896540
transform 1 0 69253 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_947
timestamp 1704896540
transform 1 0 68917 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_948
timestamp 1704896540
transform 1 0 68581 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_949
timestamp 1704896540
transform 1 0 71941 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_950
timestamp 1704896540
transform 1 0 73621 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_951
timestamp 1704896540
transform 1 0 73285 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_952
timestamp 1704896540
transform 1 0 72949 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_953
timestamp 1704896540
transform 1 0 73957 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_954
timestamp 1704896540
transform 1 0 79333 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_955
timestamp 1704896540
transform 1 0 78997 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_956
timestamp 1704896540
transform 1 0 78661 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_957
timestamp 1704896540
transform 1 0 78325 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_958
timestamp 1704896540
transform 1 0 77989 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_959
timestamp 1704896540
transform 1 0 77653 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_960
timestamp 1704896540
transform 1 0 77317 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_961
timestamp 1704896540
transform 1 0 76981 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_962
timestamp 1704896540
transform 1 0 76645 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_963
timestamp 1704896540
transform 1 0 76309 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_964
timestamp 1704896540
transform 1 0 75973 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_965
timestamp 1704896540
transform 1 0 75637 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_966
timestamp 1704896540
transform 1 0 75301 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_967
timestamp 1704896540
transform 1 0 74965 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_968
timestamp 1704896540
transform 1 0 74629 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_969
timestamp 1704896540
transform 1 0 74293 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_970
timestamp 1704896540
transform 1 0 89215 0 1 79687
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_971
timestamp 1704896540
transform 1 0 89215 0 1 79351
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_972
timestamp 1704896540
transform 1 0 89215 0 1 79015
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_973
timestamp 1704896540
transform 1 0 89215 0 1 78679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_974
timestamp 1704896540
transform 1 0 89215 0 1 78343
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_975
timestamp 1704896540
transform 1 0 89215 0 1 78007
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_976
timestamp 1704896540
transform 1 0 89215 0 1 83383
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_977
timestamp 1704896540
transform 1 0 89215 0 1 83047
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_978
timestamp 1704896540
transform 1 0 89215 0 1 82711
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_979
timestamp 1704896540
transform 1 0 89215 0 1 82375
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_980
timestamp 1704896540
transform 1 0 89215 0 1 82039
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_981
timestamp 1704896540
transform 1 0 89215 0 1 81703
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_982
timestamp 1704896540
transform 1 0 89215 0 1 81367
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_983
timestamp 1704896540
transform 1 0 89215 0 1 81031
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_984
timestamp 1704896540
transform 1 0 89215 0 1 80695
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_985
timestamp 1704896540
transform 1 0 89215 0 1 80359
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_986
timestamp 1704896540
transform 1 0 89215 0 1 80023
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_987
timestamp 1704896540
transform 1 0 79669 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_988
timestamp 1704896540
transform 1 0 81685 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_989
timestamp 1704896540
transform 1 0 81349 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_990
timestamp 1704896540
transform 1 0 81013 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_991
timestamp 1704896540
transform 1 0 80677 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_992
timestamp 1704896540
transform 1 0 80341 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_993
timestamp 1704896540
transform 1 0 80005 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_994
timestamp 1704896540
transform 1 0 85045 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_995
timestamp 1704896540
transform 1 0 84709 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_996
timestamp 1704896540
transform 1 0 84373 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_997
timestamp 1704896540
transform 1 0 84037 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_998
timestamp 1704896540
transform 1 0 83701 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_999
timestamp 1704896540
transform 1 0 83365 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_1000
timestamp 1704896540
transform 1 0 83029 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_1001
timestamp 1704896540
transform 1 0 82693 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_1002
timestamp 1704896540
transform 1 0 82357 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_1003
timestamp 1704896540
transform 1 0 82021 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_1004
timestamp 1704896540
transform 1 0 85381 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_1005
timestamp 1704896540
transform 1 0 89215 0 1 87079
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_1006
timestamp 1704896540
transform 1 0 89215 0 1 86743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_1007
timestamp 1704896540
transform 1 0 89215 0 1 86407
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_1008
timestamp 1704896540
transform 1 0 89215 0 1 86071
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_1009
timestamp 1704896540
transform 1 0 89215 0 1 85735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_1010
timestamp 1704896540
transform 1 0 89215 0 1 85399
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_1011
timestamp 1704896540
transform 1 0 89215 0 1 85063
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_1012
timestamp 1704896540
transform 1 0 89215 0 1 84727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_1013
timestamp 1704896540
transform 1 0 89215 0 1 84391
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_1014
timestamp 1704896540
transform 1 0 89215 0 1 84055
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_1015
timestamp 1704896540
transform 1 0 89215 0 1 83719
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_1016
timestamp 1704896540
transform 1 0 88741 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_1017
timestamp 1704896540
transform 1 0 88405 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_1018
timestamp 1704896540
transform 1 0 88069 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_1019
timestamp 1704896540
transform 1 0 87733 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_1020
timestamp 1704896540
transform 1 0 87397 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_1021
timestamp 1704896540
transform 1 0 87061 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_1022
timestamp 1704896540
transform 1 0 86725 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_1023
timestamp 1704896540
transform 1 0 86389 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_1024
timestamp 1704896540
transform 1 0 86053 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_1025
timestamp 1704896540
transform 1 0 85717 0 1 87463
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_0
timestamp 1704896540
transform 1 0 89212 0 1 5096
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_1
timestamp 1704896540
transform 1 0 89212 0 1 4760
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_2
timestamp 1704896540
transform 1 0 89212 0 1 4424
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_3
timestamp 1704896540
transform 1 0 89212 0 1 4088
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_4
timestamp 1704896540
transform 1 0 89212 0 1 3752
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_5
timestamp 1704896540
transform 1 0 89212 0 1 3416
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_6
timestamp 1704896540
transform 1 0 89212 0 1 3080
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_7
timestamp 1704896540
transform 1 0 89212 0 1 2744
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_8
timestamp 1704896540
transform 1 0 89212 0 1 2408
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_9
timestamp 1704896540
transform 1 0 89212 0 1 2072
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_10
timestamp 1704896540
transform 1 0 87730 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_11
timestamp 1704896540
transform 1 0 86050 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_12
timestamp 1704896540
transform 1 0 89212 0 1 5432
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_13
timestamp 1704896540
transform 1 0 84370 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_14
timestamp 1704896540
transform 1 0 82690 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_15
timestamp 1704896540
transform 1 0 81010 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_16
timestamp 1704896540
transform 1 0 89212 0 1 9464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_17
timestamp 1704896540
transform 1 0 89212 0 1 9128
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_18
timestamp 1704896540
transform 1 0 89212 0 1 8792
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_19
timestamp 1704896540
transform 1 0 89212 0 1 8456
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_20
timestamp 1704896540
transform 1 0 89212 0 1 8120
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_21
timestamp 1704896540
transform 1 0 89212 0 1 7784
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_22
timestamp 1704896540
transform 1 0 89212 0 1 7448
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_23
timestamp 1704896540
transform 1 0 89212 0 1 7112
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_24
timestamp 1704896540
transform 1 0 89212 0 1 6776
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_25
timestamp 1704896540
transform 1 0 89212 0 1 6440
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_26
timestamp 1704896540
transform 1 0 89212 0 1 6104
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_27
timestamp 1704896540
transform 1 0 89212 0 1 9800
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_28
timestamp 1704896540
transform 1 0 89212 0 1 11144
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_29
timestamp 1704896540
transform 1 0 89212 0 1 10808
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_30
timestamp 1704896540
transform 1 0 89212 0 1 10472
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_31
timestamp 1704896540
transform 1 0 89212 0 1 10136
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_32
timestamp 1704896540
transform 1 0 89212 0 1 5768
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_33
timestamp 1704896540
transform 1 0 72610 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_34
timestamp 1704896540
transform 1 0 70930 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_35
timestamp 1704896540
transform 1 0 69250 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_36
timestamp 1704896540
transform 1 0 78575 0 1 11062
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_37
timestamp 1704896540
transform 1 0 79330 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_38
timestamp 1704896540
transform 1 0 77650 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_39
timestamp 1704896540
transform 1 0 75970 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_40
timestamp 1704896540
transform 1 0 74290 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_41
timestamp 1704896540
transform 1 0 78975 0 1 17988
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_42
timestamp 1704896540
transform 1 0 79055 0 1 19546
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_43
timestamp 1704896540
transform 1 0 78655 0 1 12332
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_44
timestamp 1704896540
transform 1 0 78735 0 1 13890
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_45
timestamp 1704896540
transform 1 0 78815 0 1 15160
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_46
timestamp 1704896540
transform 1 0 78895 0 1 16718
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_47
timestamp 1704896540
transform 1 0 89212 0 1 13832
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_48
timestamp 1704896540
transform 1 0 89212 0 1 13496
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_49
timestamp 1704896540
transform 1 0 89212 0 1 13160
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_50
timestamp 1704896540
transform 1 0 89212 0 1 12824
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_51
timestamp 1704896540
transform 1 0 89212 0 1 12488
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_52
timestamp 1704896540
transform 1 0 89212 0 1 12152
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_53
timestamp 1704896540
transform 1 0 89212 0 1 11816
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_54
timestamp 1704896540
transform 1 0 89212 0 1 11480
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_55
timestamp 1704896540
transform 1 0 89212 0 1 16520
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_56
timestamp 1704896540
transform 1 0 89212 0 1 16184
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_57
timestamp 1704896540
transform 1 0 89212 0 1 15848
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_58
timestamp 1704896540
transform 1 0 89212 0 1 15512
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_59
timestamp 1704896540
transform 1 0 89212 0 1 15176
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_60
timestamp 1704896540
transform 1 0 89212 0 1 14840
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_61
timestamp 1704896540
transform 1 0 89212 0 1 14504
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_62
timestamp 1704896540
transform 1 0 89212 0 1 14168
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_63
timestamp 1704896540
transform 1 0 89212 0 1 22232
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_64
timestamp 1704896540
transform 1 0 89212 0 1 21896
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_65
timestamp 1704896540
transform 1 0 89212 0 1 21560
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_66
timestamp 1704896540
transform 1 0 89212 0 1 21224
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_67
timestamp 1704896540
transform 1 0 89212 0 1 20888
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_68
timestamp 1704896540
transform 1 0 89212 0 1 20552
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_69
timestamp 1704896540
transform 1 0 89212 0 1 20216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_70
timestamp 1704896540
transform 1 0 89212 0 1 19880
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_71
timestamp 1704896540
transform 1 0 89212 0 1 19544
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_72
timestamp 1704896540
transform 1 0 89212 0 1 19208
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_73
timestamp 1704896540
transform 1 0 89212 0 1 18872
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_74
timestamp 1704896540
transform 1 0 89212 0 1 18536
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_75
timestamp 1704896540
transform 1 0 89212 0 1 18200
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_76
timestamp 1704896540
transform 1 0 89212 0 1 17864
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_77
timestamp 1704896540
transform 1 0 89212 0 1 17528
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_78
timestamp 1704896540
transform 1 0 89212 0 1 17192
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_79
timestamp 1704896540
transform 1 0 89212 0 1 16856
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_80
timestamp 1704896540
transform 1 0 67570 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_81
timestamp 1704896540
transform 1 0 65890 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_82
timestamp 1704896540
transform 1 0 64210 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_83
timestamp 1704896540
transform 1 0 62530 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_84
timestamp 1704896540
transform 1 0 59170 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_85
timestamp 1704896540
transform 1 0 60850 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_86
timestamp 1704896540
transform 1 0 57490 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_87
timestamp 1704896540
transform 1 0 54130 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_88
timestamp 1704896540
transform 1 0 55810 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_89
timestamp 1704896540
transform 1 0 49090 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_90
timestamp 1704896540
transform 1 0 45730 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_91
timestamp 1704896540
transform 1 0 52450 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_92
timestamp 1704896540
transform 1 0 47410 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_93
timestamp 1704896540
transform 1 0 50770 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_94
timestamp 1704896540
transform 1 0 55574 0 1 13072
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_95
timestamp 1704896540
transform 1 0 50582 0 1 13072
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_96
timestamp 1704896540
transform 1 0 45590 0 1 13072
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_97
timestamp 1704896540
transform 1 0 60566 0 1 13072
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_98
timestamp 1704896540
transform 1 0 89212 0 1 22904
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_99
timestamp 1704896540
transform 1 0 89212 0 1 25256
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_100
timestamp 1704896540
transform 1 0 89212 0 1 24920
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_101
timestamp 1704896540
transform 1 0 89212 0 1 24584
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_102
timestamp 1704896540
transform 1 0 89212 0 1 24248
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_103
timestamp 1704896540
transform 1 0 89212 0 1 22568
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_104
timestamp 1704896540
transform 1 0 89212 0 1 27608
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_105
timestamp 1704896540
transform 1 0 89212 0 1 27272
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_106
timestamp 1704896540
transform 1 0 89212 0 1 26936
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_107
timestamp 1704896540
transform 1 0 89212 0 1 26600
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_108
timestamp 1704896540
transform 1 0 89212 0 1 26264
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_109
timestamp 1704896540
transform 1 0 89212 0 1 25928
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_110
timestamp 1704896540
transform 1 0 89212 0 1 23912
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_111
timestamp 1704896540
transform 1 0 89212 0 1 23576
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_112
timestamp 1704896540
transform 1 0 89212 0 1 23240
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_113
timestamp 1704896540
transform 1 0 89212 0 1 25592
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_114
timestamp 1704896540
transform 1 0 89212 0 1 29960
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_115
timestamp 1704896540
transform 1 0 89212 0 1 29624
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_116
timestamp 1704896540
transform 1 0 89212 0 1 29288
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_117
timestamp 1704896540
transform 1 0 89212 0 1 28952
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_118
timestamp 1704896540
transform 1 0 89212 0 1 28616
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_119
timestamp 1704896540
transform 1 0 89212 0 1 28280
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_120
timestamp 1704896540
transform 1 0 89212 0 1 30296
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_121
timestamp 1704896540
transform 1 0 89212 0 1 33320
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_122
timestamp 1704896540
transform 1 0 89212 0 1 32984
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_123
timestamp 1704896540
transform 1 0 89212 0 1 32648
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_124
timestamp 1704896540
transform 1 0 89212 0 1 32312
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_125
timestamp 1704896540
transform 1 0 89212 0 1 31976
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_126
timestamp 1704896540
transform 1 0 89212 0 1 31640
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_127
timestamp 1704896540
transform 1 0 89212 0 1 31304
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_128
timestamp 1704896540
transform 1 0 89212 0 1 30968
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_129
timestamp 1704896540
transform 1 0 89212 0 1 30632
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_130
timestamp 1704896540
transform 1 0 89212 0 1 27944
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_131
timestamp 1704896540
transform 1 0 89212 0 1 38360
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_132
timestamp 1704896540
transform 1 0 89212 0 1 38024
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_133
timestamp 1704896540
transform 1 0 89212 0 1 37688
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_134
timestamp 1704896540
transform 1 0 89212 0 1 37352
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_135
timestamp 1704896540
transform 1 0 89212 0 1 37016
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_136
timestamp 1704896540
transform 1 0 89212 0 1 36680
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_137
timestamp 1704896540
transform 1 0 89212 0 1 36344
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_138
timestamp 1704896540
transform 1 0 89212 0 1 36008
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_139
timestamp 1704896540
transform 1 0 89212 0 1 35672
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_140
timestamp 1704896540
transform 1 0 89212 0 1 35336
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_141
timestamp 1704896540
transform 1 0 89212 0 1 35000
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_142
timestamp 1704896540
transform 1 0 89212 0 1 34664
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_143
timestamp 1704896540
transform 1 0 89212 0 1 34328
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_144
timestamp 1704896540
transform 1 0 89212 0 1 33992
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_145
timestamp 1704896540
transform 1 0 89212 0 1 33656
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_146
timestamp 1704896540
transform 1 0 89212 0 1 39032
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_147
timestamp 1704896540
transform 1 0 89212 0 1 38696
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_148
timestamp 1704896540
transform 1 0 89212 0 1 44408
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_149
timestamp 1704896540
transform 1 0 89212 0 1 44072
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_150
timestamp 1704896540
transform 1 0 89212 0 1 43736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_151
timestamp 1704896540
transform 1 0 89212 0 1 43400
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_152
timestamp 1704896540
transform 1 0 89212 0 1 43064
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_153
timestamp 1704896540
transform 1 0 89212 0 1 42728
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_154
timestamp 1704896540
transform 1 0 89212 0 1 42392
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_155
timestamp 1704896540
transform 1 0 89212 0 1 42056
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_156
timestamp 1704896540
transform 1 0 89212 0 1 41720
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_157
timestamp 1704896540
transform 1 0 89212 0 1 41384
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_158
timestamp 1704896540
transform 1 0 89212 0 1 41048
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_159
timestamp 1704896540
transform 1 0 89212 0 1 40712
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_160
timestamp 1704896540
transform 1 0 89212 0 1 40376
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_161
timestamp 1704896540
transform 1 0 89212 0 1 40040
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_162
timestamp 1704896540
transform 1 0 89212 0 1 39704
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_163
timestamp 1704896540
transform 1 0 89212 0 1 39368
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_164
timestamp 1704896540
transform 1 0 37330 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_165
timestamp 1704896540
transform 1 0 40690 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_166
timestamp 1704896540
transform 1 0 39010 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_167
timestamp 1704896540
transform 1 0 44050 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_168
timestamp 1704896540
transform 1 0 35650 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_169
timestamp 1704896540
transform 1 0 42370 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_170
timestamp 1704896540
transform 1 0 33970 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_171
timestamp 1704896540
transform 1 0 28930 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_172
timestamp 1704896540
transform 1 0 32290 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_173
timestamp 1704896540
transform 1 0 30610 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_174
timestamp 1704896540
transform 1 0 23890 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_175
timestamp 1704896540
transform 1 0 27250 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_176
timestamp 1704896540
transform 1 0 25570 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_177
timestamp 1704896540
transform 1 0 30614 0 1 13072
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_178
timestamp 1704896540
transform 1 0 25622 0 1 13072
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_179
timestamp 1704896540
transform 1 0 40598 0 1 13072
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_180
timestamp 1704896540
transform 1 0 35606 0 1 13072
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_181
timestamp 1704896540
transform 1 0 18850 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_182
timestamp 1704896540
transform 1 0 20530 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_183
timestamp 1704896540
transform 1 0 22210 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_184
timestamp 1704896540
transform 1 0 13810 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_185
timestamp 1704896540
transform 1 0 17170 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_186
timestamp 1704896540
transform 1 0 12130 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_187
timestamp 1704896540
transform 1 0 15490 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_188
timestamp 1704896540
transform 1 0 7090 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_189
timestamp 1704896540
transform 1 0 10450 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_190
timestamp 1704896540
transform 1 0 8770 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_191
timestamp 1704896540
transform 1 0 1714 0 1 2072
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_192
timestamp 1704896540
transform 1 0 1714 0 1 5432
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_193
timestamp 1704896540
transform 1 0 1714 0 1 5096
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_194
timestamp 1704896540
transform 1 0 1714 0 1 4760
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_195
timestamp 1704896540
transform 1 0 1714 0 1 4424
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_196
timestamp 1704896540
transform 1 0 5410 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_197
timestamp 1704896540
transform 1 0 1714 0 1 4088
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_198
timestamp 1704896540
transform 1 0 3730 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_199
timestamp 1704896540
transform 1 0 1714 0 1 3752
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_200
timestamp 1704896540
transform 1 0 1714 0 1 3416
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_201
timestamp 1704896540
transform 1 0 2050 0 1 1736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_202
timestamp 1704896540
transform 1 0 1714 0 1 3080
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_203
timestamp 1704896540
transform 1 0 1714 0 1 2744
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_204
timestamp 1704896540
transform 1 0 1714 0 1 2408
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_205
timestamp 1704896540
transform 1 0 1714 0 1 11144
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_206
timestamp 1704896540
transform 1 0 1714 0 1 10808
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_207
timestamp 1704896540
transform 1 0 1714 0 1 10472
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_208
timestamp 1704896540
transform 1 0 1714 0 1 10136
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_209
timestamp 1704896540
transform 1 0 1714 0 1 9800
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_210
timestamp 1704896540
transform 1 0 1714 0 1 9464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_211
timestamp 1704896540
transform 1 0 1714 0 1 9128
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_212
timestamp 1704896540
transform 1 0 1714 0 1 8792
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_213
timestamp 1704896540
transform 1 0 1714 0 1 8456
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_214
timestamp 1704896540
transform 1 0 1714 0 1 8120
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_215
timestamp 1704896540
transform 1 0 1714 0 1 7784
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_216
timestamp 1704896540
transform 1 0 1714 0 1 7448
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_217
timestamp 1704896540
transform 1 0 1714 0 1 7112
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_218
timestamp 1704896540
transform 1 0 1714 0 1 6776
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_219
timestamp 1704896540
transform 1 0 1714 0 1 6440
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_220
timestamp 1704896540
transform 1 0 1714 0 1 6104
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_221
timestamp 1704896540
transform 1 0 1714 0 1 5768
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_222
timestamp 1704896540
transform 1 0 1714 0 1 14840
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_223
timestamp 1704896540
transform 1 0 1714 0 1 14504
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_224
timestamp 1704896540
transform 1 0 1714 0 1 12152
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_225
timestamp 1704896540
transform 1 0 1714 0 1 11816
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_226
timestamp 1704896540
transform 1 0 1714 0 1 11480
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_227
timestamp 1704896540
transform 1 0 1714 0 1 14168
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_228
timestamp 1704896540
transform 1 0 1714 0 1 13160
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_229
timestamp 1704896540
transform 1 0 1714 0 1 13832
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_230
timestamp 1704896540
transform 1 0 1714 0 1 12824
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_231
timestamp 1704896540
transform 1 0 1714 0 1 12488
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_232
timestamp 1704896540
transform 1 0 1714 0 1 16184
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_233
timestamp 1704896540
transform 1 0 1714 0 1 15848
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_234
timestamp 1704896540
transform 1 0 1714 0 1 13496
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_235
timestamp 1704896540
transform 1 0 1714 0 1 15512
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_236
timestamp 1704896540
transform 1 0 1714 0 1 15176
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_237
timestamp 1704896540
transform 1 0 1714 0 1 16520
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_238
timestamp 1704896540
transform 1 0 1714 0 1 22232
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_239
timestamp 1704896540
transform 1 0 1714 0 1 21896
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_240
timestamp 1704896540
transform 1 0 1714 0 1 21560
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_241
timestamp 1704896540
transform 1 0 1714 0 1 21224
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_242
timestamp 1704896540
transform 1 0 1714 0 1 20888
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_243
timestamp 1704896540
transform 1 0 1714 0 1 20552
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_244
timestamp 1704896540
transform 1 0 1714 0 1 20216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_245
timestamp 1704896540
transform 1 0 1714 0 1 19880
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_246
timestamp 1704896540
transform 1 0 1714 0 1 19544
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_247
timestamp 1704896540
transform 1 0 1714 0 1 19208
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_248
timestamp 1704896540
transform 1 0 1714 0 1 18872
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_249
timestamp 1704896540
transform 1 0 1714 0 1 18536
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_250
timestamp 1704896540
transform 1 0 1714 0 1 18200
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_251
timestamp 1704896540
transform 1 0 1714 0 1 17864
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_252
timestamp 1704896540
transform 1 0 1714 0 1 17528
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_253
timestamp 1704896540
transform 1 0 1714 0 1 17192
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_254
timestamp 1704896540
transform 1 0 1714 0 1 16856
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_255
timestamp 1704896540
transform 1 0 11951 0 1 30274
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_256
timestamp 1704896540
transform 1 0 11871 0 1 28716
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_257
timestamp 1704896540
transform 1 0 12111 0 1 33102
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_258
timestamp 1704896540
transform 1 0 12031 0 1 31544
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_259
timestamp 1704896540
transform 1 0 1714 0 1 24920
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_260
timestamp 1704896540
transform 1 0 1714 0 1 24584
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_261
timestamp 1704896540
transform 1 0 1714 0 1 24248
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_262
timestamp 1704896540
transform 1 0 1714 0 1 23912
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_263
timestamp 1704896540
transform 1 0 1714 0 1 23576
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_264
timestamp 1704896540
transform 1 0 1714 0 1 23240
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_265
timestamp 1704896540
transform 1 0 1714 0 1 22904
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_266
timestamp 1704896540
transform 1 0 1714 0 1 27608
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_267
timestamp 1704896540
transform 1 0 1714 0 1 27272
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_268
timestamp 1704896540
transform 1 0 1714 0 1 26936
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_269
timestamp 1704896540
transform 1 0 1714 0 1 26600
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_270
timestamp 1704896540
transform 1 0 1714 0 1 26264
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_271
timestamp 1704896540
transform 1 0 1714 0 1 25928
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_272
timestamp 1704896540
transform 1 0 1714 0 1 25592
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_273
timestamp 1704896540
transform 1 0 1714 0 1 25256
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_274
timestamp 1704896540
transform 1 0 1714 0 1 22568
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_275
timestamp 1704896540
transform 1 0 1714 0 1 30296
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_276
timestamp 1704896540
transform 1 0 1714 0 1 29960
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_277
timestamp 1704896540
transform 1 0 1714 0 1 29624
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_278
timestamp 1704896540
transform 1 0 1714 0 1 29288
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_279
timestamp 1704896540
transform 1 0 1714 0 1 28952
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_280
timestamp 1704896540
transform 1 0 1714 0 1 31640
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_281
timestamp 1704896540
transform 1 0 1714 0 1 28616
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_282
timestamp 1704896540
transform 1 0 1714 0 1 28280
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_283
timestamp 1704896540
transform 1 0 1714 0 1 31304
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_284
timestamp 1704896540
transform 1 0 1714 0 1 30968
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_285
timestamp 1704896540
transform 1 0 1714 0 1 30632
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_286
timestamp 1704896540
transform 1 0 1714 0 1 33320
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_287
timestamp 1704896540
transform 1 0 1714 0 1 32984
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_288
timestamp 1704896540
transform 1 0 1714 0 1 32648
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_289
timestamp 1704896540
transform 1 0 1714 0 1 32312
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_290
timestamp 1704896540
transform 1 0 1714 0 1 31976
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_291
timestamp 1704896540
transform 1 0 1714 0 1 27944
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_292
timestamp 1704896540
transform 1 0 1714 0 1 34328
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_293
timestamp 1704896540
transform 1 0 1714 0 1 33992
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_294
timestamp 1704896540
transform 1 0 1714 0 1 39032
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_295
timestamp 1704896540
transform 1 0 1714 0 1 38696
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_296
timestamp 1704896540
transform 1 0 1714 0 1 38360
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_297
timestamp 1704896540
transform 1 0 1714 0 1 38024
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_298
timestamp 1704896540
transform 1 0 1714 0 1 37688
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_299
timestamp 1704896540
transform 1 0 1714 0 1 37352
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_300
timestamp 1704896540
transform 1 0 1714 0 1 37016
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_301
timestamp 1704896540
transform 1 0 1714 0 1 36680
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_302
timestamp 1704896540
transform 1 0 1714 0 1 36344
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_303
timestamp 1704896540
transform 1 0 1714 0 1 36008
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_304
timestamp 1704896540
transform 1 0 1714 0 1 35672
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_305
timestamp 1704896540
transform 1 0 1714 0 1 35336
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_306
timestamp 1704896540
transform 1 0 1714 0 1 33656
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_307
timestamp 1704896540
transform 1 0 1714 0 1 35000
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_308
timestamp 1704896540
transform 1 0 1714 0 1 34664
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_309
timestamp 1704896540
transform 1 0 1714 0 1 39704
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_310
timestamp 1704896540
transform 1 0 1714 0 1 39368
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_311
timestamp 1704896540
transform 1 0 1714 0 1 44408
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_312
timestamp 1704896540
transform 1 0 1714 0 1 44072
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_313
timestamp 1704896540
transform 1 0 1714 0 1 43736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_314
timestamp 1704896540
transform 1 0 1714 0 1 43400
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_315
timestamp 1704896540
transform 1 0 1714 0 1 43064
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_316
timestamp 1704896540
transform 1 0 1714 0 1 42728
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_317
timestamp 1704896540
transform 1 0 1714 0 1 42392
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_318
timestamp 1704896540
transform 1 0 1714 0 1 42056
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_319
timestamp 1704896540
transform 1 0 1714 0 1 41720
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_320
timestamp 1704896540
transform 1 0 1714 0 1 41384
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_321
timestamp 1704896540
transform 1 0 1714 0 1 41048
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_322
timestamp 1704896540
transform 1 0 1714 0 1 40712
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_323
timestamp 1704896540
transform 1 0 1714 0 1 40376
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_324
timestamp 1704896540
transform 1 0 1714 0 1 40040
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_325
timestamp 1704896540
transform 1 0 12271 0 1 35930
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_326
timestamp 1704896540
transform 1 0 12191 0 1 34372
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_327
timestamp 1704896540
transform 1 0 12351 0 1 37200
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_328
timestamp 1704896540
transform 1 0 1714 0 1 47432
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_329
timestamp 1704896540
transform 1 0 1714 0 1 47096
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_330
timestamp 1704896540
transform 1 0 1714 0 1 46760
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_331
timestamp 1704896540
transform 1 0 1714 0 1 46424
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_332
timestamp 1704896540
transform 1 0 1714 0 1 46088
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_333
timestamp 1704896540
transform 1 0 1714 0 1 45752
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_334
timestamp 1704896540
transform 1 0 1714 0 1 45416
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_335
timestamp 1704896540
transform 1 0 1714 0 1 45080
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_336
timestamp 1704896540
transform 1 0 1714 0 1 44744
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_337
timestamp 1704896540
transform 1 0 1714 0 1 50120
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_338
timestamp 1704896540
transform 1 0 1714 0 1 49784
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_339
timestamp 1704896540
transform 1 0 1714 0 1 49448
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_340
timestamp 1704896540
transform 1 0 1714 0 1 49112
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_341
timestamp 1704896540
transform 1 0 1714 0 1 48776
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_342
timestamp 1704896540
transform 1 0 1714 0 1 48440
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_343
timestamp 1704896540
transform 1 0 1714 0 1 48104
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_344
timestamp 1704896540
transform 1 0 1714 0 1 47768
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_345
timestamp 1704896540
transform 1 0 1714 0 1 53480
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_346
timestamp 1704896540
transform 1 0 1714 0 1 53144
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_347
timestamp 1704896540
transform 1 0 1714 0 1 52808
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_348
timestamp 1704896540
transform 1 0 1714 0 1 52472
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_349
timestamp 1704896540
transform 1 0 1714 0 1 52136
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_350
timestamp 1704896540
transform 1 0 1714 0 1 51800
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_351
timestamp 1704896540
transform 1 0 1714 0 1 51464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_352
timestamp 1704896540
transform 1 0 1714 0 1 51128
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_353
timestamp 1704896540
transform 1 0 1714 0 1 50792
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_354
timestamp 1704896540
transform 1 0 1714 0 1 50456
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_355
timestamp 1704896540
transform 1 0 1714 0 1 55160
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_356
timestamp 1704896540
transform 1 0 1714 0 1 55496
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_357
timestamp 1704896540
transform 1 0 1714 0 1 53816
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_358
timestamp 1704896540
transform 1 0 1714 0 1 54488
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_359
timestamp 1704896540
transform 1 0 1714 0 1 54152
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_360
timestamp 1704896540
transform 1 0 1714 0 1 54824
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_361
timestamp 1704896540
transform 1 0 1714 0 1 57848
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_362
timestamp 1704896540
transform 1 0 1714 0 1 61208
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_363
timestamp 1704896540
transform 1 0 1714 0 1 56168
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_364
timestamp 1704896540
transform 1 0 1714 0 1 57512
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_365
timestamp 1704896540
transform 1 0 1714 0 1 57176
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_366
timestamp 1704896540
transform 1 0 1714 0 1 56840
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_367
timestamp 1704896540
transform 1 0 1714 0 1 56504
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_368
timestamp 1704896540
transform 1 0 1714 0 1 58520
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_369
timestamp 1704896540
transform 1 0 1714 0 1 58184
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_370
timestamp 1704896540
transform 1 0 1714 0 1 60872
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_371
timestamp 1704896540
transform 1 0 1714 0 1 60536
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_372
timestamp 1704896540
transform 1 0 1714 0 1 60200
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_373
timestamp 1704896540
transform 1 0 1714 0 1 55832
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_374
timestamp 1704896540
transform 1 0 1714 0 1 59864
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_375
timestamp 1704896540
transform 1 0 1714 0 1 59528
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_376
timestamp 1704896540
transform 1 0 1714 0 1 59192
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_377
timestamp 1704896540
transform 1 0 1714 0 1 58856
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_378
timestamp 1704896540
transform 1 0 1714 0 1 64904
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_379
timestamp 1704896540
transform 1 0 1714 0 1 64568
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_380
timestamp 1704896540
transform 1 0 1714 0 1 64232
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_381
timestamp 1704896540
transform 1 0 1714 0 1 63896
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_382
timestamp 1704896540
transform 1 0 1714 0 1 63560
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_383
timestamp 1704896540
transform 1 0 1714 0 1 63224
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_384
timestamp 1704896540
transform 1 0 1714 0 1 62888
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_385
timestamp 1704896540
transform 1 0 1714 0 1 62552
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_386
timestamp 1704896540
transform 1 0 1714 0 1 62216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_387
timestamp 1704896540
transform 1 0 1714 0 1 61880
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_388
timestamp 1704896540
transform 1 0 1714 0 1 61544
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_389
timestamp 1704896540
transform 1 0 1714 0 1 66584
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_390
timestamp 1704896540
transform 1 0 1714 0 1 66248
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_391
timestamp 1704896540
transform 1 0 1714 0 1 65240
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_392
timestamp 1704896540
transform 1 0 1714 0 1 65912
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_393
timestamp 1704896540
transform 1 0 1714 0 1 65576
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_394
timestamp 1704896540
transform 1 0 1714 0 1 71288
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_395
timestamp 1704896540
transform 1 0 1714 0 1 70952
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_396
timestamp 1704896540
transform 1 0 1714 0 1 70616
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_397
timestamp 1704896540
transform 1 0 1714 0 1 70280
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_398
timestamp 1704896540
transform 1 0 1714 0 1 69944
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_399
timestamp 1704896540
transform 1 0 1714 0 1 69608
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_400
timestamp 1704896540
transform 1 0 1714 0 1 69272
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_401
timestamp 1704896540
transform 1 0 1714 0 1 68936
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_402
timestamp 1704896540
transform 1 0 1714 0 1 68600
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_403
timestamp 1704896540
transform 1 0 1714 0 1 68264
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_404
timestamp 1704896540
transform 1 0 1714 0 1 67928
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_405
timestamp 1704896540
transform 1 0 1714 0 1 67592
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_406
timestamp 1704896540
transform 1 0 1714 0 1 67256
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_407
timestamp 1704896540
transform 1 0 1714 0 1 66920
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_408
timestamp 1704896540
transform 1 0 1714 0 1 72296
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_409
timestamp 1704896540
transform 1 0 1714 0 1 71960
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_410
timestamp 1704896540
transform 1 0 1714 0 1 71624
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_411
timestamp 1704896540
transform 1 0 1714 0 1 77336
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_412
timestamp 1704896540
transform 1 0 1714 0 1 77000
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_413
timestamp 1704896540
transform 1 0 1714 0 1 76664
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_414
timestamp 1704896540
transform 1 0 1714 0 1 76328
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_415
timestamp 1704896540
transform 1 0 1714 0 1 75992
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_416
timestamp 1704896540
transform 1 0 1714 0 1 75656
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_417
timestamp 1704896540
transform 1 0 1714 0 1 75320
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_418
timestamp 1704896540
transform 1 0 1714 0 1 74984
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_419
timestamp 1704896540
transform 1 0 1714 0 1 74648
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_420
timestamp 1704896540
transform 1 0 1714 0 1 74312
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_421
timestamp 1704896540
transform 1 0 1714 0 1 73976
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_422
timestamp 1704896540
transform 1 0 1714 0 1 73640
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_423
timestamp 1704896540
transform 1 0 1714 0 1 73304
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_424
timestamp 1704896540
transform 1 0 1714 0 1 72968
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_425
timestamp 1704896540
transform 1 0 1714 0 1 72632
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_426
timestamp 1704896540
transform 1 0 1714 0 1 77672
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_427
timestamp 1704896540
transform 1 0 1714 0 1 82040
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_428
timestamp 1704896540
transform 1 0 1714 0 1 81704
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_429
timestamp 1704896540
transform 1 0 1714 0 1 81368
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_430
timestamp 1704896540
transform 1 0 1714 0 1 79016
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_431
timestamp 1704896540
transform 1 0 1714 0 1 78680
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_432
timestamp 1704896540
transform 1 0 1714 0 1 78344
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_433
timestamp 1704896540
transform 1 0 1714 0 1 78008
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_434
timestamp 1704896540
transform 1 0 1714 0 1 81032
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_435
timestamp 1704896540
transform 1 0 1714 0 1 80696
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_436
timestamp 1704896540
transform 1 0 1714 0 1 80360
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_437
timestamp 1704896540
transform 1 0 1714 0 1 80024
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_438
timestamp 1704896540
transform 1 0 1714 0 1 79688
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_439
timestamp 1704896540
transform 1 0 1714 0 1 79352
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_440
timestamp 1704896540
transform 1 0 1714 0 1 83384
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_441
timestamp 1704896540
transform 1 0 1714 0 1 83048
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_442
timestamp 1704896540
transform 1 0 1714 0 1 82712
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_443
timestamp 1704896540
transform 1 0 1714 0 1 82376
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_444
timestamp 1704896540
transform 1 0 1714 0 1 87080
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_445
timestamp 1704896540
transform 1 0 1714 0 1 86744
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_446
timestamp 1704896540
transform 1 0 1714 0 1 86408
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_447
timestamp 1704896540
transform 1 0 1714 0 1 86072
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_448
timestamp 1704896540
transform 1 0 1714 0 1 85736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_449
timestamp 1704896540
transform 1 0 1714 0 1 85400
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_450
timestamp 1704896540
transform 1 0 1714 0 1 85064
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_451
timestamp 1704896540
transform 1 0 1714 0 1 84728
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_452
timestamp 1704896540
transform 1 0 1714 0 1 84392
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_453
timestamp 1704896540
transform 1 0 1714 0 1 84056
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_454
timestamp 1704896540
transform 1 0 1714 0 1 83720
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_455
timestamp 1704896540
transform 1 0 5410 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_456
timestamp 1704896540
transform 1 0 3730 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_457
timestamp 1704896540
transform 1 0 2050 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_458
timestamp 1704896540
transform 1 0 10450 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_459
timestamp 1704896540
transform 1 0 8770 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_460
timestamp 1704896540
transform 1 0 7090 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_461
timestamp 1704896540
transform 1 0 22210 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_462
timestamp 1704896540
transform 1 0 20530 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_463
timestamp 1704896540
transform 1 0 18850 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_464
timestamp 1704896540
transform 1 0 17170 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_465
timestamp 1704896540
transform 1 0 15490 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_466
timestamp 1704896540
transform 1 0 13810 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_467
timestamp 1704896540
transform 1 0 12130 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_468
timestamp 1704896540
transform 1 0 40598 0 1 77850
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_469
timestamp 1704896540
transform 1 0 35606 0 1 77850
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_470
timestamp 1704896540
transform 1 0 30614 0 1 77850
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_471
timestamp 1704896540
transform 1 0 25622 0 1 77850
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_472
timestamp 1704896540
transform 1 0 28930 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_473
timestamp 1704896540
transform 1 0 27250 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_474
timestamp 1704896540
transform 1 0 25570 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_475
timestamp 1704896540
transform 1 0 23890 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_476
timestamp 1704896540
transform 1 0 33970 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_477
timestamp 1704896540
transform 1 0 32290 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_478
timestamp 1704896540
transform 1 0 30610 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_479
timestamp 1704896540
transform 1 0 42370 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_480
timestamp 1704896540
transform 1 0 40690 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_481
timestamp 1704896540
transform 1 0 39010 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_482
timestamp 1704896540
transform 1 0 37330 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_483
timestamp 1704896540
transform 1 0 35650 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_484
timestamp 1704896540
transform 1 0 44050 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_485
timestamp 1704896540
transform 1 0 89212 0 1 47096
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_486
timestamp 1704896540
transform 1 0 89212 0 1 46760
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_487
timestamp 1704896540
transform 1 0 89212 0 1 46424
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_488
timestamp 1704896540
transform 1 0 89212 0 1 48440
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_489
timestamp 1704896540
transform 1 0 89212 0 1 48104
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_490
timestamp 1704896540
transform 1 0 89212 0 1 50120
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_491
timestamp 1704896540
transform 1 0 89212 0 1 49784
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_492
timestamp 1704896540
transform 1 0 89212 0 1 49448
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_493
timestamp 1704896540
transform 1 0 89212 0 1 46088
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_494
timestamp 1704896540
transform 1 0 89212 0 1 49112
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_495
timestamp 1704896540
transform 1 0 89212 0 1 48776
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_496
timestamp 1704896540
transform 1 0 89212 0 1 45752
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_497
timestamp 1704896540
transform 1 0 89212 0 1 45416
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_498
timestamp 1704896540
transform 1 0 89212 0 1 47768
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_499
timestamp 1704896540
transform 1 0 89212 0 1 47432
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_500
timestamp 1704896540
transform 1 0 89212 0 1 45080
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_501
timestamp 1704896540
transform 1 0 89212 0 1 44744
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_502
timestamp 1704896540
transform 1 0 89212 0 1 55496
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_503
timestamp 1704896540
transform 1 0 89212 0 1 55160
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_504
timestamp 1704896540
transform 1 0 89212 0 1 54824
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_505
timestamp 1704896540
transform 1 0 89212 0 1 54488
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_506
timestamp 1704896540
transform 1 0 89212 0 1 54152
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_507
timestamp 1704896540
transform 1 0 89212 0 1 52136
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_508
timestamp 1704896540
transform 1 0 89212 0 1 53816
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_509
timestamp 1704896540
transform 1 0 89212 0 1 53480
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_510
timestamp 1704896540
transform 1 0 89212 0 1 50456
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_511
timestamp 1704896540
transform 1 0 89212 0 1 51800
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_512
timestamp 1704896540
transform 1 0 89212 0 1 53144
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_513
timestamp 1704896540
transform 1 0 89212 0 1 51464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_514
timestamp 1704896540
transform 1 0 89212 0 1 51128
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_515
timestamp 1704896540
transform 1 0 89212 0 1 50792
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_516
timestamp 1704896540
transform 1 0 89212 0 1 52808
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_517
timestamp 1704896540
transform 1 0 89212 0 1 52472
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_518
timestamp 1704896540
transform 1 0 89212 0 1 57512
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_519
timestamp 1704896540
transform 1 0 89212 0 1 55832
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_520
timestamp 1704896540
transform 1 0 89212 0 1 57176
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_521
timestamp 1704896540
transform 1 0 89212 0 1 56840
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_522
timestamp 1704896540
transform 1 0 89212 0 1 56504
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_523
timestamp 1704896540
transform 1 0 89212 0 1 56168
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_524
timestamp 1704896540
transform 1 0 89212 0 1 61208
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_525
timestamp 1704896540
transform 1 0 89212 0 1 60872
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_526
timestamp 1704896540
transform 1 0 89212 0 1 60536
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_527
timestamp 1704896540
transform 1 0 89212 0 1 60200
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_528
timestamp 1704896540
transform 1 0 89212 0 1 59864
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_529
timestamp 1704896540
transform 1 0 89212 0 1 59528
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_530
timestamp 1704896540
transform 1 0 89212 0 1 59192
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_531
timestamp 1704896540
transform 1 0 89212 0 1 58856
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_532
timestamp 1704896540
transform 1 0 89212 0 1 58520
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_533
timestamp 1704896540
transform 1 0 89212 0 1 58184
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_534
timestamp 1704896540
transform 1 0 89212 0 1 57848
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_535
timestamp 1704896540
transform 1 0 89212 0 1 66584
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_536
timestamp 1704896540
transform 1 0 89212 0 1 66248
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_537
timestamp 1704896540
transform 1 0 89212 0 1 65912
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_538
timestamp 1704896540
transform 1 0 89212 0 1 65576
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_539
timestamp 1704896540
transform 1 0 89212 0 1 65240
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_540
timestamp 1704896540
transform 1 0 89212 0 1 64904
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_541
timestamp 1704896540
transform 1 0 89212 0 1 64568
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_542
timestamp 1704896540
transform 1 0 89212 0 1 64232
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_543
timestamp 1704896540
transform 1 0 89212 0 1 63896
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_544
timestamp 1704896540
transform 1 0 89212 0 1 63560
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_545
timestamp 1704896540
transform 1 0 89212 0 1 63224
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_546
timestamp 1704896540
transform 1 0 89212 0 1 62888
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_547
timestamp 1704896540
transform 1 0 89212 0 1 62552
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_548
timestamp 1704896540
transform 1 0 89212 0 1 62216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_549
timestamp 1704896540
transform 1 0 89212 0 1 61880
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_550
timestamp 1704896540
transform 1 0 89212 0 1 61544
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_551
timestamp 1704896540
transform 1 0 60566 0 1 77850
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_552
timestamp 1704896540
transform 1 0 50582 0 1 77850
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_553
timestamp 1704896540
transform 1 0 45590 0 1 77850
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_554
timestamp 1704896540
transform 1 0 55574 0 1 77850
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_555
timestamp 1704896540
transform 1 0 45730 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_556
timestamp 1704896540
transform 1 0 54130 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_557
timestamp 1704896540
transform 1 0 52450 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_558
timestamp 1704896540
transform 1 0 50770 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_559
timestamp 1704896540
transform 1 0 49090 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_560
timestamp 1704896540
transform 1 0 47410 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_561
timestamp 1704896540
transform 1 0 55810 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_562
timestamp 1704896540
transform 1 0 67570 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_563
timestamp 1704896540
transform 1 0 65890 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_564
timestamp 1704896540
transform 1 0 64210 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_565
timestamp 1704896540
transform 1 0 62530 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_566
timestamp 1704896540
transform 1 0 60850 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_567
timestamp 1704896540
transform 1 0 59170 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_568
timestamp 1704896540
transform 1 0 57490 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_569
timestamp 1704896540
transform 1 0 89212 0 1 70952
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_570
timestamp 1704896540
transform 1 0 89212 0 1 70616
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_571
timestamp 1704896540
transform 1 0 89212 0 1 70280
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_572
timestamp 1704896540
transform 1 0 89212 0 1 69944
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_573
timestamp 1704896540
transform 1 0 89212 0 1 69608
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_574
timestamp 1704896540
transform 1 0 89212 0 1 69272
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_575
timestamp 1704896540
transform 1 0 89212 0 1 68936
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_576
timestamp 1704896540
transform 1 0 89212 0 1 68600
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_577
timestamp 1704896540
transform 1 0 89212 0 1 71960
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_578
timestamp 1704896540
transform 1 0 89212 0 1 68264
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_579
timestamp 1704896540
transform 1 0 89212 0 1 67928
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_580
timestamp 1704896540
transform 1 0 89212 0 1 67592
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_581
timestamp 1704896540
transform 1 0 89212 0 1 67256
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_582
timestamp 1704896540
transform 1 0 89212 0 1 66920
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_583
timestamp 1704896540
transform 1 0 89212 0 1 71624
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_584
timestamp 1704896540
transform 1 0 89212 0 1 71288
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_585
timestamp 1704896540
transform 1 0 89212 0 1 72296
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_586
timestamp 1704896540
transform 1 0 89212 0 1 77672
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_587
timestamp 1704896540
transform 1 0 89212 0 1 77336
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_588
timestamp 1704896540
transform 1 0 89212 0 1 77000
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_589
timestamp 1704896540
transform 1 0 89212 0 1 76664
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_590
timestamp 1704896540
transform 1 0 89212 0 1 76328
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_591
timestamp 1704896540
transform 1 0 89212 0 1 75992
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_592
timestamp 1704896540
transform 1 0 89212 0 1 75656
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_593
timestamp 1704896540
transform 1 0 89212 0 1 75320
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_594
timestamp 1704896540
transform 1 0 89212 0 1 74984
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_595
timestamp 1704896540
transform 1 0 89212 0 1 74648
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_596
timestamp 1704896540
transform 1 0 89212 0 1 74312
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_597
timestamp 1704896540
transform 1 0 89212 0 1 73976
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_598
timestamp 1704896540
transform 1 0 89212 0 1 73640
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_599
timestamp 1704896540
transform 1 0 89212 0 1 73304
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_600
timestamp 1704896540
transform 1 0 89212 0 1 72968
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_601
timestamp 1704896540
transform 1 0 89212 0 1 72632
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_602
timestamp 1704896540
transform 1 0 70930 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_603
timestamp 1704896540
transform 1 0 69250 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_604
timestamp 1704896540
transform 1 0 72610 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_605
timestamp 1704896540
transform 1 0 79330 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_606
timestamp 1704896540
transform 1 0 77650 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_607
timestamp 1704896540
transform 1 0 75970 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_608
timestamp 1704896540
transform 1 0 74290 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_609
timestamp 1704896540
transform 1 0 89212 0 1 79352
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_610
timestamp 1704896540
transform 1 0 89212 0 1 79016
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_611
timestamp 1704896540
transform 1 0 89212 0 1 78680
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_612
timestamp 1704896540
transform 1 0 89212 0 1 78344
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_613
timestamp 1704896540
transform 1 0 89212 0 1 78008
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_614
timestamp 1704896540
transform 1 0 89212 0 1 83384
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_615
timestamp 1704896540
transform 1 0 89212 0 1 83048
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_616
timestamp 1704896540
transform 1 0 89212 0 1 82712
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_617
timestamp 1704896540
transform 1 0 89212 0 1 82376
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_618
timestamp 1704896540
transform 1 0 89212 0 1 82040
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_619
timestamp 1704896540
transform 1 0 89212 0 1 81704
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_620
timestamp 1704896540
transform 1 0 89212 0 1 81368
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_621
timestamp 1704896540
transform 1 0 89212 0 1 81032
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_622
timestamp 1704896540
transform 1 0 89212 0 1 80696
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_623
timestamp 1704896540
transform 1 0 89212 0 1 80360
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_624
timestamp 1704896540
transform 1 0 89212 0 1 80024
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_625
timestamp 1704896540
transform 1 0 89212 0 1 79688
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_626
timestamp 1704896540
transform 1 0 81010 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_627
timestamp 1704896540
transform 1 0 84370 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_628
timestamp 1704896540
transform 1 0 82690 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_629
timestamp 1704896540
transform 1 0 89212 0 1 87080
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_630
timestamp 1704896540
transform 1 0 89212 0 1 86744
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_631
timestamp 1704896540
transform 1 0 89212 0 1 86408
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_632
timestamp 1704896540
transform 1 0 89212 0 1 86072
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_633
timestamp 1704896540
transform 1 0 89212 0 1 85736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_634
timestamp 1704896540
transform 1 0 89212 0 1 85400
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_635
timestamp 1704896540
transform 1 0 89212 0 1 85064
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_636
timestamp 1704896540
transform 1 0 89212 0 1 84728
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_637
timestamp 1704896540
transform 1 0 89212 0 1 84392
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_638
timestamp 1704896540
transform 1 0 89212 0 1 84056
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_639
timestamp 1704896540
transform 1 0 89212 0 1 83720
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_640
timestamp 1704896540
transform 1 0 87730 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_641
timestamp 1704896540
transform 1 0 86050 0 1 87464
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_32  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_32_0
timestamp 1704896540
transform 1 0 79255 0 1 19868
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_32  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_32_1
timestamp 1704896540
transform 1 0 11753 0 1 2711
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_32  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_32_2
timestamp 1704896540
transform 1 0 11753 0 1 28384
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_32  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_32_3
timestamp 1704896540
transform 1 0 79255 0 1 86479
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_0
timestamp 1704896540
transform 1 0 89760 0 1 2045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1
timestamp 1704896540
transform 1 0 87584 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2
timestamp 1704896540
transform 1 0 87584 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_3
timestamp 1704896540
transform 1 0 86088 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_4
timestamp 1704896540
transform 1 0 86088 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_5
timestamp 1704896540
transform 1 0 89760 0 1 3677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_6
timestamp 1704896540
transform 1 0 89760 0 1 5309
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_7
timestamp 1704896540
transform 1 0 84320 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_8
timestamp 1704896540
transform 1 0 82824 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_9
timestamp 1704896540
transform 1 0 82824 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_10
timestamp 1704896540
transform 1 0 80920 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_11
timestamp 1704896540
transform 1 0 80920 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_12
timestamp 1704896540
transform 1 0 84320 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_13
timestamp 1704896540
transform 1 0 79832 0 1 10341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_14
timestamp 1704896540
transform 1 0 89760 0 1 10341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_15
timestamp 1704896540
transform 1 0 89760 0 1 7213
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_16
timestamp 1704896540
transform 1 0 89760 0 1 8709
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_17
timestamp 1704896540
transform 1 0 70856 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_18
timestamp 1704896540
transform 1 0 70856 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_19
timestamp 1704896540
transform 1 0 69360 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_20
timestamp 1704896540
transform 1 0 75888 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_21
timestamp 1704896540
transform 1 0 75888 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_22
timestamp 1704896540
transform 1 0 74392 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_23
timestamp 1704896540
transform 1 0 79288 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_24
timestamp 1704896540
transform 1 0 79288 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_25
timestamp 1704896540
transform 1 0 69360 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_26
timestamp 1704896540
transform 1 0 77656 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_27
timestamp 1704896540
transform 1 0 74392 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_28
timestamp 1704896540
transform 1 0 72624 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_29
timestamp 1704896540
transform 1 0 72624 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_30
timestamp 1704896540
transform 1 0 77656 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_31
timestamp 1704896540
transform 1 0 72896 0 1 21493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_32
timestamp 1704896540
transform 1 0 73032 0 1 21085
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_33
timestamp 1704896540
transform 1 0 73032 0 1 21357
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_34
timestamp 1704896540
transform 1 0 74800 0 1 21221
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_35
timestamp 1704896540
transform 1 0 71672 0 1 22173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_36
timestamp 1704896540
transform 1 0 71808 0 1 20949
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_37
timestamp 1704896540
transform 1 0 77112 0 1 20541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_38
timestamp 1704896540
transform 1 0 71400 0 1 20949
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_39
timestamp 1704896540
transform 1 0 75888 0 1 20677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_40
timestamp 1704896540
transform 1 0 75888 0 1 21357
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_41
timestamp 1704896540
transform 1 0 75072 0 1 21493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_42
timestamp 1704896540
transform 1 0 75072 0 1 21221
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_43
timestamp 1704896540
transform 1 0 75072 0 1 20677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_44
timestamp 1704896540
transform 1 0 72080 0 1 22037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_45
timestamp 1704896540
transform 1 0 72080 0 1 21765
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_46
timestamp 1704896540
transform 1 0 71400 0 1 20677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_47
timestamp 1704896540
transform 1 0 75480 0 1 20677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_48
timestamp 1704896540
transform 1 0 75480 0 1 21357
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_49
timestamp 1704896540
transform 1 0 74800 0 1 20677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_50
timestamp 1704896540
transform 1 0 71264 0 1 22173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_51
timestamp 1704896540
transform 1 0 77112 0 1 18909
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_52
timestamp 1704896540
transform 1 0 71808 0 1 20677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_53
timestamp 1704896540
transform 1 0 75480 0 1 21493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_54
timestamp 1704896540
transform 1 0 72216 0 1 21085
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_55
timestamp 1704896540
transform 1 0 72216 0 1 21357
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_56
timestamp 1704896540
transform 1 0 72896 0 1 22309
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_57
timestamp 1704896540
transform 1 0 73032 0 1 20677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_58
timestamp 1704896540
transform 1 0 73032 0 1 20949
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_59
timestamp 1704896540
transform 1 0 72896 0 1 21765
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_60
timestamp 1704896540
transform 1 0 89760 0 1 15509
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_61
timestamp 1704896540
transform 1 0 89760 0 1 12245
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_62
timestamp 1704896540
transform 1 0 89760 0 1 13877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_63
timestamp 1704896540
transform 1 0 79968 0 1 14557
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_64
timestamp 1704896540
transform 1 0 79832 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_65
timestamp 1704896540
transform 1 0 79832 0 1 13061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_66
timestamp 1704896540
transform 1 0 79968 0 1 14421
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_67
timestamp 1704896540
transform 1 0 79968 0 1 11837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_68
timestamp 1704896540
transform 1 0 79832 0 1 13197
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_69
timestamp 1704896540
transform 1 0 79832 0 1 15917
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_70
timestamp 1704896540
transform 1 0 79968 0 1 17277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_71
timestamp 1704896540
transform 1 0 79968 0 1 17413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_72
timestamp 1704896540
transform 1 0 79968 0 1 20133
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_73
timestamp 1704896540
transform 1 0 79832 0 1 20269
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_74
timestamp 1704896540
transform 1 0 79832 0 1 20541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_75
timestamp 1704896540
transform 1 0 79832 0 1 18637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_76
timestamp 1704896540
transform 1 0 89760 0 1 22173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_77
timestamp 1704896540
transform 1 0 89760 0 1 20541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_78
timestamp 1704896540
transform 1 0 89760 0 1 18773
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_79
timestamp 1704896540
transform 1 0 89760 0 1 17141
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_80
timestamp 1704896540
transform 1 0 57392 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_81
timestamp 1704896540
transform 1 0 57392 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_82
timestamp 1704896540
transform 1 0 62424 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_83
timestamp 1704896540
transform 1 0 62424 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_84
timestamp 1704896540
transform 1 0 59296 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_85
timestamp 1704896540
transform 1 0 59296 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_86
timestamp 1704896540
transform 1 0 60792 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_87
timestamp 1704896540
transform 1 0 60792 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_88
timestamp 1704896540
transform 1 0 65280 0 1 10477
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_89
timestamp 1704896540
transform 1 0 67592 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_90
timestamp 1704896540
transform 1 0 65280 0 1 10885
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_91
timestamp 1704896540
transform 1 0 67592 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_92
timestamp 1704896540
transform 1 0 65416 0 1 9389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_93
timestamp 1704896540
transform 1 0 60792 0 1 10885
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_94
timestamp 1704896540
transform 1 0 64328 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_95
timestamp 1704896540
transform 1 0 64328 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_96
timestamp 1704896540
transform 1 0 65824 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_97
timestamp 1704896540
transform 1 0 65824 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_98
timestamp 1704896540
transform 1 0 54128 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_99
timestamp 1704896540
transform 1 0 54128 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_100
timestamp 1704896540
transform 1 0 52360 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_101
timestamp 1704896540
transform 1 0 52360 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_102
timestamp 1704896540
transform 1 0 50864 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_103
timestamp 1704896540
transform 1 0 50864 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_104
timestamp 1704896540
transform 1 0 50728 0 1 10885
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_105
timestamp 1704896540
transform 1 0 49096 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_106
timestamp 1704896540
transform 1 0 49096 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_107
timestamp 1704896540
transform 1 0 47328 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_108
timestamp 1704896540
transform 1 0 47328 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_109
timestamp 1704896540
transform 1 0 45832 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_110
timestamp 1704896540
transform 1 0 45832 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_111
timestamp 1704896540
transform 1 0 45696 0 1 10885
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_112
timestamp 1704896540
transform 1 0 55760 0 1 10885
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_113
timestamp 1704896540
transform 1 0 55896 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_114
timestamp 1704896540
transform 1 0 55896 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_115
timestamp 1704896540
transform 1 0 54128 0 1 19589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_116
timestamp 1704896540
transform 1 0 54128 0 1 19045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_117
timestamp 1704896540
transform 1 0 53176 0 1 19589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_118
timestamp 1704896540
transform 1 0 53176 0 1 19045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_119
timestamp 1704896540
transform 1 0 51000 0 1 13197
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_120
timestamp 1704896540
transform 1 0 51952 0 1 19589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_121
timestamp 1704896540
transform 1 0 51952 0 1 19045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_122
timestamp 1704896540
transform 1 0 50728 0 1 12789
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_123
timestamp 1704896540
transform 1 0 51408 0 1 18909
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_124
timestamp 1704896540
transform 1 0 51408 0 1 14285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_125
timestamp 1704896540
transform 1 0 50728 0 1 13469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_126
timestamp 1704896540
transform 1 0 50728 0 1 14149
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_127
timestamp 1704896540
transform 1 0 50864 0 1 13333
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_128
timestamp 1704896540
transform 1 0 50864 0 1 11837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_129
timestamp 1704896540
transform 1 0 50728 0 1 11701
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_130
timestamp 1704896540
transform 1 0 50728 0 1 19589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_131
timestamp 1704896540
transform 1 0 50728 0 1 19045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_132
timestamp 1704896540
transform 1 0 50184 0 1 19045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_133
timestamp 1704896540
transform 1 0 50184 0 1 19589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_134
timestamp 1704896540
transform 1 0 49368 0 1 19589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_135
timestamp 1704896540
transform 1 0 49368 0 1 19045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_136
timestamp 1704896540
transform 1 0 47872 0 1 19589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_137
timestamp 1704896540
transform 1 0 47872 0 1 19045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_138
timestamp 1704896540
transform 1 0 46920 0 1 19589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_139
timestamp 1704896540
transform 1 0 46920 0 1 19045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_140
timestamp 1704896540
transform 1 0 45968 0 1 13469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_141
timestamp 1704896540
transform 1 0 45968 0 1 14149
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_142
timestamp 1704896540
transform 1 0 45696 0 1 13333
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_143
timestamp 1704896540
transform 1 0 45696 0 1 11837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_144
timestamp 1704896540
transform 1 0 45696 0 1 11701
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_145
timestamp 1704896540
transform 1 0 45696 0 1 14285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_146
timestamp 1704896540
transform 1 0 45696 0 1 18909
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_147
timestamp 1704896540
transform 1 0 45560 0 1 19045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_148
timestamp 1704896540
transform 1 0 45560 0 1 19589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_149
timestamp 1704896540
transform 1 0 50728 0 1 12381
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_150
timestamp 1704896540
transform 1 0 55488 0 1 12925
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_151
timestamp 1704896540
transform 1 0 50456 0 1 12925
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_152
timestamp 1704896540
transform 1 0 45560 0 1 12925
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_153
timestamp 1704896540
transform 1 0 51000 0 1 11565
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_154
timestamp 1704896540
transform 1 0 51000 0 1 12245
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_155
timestamp 1704896540
transform 1 0 45968 0 1 17413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_156
timestamp 1704896540
transform 1 0 45968 0 1 14965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_157
timestamp 1704896540
transform 1 0 55760 0 1 13469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_158
timestamp 1704896540
transform 1 0 55760 0 1 14149
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_159
timestamp 1704896540
transform 1 0 45832 0 1 14965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_160
timestamp 1704896540
transform 1 0 45832 0 1 13197
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_161
timestamp 1704896540
transform 1 0 45832 0 1 12925
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_162
timestamp 1704896540
transform 1 0 45832 0 1 12381
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_163
timestamp 1704896540
transform 1 0 45832 0 1 11565
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_164
timestamp 1704896540
transform 1 0 45832 0 1 12245
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_165
timestamp 1704896540
transform 1 0 55896 0 1 13333
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_166
timestamp 1704896540
transform 1 0 55896 0 1 11837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_167
timestamp 1704896540
transform 1 0 55760 0 1 11701
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_168
timestamp 1704896540
transform 1 0 55760 0 1 14285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_169
timestamp 1704896540
transform 1 0 55760 0 1 18909
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_170
timestamp 1704896540
transform 1 0 55760 0 1 19589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_171
timestamp 1704896540
transform 1 0 55760 0 1 19045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_172
timestamp 1704896540
transform 1 0 56168 0 1 17413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_173
timestamp 1704896540
transform 1 0 56168 0 1 14965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_174
timestamp 1704896540
transform 1 0 56032 0 1 14965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_175
timestamp 1704896540
transform 1 0 56032 0 1 13197
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_176
timestamp 1704896540
transform 1 0 55760 0 1 12789
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_177
timestamp 1704896540
transform 1 0 55760 0 1 12381
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_178
timestamp 1704896540
transform 1 0 56032 0 1 11565
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_179
timestamp 1704896540
transform 1 0 56032 0 1 12245
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_180
timestamp 1704896540
transform 1 0 51136 0 1 17413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_181
timestamp 1704896540
transform 1 0 51136 0 1 14965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_182
timestamp 1704896540
transform 1 0 51000 0 1 14965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_183
timestamp 1704896540
transform 1 0 56984 0 1 19589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_184
timestamp 1704896540
transform 1 0 56984 0 1 19045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_185
timestamp 1704896540
transform 1 0 60520 0 1 12925
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_186
timestamp 1704896540
transform 1 0 66368 0 1 21629
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_187
timestamp 1704896540
transform 1 0 66368 0 1 21901
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_188
timestamp 1704896540
transform 1 0 66504 0 1 21493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_189
timestamp 1704896540
transform 1 0 66504 0 1 21221
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_190
timestamp 1704896540
transform 1 0 66504 0 1 20813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_191
timestamp 1704896540
transform 1 0 66504 0 1 21085
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_192
timestamp 1704896540
transform 1 0 66368 0 1 20133
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_193
timestamp 1704896540
transform 1 0 66368 0 1 17549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_194
timestamp 1704896540
transform 1 0 60928 0 1 17413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_195
timestamp 1704896540
transform 1 0 60928 0 1 14965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_196
timestamp 1704896540
transform 1 0 61064 0 1 14965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_197
timestamp 1704896540
transform 1 0 61064 0 1 13197
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_198
timestamp 1704896540
transform 1 0 65416 0 1 11429
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_199
timestamp 1704896540
transform 1 0 60792 0 1 12789
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_200
timestamp 1704896540
transform 1 0 60792 0 1 12381
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_201
timestamp 1704896540
transform 1 0 60656 0 1 11565
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_202
timestamp 1704896540
transform 1 0 60656 0 1 12245
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_203
timestamp 1704896540
transform 1 0 65688 0 1 19589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_204
timestamp 1704896540
transform 1 0 65688 0 1 19045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_205
timestamp 1704896540
transform 1 0 63920 0 1 19045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_206
timestamp 1704896540
transform 1 0 63920 0 1 19589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_207
timestamp 1704896540
transform 1 0 62832 0 1 19589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_208
timestamp 1704896540
transform 1 0 62832 0 1 19045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_209
timestamp 1704896540
transform 1 0 61880 0 1 19589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_210
timestamp 1704896540
transform 1 0 61880 0 1 19045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_211
timestamp 1704896540
transform 1 0 61472 0 1 18909
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_212
timestamp 1704896540
transform 1 0 61472 0 1 14285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_213
timestamp 1704896540
transform 1 0 60792 0 1 13469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_214
timestamp 1704896540
transform 1 0 60792 0 1 14149
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_215
timestamp 1704896540
transform 1 0 60928 0 1 13333
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_216
timestamp 1704896540
transform 1 0 60928 0 1 11837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_217
timestamp 1704896540
transform 1 0 60792 0 1 11701
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_218
timestamp 1704896540
transform 1 0 60656 0 1 19589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_219
timestamp 1704896540
transform 1 0 60656 0 1 19045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_220
timestamp 1704896540
transform 1 0 60112 0 1 19045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_221
timestamp 1704896540
transform 1 0 60112 0 1 19589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_222
timestamp 1704896540
transform 1 0 59432 0 1 19589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_223
timestamp 1704896540
transform 1 0 59432 0 1 19045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_224
timestamp 1704896540
transform 1 0 58888 0 1 19045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_225
timestamp 1704896540
transform 1 0 58888 0 1 19589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_226
timestamp 1704896540
transform 1 0 58208 0 1 19589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_227
timestamp 1704896540
transform 1 0 58208 0 1 19045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_228
timestamp 1704896540
transform 1 0 66368 0 1 25573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_229
timestamp 1704896540
transform 1 0 66368 0 1 29925
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_230
timestamp 1704896540
transform 1 0 66368 0 1 25029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_231
timestamp 1704896540
transform 1 0 66368 0 1 24757
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_232
timestamp 1704896540
transform 1 0 66368 0 1 30197
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_233
timestamp 1704896540
transform 1 0 66504 0 1 38085
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_234
timestamp 1704896540
transform 1 0 66368 0 1 41621
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_235
timestamp 1704896540
transform 1 0 66368 0 1 41349
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_236
timestamp 1704896540
transform 1 0 66504 0 1 37677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_237
timestamp 1704896540
transform 1 0 66504 0 1 29517
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_238
timestamp 1704896540
transform 1 0 66504 0 1 29789
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_239
timestamp 1704896540
transform 1 0 66368 0 1 36589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_240
timestamp 1704896540
transform 1 0 66368 0 1 36861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_241
timestamp 1704896540
transform 1 0 66504 0 1 42165
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_242
timestamp 1704896540
transform 1 0 66504 0 1 42437
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_243
timestamp 1704896540
transform 1 0 66368 0 1 25845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_244
timestamp 1704896540
transform 1 0 66368 0 1 33733
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_245
timestamp 1704896540
transform 1 0 66368 0 1 33461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_246
timestamp 1704896540
transform 1 0 66504 0 1 33869
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_247
timestamp 1704896540
transform 1 0 66504 0 1 34141
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_248
timestamp 1704896540
transform 1 0 66368 0 1 32917
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_249
timestamp 1704896540
transform 1 0 66504 0 1 38765
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_250
timestamp 1704896540
transform 1 0 66504 0 1 38493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_251
timestamp 1704896540
transform 1 0 66368 0 1 32645
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_252
timestamp 1704896540
transform 1 0 66368 0 1 37813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_253
timestamp 1704896540
transform 1 0 66368 0 1 38085
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_254
timestamp 1704896540
transform 1 0 66504 0 1 28973
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_255
timestamp 1704896540
transform 1 0 66504 0 1 28701
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_256
timestamp 1704896540
transform 1 0 66368 0 1 39309
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_257
timestamp 1704896540
transform 1 0 66368 0 1 39037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_258
timestamp 1704896540
transform 1 0 66368 0 1 41893
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_259
timestamp 1704896540
transform 1 0 66368 0 1 42165
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_260
timestamp 1704896540
transform 1 0 89760 0 1 25573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_261
timestamp 1704896540
transform 1 0 89760 0 1 23805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_262
timestamp 1704896540
transform 1 0 89760 0 1 27341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_263
timestamp 1704896540
transform 1 0 89760 0 1 30605
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_264
timestamp 1704896540
transform 1 0 89760 0 1 28973
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_265
timestamp 1704896540
transform 1 0 89760 0 1 32373
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_266
timestamp 1704896540
transform 1 0 74800 0 1 27613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_267
timestamp 1704896540
transform 1 0 74664 0 1 23805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_268
timestamp 1704896540
transform 1 0 74664 0 1 23669
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_269
timestamp 1704896540
transform 1 0 74664 0 1 22989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_270
timestamp 1704896540
transform 1 0 75072 0 1 23805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_271
timestamp 1704896540
transform 1 0 75072 0 1 24077
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_272
timestamp 1704896540
transform 1 0 74664 0 1 25301
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_273
timestamp 1704896540
transform 1 0 77384 0 1 25437
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_274
timestamp 1704896540
transform 1 0 77384 0 1 25845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_275
timestamp 1704896540
transform 1 0 74664 0 1 25437
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_276
timestamp 1704896540
transform 1 0 76024 0 1 26797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_277
timestamp 1704896540
transform 1 0 76432 0 1 26933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_278
timestamp 1704896540
transform 1 0 76432 0 1 27613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_279
timestamp 1704896540
transform 1 0 76432 0 1 25437
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_280
timestamp 1704896540
transform 1 0 76432 0 1 25981
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_281
timestamp 1704896540
transform 1 0 76296 0 1 26797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_282
timestamp 1704896540
transform 1 0 76296 0 1 26253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_283
timestamp 1704896540
transform 1 0 76296 0 1 25301
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_284
timestamp 1704896540
transform 1 0 76296 0 1 23805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_285
timestamp 1704896540
transform 1 0 76024 0 1 23669
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_286
timestamp 1704896540
transform 1 0 76024 0 1 22989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_287
timestamp 1704896540
transform 1 0 76296 0 1 25981
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_288
timestamp 1704896540
transform 1 0 76296 0 1 25573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_289
timestamp 1704896540
transform 1 0 75072 0 1 22853
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_290
timestamp 1704896540
transform 1 0 75072 0 1 25437
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_291
timestamp 1704896540
transform 1 0 75072 0 1 25981
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_292
timestamp 1704896540
transform 1 0 75208 0 1 26117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_293
timestamp 1704896540
transform 1 0 75208 0 1 26797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_294
timestamp 1704896540
transform 1 0 75208 0 1 26933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_295
timestamp 1704896540
transform 1 0 75208 0 1 27613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_296
timestamp 1704896540
transform 1 0 74664 0 1 26117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_297
timestamp 1704896540
transform 1 0 74664 0 1 26389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_298
timestamp 1704896540
transform 1 0 74664 0 1 25981
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_299
timestamp 1704896540
transform 1 0 76024 0 1 26253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_300
timestamp 1704896540
transform 1 0 75752 0 1 25437
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_301
timestamp 1704896540
transform 1 0 75752 0 1 25981
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_302
timestamp 1704896540
transform 1 0 75480 0 1 23669
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_303
timestamp 1704896540
transform 1 0 75480 0 1 22989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_304
timestamp 1704896540
transform 1 0 75480 0 1 22853
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_305
timestamp 1704896540
transform 1 0 74800 0 1 26933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_306
timestamp 1704896540
transform 1 0 71264 0 1 27749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_307
timestamp 1704896540
transform 1 0 71264 0 1 27341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_308
timestamp 1704896540
transform 1 0 71264 0 1 27613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_309
timestamp 1704896540
transform 1 0 71264 0 1 26797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_310
timestamp 1704896540
transform 1 0 71672 0 1 22989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_311
timestamp 1704896540
transform 1 0 71400 0 1 24077
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_312
timestamp 1704896540
transform 1 0 71400 0 1 23805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_313
timestamp 1704896540
transform 1 0 71264 0 1 23669
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_314
timestamp 1704896540
transform 1 0 71400 0 1 24621
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_315
timestamp 1704896540
transform 1 0 71400 0 1 24893
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_316
timestamp 1704896540
transform 1 0 72080 0 1 23261
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_317
timestamp 1704896540
transform 1 0 72080 0 1 22989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_318
timestamp 1704896540
transform 1 0 72080 0 1 22581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_319
timestamp 1704896540
transform 1 0 72080 0 1 22853
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_320
timestamp 1704896540
transform 1 0 72216 0 1 25029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_321
timestamp 1704896540
transform 1 0 72216 0 1 25301
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_322
timestamp 1704896540
transform 1 0 71672 0 1 23805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_323
timestamp 1704896540
transform 1 0 71808 0 1 26797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_324
timestamp 1704896540
transform 1 0 71808 0 1 26525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_325
timestamp 1704896540
transform 1 0 71264 0 1 23397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_326
timestamp 1704896540
transform 1 0 71264 0 1 22989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_327
timestamp 1704896540
transform 1 0 72896 0 1 22581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_328
timestamp 1704896540
transform 1 0 71672 0 1 23261
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_329
timestamp 1704896540
transform 1 0 71672 0 1 24077
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_330
timestamp 1704896540
transform 1 0 71400 0 1 25301
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_331
timestamp 1704896540
transform 1 0 71400 0 1 25029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_332
timestamp 1704896540
transform 1 0 72624 0 1 27341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_333
timestamp 1704896540
transform 1 0 72624 0 1 27613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_334
timestamp 1704896540
transform 1 0 72216 0 1 25981
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_335
timestamp 1704896540
transform 1 0 73032 0 1 26253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_336
timestamp 1704896540
transform 1 0 73032 0 1 26525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_337
timestamp 1704896540
transform 1 0 72216 0 1 25709
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_338
timestamp 1704896540
transform 1 0 72488 0 1 22853
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_339
timestamp 1704896540
transform 1 0 71672 0 1 26933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_340
timestamp 1704896540
transform 1 0 71672 0 1 27205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_341
timestamp 1704896540
transform 1 0 71808 0 1 22853
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_342
timestamp 1704896540
transform 1 0 71808 0 1 22581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_343
timestamp 1704896540
transform 1 0 71264 0 1 24213
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_344
timestamp 1704896540
transform 1 0 71264 0 1 24485
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_345
timestamp 1704896540
transform 1 0 73032 0 1 23669
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_346
timestamp 1704896540
transform 1 0 73032 0 1 23397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_347
timestamp 1704896540
transform 1 0 72896 0 1 23261
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_348
timestamp 1704896540
transform 1 0 72896 0 1 22989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_349
timestamp 1704896540
transform 1 0 72896 0 1 25301
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_350
timestamp 1704896540
transform 1 0 72080 0 1 23805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_351
timestamp 1704896540
transform 1 0 72896 0 1 25029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_352
timestamp 1704896540
transform 1 0 72488 0 1 22581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_353
timestamp 1704896540
transform 1 0 73032 0 1 25437
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_354
timestamp 1704896540
transform 1 0 73032 0 1 25709
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_355
timestamp 1704896540
transform 1 0 72080 0 1 24077
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_356
timestamp 1704896540
transform 1 0 71672 0 1 27749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_357
timestamp 1704896540
transform 1 0 71672 0 1 27341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_358
timestamp 1704896540
transform 1 0 71672 0 1 27613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_359
timestamp 1704896540
transform 1 0 71264 0 1 23261
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_360
timestamp 1704896540
transform 1 0 72216 0 1 27749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_361
timestamp 1704896540
transform 1 0 72624 0 1 24213
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_362
timestamp 1704896540
transform 1 0 71672 0 1 26389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_363
timestamp 1704896540
transform 1 0 71672 0 1 26117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_364
timestamp 1704896540
transform 1 0 72624 0 1 24485
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_365
timestamp 1704896540
transform 1 0 72896 0 1 27749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_366
timestamp 1704896540
transform 1 0 71672 0 1 23669
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_367
timestamp 1704896540
transform 1 0 72080 0 1 23397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_368
timestamp 1704896540
transform 1 0 72080 0 1 23669
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_369
timestamp 1704896540
transform 1 0 71672 0 1 23397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_370
timestamp 1704896540
transform 1 0 71672 0 1 24213
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_371
timestamp 1704896540
transform 1 0 72896 0 1 23805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_372
timestamp 1704896540
transform 1 0 72896 0 1 24077
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_373
timestamp 1704896540
transform 1 0 72488 0 1 24077
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_374
timestamp 1704896540
transform 1 0 72488 0 1 23805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_375
timestamp 1704896540
transform 1 0 72352 0 1 26525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_376
timestamp 1704896540
transform 1 0 72352 0 1 26797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_377
timestamp 1704896540
transform 1 0 72488 0 1 27205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_378
timestamp 1704896540
transform 1 0 72488 0 1 26933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_379
timestamp 1704896540
transform 1 0 71264 0 1 26117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_380
timestamp 1704896540
transform 1 0 71264 0 1 26389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_381
timestamp 1704896540
transform 1 0 71672 0 1 24485
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_382
timestamp 1704896540
transform 1 0 71672 0 1 24893
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_383
timestamp 1704896540
transform 1 0 71672 0 1 24621
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_384
timestamp 1704896540
transform 1 0 71400 0 1 27205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_385
timestamp 1704896540
transform 1 0 71400 0 1 26933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_386
timestamp 1704896540
transform 1 0 71264 0 1 26525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_387
timestamp 1704896540
transform 1 0 71672 0 1 25301
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_388
timestamp 1704896540
transform 1 0 71672 0 1 25029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_389
timestamp 1704896540
transform 1 0 72216 0 1 24893
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_390
timestamp 1704896540
transform 1 0 72216 0 1 24621
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_391
timestamp 1704896540
transform 1 0 73032 0 1 24213
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_392
timestamp 1704896540
transform 1 0 71400 0 1 22853
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_393
timestamp 1704896540
transform 1 0 71400 0 1 22581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_394
timestamp 1704896540
transform 1 0 73032 0 1 24485
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_395
timestamp 1704896540
transform 1 0 73032 0 1 24893
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_396
timestamp 1704896540
transform 1 0 73032 0 1 24621
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_397
timestamp 1704896540
transform 1 0 72896 0 1 27205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_398
timestamp 1704896540
transform 1 0 72896 0 1 26933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_399
timestamp 1704896540
transform 1 0 71808 0 1 30469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_400
timestamp 1704896540
transform 1 0 72216 0 1 29789
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_401
timestamp 1704896540
transform 1 0 72216 0 1 30061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_402
timestamp 1704896540
transform 1 0 71808 0 1 30741
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_403
timestamp 1704896540
transform 1 0 71808 0 1 31149
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_404
timestamp 1704896540
transform 1 0 71808 0 1 30877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_405
timestamp 1704896540
transform 1 0 71808 0 1 33325
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_406
timestamp 1704896540
transform 1 0 72488 0 1 28157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_407
timestamp 1704896540
transform 1 0 71672 0 1 28157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_408
timestamp 1704896540
transform 1 0 71672 0 1 28429
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_409
timestamp 1704896540
transform 1 0 71808 0 1 28837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_410
timestamp 1704896540
transform 1 0 71808 0 1 28565
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_411
timestamp 1704896540
transform 1 0 71400 0 1 28973
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_412
timestamp 1704896540
transform 1 0 71400 0 1 29245
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_413
timestamp 1704896540
transform 1 0 71672 0 1 32509
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_414
timestamp 1704896540
transform 1 0 71672 0 1 32781
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_415
timestamp 1704896540
transform 1 0 73032 0 1 29245
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_416
timestamp 1704896540
transform 1 0 73032 0 1 28973
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_417
timestamp 1704896540
transform 1 0 71808 0 1 33189
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_418
timestamp 1704896540
transform 1 0 71808 0 1 32917
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_419
timestamp 1704896540
transform 1 0 71672 0 1 31285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_420
timestamp 1704896540
transform 1 0 71672 0 1 31557
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_421
timestamp 1704896540
transform 1 0 72080 0 1 30741
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_422
timestamp 1704896540
transform 1 0 72080 0 1 30469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_423
timestamp 1704896540
transform 1 0 72624 0 1 29789
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_424
timestamp 1704896540
transform 1 0 72080 0 1 31285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_425
timestamp 1704896540
transform 1 0 73032 0 1 29381
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_426
timestamp 1704896540
transform 1 0 73032 0 1 29653
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_427
timestamp 1704896540
transform 1 0 72080 0 1 31557
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_428
timestamp 1704896540
transform 1 0 72624 0 1 30061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_429
timestamp 1704896540
transform 1 0 72624 0 1 32373
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_430
timestamp 1704896540
transform 1 0 72624 0 1 32101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_431
timestamp 1704896540
transform 1 0 72488 0 1 31965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_432
timestamp 1704896540
transform 1 0 72488 0 1 31693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_433
timestamp 1704896540
transform 1 0 72216 0 1 28021
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_434
timestamp 1704896540
transform 1 0 72896 0 1 28021
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_435
timestamp 1704896540
transform 1 0 71400 0 1 31965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_436
timestamp 1704896540
transform 1 0 71400 0 1 31693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_437
timestamp 1704896540
transform 1 0 71400 0 1 30741
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_438
timestamp 1704896540
transform 1 0 71400 0 1 30469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_439
timestamp 1704896540
transform 1 0 73032 0 1 28837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_440
timestamp 1704896540
transform 1 0 73032 0 1 28565
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_441
timestamp 1704896540
transform 1 0 72896 0 1 28157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_442
timestamp 1704896540
transform 1 0 72896 0 1 28429
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_443
timestamp 1704896540
transform 1 0 71808 0 1 32373
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_444
timestamp 1704896540
transform 1 0 71808 0 1 32101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_445
timestamp 1704896540
transform 1 0 71672 0 1 31693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_446
timestamp 1704896540
transform 1 0 71672 0 1 31965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_447
timestamp 1704896540
transform 1 0 72896 0 1 33325
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_448
timestamp 1704896540
transform 1 0 72624 0 1 32917
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_449
timestamp 1704896540
transform 1 0 71400 0 1 32781
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_450
timestamp 1704896540
transform 1 0 71400 0 1 32509
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_451
timestamp 1704896540
transform 1 0 71400 0 1 32101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_452
timestamp 1704896540
transform 1 0 71400 0 1 32373
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_453
timestamp 1704896540
transform 1 0 72624 0 1 33189
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_454
timestamp 1704896540
transform 1 0 72080 0 1 28157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_455
timestamp 1704896540
transform 1 0 72080 0 1 28429
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_456
timestamp 1704896540
transform 1 0 72896 0 1 30469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_457
timestamp 1704896540
transform 1 0 72896 0 1 30197
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_458
timestamp 1704896540
transform 1 0 73032 0 1 29789
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_459
timestamp 1704896540
transform 1 0 73032 0 1 30061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_460
timestamp 1704896540
transform 1 0 72080 0 1 32101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_461
timestamp 1704896540
transform 1 0 72896 0 1 32509
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_462
timestamp 1704896540
transform 1 0 72896 0 1 32781
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_463
timestamp 1704896540
transform 1 0 73032 0 1 33189
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_464
timestamp 1704896540
transform 1 0 73032 0 1 32917
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_465
timestamp 1704896540
transform 1 0 71400 0 1 33325
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_466
timestamp 1704896540
transform 1 0 71264 0 1 30877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_467
timestamp 1704896540
transform 1 0 71400 0 1 28157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_468
timestamp 1704896540
transform 1 0 71400 0 1 28429
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_469
timestamp 1704896540
transform 1 0 71264 0 1 31149
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_470
timestamp 1704896540
transform 1 0 71400 0 1 31557
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_471
timestamp 1704896540
transform 1 0 71400 0 1 31285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_472
timestamp 1704896540
transform 1 0 72080 0 1 32373
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_473
timestamp 1704896540
transform 1 0 72352 0 1 32509
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_474
timestamp 1704896540
transform 1 0 72352 0 1 32781
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_475
timestamp 1704896540
transform 1 0 71264 0 1 28837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_476
timestamp 1704896540
transform 1 0 71264 0 1 28565
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_477
timestamp 1704896540
transform 1 0 71264 0 1 33189
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_478
timestamp 1704896540
transform 1 0 71264 0 1 32917
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_479
timestamp 1704896540
transform 1 0 72352 0 1 33461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_480
timestamp 1704896540
transform 1 0 72352 0 1 33189
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_481
timestamp 1704896540
transform 1 0 73032 0 1 32373
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_482
timestamp 1704896540
transform 1 0 73032 0 1 32101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_483
timestamp 1704896540
transform 1 0 73032 0 1 31693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_484
timestamp 1704896540
transform 1 0 73032 0 1 31965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_485
timestamp 1704896540
transform 1 0 71672 0 1 28021
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_486
timestamp 1704896540
transform 1 0 71808 0 1 28973
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_487
timestamp 1704896540
transform 1 0 71808 0 1 29245
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_488
timestamp 1704896540
transform 1 0 72488 0 1 28837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_489
timestamp 1704896540
transform 1 0 72488 0 1 28565
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_490
timestamp 1704896540
transform 1 0 72488 0 1 28429
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_491
timestamp 1704896540
transform 1 0 71264 0 1 28021
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_492
timestamp 1704896540
transform 1 0 72080 0 1 36453
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_493
timestamp 1704896540
transform 1 0 72080 0 1 36725
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_494
timestamp 1704896540
transform 1 0 71400 0 1 37133
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_495
timestamp 1704896540
transform 1 0 72488 0 1 36317
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_496
timestamp 1704896540
transform 1 0 71400 0 1 33597
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_497
timestamp 1704896540
transform 1 0 71264 0 1 37541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_498
timestamp 1704896540
transform 1 0 71264 0 1 37269
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_499
timestamp 1704896540
transform 1 0 71672 0 1 37269
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_500
timestamp 1704896540
transform 1 0 72216 0 1 38629
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_501
timestamp 1704896540
transform 1 0 72216 0 1 38357
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_502
timestamp 1704896540
transform 1 0 72080 0 1 37677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_503
timestamp 1704896540
transform 1 0 72080 0 1 37949
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_504
timestamp 1704896540
transform 1 0 72352 0 1 35501
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_505
timestamp 1704896540
transform 1 0 72352 0 1 35229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_506
timestamp 1704896540
transform 1 0 72216 0 1 35501
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_507
timestamp 1704896540
transform 1 0 73032 0 1 36725
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_508
timestamp 1704896540
transform 1 0 73032 0 1 36453
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_509
timestamp 1704896540
transform 1 0 73032 0 1 34413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_510
timestamp 1704896540
transform 1 0 73032 0 1 34141
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_511
timestamp 1704896540
transform 1 0 72216 0 1 35229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_512
timestamp 1704896540
transform 1 0 72488 0 1 36045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_513
timestamp 1704896540
transform 1 0 72488 0 1 36861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_514
timestamp 1704896540
transform 1 0 71672 0 1 34685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_515
timestamp 1704896540
transform 1 0 71672 0 1 34413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_516
timestamp 1704896540
transform 1 0 71264 0 1 34685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_517
timestamp 1704896540
transform 1 0 71264 0 1 34413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_518
timestamp 1704896540
transform 1 0 71264 0 1 36045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_519
timestamp 1704896540
transform 1 0 71264 0 1 36317
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_520
timestamp 1704896540
transform 1 0 71264 0 1 38765
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_521
timestamp 1704896540
transform 1 0 71808 0 1 33597
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_522
timestamp 1704896540
transform 1 0 72352 0 1 36453
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_523
timestamp 1704896540
transform 1 0 71808 0 1 38765
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_524
timestamp 1704896540
transform 1 0 71264 0 1 36725
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_525
timestamp 1704896540
transform 1 0 71264 0 1 36453
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_526
timestamp 1704896540
transform 1 0 72896 0 1 36317
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_527
timestamp 1704896540
transform 1 0 72896 0 1 36045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_528
timestamp 1704896540
transform 1 0 71400 0 1 35909
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_529
timestamp 1704896540
transform 1 0 71400 0 1 35637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_530
timestamp 1704896540
transform 1 0 71264 0 1 35229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_531
timestamp 1704896540
transform 1 0 71264 0 1 35501
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_532
timestamp 1704896540
transform 1 0 72488 0 1 37133
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_533
timestamp 1704896540
transform 1 0 72896 0 1 35637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_534
timestamp 1704896540
transform 1 0 72080 0 1 35637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_535
timestamp 1704896540
transform 1 0 72896 0 1 35909
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_536
timestamp 1704896540
transform 1 0 71672 0 1 37541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_537
timestamp 1704896540
transform 1 0 72624 0 1 34005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_538
timestamp 1704896540
transform 1 0 72624 0 1 33733
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_539
timestamp 1704896540
transform 1 0 72896 0 1 36861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_540
timestamp 1704896540
transform 1 0 72896 0 1 37133
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_541
timestamp 1704896540
transform 1 0 73032 0 1 37541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_542
timestamp 1704896540
transform 1 0 73032 0 1 37269
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_543
timestamp 1704896540
transform 1 0 72896 0 1 37677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_544
timestamp 1704896540
transform 1 0 72896 0 1 37949
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_545
timestamp 1704896540
transform 1 0 72896 0 1 38357
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_546
timestamp 1704896540
transform 1 0 72896 0 1 38085
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_547
timestamp 1704896540
transform 1 0 72352 0 1 36725
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_548
timestamp 1704896540
transform 1 0 71264 0 1 34821
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_549
timestamp 1704896540
transform 1 0 72896 0 1 34005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_550
timestamp 1704896540
transform 1 0 72896 0 1 33733
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_551
timestamp 1704896540
transform 1 0 72896 0 1 33597
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_552
timestamp 1704896540
transform 1 0 71264 0 1 35093
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_553
timestamp 1704896540
transform 1 0 71808 0 1 35501
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_554
timestamp 1704896540
transform 1 0 71808 0 1 35229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_555
timestamp 1704896540
transform 1 0 71808 0 1 34821
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_556
timestamp 1704896540
transform 1 0 71808 0 1 35093
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_557
timestamp 1704896540
transform 1 0 71672 0 1 36725
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_558
timestamp 1704896540
transform 1 0 71672 0 1 36453
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_559
timestamp 1704896540
transform 1 0 71672 0 1 35637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_560
timestamp 1704896540
transform 1 0 71672 0 1 35909
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_561
timestamp 1704896540
transform 1 0 71672 0 1 36317
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_562
timestamp 1704896540
transform 1 0 71672 0 1 36045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_563
timestamp 1704896540
transform 1 0 72080 0 1 35909
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_564
timestamp 1704896540
transform 1 0 72352 0 1 35909
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_565
timestamp 1704896540
transform 1 0 72352 0 1 35637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_566
timestamp 1704896540
transform 1 0 72216 0 1 34685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_567
timestamp 1704896540
transform 1 0 71672 0 1 36861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_568
timestamp 1704896540
transform 1 0 71672 0 1 37133
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_569
timestamp 1704896540
transform 1 0 72216 0 1 34413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_570
timestamp 1704896540
transform 1 0 71400 0 1 36861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_571
timestamp 1704896540
transform 1 0 72488 0 1 40397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_572
timestamp 1704896540
transform 1 0 72352 0 1 43389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_573
timestamp 1704896540
transform 1 0 72352 0 1 43117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_574
timestamp 1704896540
transform 1 0 72216 0 1 43389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_575
timestamp 1704896540
transform 1 0 72216 0 1 43117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_576
timestamp 1704896540
transform 1 0 72080 0 1 42573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_577
timestamp 1704896540
transform 1 0 72080 0 1 42301
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_578
timestamp 1704896540
transform 1 0 72896 0 1 40805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_579
timestamp 1704896540
transform 1 0 72896 0 1 41077
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_580
timestamp 1704896540
transform 1 0 72080 0 1 39989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_581
timestamp 1704896540
transform 1 0 72080 0 1 40261
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_582
timestamp 1704896540
transform 1 0 71264 0 1 39173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_583
timestamp 1704896540
transform 1 0 71264 0 1 39445
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_584
timestamp 1704896540
transform 1 0 73032 0 1 39853
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_585
timestamp 1704896540
transform 1 0 73032 0 1 39581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_586
timestamp 1704896540
transform 1 0 72624 0 1 43525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_587
timestamp 1704896540
transform 1 0 72624 0 1 43797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_588
timestamp 1704896540
transform 1 0 72352 0 1 44341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_589
timestamp 1704896540
transform 1 0 71672 0 1 43933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_590
timestamp 1704896540
transform 1 0 71672 0 1 44205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_591
timestamp 1704896540
transform 1 0 71808 0 1 44341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_592
timestamp 1704896540
transform 1 0 72896 0 1 44341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_593
timestamp 1704896540
transform 1 0 71808 0 1 42981
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_594
timestamp 1704896540
transform 1 0 71808 0 1 42709
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_595
timestamp 1704896540
transform 1 0 72080 0 1 44341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_596
timestamp 1704896540
transform 1 0 73032 0 1 41893
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_597
timestamp 1704896540
transform 1 0 73032 0 1 41621
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_598
timestamp 1704896540
transform 1 0 72896 0 1 41213
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_599
timestamp 1704896540
transform 1 0 72896 0 1 41485
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_600
timestamp 1704896540
transform 1 0 72352 0 1 40261
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_601
timestamp 1704896540
transform 1 0 72352 0 1 39989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_602
timestamp 1704896540
transform 1 0 72896 0 1 40669
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_603
timestamp 1704896540
transform 1 0 72896 0 1 40397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_604
timestamp 1704896540
transform 1 0 72896 0 1 39989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_605
timestamp 1704896540
transform 1 0 72896 0 1 40261
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_606
timestamp 1704896540
transform 1 0 73032 0 1 43525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_607
timestamp 1704896540
transform 1 0 73032 0 1 43797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_608
timestamp 1704896540
transform 1 0 71400 0 1 43117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_609
timestamp 1704896540
transform 1 0 71400 0 1 43389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_610
timestamp 1704896540
transform 1 0 71264 0 1 43525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_611
timestamp 1704896540
transform 1 0 71264 0 1 43797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_612
timestamp 1704896540
transform 1 0 72352 0 1 39581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_613
timestamp 1704896540
transform 1 0 72352 0 1 39853
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_614
timestamp 1704896540
transform 1 0 72216 0 1 39581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_615
timestamp 1704896540
transform 1 0 72216 0 1 39853
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_616
timestamp 1704896540
transform 1 0 72080 0 1 39445
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_617
timestamp 1704896540
transform 1 0 72080 0 1 39173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_618
timestamp 1704896540
transform 1 0 71808 0 1 41485
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_619
timestamp 1704896540
transform 1 0 71808 0 1 41213
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_620
timestamp 1704896540
transform 1 0 71808 0 1 40805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_621
timestamp 1704896540
transform 1 0 71808 0 1 41077
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_622
timestamp 1704896540
transform 1 0 71672 0 1 41621
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_623
timestamp 1704896540
transform 1 0 71672 0 1 41893
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_624
timestamp 1704896540
transform 1 0 72896 0 1 42029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_625
timestamp 1704896540
transform 1 0 72896 0 1 42301
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_626
timestamp 1704896540
transform 1 0 71400 0 1 44341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_627
timestamp 1704896540
transform 1 0 71264 0 1 43933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_628
timestamp 1704896540
transform 1 0 71264 0 1 44205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_629
timestamp 1704896540
transform 1 0 71400 0 1 41485
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_630
timestamp 1704896540
transform 1 0 71400 0 1 41213
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_631
timestamp 1704896540
transform 1 0 71400 0 1 40805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_632
timestamp 1704896540
transform 1 0 73032 0 1 42845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_633
timestamp 1704896540
transform 1 0 73032 0 1 43117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_634
timestamp 1704896540
transform 1 0 71400 0 1 41077
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_635
timestamp 1704896540
transform 1 0 71264 0 1 39581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_636
timestamp 1704896540
transform 1 0 71264 0 1 39853
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_637
timestamp 1704896540
transform 1 0 71264 0 1 42981
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_638
timestamp 1704896540
transform 1 0 71264 0 1 42709
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_639
timestamp 1704896540
transform 1 0 71400 0 1 40669
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_640
timestamp 1704896540
transform 1 0 71400 0 1 40397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_641
timestamp 1704896540
transform 1 0 71400 0 1 39989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_642
timestamp 1704896540
transform 1 0 71400 0 1 40261
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_643
timestamp 1704896540
transform 1 0 71672 0 1 40397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_644
timestamp 1704896540
transform 1 0 72216 0 1 44205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_645
timestamp 1704896540
transform 1 0 71672 0 1 39989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_646
timestamp 1704896540
transform 1 0 71672 0 1 40261
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_647
timestamp 1704896540
transform 1 0 71264 0 1 41621
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_648
timestamp 1704896540
transform 1 0 71264 0 1 41893
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_649
timestamp 1704896540
transform 1 0 72216 0 1 43933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_650
timestamp 1704896540
transform 1 0 71808 0 1 39853
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_651
timestamp 1704896540
transform 1 0 71808 0 1 39581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_652
timestamp 1704896540
transform 1 0 72080 0 1 40805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_653
timestamp 1704896540
transform 1 0 71672 0 1 40669
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_654
timestamp 1704896540
transform 1 0 71808 0 1 39445
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_655
timestamp 1704896540
transform 1 0 71808 0 1 39173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_656
timestamp 1704896540
transform 1 0 72080 0 1 41077
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_657
timestamp 1704896540
transform 1 0 72624 0 1 41621
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_658
timestamp 1704896540
transform 1 0 72624 0 1 41893
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_659
timestamp 1704896540
transform 1 0 72488 0 1 40669
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_660
timestamp 1704896540
transform 1 0 71808 0 1 43117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_661
timestamp 1704896540
transform 1 0 71808 0 1 43389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_662
timestamp 1704896540
transform 1 0 71672 0 1 43797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_663
timestamp 1704896540
transform 1 0 71672 0 1 43525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_664
timestamp 1704896540
transform 1 0 71264 0 1 39037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_665
timestamp 1704896540
transform 1 0 71808 0 1 39037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_666
timestamp 1704896540
transform 1 0 89760 0 1 35637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_667
timestamp 1704896540
transform 1 0 89760 0 1 37269
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_668
timestamp 1704896540
transform 1 0 89760 0 1 34005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_669
timestamp 1704896540
transform 1 0 89760 0 1 39173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_670
timestamp 1704896540
transform 1 0 89760 0 1 42301
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_671
timestamp 1704896540
transform 1 0 89760 0 1 40805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_672
timestamp 1704896540
transform 1 0 89760 0 1 43933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_673
timestamp 1704896540
transform 1 0 71672 0 1 22445
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_674
timestamp 1704896540
transform 1 0 71264 0 1 22445
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_675
timestamp 1704896540
transform 1 0 42296 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_676
timestamp 1704896540
transform 1 0 42296 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_677
timestamp 1704896540
transform 1 0 38896 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_678
timestamp 1704896540
transform 1 0 38896 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_679
timestamp 1704896540
transform 1 0 43928 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_680
timestamp 1704896540
transform 1 0 40800 0 1 10885
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_681
timestamp 1704896540
transform 1 0 43928 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_682
timestamp 1704896540
transform 1 0 40800 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_683
timestamp 1704896540
transform 1 0 40800 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_684
timestamp 1704896540
transform 1 0 37400 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_685
timestamp 1704896540
transform 1 0 37400 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_686
timestamp 1704896540
transform 1 0 35632 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_687
timestamp 1704896540
transform 1 0 35632 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_688
timestamp 1704896540
transform 1 0 35768 0 1 10885
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_689
timestamp 1704896540
transform 1 0 30736 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_690
timestamp 1704896540
transform 1 0 30736 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_691
timestamp 1704896540
transform 1 0 28832 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_692
timestamp 1704896540
transform 1 0 28832 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_693
timestamp 1704896540
transform 1 0 32368 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_694
timestamp 1704896540
transform 1 0 32368 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_695
timestamp 1704896540
transform 1 0 33864 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_696
timestamp 1704896540
transform 1 0 33864 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_697
timestamp 1704896540
transform 1 0 25160 0 1 3677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_698
timestamp 1704896540
transform 1 0 25568 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_699
timestamp 1704896540
transform 1 0 25568 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_700
timestamp 1704896540
transform 1 0 27336 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_701
timestamp 1704896540
transform 1 0 25160 0 1 1773
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_702
timestamp 1704896540
transform 1 0 27336 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_703
timestamp 1704896540
transform 1 0 25704 0 1 2861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_704
timestamp 1704896540
transform 1 0 24752 0 1 2861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_705
timestamp 1704896540
transform 1 0 23392 0 1 2861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_706
timestamp 1704896540
transform 1 0 23800 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_707
timestamp 1704896540
transform 1 0 23800 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_708
timestamp 1704896540
transform 1 0 25568 0 1 10885
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_709
timestamp 1704896540
transform 1 0 25568 0 1 10477
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_710
timestamp 1704896540
transform 1 0 25160 0 1 11157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_711
timestamp 1704896540
transform 1 0 25160 0 1 9389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_712
timestamp 1704896540
transform 1 0 25704 0 1 10885
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_713
timestamp 1704896540
transform 1 0 30872 0 1 10885
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_714
timestamp 1704896540
transform 1 0 25976 0 1 14965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_715
timestamp 1704896540
transform 1 0 31960 0 1 19045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_716
timestamp 1704896540
transform 1 0 26112 0 1 14965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_717
timestamp 1704896540
transform 1 0 26112 0 1 13197
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_718
timestamp 1704896540
transform 1 0 25840 0 1 12789
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_719
timestamp 1704896540
transform 1 0 25840 0 1 12381
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_720
timestamp 1704896540
transform 1 0 25840 0 1 11565
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_721
timestamp 1704896540
transform 1 0 25840 0 1 12245
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_722
timestamp 1704896540
transform 1 0 25976 0 1 11837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_723
timestamp 1704896540
transform 1 0 31008 0 1 12925
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_724
timestamp 1704896540
transform 1 0 31552 0 1 19045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_725
timestamp 1704896540
transform 1 0 31552 0 1 19589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_726
timestamp 1704896540
transform 1 0 30736 0 1 13469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_727
timestamp 1704896540
transform 1 0 30736 0 1 14149
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_728
timestamp 1704896540
transform 1 0 31008 0 1 12381
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_729
timestamp 1704896540
transform 1 0 24480 0 1 21629
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_730
timestamp 1704896540
transform 1 0 24480 0 1 21221
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_731
timestamp 1704896540
transform 1 0 30736 0 1 11565
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_732
timestamp 1704896540
transform 1 0 30736 0 1 12245
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_733
timestamp 1704896540
transform 1 0 30464 0 1 12925
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_734
timestamp 1704896540
transform 1 0 25296 0 1 12925
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_735
timestamp 1704896540
transform 1 0 24344 0 1 21901
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_736
timestamp 1704896540
transform 1 0 24344 0 1 21629
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_737
timestamp 1704896540
transform 1 0 24616 0 1 21221
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_738
timestamp 1704896540
transform 1 0 24616 0 1 21493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_739
timestamp 1704896540
transform 1 0 31960 0 1 19589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_740
timestamp 1704896540
transform 1 0 25976 0 1 17413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_741
timestamp 1704896540
transform 1 0 30872 0 1 13333
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_742
timestamp 1704896540
transform 1 0 30872 0 1 11837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_743
timestamp 1704896540
transform 1 0 30872 0 1 11701
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_744
timestamp 1704896540
transform 1 0 30736 0 1 14285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_745
timestamp 1704896540
transform 1 0 30736 0 1 18909
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_746
timestamp 1704896540
transform 1 0 31144 0 1 17413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_747
timestamp 1704896540
transform 1 0 31144 0 1 14965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_748
timestamp 1704896540
transform 1 0 31008 0 1 14965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_749
timestamp 1704896540
transform 1 0 25296 0 1 19045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_750
timestamp 1704896540
transform 1 0 25296 0 1 19589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_751
timestamp 1704896540
transform 1 0 26520 0 1 19045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_752
timestamp 1704896540
transform 1 0 26520 0 1 19589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_753
timestamp 1704896540
transform 1 0 30328 0 1 19589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_754
timestamp 1704896540
transform 1 0 30328 0 1 19045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_755
timestamp 1704896540
transform 1 0 31008 0 1 13197
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_756
timestamp 1704896540
transform 1 0 25704 0 1 11701
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_757
timestamp 1704896540
transform 1 0 29648 0 1 19045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_758
timestamp 1704896540
transform 1 0 29648 0 1 19589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_759
timestamp 1704896540
transform 1 0 26792 0 1 18909
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_760
timestamp 1704896540
transform 1 0 26792 0 1 14285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_761
timestamp 1704896540
transform 1 0 29512 0 1 19589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_762
timestamp 1704896540
transform 1 0 29512 0 1 19045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_763
timestamp 1704896540
transform 1 0 28152 0 1 19589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_764
timestamp 1704896540
transform 1 0 28152 0 1 19045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_765
timestamp 1704896540
transform 1 0 33184 0 1 19589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_766
timestamp 1704896540
transform 1 0 33184 0 1 19045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_767
timestamp 1704896540
transform 1 0 32640 0 1 19045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_768
timestamp 1704896540
transform 1 0 32640 0 1 19589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_769
timestamp 1704896540
transform 1 0 25976 0 1 13469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_770
timestamp 1704896540
transform 1 0 25976 0 1 14149
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_771
timestamp 1704896540
transform 1 0 25976 0 1 13333
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_772
timestamp 1704896540
transform 1 0 44472 0 1 19589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_773
timestamp 1704896540
transform 1 0 44472 0 1 19045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_774
timestamp 1704896540
transform 1 0 43928 0 1 19045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_775
timestamp 1704896540
transform 1 0 43928 0 1 19589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_776
timestamp 1704896540
transform 1 0 40528 0 1 12925
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_777
timestamp 1704896540
transform 1 0 35496 0 1 12925
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_778
timestamp 1704896540
transform 1 0 42704 0 1 19045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_779
timestamp 1704896540
transform 1 0 42704 0 1 19589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_780
timestamp 1704896540
transform 1 0 41480 0 1 19045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_781
timestamp 1704896540
transform 1 0 41480 0 1 19589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_782
timestamp 1704896540
transform 1 0 41480 0 1 18909
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_783
timestamp 1704896540
transform 1 0 41480 0 1 14285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_784
timestamp 1704896540
transform 1 0 40936 0 1 13469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_785
timestamp 1704896540
transform 1 0 40936 0 1 14149
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_786
timestamp 1704896540
transform 1 0 40936 0 1 13333
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_787
timestamp 1704896540
transform 1 0 40936 0 1 11837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_788
timestamp 1704896540
transform 1 0 40800 0 1 11701
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_789
timestamp 1704896540
transform 1 0 40800 0 1 19589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_790
timestamp 1704896540
transform 1 0 40800 0 1 19045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_791
timestamp 1704896540
transform 1 0 38352 0 1 19045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_792
timestamp 1704896540
transform 1 0 38352 0 1 19589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_793
timestamp 1704896540
transform 1 0 36448 0 1 19045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_794
timestamp 1704896540
transform 1 0 36448 0 1 19589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_795
timestamp 1704896540
transform 1 0 36448 0 1 18909
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_796
timestamp 1704896540
transform 1 0 36448 0 1 14285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_797
timestamp 1704896540
transform 1 0 35768 0 1 13469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_798
timestamp 1704896540
transform 1 0 35768 0 1 14149
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_799
timestamp 1704896540
transform 1 0 35904 0 1 13333
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_800
timestamp 1704896540
transform 1 0 35904 0 1 11837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_801
timestamp 1704896540
transform 1 0 35768 0 1 11701
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_802
timestamp 1704896540
transform 1 0 35768 0 1 19589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_803
timestamp 1704896540
transform 1 0 35768 0 1 19045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_804
timestamp 1704896540
transform 1 0 35224 0 1 19045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_805
timestamp 1704896540
transform 1 0 35224 0 1 19589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_806
timestamp 1704896540
transform 1 0 34544 0 1 19589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_807
timestamp 1704896540
transform 1 0 34544 0 1 19045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_808
timestamp 1704896540
transform 1 0 40936 0 1 17413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_809
timestamp 1704896540
transform 1 0 40936 0 1 14965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_810
timestamp 1704896540
transform 1 0 41072 0 1 14965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_811
timestamp 1704896540
transform 1 0 41072 0 1 13197
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_812
timestamp 1704896540
transform 1 0 40800 0 1 12789
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_813
timestamp 1704896540
transform 1 0 40800 0 1 12381
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_814
timestamp 1704896540
transform 1 0 41072 0 1 11565
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_815
timestamp 1704896540
transform 1 0 41072 0 1 12245
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_816
timestamp 1704896540
transform 1 0 36176 0 1 17413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_817
timestamp 1704896540
transform 1 0 36176 0 1 14965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_818
timestamp 1704896540
transform 1 0 36040 0 1 14965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_819
timestamp 1704896540
transform 1 0 36040 0 1 13197
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_820
timestamp 1704896540
transform 1 0 35768 0 1 12789
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_821
timestamp 1704896540
transform 1 0 35768 0 1 12381
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_822
timestamp 1704896540
transform 1 0 35632 0 1 11565
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_823
timestamp 1704896540
transform 1 0 35632 0 1 12245
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_824
timestamp 1704896540
transform 1 0 19992 0 1 2861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_825
timestamp 1704896540
transform 1 0 18904 0 1 2861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_826
timestamp 1704896540
transform 1 0 17680 0 1 2861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_827
timestamp 1704896540
transform 1 0 22304 0 1 2861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_828
timestamp 1704896540
transform 1 0 20400 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_829
timestamp 1704896540
transform 1 0 18768 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_830
timestamp 1704896540
transform 1 0 18768 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_831
timestamp 1704896540
transform 1 0 21080 0 1 2861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_832
timestamp 1704896540
transform 1 0 20400 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_833
timestamp 1704896540
transform 1 0 22168 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_834
timestamp 1704896540
transform 1 0 22168 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_835
timestamp 1704896540
transform 1 0 13872 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_836
timestamp 1704896540
transform 1 0 13872 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_837
timestamp 1704896540
transform 1 0 12104 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_838
timestamp 1704896540
transform 1 0 13328 0 1 549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_839
timestamp 1704896540
transform 1 0 12104 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_840
timestamp 1704896540
transform 1 0 13328 0 1 2317
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_841
timestamp 1704896540
transform 1 0 12920 0 1 2861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_842
timestamp 1704896540
transform 1 0 15368 0 1 2861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_843
timestamp 1704896540
transform 1 0 14280 0 1 2861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_844
timestamp 1704896540
transform 1 0 16456 0 1 3949
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_845
timestamp 1704896540
transform 1 0 15504 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_846
timestamp 1704896540
transform 1 0 15504 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_847
timestamp 1704896540
transform 1 0 16456 0 1 2861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_848
timestamp 1704896540
transform 1 0 17136 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_849
timestamp 1704896540
transform 1 0 17136 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_850
timestamp 1704896540
transform 1 0 16592 0 1 6397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_851
timestamp 1704896540
transform 1 0 11696 0 1 10885
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_852
timestamp 1704896540
transform 1 0 16456 0 1 7621
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_853
timestamp 1704896540
transform 1 0 11696 0 1 10749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_854
timestamp 1704896540
transform 1 0 16456 0 1 10477
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_855
timestamp 1704896540
transform 1 0 11696 0 1 8029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_856
timestamp 1704896540
transform 1 0 16592 0 1 9117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_857
timestamp 1704896540
transform 1 0 16456 0 1 7757
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_858
timestamp 1704896540
transform 1 0 16592 0 1 9253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_859
timestamp 1704896540
transform 1 0 17952 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_860
timestamp 1704896540
transform 1 0 10336 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_861
timestamp 1704896540
transform 1 0 8840 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_862
timestamp 1704896540
transform 1 0 7072 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_863
timestamp 1704896540
transform 1 0 7072 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_864
timestamp 1704896540
transform 1 0 8840 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_865
timestamp 1704896540
transform 1 0 10336 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_866
timestamp 1704896540
transform 1 0 1904 0 1 1773
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_867
timestamp 1704896540
transform 1 0 1904 0 1 2045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_868
timestamp 1704896540
transform 1 0 1224 0 1 3677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_869
timestamp 1704896540
transform 1 0 1224 0 1 5309
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_870
timestamp 1704896540
transform 1 0 5304 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_871
timestamp 1704896540
transform 1 0 5304 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_872
timestamp 1704896540
transform 1 0 3672 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_873
timestamp 1704896540
transform 1 0 3672 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_874
timestamp 1704896540
transform 1 0 1904 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_875
timestamp 1704896540
transform 1 0 1904 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_876
timestamp 1704896540
transform 1 0 544 0 1 10885
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_877
timestamp 1704896540
transform 1 0 544 0 1 7893
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_878
timestamp 1704896540
transform 1 0 1224 0 1 7077
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_879
timestamp 1704896540
transform 1 0 2856 0 1 8301
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_880
timestamp 1704896540
transform 1 0 2856 0 1 8573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_881
timestamp 1704896540
transform 1 0 1224 0 1 10477
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_882
timestamp 1704896540
transform 1 0 1224 0 1 8845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_883
timestamp 1704896540
transform 1 0 2448 0 1 9253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_884
timestamp 1704896540
transform 1 0 2448 0 1 8845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_885
timestamp 1704896540
transform 1 0 11424 0 1 13741
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_886
timestamp 1704896540
transform 1 0 11424 0 1 16325
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_887
timestamp 1704896540
transform 1 0 2448 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_888
timestamp 1704896540
transform 1 0 1224 0 1 15645
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_889
timestamp 1704896540
transform 1 0 1224 0 1 12245
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_890
timestamp 1704896540
transform 1 0 544 0 1 15101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_891
timestamp 1704896540
transform 1 0 1224 0 1 13741
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_892
timestamp 1704896540
transform 1 0 1224 0 1 17141
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_893
timestamp 1704896540
transform 1 0 2448 0 1 17141
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_894
timestamp 1704896540
transform 1 0 1224 0 1 22173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_895
timestamp 1704896540
transform 1 0 1224 0 1 18773
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_896
timestamp 1704896540
transform 1 0 3128 0 1 19181
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_897
timestamp 1704896540
transform 1 0 3128 0 1 18909
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_898
timestamp 1704896540
transform 1 0 1224 0 1 20405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_899
timestamp 1704896540
transform 1 0 2455 0 1 18260
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_900
timestamp 1704896540
transform 1 0 3944 0 1 20541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_901
timestamp 1704896540
transform 1 0 544 0 1 20813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_902
timestamp 1704896540
transform 1 0 3672 0 1 20813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_903
timestamp 1704896540
transform 1 0 3944 0 1 17957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_904
timestamp 1704896540
transform 1 0 19584 0 1 20677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_905
timestamp 1704896540
transform 1 0 19584 0 1 20949
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_906
timestamp 1704896540
transform 1 0 17816 0 1 21493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_907
timestamp 1704896540
transform 1 0 19448 0 1 22173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_908
timestamp 1704896540
transform 1 0 17816 0 1 21765
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_909
timestamp 1704896540
transform 1 0 17952 0 1 20677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_910
timestamp 1704896540
transform 1 0 17952 0 1 20949
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_911
timestamp 1704896540
transform 1 0 17952 0 1 21357
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_912
timestamp 1704896540
transform 1 0 17952 0 1 21085
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_913
timestamp 1704896540
transform 1 0 18768 0 1 22037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_914
timestamp 1704896540
transform 1 0 18768 0 1 21765
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_915
timestamp 1704896540
transform 1 0 17952 0 1 22309
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_916
timestamp 1704896540
transform 1 0 18904 0 1 21085
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_917
timestamp 1704896540
transform 1 0 18904 0 1 21357
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_918
timestamp 1704896540
transform 1 0 16592 0 1 17549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_919
timestamp 1704896540
transform 1 0 16592 0 1 14829
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_920
timestamp 1704896540
transform 1 0 16592 0 1 11837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_921
timestamp 1704896540
transform 1 0 16592 0 1 14693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_922
timestamp 1704896540
transform 1 0 16592 0 1 12109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_923
timestamp 1704896540
transform 1 0 15776 0 1 20677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_924
timestamp 1704896540
transform 1 0 15776 0 1 21221
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_925
timestamp 1704896540
transform 1 0 15096 0 1 21493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_926
timestamp 1704896540
transform 1 0 11696 0 1 13469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_927
timestamp 1704896540
transform 1 0 13600 0 1 20541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_928
timestamp 1704896540
transform 1 0 13600 0 1 19317
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_929
timestamp 1704896540
transform 1 0 19040 0 1 20677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_930
timestamp 1704896540
transform 1 0 19040 0 1 20949
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_931
timestamp 1704896540
transform 1 0 18360 0 1 22037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_932
timestamp 1704896540
transform 1 0 18360 0 1 21765
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_933
timestamp 1704896540
transform 1 0 18496 0 1 20813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_934
timestamp 1704896540
transform 1 0 18496 0 1 20541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_935
timestamp 1704896540
transform 1 0 19040 0 1 22173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_936
timestamp 1704896540
transform 1 0 19176 0 1 19861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_937
timestamp 1704896540
transform 1 0 19176 0 1 16325
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_938
timestamp 1704896540
transform 1 0 17952 0 1 13333
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_939
timestamp 1704896540
transform 1 0 16456 0 1 16189
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_940
timestamp 1704896540
transform 1 0 16456 0 1 13469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_941
timestamp 1704896540
transform 1 0 16184 0 1 20677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_942
timestamp 1704896540
transform 1 0 16184 0 1 21221
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_943
timestamp 1704896540
transform 1 0 15232 0 1 21493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_944
timestamp 1704896540
transform 1 0 19448 0 1 20133
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_945
timestamp 1704896540
transform 1 0 19040 0 1 20541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_946
timestamp 1704896540
transform 1 0 14008 0 1 20541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_947
timestamp 1704896540
transform 1 0 14008 0 1 17957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_948
timestamp 1704896540
transform 1 0 11696 0 1 15101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_949
timestamp 1704896540
transform 1 0 11696 0 1 17821
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_950
timestamp 1704896540
transform 1 0 19040 0 1 17685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_951
timestamp 1704896540
transform 1 0 19448 0 1 20541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_952
timestamp 1704896540
transform 1 0 11560 0 1 19181
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_953
timestamp 1704896540
transform 1 0 11560 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_954
timestamp 1704896540
transform 1 0 11560 0 1 14965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_955
timestamp 1704896540
transform 1 0 11560 0 1 12245
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_956
timestamp 1704896540
transform 1 0 11560 0 1 12109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_957
timestamp 1704896540
transform 1 0 11560 0 1 9389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_958
timestamp 1704896540
transform 1 0 17952 0 1 25709
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_959
timestamp 1704896540
transform 1 0 17952 0 1 25437
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_960
timestamp 1704896540
transform 1 0 17952 0 1 24213
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_961
timestamp 1704896540
transform 1 0 19448 0 1 27341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_962
timestamp 1704896540
transform 1 0 17680 0 1 25573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_963
timestamp 1704896540
transform 1 0 17816 0 1 27749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_964
timestamp 1704896540
transform 1 0 18496 0 1 23805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_965
timestamp 1704896540
transform 1 0 18496 0 1 24077
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_966
timestamp 1704896540
transform 1 0 18360 0 1 23805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_967
timestamp 1704896540
transform 1 0 18496 0 1 25301
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_968
timestamp 1704896540
transform 1 0 19584 0 1 27749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_969
timestamp 1704896540
transform 1 0 18496 0 1 25029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_970
timestamp 1704896540
transform 1 0 19584 0 1 22853
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_971
timestamp 1704896540
transform 1 0 19584 0 1 22581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_972
timestamp 1704896540
transform 1 0 19176 0 1 24621
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_973
timestamp 1704896540
transform 1 0 19584 0 1 27205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_974
timestamp 1704896540
transform 1 0 19584 0 1 26933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_975
timestamp 1704896540
transform 1 0 19448 0 1 26525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_976
timestamp 1704896540
transform 1 0 19448 0 1 26797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_977
timestamp 1704896540
transform 1 0 19176 0 1 24893
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_978
timestamp 1704896540
transform 1 0 18360 0 1 24077
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_979
timestamp 1704896540
transform 1 0 19176 0 1 26933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_980
timestamp 1704896540
transform 1 0 19448 0 1 24893
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_981
timestamp 1704896540
transform 1 0 19448 0 1 24621
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_982
timestamp 1704896540
transform 1 0 19176 0 1 27205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_983
timestamp 1704896540
transform 1 0 19176 0 1 23397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_984
timestamp 1704896540
transform 1 0 19176 0 1 23669
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_985
timestamp 1704896540
transform 1 0 19176 0 1 26389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_986
timestamp 1704896540
transform 1 0 18496 0 1 26525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_987
timestamp 1704896540
transform 1 0 18496 0 1 26797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_988
timestamp 1704896540
transform 1 0 19176 0 1 26117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_989
timestamp 1704896540
transform 1 0 18496 0 1 23261
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_990
timestamp 1704896540
transform 1 0 19448 0 1 23805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_991
timestamp 1704896540
transform 1 0 19448 0 1 24077
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_992
timestamp 1704896540
transform 1 0 19584 0 1 24485
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_993
timestamp 1704896540
transform 1 0 19584 0 1 24213
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_994
timestamp 1704896540
transform 1 0 18496 0 1 22989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_995
timestamp 1704896540
transform 1 0 18224 0 1 24485
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_996
timestamp 1704896540
transform 1 0 18224 0 1 24213
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_997
timestamp 1704896540
transform 1 0 17680 0 1 25981
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_998
timestamp 1704896540
transform 1 0 19448 0 1 23669
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_999
timestamp 1704896540
transform 1 0 19448 0 1 23397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1000
timestamp 1704896540
transform 1 0 19584 0 1 22989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1001
timestamp 1704896540
transform 1 0 19584 0 1 23261
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1002
timestamp 1704896540
transform 1 0 19448 0 1 26389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1003
timestamp 1704896540
transform 1 0 19448 0 1 26117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1004
timestamp 1704896540
transform 1 0 18768 0 1 27749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1005
timestamp 1704896540
transform 1 0 17816 0 1 23669
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1006
timestamp 1704896540
transform 1 0 18496 0 1 27613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1007
timestamp 1704896540
transform 1 0 18496 0 1 27341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1008
timestamp 1704896540
transform 1 0 18632 0 1 25709
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1009
timestamp 1704896540
transform 1 0 18632 0 1 25981
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1010
timestamp 1704896540
transform 1 0 17816 0 1 23397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1011
timestamp 1704896540
transform 1 0 19040 0 1 27749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1012
timestamp 1704896540
transform 1 0 19040 0 1 27341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1013
timestamp 1704896540
transform 1 0 19040 0 1 26525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1014
timestamp 1704896540
transform 1 0 19040 0 1 26797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1015
timestamp 1704896540
transform 1 0 19040 0 1 27613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1016
timestamp 1704896540
transform 1 0 19040 0 1 25029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1017
timestamp 1704896540
transform 1 0 19040 0 1 25301
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1018
timestamp 1704896540
transform 1 0 19176 0 1 23805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1019
timestamp 1704896540
transform 1 0 19176 0 1 24077
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1020
timestamp 1704896540
transform 1 0 18768 0 1 24893
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1021
timestamp 1704896540
transform 1 0 18768 0 1 24621
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1022
timestamp 1704896540
transform 1 0 18632 0 1 24213
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1023
timestamp 1704896540
transform 1 0 18632 0 1 24485
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1024
timestamp 1704896540
transform 1 0 17816 0 1 25301
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1025
timestamp 1704896540
transform 1 0 17952 0 1 26253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1026
timestamp 1704896540
transform 1 0 17952 0 1 26525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1027
timestamp 1704896540
transform 1 0 17816 0 1 26933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1028
timestamp 1704896540
transform 1 0 18224 0 1 25029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1029
timestamp 1704896540
transform 1 0 18224 0 1 25301
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1030
timestamp 1704896540
transform 1 0 17816 0 1 27205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1031
timestamp 1704896540
transform 1 0 19448 0 1 27613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1032
timestamp 1704896540
transform 1 0 18768 0 1 27613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1033
timestamp 1704896540
transform 1 0 18768 0 1 27341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1034
timestamp 1704896540
transform 1 0 18904 0 1 26525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1035
timestamp 1704896540
transform 1 0 18904 0 1 26797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1036
timestamp 1704896540
transform 1 0 18632 0 1 27205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1037
timestamp 1704896540
transform 1 0 18632 0 1 26933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1038
timestamp 1704896540
transform 1 0 19176 0 1 22581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1039
timestamp 1704896540
transform 1 0 19176 0 1 22853
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1040
timestamp 1704896540
transform 1 0 19176 0 1 23261
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1041
timestamp 1704896540
transform 1 0 19176 0 1 22989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1042
timestamp 1704896540
transform 1 0 17816 0 1 23805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1043
timestamp 1704896540
transform 1 0 17816 0 1 24077
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1044
timestamp 1704896540
transform 1 0 17816 0 1 22989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1045
timestamp 1704896540
transform 1 0 17816 0 1 23261
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1046
timestamp 1704896540
transform 1 0 17816 0 1 24893
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1047
timestamp 1704896540
transform 1 0 19584 0 1 25029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1048
timestamp 1704896540
transform 1 0 17952 0 1 24485
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1049
timestamp 1704896540
transform 1 0 19040 0 1 24485
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1050
timestamp 1704896540
transform 1 0 19040 0 1 24213
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1051
timestamp 1704896540
transform 1 0 18224 0 1 27749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1052
timestamp 1704896540
transform 1 0 17952 0 1 22581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1053
timestamp 1704896540
transform 1 0 18224 0 1 23669
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1054
timestamp 1704896540
transform 1 0 18224 0 1 23397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1055
timestamp 1704896540
transform 1 0 19584 0 1 25301
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1056
timestamp 1704896540
transform 1 0 17816 0 1 25029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1057
timestamp 1704896540
transform 1 0 17816 0 1 24621
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1058
timestamp 1704896540
transform 1 0 15096 0 1 25437
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1059
timestamp 1704896540
transform 1 0 15776 0 1 27613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1060
timestamp 1704896540
transform 1 0 15776 0 1 26933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1061
timestamp 1704896540
transform 1 0 15096 0 1 25981
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1062
timestamp 1704896540
transform 1 0 15096 0 1 26797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1063
timestamp 1704896540
transform 1 0 15096 0 1 26253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1064
timestamp 1704896540
transform 1 0 15232 0 1 23805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1065
timestamp 1704896540
transform 1 0 14416 0 1 25437
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1066
timestamp 1704896540
transform 1 0 15640 0 1 22853
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1067
timestamp 1704896540
transform 1 0 15232 0 1 25165
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1068
timestamp 1704896540
transform 1 0 15640 0 1 22581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1069
timestamp 1704896540
transform 1 0 15096 0 1 22581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1070
timestamp 1704896540
transform 1 0 12920 0 1 25437
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1071
timestamp 1704896540
transform 1 0 16184 0 1 26117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1072
timestamp 1704896540
transform 1 0 14688 0 1 23805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1073
timestamp 1704896540
transform 1 0 14416 0 1 25981
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1074
timestamp 1704896540
transform 1 0 16048 0 1 25981
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1075
timestamp 1704896540
transform 1 0 14824 0 1 25981
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1076
timestamp 1704896540
transform 1 0 14824 0 1 25573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1077
timestamp 1704896540
transform 1 0 16048 0 1 25437
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1078
timestamp 1704896540
transform 1 0 15640 0 1 26117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1079
timestamp 1704896540
transform 1 0 15912 0 1 26253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1080
timestamp 1704896540
transform 1 0 15912 0 1 25437
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1081
timestamp 1704896540
transform 1 0 15776 0 1 25437
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1082
timestamp 1704896540
transform 1 0 15232 0 1 22853
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1083
timestamp 1704896540
transform 1 0 15232 0 1 22989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1084
timestamp 1704896540
transform 1 0 15776 0 1 25981
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1085
timestamp 1704896540
transform 1 0 14824 0 1 27749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1086
timestamp 1704896540
transform 1 0 15232 0 1 23669
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1087
timestamp 1704896540
transform 1 0 15776 0 1 22989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1088
timestamp 1704896540
transform 1 0 15776 0 1 23669
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1089
timestamp 1704896540
transform 1 0 15640 0 1 26797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1090
timestamp 1704896540
transform 1 0 16184 0 1 22989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1091
timestamp 1704896540
transform 1 0 14688 0 1 25301
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1092
timestamp 1704896540
transform 1 0 14552 0 1 26933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1093
timestamp 1704896540
transform 1 0 14552 0 1 27613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1094
timestamp 1704896540
transform 1 0 14416 0 1 26797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1095
timestamp 1704896540
transform 1 0 16184 0 1 23669
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1096
timestamp 1704896540
transform 1 0 16184 0 1 26797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1097
timestamp 1704896540
transform 1 0 14416 0 1 26253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1098
timestamp 1704896540
transform 1 0 15368 0 1 26933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1099
timestamp 1704896540
transform 1 0 15368 0 1 27613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1100
timestamp 1704896540
transform 1 0 12920 0 1 28021
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1101
timestamp 1704896540
transform 1 0 14824 0 1 29381
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1102
timestamp 1704896540
transform 1 0 19176 0 1 28157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1103
timestamp 1704896540
transform 1 0 17816 0 1 28157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1104
timestamp 1704896540
transform 1 0 19584 0 1 33325
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1105
timestamp 1704896540
transform 1 0 17816 0 1 28429
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1106
timestamp 1704896540
transform 1 0 19584 0 1 28429
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1107
timestamp 1704896540
transform 1 0 19584 0 1 28157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1108
timestamp 1704896540
transform 1 0 19584 0 1 28021
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1109
timestamp 1704896540
transform 1 0 19448 0 1 28973
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1110
timestamp 1704896540
transform 1 0 19448 0 1 29245
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1111
timestamp 1704896540
transform 1 0 19584 0 1 33189
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1112
timestamp 1704896540
transform 1 0 19584 0 1 32917
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1113
timestamp 1704896540
transform 1 0 19448 0 1 32509
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1114
timestamp 1704896540
transform 1 0 19448 0 1 32781
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1115
timestamp 1704896540
transform 1 0 19448 0 1 31965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1116
timestamp 1704896540
transform 1 0 19448 0 1 31693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1117
timestamp 1704896540
transform 1 0 19448 0 1 31285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1118
timestamp 1704896540
transform 1 0 19448 0 1 31557
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1119
timestamp 1704896540
transform 1 0 17816 0 1 29789
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1120
timestamp 1704896540
transform 1 0 17816 0 1 30061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1121
timestamp 1704896540
transform 1 0 18768 0 1 28021
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1122
timestamp 1704896540
transform 1 0 18632 0 1 30061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1123
timestamp 1704896540
transform 1 0 18632 0 1 29789
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1124
timestamp 1704896540
transform 1 0 18632 0 1 33189
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1125
timestamp 1704896540
transform 1 0 18632 0 1 32917
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1126
timestamp 1704896540
transform 1 0 19176 0 1 32781
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1127
timestamp 1704896540
transform 1 0 18768 0 1 29245
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1128
timestamp 1704896540
transform 1 0 18768 0 1 28973
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1129
timestamp 1704896540
transform 1 0 19176 0 1 32509
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1130
timestamp 1704896540
transform 1 0 19176 0 1 32101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1131
timestamp 1704896540
transform 1 0 19176 0 1 32373
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1132
timestamp 1704896540
transform 1 0 18768 0 1 32101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1133
timestamp 1704896540
transform 1 0 18768 0 1 32373
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1134
timestamp 1704896540
transform 1 0 19176 0 1 30741
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1135
timestamp 1704896540
transform 1 0 19176 0 1 30469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1136
timestamp 1704896540
transform 1 0 18496 0 1 33325
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1137
timestamp 1704896540
transform 1 0 18496 0 1 31965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1138
timestamp 1704896540
transform 1 0 18496 0 1 31693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1139
timestamp 1704896540
transform 1 0 19040 0 1 28565
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1140
timestamp 1704896540
transform 1 0 19040 0 1 28837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1141
timestamp 1704896540
transform 1 0 19040 0 1 29245
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1142
timestamp 1704896540
transform 1 0 19040 0 1 28973
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1143
timestamp 1704896540
transform 1 0 19040 0 1 28021
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1144
timestamp 1704896540
transform 1 0 18496 0 1 30741
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1145
timestamp 1704896540
transform 1 0 18496 0 1 30469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1146
timestamp 1704896540
transform 1 0 19176 0 1 31557
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1147
timestamp 1704896540
transform 1 0 19176 0 1 31285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1148
timestamp 1704896540
transform 1 0 19040 0 1 30877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1149
timestamp 1704896540
transform 1 0 19040 0 1 31149
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1150
timestamp 1704896540
transform 1 0 17816 0 1 28565
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1151
timestamp 1704896540
transform 1 0 17816 0 1 28837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1152
timestamp 1704896540
transform 1 0 18360 0 1 32101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1153
timestamp 1704896540
transform 1 0 18360 0 1 32373
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1154
timestamp 1704896540
transform 1 0 18360 0 1 32509
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1155
timestamp 1704896540
transform 1 0 18360 0 1 32781
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1156
timestamp 1704896540
transform 1 0 17816 0 1 29653
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1157
timestamp 1704896540
transform 1 0 17816 0 1 29381
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1158
timestamp 1704896540
transform 1 0 18496 0 1 28837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1159
timestamp 1704896540
transform 1 0 18496 0 1 28565
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1160
timestamp 1704896540
transform 1 0 18224 0 1 28837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1161
timestamp 1704896540
transform 1 0 17816 0 1 28973
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1162
timestamp 1704896540
transform 1 0 19584 0 1 32101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1163
timestamp 1704896540
transform 1 0 18224 0 1 28565
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1164
timestamp 1704896540
transform 1 0 18360 0 1 28157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1165
timestamp 1704896540
transform 1 0 19584 0 1 32373
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1166
timestamp 1704896540
transform 1 0 19584 0 1 28837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1167
timestamp 1704896540
transform 1 0 19584 0 1 28565
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1168
timestamp 1704896540
transform 1 0 17816 0 1 29245
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1169
timestamp 1704896540
transform 1 0 18360 0 1 28429
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1170
timestamp 1704896540
transform 1 0 19176 0 1 33325
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1171
timestamp 1704896540
transform 1 0 17816 0 1 33325
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1172
timestamp 1704896540
transform 1 0 17952 0 1 31693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1173
timestamp 1704896540
transform 1 0 17952 0 1 31965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1174
timestamp 1704896540
transform 1 0 17816 0 1 30197
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1175
timestamp 1704896540
transform 1 0 17816 0 1 30469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1176
timestamp 1704896540
transform 1 0 17816 0 1 28021
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1177
timestamp 1704896540
transform 1 0 18360 0 1 31557
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1178
timestamp 1704896540
transform 1 0 17952 0 1 32101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1179
timestamp 1704896540
transform 1 0 17952 0 1 32373
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1180
timestamp 1704896540
transform 1 0 19448 0 1 30877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1181
timestamp 1704896540
transform 1 0 19448 0 1 31149
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1182
timestamp 1704896540
transform 1 0 19584 0 1 30469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1183
timestamp 1704896540
transform 1 0 18360 0 1 31285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1184
timestamp 1704896540
transform 1 0 17816 0 1 32509
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1185
timestamp 1704896540
transform 1 0 17816 0 1 32781
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1186
timestamp 1704896540
transform 1 0 17952 0 1 33189
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1187
timestamp 1704896540
transform 1 0 17952 0 1 32917
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1188
timestamp 1704896540
transform 1 0 18224 0 1 28021
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1189
timestamp 1704896540
transform 1 0 19584 0 1 30741
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1190
timestamp 1704896540
transform 1 0 19040 0 1 31693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1191
timestamp 1704896540
transform 1 0 19040 0 1 31965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1192
timestamp 1704896540
transform 1 0 19040 0 1 32917
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1193
timestamp 1704896540
transform 1 0 19040 0 1 33189
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1194
timestamp 1704896540
transform 1 0 19176 0 1 28429
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1195
timestamp 1704896540
transform 1 0 3672 0 1 23397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1196
timestamp 1704896540
transform 1 0 1224 0 1 25573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1197
timestamp 1704896540
transform 1 0 2176 0 1 25029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1198
timestamp 1704896540
transform 1 0 2176 0 1 25573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1199
timestamp 1704896540
transform 1 0 1224 0 1 27205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1200
timestamp 1704896540
transform 1 0 2455 0 1 25667
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1201
timestamp 1704896540
transform 1 0 1224 0 1 23805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1202
timestamp 1704896540
transform 1 0 544 0 1 26253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1203
timestamp 1704896540
transform 1 0 1224 0 1 28837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1204
timestamp 1704896540
transform 1 0 1224 0 1 30741
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1205
timestamp 1704896540
transform 1 0 1224 0 1 32237
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1206
timestamp 1704896540
transform 1 0 11016 0 1 32373
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1207
timestamp 1704896540
transform 1 0 11016 0 1 29517
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1208
timestamp 1704896540
transform 1 0 11016 0 1 32237
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1209
timestamp 1704896540
transform 1 0 11152 0 1 31013
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1210
timestamp 1704896540
transform 1 0 11152 0 1 30877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1211
timestamp 1704896540
transform 1 0 11152 0 1 28157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1212
timestamp 1704896540
transform 1 0 11152 0 1 35229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1213
timestamp 1704896540
transform 1 0 11152 0 1 37949
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1214
timestamp 1704896540
transform 1 0 11016 0 1 35093
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1215
timestamp 1704896540
transform 1 0 11288 0 1 33869
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1216
timestamp 1704896540
transform 1 0 11152 0 1 33597
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1217
timestamp 1704896540
transform 1 0 11288 0 1 36453
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1218
timestamp 1704896540
transform 1 0 1224 0 1 34005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1219
timestamp 1704896540
transform 1 0 1224 0 1 35637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1220
timestamp 1704896540
transform 1 0 1224 0 1 37269
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1221
timestamp 1704896540
transform 1 0 1224 0 1 44205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1222
timestamp 1704896540
transform 1 0 1224 0 1 40669
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1223
timestamp 1704896540
transform 1 0 1224 0 1 42301
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1224
timestamp 1704896540
transform 1 0 1224 0 1 39173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1225
timestamp 1704896540
transform 1 0 17816 0 1 36317
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1226
timestamp 1704896540
transform 1 0 17816 0 1 36045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1227
timestamp 1704896540
transform 1 0 17816 0 1 35637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1228
timestamp 1704896540
transform 1 0 19040 0 1 38765
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1229
timestamp 1704896540
transform 1 0 17816 0 1 35909
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1230
timestamp 1704896540
transform 1 0 17816 0 1 34005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1231
timestamp 1704896540
transform 1 0 19584 0 1 33597
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1232
timestamp 1704896540
transform 1 0 19584 0 1 36453
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1233
timestamp 1704896540
transform 1 0 17816 0 1 33733
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1234
timestamp 1704896540
transform 1 0 19448 0 1 37133
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1235
timestamp 1704896540
transform 1 0 19448 0 1 35637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1236
timestamp 1704896540
transform 1 0 19448 0 1 35909
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1237
timestamp 1704896540
transform 1 0 19448 0 1 36317
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1238
timestamp 1704896540
transform 1 0 18904 0 1 36725
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1239
timestamp 1704896540
transform 1 0 18904 0 1 36453
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1240
timestamp 1704896540
transform 1 0 18904 0 1 35229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1241
timestamp 1704896540
transform 1 0 18904 0 1 35501
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1242
timestamp 1704896540
transform 1 0 19448 0 1 36045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1243
timestamp 1704896540
transform 1 0 19584 0 1 35501
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1244
timestamp 1704896540
transform 1 0 19584 0 1 35229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1245
timestamp 1704896540
transform 1 0 17816 0 1 37133
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1246
timestamp 1704896540
transform 1 0 18904 0 1 35637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1247
timestamp 1704896540
transform 1 0 18904 0 1 35909
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1248
timestamp 1704896540
transform 1 0 17952 0 1 37541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1249
timestamp 1704896540
transform 1 0 19448 0 1 34413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1250
timestamp 1704896540
transform 1 0 19448 0 1 34685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1251
timestamp 1704896540
transform 1 0 19448 0 1 35093
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1252
timestamp 1704896540
transform 1 0 18632 0 1 34005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1253
timestamp 1704896540
transform 1 0 18632 0 1 33733
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1254
timestamp 1704896540
transform 1 0 18904 0 1 38629
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1255
timestamp 1704896540
transform 1 0 18904 0 1 38357
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1256
timestamp 1704896540
transform 1 0 18632 0 1 34413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1257
timestamp 1704896540
transform 1 0 18632 0 1 34685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1258
timestamp 1704896540
transform 1 0 19448 0 1 34821
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1259
timestamp 1704896540
transform 1 0 19040 0 1 36045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1260
timestamp 1704896540
transform 1 0 19040 0 1 36317
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1261
timestamp 1704896540
transform 1 0 19040 0 1 34685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1262
timestamp 1704896540
transform 1 0 18496 0 1 33597
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1263
timestamp 1704896540
transform 1 0 18224 0 1 33733
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1264
timestamp 1704896540
transform 1 0 18224 0 1 34005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1265
timestamp 1704896540
transform 1 0 18496 0 1 35229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1266
timestamp 1704896540
transform 1 0 18496 0 1 35501
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1267
timestamp 1704896540
transform 1 0 19584 0 1 36725
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1268
timestamp 1704896540
transform 1 0 18496 0 1 37677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1269
timestamp 1704896540
transform 1 0 18496 0 1 37949
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1270
timestamp 1704896540
transform 1 0 19040 0 1 34413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1271
timestamp 1704896540
transform 1 0 17816 0 1 33597
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1272
timestamp 1704896540
transform 1 0 19176 0 1 35909
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1273
timestamp 1704896540
transform 1 0 19176 0 1 35637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1274
timestamp 1704896540
transform 1 0 17952 0 1 37269
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1275
timestamp 1704896540
transform 1 0 19448 0 1 38765
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1276
timestamp 1704896540
transform 1 0 19176 0 1 33597
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1277
timestamp 1704896540
transform 1 0 17952 0 1 36453
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1278
timestamp 1704896540
transform 1 0 17952 0 1 36725
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1279
timestamp 1704896540
transform 1 0 18360 0 1 36861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1280
timestamp 1704896540
transform 1 0 18360 0 1 37133
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1281
timestamp 1704896540
transform 1 0 17816 0 1 36861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1282
timestamp 1704896540
transform 1 0 19176 0 1 36453
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1283
timestamp 1704896540
transform 1 0 19176 0 1 36725
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1284
timestamp 1704896540
transform 1 0 19176 0 1 37133
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1285
timestamp 1704896540
transform 1 0 19176 0 1 36861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1286
timestamp 1704896540
transform 1 0 17816 0 1 38357
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1287
timestamp 1704896540
transform 1 0 17816 0 1 38085
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1288
timestamp 1704896540
transform 1 0 17816 0 1 37949
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1289
timestamp 1704896540
transform 1 0 17816 0 1 37677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1290
timestamp 1704896540
transform 1 0 18224 0 1 36725
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1291
timestamp 1704896540
transform 1 0 18224 0 1 36453
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1292
timestamp 1704896540
transform 1 0 17952 0 1 34413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1293
timestamp 1704896540
transform 1 0 17952 0 1 34141
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1294
timestamp 1704896540
transform 1 0 19040 0 1 34821
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1295
timestamp 1704896540
transform 1 0 19040 0 1 35093
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1296
timestamp 1704896540
transform 1 0 19040 0 1 35501
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1297
timestamp 1704896540
transform 1 0 19040 0 1 35229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1298
timestamp 1704896540
transform 1 0 19040 0 1 37269
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1299
timestamp 1704896540
transform 1 0 19584 0 1 37541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1300
timestamp 1704896540
transform 1 0 19040 0 1 37541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1301
timestamp 1704896540
transform 1 0 19584 0 1 37269
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1302
timestamp 1704896540
transform 1 0 19448 0 1 36861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1303
timestamp 1704896540
transform 1 0 19448 0 1 40397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1304
timestamp 1704896540
transform 1 0 19448 0 1 40669
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1305
timestamp 1704896540
transform 1 0 19448 0 1 41077
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1306
timestamp 1704896540
transform 1 0 19448 0 1 40805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1307
timestamp 1704896540
transform 1 0 19448 0 1 41621
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1308
timestamp 1704896540
transform 1 0 19448 0 1 41893
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1309
timestamp 1704896540
transform 1 0 19584 0 1 44341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1310
timestamp 1704896540
transform 1 0 19584 0 1 43525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1311
timestamp 1704896540
transform 1 0 19584 0 1 43797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1312
timestamp 1704896540
transform 1 0 19584 0 1 44205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1313
timestamp 1704896540
transform 1 0 19584 0 1 43933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1314
timestamp 1704896540
transform 1 0 18904 0 1 39581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1315
timestamp 1704896540
transform 1 0 18904 0 1 39853
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1316
timestamp 1704896540
transform 1 0 18632 0 1 40261
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1317
timestamp 1704896540
transform 1 0 18632 0 1 39989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1318
timestamp 1704896540
transform 1 0 18768 0 1 39445
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1319
timestamp 1704896540
transform 1 0 18768 0 1 39173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1320
timestamp 1704896540
transform 1 0 18904 0 1 43389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1321
timestamp 1704896540
transform 1 0 18904 0 1 43117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1322
timestamp 1704896540
transform 1 0 18904 0 1 43933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1323
timestamp 1704896540
transform 1 0 18904 0 1 44205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1324
timestamp 1704896540
transform 1 0 18632 0 1 44341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1325
timestamp 1704896540
transform 1 0 19448 0 1 39445
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1326
timestamp 1704896540
transform 1 0 18360 0 1 42573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1327
timestamp 1704896540
transform 1 0 18360 0 1 42301
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1328
timestamp 1704896540
transform 1 0 19448 0 1 42709
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1329
timestamp 1704896540
transform 1 0 18496 0 1 39445
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1330
timestamp 1704896540
transform 1 0 18496 0 1 39173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1331
timestamp 1704896540
transform 1 0 18360 0 1 39445
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1332
timestamp 1704896540
transform 1 0 18360 0 1 39173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1333
timestamp 1704896540
transform 1 0 18496 0 1 41349
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1334
timestamp 1704896540
transform 1 0 18496 0 1 41077
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1335
timestamp 1704896540
transform 1 0 18224 0 1 39581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1336
timestamp 1704896540
transform 1 0 18224 0 1 39853
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1337
timestamp 1704896540
transform 1 0 18224 0 1 41621
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1338
timestamp 1704896540
transform 1 0 18224 0 1 41893
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1339
timestamp 1704896540
transform 1 0 19448 0 1 42981
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1340
timestamp 1704896540
transform 1 0 19448 0 1 43389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1341
timestamp 1704896540
transform 1 0 19448 0 1 43117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1342
timestamp 1704896540
transform 1 0 18224 0 1 44205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1343
timestamp 1704896540
transform 1 0 18224 0 1 43933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1344
timestamp 1704896540
transform 1 0 18360 0 1 43797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1345
timestamp 1704896540
transform 1 0 18360 0 1 43525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1346
timestamp 1704896540
transform 1 0 18496 0 1 40669
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1347
timestamp 1704896540
transform 1 0 18496 0 1 40397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1348
timestamp 1704896540
transform 1 0 18360 0 1 40669
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1349
timestamp 1704896540
transform 1 0 18360 0 1 40397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1350
timestamp 1704896540
transform 1 0 19584 0 1 41485
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1351
timestamp 1704896540
transform 1 0 19584 0 1 41213
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1352
timestamp 1704896540
transform 1 0 19176 0 1 44341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1353
timestamp 1704896540
transform 1 0 19176 0 1 41893
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1354
timestamp 1704896540
transform 1 0 19176 0 1 41621
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1355
timestamp 1704896540
transform 1 0 19176 0 1 40805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1356
timestamp 1704896540
transform 1 0 19176 0 1 41077
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1357
timestamp 1704896540
transform 1 0 19176 0 1 41485
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1358
timestamp 1704896540
transform 1 0 19176 0 1 41213
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1359
timestamp 1704896540
transform 1 0 19176 0 1 39445
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1360
timestamp 1704896540
transform 1 0 19176 0 1 39173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1361
timestamp 1704896540
transform 1 0 19040 0 1 44205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1362
timestamp 1704896540
transform 1 0 19040 0 1 43933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1363
timestamp 1704896540
transform 1 0 19040 0 1 43525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1364
timestamp 1704896540
transform 1 0 19040 0 1 43797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1365
timestamp 1704896540
transform 1 0 19040 0 1 39581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1366
timestamp 1704896540
transform 1 0 19040 0 1 39853
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1367
timestamp 1704896540
transform 1 0 19448 0 1 39173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1368
timestamp 1704896540
transform 1 0 19040 0 1 43389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1369
timestamp 1704896540
transform 1 0 19040 0 1 43117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1370
timestamp 1704896540
transform 1 0 19040 0 1 42709
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1371
timestamp 1704896540
transform 1 0 19040 0 1 42981
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1372
timestamp 1704896540
transform 1 0 19176 0 1 40669
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1373
timestamp 1704896540
transform 1 0 19176 0 1 40397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1374
timestamp 1704896540
transform 1 0 19176 0 1 39989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1375
timestamp 1704896540
transform 1 0 19176 0 1 40261
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1376
timestamp 1704896540
transform 1 0 17816 0 1 40397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1377
timestamp 1704896540
transform 1 0 17816 0 1 40669
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1378
timestamp 1704896540
transform 1 0 17816 0 1 44341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1379
timestamp 1704896540
transform 1 0 19040 0 1 41213
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1380
timestamp 1704896540
transform 1 0 19040 0 1 41757
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1381
timestamp 1704896540
transform 1 0 17952 0 1 40805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1382
timestamp 1704896540
transform 1 0 17952 0 1 41077
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1383
timestamp 1704896540
transform 1 0 17952 0 1 41485
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1384
timestamp 1704896540
transform 1 0 17952 0 1 41213
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1385
timestamp 1704896540
transform 1 0 17816 0 1 42301
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1386
timestamp 1704896540
transform 1 0 17816 0 1 42029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1387
timestamp 1704896540
transform 1 0 17816 0 1 41621
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1388
timestamp 1704896540
transform 1 0 17816 0 1 41893
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1389
timestamp 1704896540
transform 1 0 17816 0 1 39581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1390
timestamp 1704896540
transform 1 0 17816 0 1 39853
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1391
timestamp 1704896540
transform 1 0 17952 0 1 40261
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1392
timestamp 1704896540
transform 1 0 17952 0 1 39989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1393
timestamp 1704896540
transform 1 0 17952 0 1 43525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1394
timestamp 1704896540
transform 1 0 17952 0 1 43797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1395
timestamp 1704896540
transform 1 0 17816 0 1 43117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1396
timestamp 1704896540
transform 1 0 17816 0 1 42845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1397
timestamp 1704896540
transform 1 0 19584 0 1 40261
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1398
timestamp 1704896540
transform 1 0 19584 0 1 39989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1399
timestamp 1704896540
transform 1 0 19584 0 1 39853
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1400
timestamp 1704896540
transform 1 0 19584 0 1 39581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1401
timestamp 1704896540
transform 1 0 19448 0 1 39037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1402
timestamp 1704896540
transform 1 0 19040 0 1 39037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1403
timestamp 1704896540
transform 1 0 24616 0 1 34549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1404
timestamp 1704896540
transform 1 0 24616 0 1 24757
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1405
timestamp 1704896540
transform 1 0 24616 0 1 25029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1406
timestamp 1704896540
transform 1 0 24616 0 1 37813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1407
timestamp 1704896540
transform 1 0 24616 0 1 38085
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1408
timestamp 1704896540
transform 1 0 24480 0 1 33733
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1409
timestamp 1704896540
transform 1 0 24480 0 1 33461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1410
timestamp 1704896540
transform 1 0 24616 0 1 36589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1411
timestamp 1704896540
transform 1 0 24616 0 1 36861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1412
timestamp 1704896540
transform 1 0 24616 0 1 34141
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1413
timestamp 1704896540
transform 1 0 24616 0 1 33733
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1414
timestamp 1704896540
transform 1 0 24344 0 1 42709
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1415
timestamp 1704896540
transform 1 0 24344 0 1 42437
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1416
timestamp 1704896540
transform 1 0 24480 0 1 30197
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1417
timestamp 1704896540
transform 1 0 24480 0 1 29925
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1418
timestamp 1704896540
transform 1 0 24616 0 1 25573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1419
timestamp 1704896540
transform 1 0 24616 0 1 25845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1420
timestamp 1704896540
transform 1 0 24480 0 1 31421
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1421
timestamp 1704896540
transform 1 0 24480 0 1 31149
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1422
timestamp 1704896540
transform 1 0 24616 0 1 42165
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1423
timestamp 1704896540
transform 1 0 24616 0 1 42437
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1424
timestamp 1704896540
transform 1 0 24344 0 1 39309
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1425
timestamp 1704896540
transform 1 0 24344 0 1 39037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1426
timestamp 1704896540
transform 1 0 24616 0 1 30333
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1427
timestamp 1704896540
transform 1 0 24616 0 1 30605
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1428
timestamp 1704896540
transform 1 0 24616 0 1 34277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1429
timestamp 1704896540
transform 1 0 19448 0 1 22445
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1430
timestamp 1704896540
transform 1 0 19040 0 1 22445
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1431
timestamp 1704896540
transform 1 0 24480 0 1 45837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1432
timestamp 1704896540
transform 1 0 24480 0 1 46109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1433
timestamp 1704896540
transform 1 0 24344 0 1 58621
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1434
timestamp 1704896540
transform 1 0 24480 0 1 63789
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1435
timestamp 1704896540
transform 1 0 24480 0 1 63517
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1436
timestamp 1704896540
transform 1 0 24344 0 1 58349
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1437
timestamp 1704896540
transform 1 0 24344 0 1 62973
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1438
timestamp 1704896540
transform 1 0 24616 0 1 66645
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1439
timestamp 1704896540
transform 1 0 24344 0 1 62701
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1440
timestamp 1704896540
transform 1 0 24480 0 1 46789
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1441
timestamp 1704896540
transform 1 0 24480 0 1 46517
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1442
timestamp 1704896540
transform 1 0 24344 0 1 45565
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1443
timestamp 1704896540
transform 1 0 24344 0 1 45293
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1444
timestamp 1704896540
transform 1 0 24616 0 1 59573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1445
timestamp 1704896540
transform 1 0 24616 0 1 59845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1446
timestamp 1704896540
transform 1 0 24480 0 1 50869
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1447
timestamp 1704896540
transform 1 0 24480 0 1 50461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1448
timestamp 1704896540
transform 1 0 24616 0 1 54677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1449
timestamp 1704896540
transform 1 0 24616 0 1 54405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1450
timestamp 1704896540
transform 1 0 24344 0 1 54269
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1451
timestamp 1704896540
transform 1 0 24344 0 1 53997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1452
timestamp 1704896540
transform 1 0 24616 0 1 63381
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1453
timestamp 1704896540
transform 1 0 24616 0 1 63109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1454
timestamp 1704896540
transform 1 0 24616 0 1 50869
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1455
timestamp 1704896540
transform 1 0 24616 0 1 51141
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1456
timestamp 1704896540
transform 1 0 24616 0 1 65829
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1457
timestamp 1704896540
transform 1 0 24616 0 1 66101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1458
timestamp 1704896540
transform 1 0 19176 0 1 47741
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1459
timestamp 1704896540
transform 1 0 17952 0 1 48965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1460
timestamp 1704896540
transform 1 0 19040 0 1 47061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1461
timestamp 1704896540
transform 1 0 19040 0 1 47333
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1462
timestamp 1704896540
transform 1 0 19176 0 1 49509
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1463
timestamp 1704896540
transform 1 0 17952 0 1 45429
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1464
timestamp 1704896540
transform 1 0 18224 0 1 48557
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1465
timestamp 1704896540
transform 1 0 19176 0 1 49781
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1466
timestamp 1704896540
transform 1 0 18768 0 1 49509
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1467
timestamp 1704896540
transform 1 0 18632 0 1 48693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1468
timestamp 1704896540
transform 1 0 17952 0 1 48693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1469
timestamp 1704896540
transform 1 0 17816 0 1 48285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1470
timestamp 1704896540
transform 1 0 19584 0 1 48557
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1471
timestamp 1704896540
transform 1 0 19584 0 1 48285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1472
timestamp 1704896540
transform 1 0 17816 0 1 48557
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1473
timestamp 1704896540
transform 1 0 18768 0 1 46381
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1474
timestamp 1704896540
transform 1 0 18224 0 1 48285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1475
timestamp 1704896540
transform 1 0 17952 0 1 45837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1476
timestamp 1704896540
transform 1 0 19040 0 1 44749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1477
timestamp 1704896540
transform 1 0 19448 0 1 45021
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1478
timestamp 1704896540
transform 1 0 19176 0 1 45837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1479
timestamp 1704896540
transform 1 0 19176 0 1 45565
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1480
timestamp 1704896540
transform 1 0 19040 0 1 48557
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1481
timestamp 1704896540
transform 1 0 19040 0 1 48285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1482
timestamp 1704896540
transform 1 0 19040 0 1 47877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1483
timestamp 1704896540
transform 1 0 19448 0 1 44749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1484
timestamp 1704896540
transform 1 0 19040 0 1 45021
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1485
timestamp 1704896540
transform 1 0 19448 0 1 48693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1486
timestamp 1704896540
transform 1 0 19448 0 1 45565
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1487
timestamp 1704896540
transform 1 0 19448 0 1 45837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1488
timestamp 1704896540
transform 1 0 19584 0 1 47333
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1489
timestamp 1704896540
transform 1 0 19584 0 1 47061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1490
timestamp 1704896540
transform 1 0 19448 0 1 48965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1491
timestamp 1704896540
transform 1 0 19040 0 1 48149
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1492
timestamp 1704896540
transform 1 0 19584 0 1 49781
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1493
timestamp 1704896540
transform 1 0 19584 0 1 49509
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1494
timestamp 1704896540
transform 1 0 17952 0 1 46245
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1495
timestamp 1704896540
transform 1 0 19176 0 1 49373
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1496
timestamp 1704896540
transform 1 0 19448 0 1 45429
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1497
timestamp 1704896540
transform 1 0 19448 0 1 45157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1498
timestamp 1704896540
transform 1 0 19176 0 1 49101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1499
timestamp 1704896540
transform 1 0 19176 0 1 48693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1500
timestamp 1704896540
transform 1 0 19176 0 1 48965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1501
timestamp 1704896540
transform 1 0 17952 0 1 45973
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1502
timestamp 1704896540
transform 1 0 19448 0 1 49373
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1503
timestamp 1704896540
transform 1 0 18224 0 1 47877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1504
timestamp 1704896540
transform 1 0 18224 0 1 48149
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1505
timestamp 1704896540
transform 1 0 19448 0 1 49101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1506
timestamp 1704896540
transform 1 0 18768 0 1 46653
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1507
timestamp 1704896540
transform 1 0 19040 0 1 45429
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1508
timestamp 1704896540
transform 1 0 18496 0 1 45837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1509
timestamp 1704896540
transform 1 0 18496 0 1 45565
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1510
timestamp 1704896540
transform 1 0 17952 0 1 45565
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1511
timestamp 1704896540
transform 1 0 18768 0 1 49373
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1512
timestamp 1704896540
transform 1 0 19040 0 1 45157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1513
timestamp 1704896540
transform 1 0 18360 0 1 45565
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1514
timestamp 1704896540
transform 1 0 18360 0 1 45021
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1515
timestamp 1704896540
transform 1 0 18360 0 1 44749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1516
timestamp 1704896540
transform 1 0 18360 0 1 45837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1517
timestamp 1704896540
transform 1 0 18224 0 1 49781
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1518
timestamp 1704896540
transform 1 0 19448 0 1 47469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1519
timestamp 1704896540
transform 1 0 19448 0 1 47741
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1520
timestamp 1704896540
transform 1 0 19448 0 1 48149
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1521
timestamp 1704896540
transform 1 0 19448 0 1 47877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1522
timestamp 1704896540
transform 1 0 18224 0 1 49509
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1523
timestamp 1704896540
transform 1 0 18768 0 1 49101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1524
timestamp 1704896540
transform 1 0 18904 0 1 47061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1525
timestamp 1704896540
transform 1 0 17816 0 1 44749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1526
timestamp 1704896540
transform 1 0 17816 0 1 45021
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1527
timestamp 1704896540
transform 1 0 17952 0 1 49509
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1528
timestamp 1704896540
transform 1 0 17952 0 1 49781
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1529
timestamp 1704896540
transform 1 0 17952 0 1 46789
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1530
timestamp 1704896540
transform 1 0 17816 0 1 46653
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1531
timestamp 1704896540
transform 1 0 18496 0 1 46925
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1532
timestamp 1704896540
transform 1 0 17952 0 1 47061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1533
timestamp 1704896540
transform 1 0 17816 0 1 49373
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1534
timestamp 1704896540
transform 1 0 18496 0 1 46653
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1535
timestamp 1704896540
transform 1 0 17816 0 1 46381
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1536
timestamp 1704896540
transform 1 0 18904 0 1 48285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1537
timestamp 1704896540
transform 1 0 18904 0 1 48557
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1538
timestamp 1704896540
transform 1 0 17816 0 1 49101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1539
timestamp 1704896540
transform 1 0 18904 0 1 47333
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1540
timestamp 1704896540
transform 1 0 17952 0 1 49917
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1541
timestamp 1704896540
transform 1 0 19176 0 1 47469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1542
timestamp 1704896540
transform 1 0 18632 0 1 48965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1543
timestamp 1704896540
transform 1 0 17952 0 1 45157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1544
timestamp 1704896540
transform 1 0 18768 0 1 49781
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1545
timestamp 1704896540
transform 1 0 18360 0 1 54541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1546
timestamp 1704896540
transform 1 0 18224 0 1 52637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1547
timestamp 1704896540
transform 1 0 18224 0 1 52909
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1548
timestamp 1704896540
transform 1 0 19176 0 1 51821
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1549
timestamp 1704896540
transform 1 0 19176 0 1 52093
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1550
timestamp 1704896540
transform 1 0 19584 0 1 52229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1551
timestamp 1704896540
transform 1 0 19584 0 1 52501
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1552
timestamp 1704896540
transform 1 0 19176 0 1 53725
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1553
timestamp 1704896540
transform 1 0 19176 0 1 53453
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1554
timestamp 1704896540
transform 1 0 19040 0 1 52229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1555
timestamp 1704896540
transform 1 0 19448 0 1 52637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1556
timestamp 1704896540
transform 1 0 19448 0 1 52909
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1557
timestamp 1704896540
transform 1 0 19040 0 1 52501
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1558
timestamp 1704896540
transform 1 0 17816 0 1 52501
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1559
timestamp 1704896540
transform 1 0 17816 0 1 52637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1560
timestamp 1704896540
transform 1 0 17816 0 1 52909
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1561
timestamp 1704896540
transform 1 0 17816 0 1 52229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1562
timestamp 1704896540
transform 1 0 19040 0 1 51685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1563
timestamp 1704896540
transform 1 0 19040 0 1 51413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1564
timestamp 1704896540
transform 1 0 19176 0 1 51277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1565
timestamp 1704896540
transform 1 0 19176 0 1 51005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1566
timestamp 1704896540
transform 1 0 19176 0 1 53861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1567
timestamp 1704896540
transform 1 0 19448 0 1 52093
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1568
timestamp 1704896540
transform 1 0 19448 0 1 51821
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1569
timestamp 1704896540
transform 1 0 19176 0 1 54133
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1570
timestamp 1704896540
transform 1 0 19176 0 1 53317
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1571
timestamp 1704896540
transform 1 0 19176 0 1 53045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1572
timestamp 1704896540
transform 1 0 19040 0 1 52637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1573
timestamp 1704896540
transform 1 0 19448 0 1 51005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1574
timestamp 1704896540
transform 1 0 19448 0 1 51277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1575
timestamp 1704896540
transform 1 0 19584 0 1 51685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1576
timestamp 1704896540
transform 1 0 19584 0 1 51413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1577
timestamp 1704896540
transform 1 0 19040 0 1 52909
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1578
timestamp 1704896540
transform 1 0 19448 0 1 54133
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1579
timestamp 1704896540
transform 1 0 19448 0 1 53861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1580
timestamp 1704896540
transform 1 0 19448 0 1 53045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1581
timestamp 1704896540
transform 1 0 19448 0 1 53317
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1582
timestamp 1704896540
transform 1 0 19448 0 1 53725
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1583
timestamp 1704896540
transform 1 0 19448 0 1 53453
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1584
timestamp 1704896540
transform 1 0 18360 0 1 54269
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1585
timestamp 1704896540
transform 1 0 19584 0 1 55629
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1586
timestamp 1704896540
transform 1 0 19584 0 1 55357
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1587
timestamp 1704896540
transform 1 0 17816 0 1 53045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1588
timestamp 1704896540
transform 1 0 17816 0 1 53317
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1589
timestamp 1704896540
transform 1 0 17816 0 1 53725
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1590
timestamp 1704896540
transform 1 0 17816 0 1 53453
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1591
timestamp 1704896540
transform 1 0 17952 0 1 53861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1592
timestamp 1704896540
transform 1 0 17952 0 1 54133
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1593
timestamp 1704896540
transform 1 0 18496 0 1 51005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1594
timestamp 1704896540
transform 1 0 18496 0 1 51277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1595
timestamp 1704896540
transform 1 0 17816 0 1 51005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1596
timestamp 1704896540
transform 1 0 18496 0 1 52501
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1597
timestamp 1704896540
transform 1 0 18496 0 1 52229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1598
timestamp 1704896540
transform 1 0 18360 0 1 52501
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1599
timestamp 1704896540
transform 1 0 18360 0 1 52229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1600
timestamp 1704896540
transform 1 0 17816 0 1 50733
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1601
timestamp 1704896540
transform 1 0 17952 0 1 50597
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1602
timestamp 1704896540
transform 1 0 17952 0 1 50325
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1603
timestamp 1704896540
transform 1 0 19176 0 1 55629
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1604
timestamp 1704896540
transform 1 0 19176 0 1 55357
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1605
timestamp 1704896540
transform 1 0 18904 0 1 52093
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1606
timestamp 1704896540
transform 1 0 18904 0 1 51821
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1607
timestamp 1704896540
transform 1 0 18496 0 1 53045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1608
timestamp 1704896540
transform 1 0 18496 0 1 53317
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1609
timestamp 1704896540
transform 1 0 18904 0 1 51141
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1610
timestamp 1704896540
transform 1 0 18904 0 1 50733
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1611
timestamp 1704896540
transform 1 0 18632 0 1 50325
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1612
timestamp 1704896540
transform 1 0 18632 0 1 50597
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1613
timestamp 1704896540
transform 1 0 17952 0 1 54949
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1614
timestamp 1704896540
transform 1 0 18632 0 1 55221
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1615
timestamp 1704896540
transform 1 0 18632 0 1 54949
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1616
timestamp 1704896540
transform 1 0 17952 0 1 54677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1617
timestamp 1704896540
transform 1 0 18904 0 1 52637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1618
timestamp 1704896540
transform 1 0 18904 0 1 52909
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1619
timestamp 1704896540
transform 1 0 17816 0 1 54269
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1620
timestamp 1704896540
transform 1 0 17816 0 1 54541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1621
timestamp 1704896540
transform 1 0 18496 0 1 54269
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1622
timestamp 1704896540
transform 1 0 18496 0 1 54541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1623
timestamp 1704896540
transform 1 0 17952 0 1 50189
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1624
timestamp 1704896540
transform 1 0 1224 0 1 47333
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1625
timestamp 1704896540
transform 1 0 1224 0 1 48965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1626
timestamp 1704896540
transform 1 0 1224 0 1 45701
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1627
timestamp 1704896540
transform 1 0 1224 0 1 54133
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1628
timestamp 1704896540
transform 1 0 1224 0 1 52501
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1629
timestamp 1704896540
transform 1 0 1224 0 1 50733
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1630
timestamp 1704896540
transform 1 0 1224 0 1 60797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1631
timestamp 1704896540
transform 1 0 1224 0 1 55765
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1632
timestamp 1704896540
transform 1 0 1224 0 1 59165
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1633
timestamp 1704896540
transform 1 0 1224 0 1 57397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1634
timestamp 1704896540
transform 1 0 1224 0 1 64197
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1635
timestamp 1704896540
transform 1 0 1224 0 1 65829
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1636
timestamp 1704896540
transform 1 0 1224 0 1 62429
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1637
timestamp 1704896540
transform 1 0 18768 0 1 59981
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1638
timestamp 1704896540
transform 1 0 18768 0 1 59709
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1639
timestamp 1704896540
transform 1 0 19176 0 1 59709
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1640
timestamp 1704896540
transform 1 0 19176 0 1 59981
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1641
timestamp 1704896540
transform 1 0 18496 0 1 59709
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1642
timestamp 1704896540
transform 1 0 18496 0 1 59981
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1643
timestamp 1704896540
transform 1 0 18360 0 1 59709
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1644
timestamp 1704896540
transform 1 0 18360 0 1 59981
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1645
timestamp 1704896540
transform 1 0 18360 0 1 61205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1646
timestamp 1704896540
transform 1 0 18360 0 1 60933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1647
timestamp 1704896540
transform 1 0 19040 0 1 60797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1648
timestamp 1704896540
transform 1 0 19040 0 1 60525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1649
timestamp 1704896540
transform 1 0 17952 0 1 56581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1650
timestamp 1704896540
transform 1 0 17952 0 1 56853
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1651
timestamp 1704896540
transform 1 0 17816 0 1 56445
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1652
timestamp 1704896540
transform 1 0 17816 0 1 56173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1653
timestamp 1704896540
transform 1 0 18496 0 1 58757
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1654
timestamp 1704896540
transform 1 0 18496 0 1 58485
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1655
timestamp 1704896540
transform 1 0 17816 0 1 58485
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1656
timestamp 1704896540
transform 1 0 19176 0 1 56173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1657
timestamp 1704896540
transform 1 0 19176 0 1 56445
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1658
timestamp 1704896540
transform 1 0 19176 0 1 56853
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1659
timestamp 1704896540
transform 1 0 18496 0 1 56853
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1660
timestamp 1704896540
transform 1 0 18496 0 1 56581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1661
timestamp 1704896540
transform 1 0 18496 0 1 56173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1662
timestamp 1704896540
transform 1 0 18496 0 1 56445
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1663
timestamp 1704896540
transform 1 0 18360 0 1 56853
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1664
timestamp 1704896540
transform 1 0 18360 0 1 56581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1665
timestamp 1704896540
transform 1 0 18360 0 1 56173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1666
timestamp 1704896540
transform 1 0 18360 0 1 56445
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1667
timestamp 1704896540
transform 1 0 18224 0 1 56989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1668
timestamp 1704896540
transform 1 0 18224 0 1 57261
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1669
timestamp 1704896540
transform 1 0 19176 0 1 56581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1670
timestamp 1704896540
transform 1 0 17816 0 1 58213
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1671
timestamp 1704896540
transform 1 0 18224 0 1 60117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1672
timestamp 1704896540
transform 1 0 18224 0 1 60389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1673
timestamp 1704896540
transform 1 0 17816 0 1 56989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1674
timestamp 1704896540
transform 1 0 19176 0 1 57669
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1675
timestamp 1704896540
transform 1 0 19176 0 1 57397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1676
timestamp 1704896540
transform 1 0 19040 0 1 56989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1677
timestamp 1704896540
transform 1 0 19448 0 1 57397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1678
timestamp 1704896540
transform 1 0 19448 0 1 57669
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1679
timestamp 1704896540
transform 1 0 19448 0 1 58077
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1680
timestamp 1704896540
transform 1 0 19448 0 1 57805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1681
timestamp 1704896540
transform 1 0 19040 0 1 57261
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1682
timestamp 1704896540
transform 1 0 19040 0 1 56037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1683
timestamp 1704896540
transform 1 0 19040 0 1 55765
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1684
timestamp 1704896540
transform 1 0 19040 0 1 57805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1685
timestamp 1704896540
transform 1 0 19584 0 1 56173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1686
timestamp 1704896540
transform 1 0 19584 0 1 56445
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1687
timestamp 1704896540
transform 1 0 19040 0 1 58077
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1688
timestamp 1704896540
transform 1 0 17816 0 1 57261
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1689
timestamp 1704896540
transform 1 0 19448 0 1 59709
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1690
timestamp 1704896540
transform 1 0 19448 0 1 59981
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1691
timestamp 1704896540
transform 1 0 17816 0 1 59437
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1692
timestamp 1704896540
transform 1 0 19040 0 1 60933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1693
timestamp 1704896540
transform 1 0 19584 0 1 57261
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1694
timestamp 1704896540
transform 1 0 19584 0 1 56989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1695
timestamp 1704896540
transform 1 0 19584 0 1 56581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1696
timestamp 1704896540
transform 1 0 19584 0 1 56853
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1697
timestamp 1704896540
transform 1 0 19040 0 1 61205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1698
timestamp 1704896540
transform 1 0 17816 0 1 59709
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1699
timestamp 1704896540
transform 1 0 19584 0 1 60933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1700
timestamp 1704896540
transform 1 0 19584 0 1 61205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1701
timestamp 1704896540
transform 1 0 17816 0 1 58621
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1702
timestamp 1704896540
transform 1 0 17816 0 1 58893
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1703
timestamp 1704896540
transform 1 0 19584 0 1 56037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1704
timestamp 1704896540
transform 1 0 19584 0 1 55765
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1705
timestamp 1704896540
transform 1 0 18632 0 1 60525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1706
timestamp 1704896540
transform 1 0 18632 0 1 60797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1707
timestamp 1704896540
transform 1 0 18768 0 1 61205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1708
timestamp 1704896540
transform 1 0 17816 0 1 57397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1709
timestamp 1704896540
transform 1 0 17816 0 1 57669
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1710
timestamp 1704896540
transform 1 0 17952 0 1 60117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1711
timestamp 1704896540
transform 1 0 17952 0 1 61205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1712
timestamp 1704896540
transform 1 0 17952 0 1 60933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1713
timestamp 1704896540
transform 1 0 19584 0 1 59573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1714
timestamp 1704896540
transform 1 0 19584 0 1 59301
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1715
timestamp 1704896540
transform 1 0 19448 0 1 60797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1716
timestamp 1704896540
transform 1 0 19448 0 1 60525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1717
timestamp 1704896540
transform 1 0 19448 0 1 60117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1718
timestamp 1704896540
transform 1 0 19448 0 1 60389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1719
timestamp 1704896540
transform 1 0 18768 0 1 58213
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1720
timestamp 1704896540
transform 1 0 18768 0 1 58485
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1721
timestamp 1704896540
transform 1 0 17952 0 1 60389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1722
timestamp 1704896540
transform 1 0 17816 0 1 58077
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1723
timestamp 1704896540
transform 1 0 18632 0 1 57669
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1724
timestamp 1704896540
transform 1 0 18632 0 1 57397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1725
timestamp 1704896540
transform 1 0 17816 0 1 57805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1726
timestamp 1704896540
transform 1 0 19176 0 1 59301
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1727
timestamp 1704896540
transform 1 0 18904 0 1 58893
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1728
timestamp 1704896540
transform 1 0 18904 0 1 59165
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1729
timestamp 1704896540
transform 1 0 18904 0 1 60389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1730
timestamp 1704896540
transform 1 0 18904 0 1 60117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1731
timestamp 1704896540
transform 1 0 18904 0 1 55765
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1732
timestamp 1704896540
transform 1 0 18904 0 1 56037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1733
timestamp 1704896540
transform 1 0 19176 0 1 59573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1734
timestamp 1704896540
transform 1 0 18768 0 1 60933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1735
timestamp 1704896540
transform 1 0 19040 0 1 60389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1736
timestamp 1704896540
transform 1 0 19040 0 1 60117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1737
timestamp 1704896540
transform 1 0 18904 0 1 66101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1738
timestamp 1704896540
transform 1 0 18904 0 1 66373
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1739
timestamp 1704896540
transform 1 0 18496 0 1 65557
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1740
timestamp 1704896540
transform 1 0 18496 0 1 65285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1741
timestamp 1704896540
transform 1 0 18224 0 1 65285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1742
timestamp 1704896540
transform 1 0 18224 0 1 65557
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1743
timestamp 1704896540
transform 1 0 18224 0 1 65693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1744
timestamp 1704896540
transform 1 0 18224 0 1 65965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1745
timestamp 1704896540
transform 1 0 18224 0 1 61341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1746
timestamp 1704896540
transform 1 0 18224 0 1 61613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1747
timestamp 1704896540
transform 1 0 18224 0 1 64469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1748
timestamp 1704896540
transform 1 0 18224 0 1 64741
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1749
timestamp 1704896540
transform 1 0 18496 0 1 62973
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1750
timestamp 1704896540
transform 1 0 18496 0 1 63245
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1751
timestamp 1704896540
transform 1 0 18360 0 1 62429
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1752
timestamp 1704896540
transform 1 0 18360 0 1 62157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1753
timestamp 1704896540
transform 1 0 18360 0 1 64333
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1754
timestamp 1704896540
transform 1 0 18360 0 1 64061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1755
timestamp 1704896540
transform 1 0 19448 0 1 64877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1756
timestamp 1704896540
transform 1 0 19448 0 1 65149
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1757
timestamp 1704896540
transform 1 0 19448 0 1 65557
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1758
timestamp 1704896540
transform 1 0 19448 0 1 65285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1759
timestamp 1704896540
transform 1 0 19584 0 1 64741
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1760
timestamp 1704896540
transform 1 0 19584 0 1 64469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1761
timestamp 1704896540
transform 1 0 19448 0 1 65693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1762
timestamp 1704896540
transform 1 0 19448 0 1 65965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1763
timestamp 1704896540
transform 1 0 19448 0 1 66101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1764
timestamp 1704896540
transform 1 0 19448 0 1 66373
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1765
timestamp 1704896540
transform 1 0 19448 0 1 61341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1766
timestamp 1704896540
transform 1 0 19448 0 1 61613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1767
timestamp 1704896540
transform 1 0 19448 0 1 61749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1768
timestamp 1704896540
transform 1 0 19448 0 1 62021
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1769
timestamp 1704896540
transform 1 0 19584 0 1 62157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1770
timestamp 1704896540
transform 1 0 19584 0 1 62429
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1771
timestamp 1704896540
transform 1 0 19584 0 1 63653
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1772
timestamp 1704896540
transform 1 0 19584 0 1 63925
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1773
timestamp 1704896540
transform 1 0 19584 0 1 64333
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1774
timestamp 1704896540
transform 1 0 19584 0 1 64061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1775
timestamp 1704896540
transform 1 0 18904 0 1 64469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1776
timestamp 1704896540
transform 1 0 18904 0 1 64741
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1777
timestamp 1704896540
transform 1 0 18904 0 1 63653
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1778
timestamp 1704896540
transform 1 0 18904 0 1 63925
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1779
timestamp 1704896540
transform 1 0 18768 0 1 61613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1780
timestamp 1704896540
transform 1 0 18768 0 1 61341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1781
timestamp 1704896540
transform 1 0 19176 0 1 62021
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1782
timestamp 1704896540
transform 1 0 19176 0 1 61749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1783
timestamp 1704896540
transform 1 0 18632 0 1 64877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1784
timestamp 1704896540
transform 1 0 18632 0 1 65149
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1785
timestamp 1704896540
transform 1 0 18904 0 1 61749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1786
timestamp 1704896540
transform 1 0 19176 0 1 66373
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1787
timestamp 1704896540
transform 1 0 19176 0 1 66101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1788
timestamp 1704896540
transform 1 0 19176 0 1 64877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1789
timestamp 1704896540
transform 1 0 19176 0 1 65149
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1790
timestamp 1704896540
transform 1 0 19176 0 1 63653
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1791
timestamp 1704896540
transform 1 0 19176 0 1 63925
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1792
timestamp 1704896540
transform 1 0 19040 0 1 61613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1793
timestamp 1704896540
transform 1 0 19040 0 1 61341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1794
timestamp 1704896540
transform 1 0 19040 0 1 62157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1795
timestamp 1704896540
transform 1 0 19040 0 1 62429
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1796
timestamp 1704896540
transform 1 0 18904 0 1 62021
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1797
timestamp 1704896540
transform 1 0 19040 0 1 65965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1798
timestamp 1704896540
transform 1 0 19040 0 1 65693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1799
timestamp 1704896540
transform 1 0 19040 0 1 65285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1800
timestamp 1704896540
transform 1 0 19040 0 1 65557
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1801
timestamp 1704896540
transform 1 0 19040 0 1 64741
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1802
timestamp 1704896540
transform 1 0 19040 0 1 64469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1803
timestamp 1704896540
transform 1 0 19176 0 1 64061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1804
timestamp 1704896540
transform 1 0 19176 0 1 64333
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1805
timestamp 1704896540
transform 1 0 17816 0 1 65557
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1806
timestamp 1704896540
transform 1 0 17816 0 1 65285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1807
timestamp 1704896540
transform 1 0 17952 0 1 63245
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1808
timestamp 1704896540
transform 1 0 17952 0 1 62973
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1809
timestamp 1704896540
transform 1 0 17952 0 1 62565
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1810
timestamp 1704896540
transform 1 0 17952 0 1 62837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1811
timestamp 1704896540
transform 1 0 17816 0 1 63381
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1812
timestamp 1704896540
transform 1 0 17816 0 1 63653
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1813
timestamp 1704896540
transform 1 0 17952 0 1 64333
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1814
timestamp 1704896540
transform 1 0 17952 0 1 64061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1815
timestamp 1704896540
transform 1 0 17816 0 1 65693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1816
timestamp 1704896540
transform 1 0 17816 0 1 65965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1817
timestamp 1704896540
transform 1 0 17952 0 1 66373
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1818
timestamp 1704896540
transform 1 0 17952 0 1 66101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1819
timestamp 1704896540
transform 1 0 17816 0 1 66509
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1820
timestamp 1704896540
transform 1 0 17816 0 1 61341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1821
timestamp 1704896540
transform 1 0 17816 0 1 61613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1822
timestamp 1704896540
transform 1 0 17816 0 1 65149
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1823
timestamp 1704896540
transform 1 0 17816 0 1 64877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1824
timestamp 1704896540
transform 1 0 17816 0 1 62429
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1825
timestamp 1704896540
transform 1 0 17816 0 1 62157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1826
timestamp 1704896540
transform 1 0 17816 0 1 61749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1827
timestamp 1704896540
transform 1 0 17816 0 1 62021
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1828
timestamp 1704896540
transform 1 0 18768 0 1 65965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1829
timestamp 1704896540
transform 1 0 18768 0 1 65693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1830
timestamp 1704896540
transform 1 0 19584 0 1 69637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1831
timestamp 1704896540
transform 1 0 19584 0 1 69909
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1832
timestamp 1704896540
transform 1 0 19584 0 1 70317
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1833
timestamp 1704896540
transform 1 0 19584 0 1 70045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1834
timestamp 1704896540
transform 1 0 19448 0 1 67869
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1835
timestamp 1704896540
transform 1 0 19448 0 1 67597
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1836
timestamp 1704896540
transform 1 0 19176 0 1 68413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1837
timestamp 1704896540
transform 1 0 19176 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1838
timestamp 1704896540
transform 1 0 18904 0 1 70045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1839
timestamp 1704896540
transform 1 0 18904 0 1 70317
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1840
timestamp 1704896540
transform 1 0 18496 0 1 67869
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1841
timestamp 1704896540
transform 1 0 18496 0 1 67597
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1842
timestamp 1704896540
transform 1 0 18496 0 1 66917
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1843
timestamp 1704896540
transform 1 0 18496 0 1 67189
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1844
timestamp 1704896540
transform 1 0 18224 0 1 69637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1845
timestamp 1704896540
transform 1 0 18224 0 1 69909
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1846
timestamp 1704896540
transform 1 0 18496 0 1 69093
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1847
timestamp 1704896540
transform 1 0 18496 0 1 68821
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1848
timestamp 1704896540
transform 1 0 18224 0 1 70045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1849
timestamp 1704896540
transform 1 0 18224 0 1 70317
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1850
timestamp 1704896540
transform 1 0 18224 0 1 69501
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1851
timestamp 1704896540
transform 1 0 18224 0 1 69229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1852
timestamp 1704896540
transform 1 0 18224 0 1 68821
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1853
timestamp 1704896540
transform 1 0 18224 0 1 69093
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1854
timestamp 1704896540
transform 1 0 18496 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1855
timestamp 1704896540
transform 1 0 18496 0 1 68413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1856
timestamp 1704896540
transform 1 0 18360 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1857
timestamp 1704896540
transform 1 0 18360 0 1 68413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1858
timestamp 1704896540
transform 1 0 19040 0 1 69093
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1859
timestamp 1704896540
transform 1 0 19040 0 1 68821
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1860
timestamp 1704896540
transform 1 0 19176 0 1 69909
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1861
timestamp 1704896540
transform 1 0 19176 0 1 69637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1862
timestamp 1704896540
transform 1 0 19176 0 1 69229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1863
timestamp 1704896540
transform 1 0 19176 0 1 69501
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1864
timestamp 1704896540
transform 1 0 19040 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1865
timestamp 1704896540
transform 1 0 19040 0 1 68005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1866
timestamp 1704896540
transform 1 0 19040 0 1 67597
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1867
timestamp 1704896540
transform 1 0 19040 0 1 67869
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1868
timestamp 1704896540
transform 1 0 17952 0 1 70317
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1869
timestamp 1704896540
transform 1 0 17816 0 1 67325
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1870
timestamp 1704896540
transform 1 0 17816 0 1 67597
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1871
timestamp 1704896540
transform 1 0 17816 0 1 69501
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1872
timestamp 1704896540
transform 1 0 17816 0 1 69229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1873
timestamp 1704896540
transform 1 0 17816 0 1 68821
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1874
timestamp 1704896540
transform 1 0 17816 0 1 69093
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1875
timestamp 1704896540
transform 1 0 17816 0 1 67189
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1876
timestamp 1704896540
transform 1 0 17816 0 1 66917
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1877
timestamp 1704896540
transform 1 0 17952 0 1 70045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1878
timestamp 1704896540
transform 1 0 17952 0 1 69637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1879
timestamp 1704896540
transform 1 0 19040 0 1 70317
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1880
timestamp 1704896540
transform 1 0 19040 0 1 70045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1881
timestamp 1704896540
transform 1 0 17952 0 1 69909
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1882
timestamp 1704896540
transform 1 0 19448 0 1 69229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1883
timestamp 1704896540
transform 1 0 19448 0 1 69501
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1884
timestamp 1704896540
transform 1 0 19584 0 1 68005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1885
timestamp 1704896540
transform 1 0 19584 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1886
timestamp 1704896540
transform 1 0 19584 0 1 69093
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1887
timestamp 1704896540
transform 1 0 19584 0 1 68821
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1888
timestamp 1704896540
transform 1 0 19448 0 1 68413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1889
timestamp 1704896540
transform 1 0 19448 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1890
timestamp 1704896540
transform 1 0 1224 0 1 69229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1891
timestamp 1704896540
transform 1 0 1224 0 1 70997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1892
timestamp 1704896540
transform 1 0 1224 0 1 67733
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1893
timestamp 1704896540
transform 1 0 1224 0 1 77661
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1894
timestamp 1704896540
transform 1 0 1224 0 1 75893
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1895
timestamp 1704896540
transform 1 0 1224 0 1 72629
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1896
timestamp 1704896540
transform 1 0 1224 0 1 74261
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1897
timestamp 1704896540
transform 1 0 1224 0 1 82693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1898
timestamp 1704896540
transform 1 0 1224 0 1 80925
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1899
timestamp 1704896540
transform 1 0 1224 0 1 79293
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1900
timestamp 1704896540
transform 1 0 5304 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1901
timestamp 1704896540
transform 1 0 5304 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1902
timestamp 1704896540
transform 1 0 3808 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1903
timestamp 1704896540
transform 1 0 3808 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1904
timestamp 1704896540
transform 1 0 2176 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1905
timestamp 1704896540
transform 1 0 2176 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1906
timestamp 1704896540
transform 1 0 1224 0 1 85957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1907
timestamp 1704896540
transform 1 0 1224 0 1 84325
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1908
timestamp 1704896540
transform 1 0 10336 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1909
timestamp 1704896540
transform 1 0 10336 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1910
timestamp 1704896540
transform 1 0 8840 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1911
timestamp 1704896540
transform 1 0 8840 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1912
timestamp 1704896540
transform 1 0 7072 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1913
timestamp 1704896540
transform 1 0 7072 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1914
timestamp 1704896540
transform 1 0 22168 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1915
timestamp 1704896540
transform 1 0 22168 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1916
timestamp 1704896540
transform 1 0 20536 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1917
timestamp 1704896540
transform 1 0 20536 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1918
timestamp 1704896540
transform 1 0 18904 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1919
timestamp 1704896540
transform 1 0 18904 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1920
timestamp 1704896540
transform 1 0 17272 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1921
timestamp 1704896540
transform 1 0 17272 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1922
timestamp 1704896540
transform 1 0 15368 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1923
timestamp 1704896540
transform 1 0 15368 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1924
timestamp 1704896540
transform 1 0 13872 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1925
timestamp 1704896540
transform 1 0 13872 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1926
timestamp 1704896540
transform 1 0 12104 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1927
timestamp 1704896540
transform 1 0 12104 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1928
timestamp 1704896540
transform 1 0 43248 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1929
timestamp 1704896540
transform 1 0 43248 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1930
timestamp 1704896540
transform 1 0 41072 0 1 73581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1931
timestamp 1704896540
transform 1 0 40936 0 1 76029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1932
timestamp 1704896540
transform 1 0 41072 0 1 76029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1933
timestamp 1704896540
transform 1 0 41072 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1934
timestamp 1704896540
transform 1 0 36040 0 1 73581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1935
timestamp 1704896540
transform 1 0 36040 0 1 76029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1936
timestamp 1704896540
transform 1 0 35904 0 1 76029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1937
timestamp 1704896540
transform 1 0 35904 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1938
timestamp 1704896540
transform 1 0 42704 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1939
timestamp 1704896540
transform 1 0 42704 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1940
timestamp 1704896540
transform 1 0 35768 0 1 77525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1941
timestamp 1704896540
transform 1 0 35768 0 1 76845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1942
timestamp 1704896540
transform 1 0 41616 0 1 71269
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1943
timestamp 1704896540
transform 1 0 41616 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1944
timestamp 1704896540
transform 1 0 40936 0 1 77525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1945
timestamp 1704896540
transform 1 0 40936 0 1 76845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1946
timestamp 1704896540
transform 1 0 35768 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1947
timestamp 1704896540
transform 1 0 35768 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1948
timestamp 1704896540
transform 1 0 40800 0 1 76573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1949
timestamp 1704896540
transform 1 0 40800 0 1 71949
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1950
timestamp 1704896540
transform 1 0 40664 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1951
timestamp 1704896540
transform 1 0 40664 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1952
timestamp 1704896540
transform 1 0 40256 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1953
timestamp 1704896540
transform 1 0 40256 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1954
timestamp 1704896540
transform 1 0 39440 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1955
timestamp 1704896540
transform 1 0 39440 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1956
timestamp 1704896540
transform 1 0 34408 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1957
timestamp 1704896540
transform 1 0 34408 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1958
timestamp 1704896540
transform 1 0 38216 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1959
timestamp 1704896540
transform 1 0 38216 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1960
timestamp 1704896540
transform 1 0 37672 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1961
timestamp 1704896540
transform 1 0 37672 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1962
timestamp 1704896540
transform 1 0 35224 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1963
timestamp 1704896540
transform 1 0 35224 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1964
timestamp 1704896540
transform 1 0 36992 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1965
timestamp 1704896540
transform 1 0 36992 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1966
timestamp 1704896540
transform 1 0 36448 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1967
timestamp 1704896540
transform 1 0 36448 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1968
timestamp 1704896540
transform 1 0 45152 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1969
timestamp 1704896540
transform 1 0 45152 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1970
timestamp 1704896540
transform 1 0 36856 0 1 71949
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1971
timestamp 1704896540
transform 1 0 36856 0 1 76573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1972
timestamp 1704896540
transform 1 0 43928 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1973
timestamp 1704896540
transform 1 0 43928 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1974
timestamp 1704896540
transform 1 0 34000 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1975
timestamp 1704896540
transform 1 0 34000 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1976
timestamp 1704896540
transform 1 0 33048 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1977
timestamp 1704896540
transform 1 0 33048 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1978
timestamp 1704896540
transform 1 0 26792 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1979
timestamp 1704896540
transform 1 0 31008 0 1 73581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1980
timestamp 1704896540
transform 1 0 31008 0 1 76029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1981
timestamp 1704896540
transform 1 0 30872 0 1 76029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1982
timestamp 1704896540
transform 1 0 30872 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1983
timestamp 1704896540
transform 1 0 26112 0 1 73581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1984
timestamp 1704896540
transform 1 0 26112 0 1 76029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1985
timestamp 1704896540
transform 1 0 25976 0 1 76029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1986
timestamp 1704896540
transform 1 0 25976 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1987
timestamp 1704896540
transform 1 0 24344 0 1 67325
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1988
timestamp 1704896540
transform 1 0 24344 0 1 67053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1989
timestamp 1704896540
transform 1 0 24616 0 1 66917
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1990
timestamp 1704896540
transform 1 0 25976 0 1 73309
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1991
timestamp 1704896540
transform 1 0 25976 0 1 70861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1992
timestamp 1704896540
transform 1 0 26792 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1993
timestamp 1704896540
transform 1 0 32504 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1994
timestamp 1704896540
transform 1 0 32504 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1995
timestamp 1704896540
transform 1 0 31960 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1996
timestamp 1704896540
transform 1 0 31960 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1997
timestamp 1704896540
transform 1 0 31416 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1998
timestamp 1704896540
transform 1 0 31416 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_1999
timestamp 1704896540
transform 1 0 30736 0 1 77525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2000
timestamp 1704896540
transform 1 0 30736 0 1 76845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2001
timestamp 1704896540
transform 1 0 30736 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2002
timestamp 1704896540
transform 1 0 30736 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2003
timestamp 1704896540
transform 1 0 25840 0 1 77525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2004
timestamp 1704896540
transform 1 0 25840 0 1 76845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2005
timestamp 1704896540
transform 1 0 30328 0 1 76573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2006
timestamp 1704896540
transform 1 0 30328 0 1 71949
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2007
timestamp 1704896540
transform 1 0 29512 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2008
timestamp 1704896540
transform 1 0 29512 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2009
timestamp 1704896540
transform 1 0 25840 0 1 76573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2010
timestamp 1704896540
transform 1 0 25840 0 1 71949
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2011
timestamp 1704896540
transform 1 0 28968 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2012
timestamp 1704896540
transform 1 0 28968 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2013
timestamp 1704896540
transform 1 0 27744 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2014
timestamp 1704896540
transform 1 0 27744 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2015
timestamp 1704896540
transform 1 0 25568 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2016
timestamp 1704896540
transform 1 0 25568 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2017
timestamp 1704896540
transform 1 0 27608 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2018
timestamp 1704896540
transform 1 0 27608 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2019
timestamp 1704896540
transform 1 0 23936 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2020
timestamp 1704896540
transform 1 0 32368 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2021
timestamp 1704896540
transform 1 0 32368 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2022
timestamp 1704896540
transform 1 0 30600 0 1 77933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2023
timestamp 1704896540
transform 1 0 25568 0 1 77933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2024
timestamp 1704896540
transform 1 0 30464 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2025
timestamp 1704896540
transform 1 0 30464 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2026
timestamp 1704896540
transform 1 0 28832 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2027
timestamp 1704896540
transform 1 0 28832 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2028
timestamp 1704896540
transform 1 0 27336 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2029
timestamp 1704896540
transform 1 0 27336 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2030
timestamp 1704896540
transform 1 0 25432 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2031
timestamp 1704896540
transform 1 0 25432 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2032
timestamp 1704896540
transform 1 0 23936 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2033
timestamp 1704896540
transform 1 0 33864 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2034
timestamp 1704896540
transform 1 0 33864 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2035
timestamp 1704896540
transform 1 0 40664 0 1 77933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2036
timestamp 1704896540
transform 1 0 35632 0 1 77933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2037
timestamp 1704896540
transform 1 0 43928 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2038
timestamp 1704896540
transform 1 0 43928 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2039
timestamp 1704896540
transform 1 0 42432 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2040
timestamp 1704896540
transform 1 0 42432 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2041
timestamp 1704896540
transform 1 0 40936 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2042
timestamp 1704896540
transform 1 0 40936 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2043
timestamp 1704896540
transform 1 0 39032 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2044
timestamp 1704896540
transform 1 0 39032 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2045
timestamp 1704896540
transform 1 0 37400 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2046
timestamp 1704896540
transform 1 0 37400 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2047
timestamp 1704896540
transform 1 0 35904 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2048
timestamp 1704896540
transform 1 0 35904 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2049
timestamp 1704896540
transform 1 0 22848 0 1 46109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2050
timestamp 1704896540
transform 1 0 22848 0 1 45565
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2051
timestamp 1704896540
transform 1 0 17816 0 1 66781
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2052
timestamp 1704896540
transform 1 0 89760 0 1 47333
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2053
timestamp 1704896540
transform 1 0 89760 0 1 49101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2054
timestamp 1704896540
transform 1 0 89760 0 1 45701
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2055
timestamp 1704896540
transform 1 0 89760 0 1 52365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2056
timestamp 1704896540
transform 1 0 89760 0 1 54133
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2057
timestamp 1704896540
transform 1 0 89760 0 1 50733
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2058
timestamp 1704896540
transform 1 0 70720 0 1 45429
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2059
timestamp 1704896540
transform 1 0 69360 0 1 45973
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2060
timestamp 1704896540
transform 1 0 72080 0 1 45837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2061
timestamp 1704896540
transform 1 0 71672 0 1 45429
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2062
timestamp 1704896540
transform 1 0 71672 0 1 45157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2063
timestamp 1704896540
transform 1 0 71264 0 1 49101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2064
timestamp 1704896540
transform 1 0 71264 0 1 48149
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2065
timestamp 1704896540
transform 1 0 71264 0 1 49373
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2066
timestamp 1704896540
transform 1 0 72352 0 1 45429
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2067
timestamp 1704896540
transform 1 0 72352 0 1 45157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2068
timestamp 1704896540
transform 1 0 72216 0 1 45429
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2069
timestamp 1704896540
transform 1 0 71808 0 1 47469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2070
timestamp 1704896540
transform 1 0 71808 0 1 47741
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2071
timestamp 1704896540
transform 1 0 72216 0 1 45157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2072
timestamp 1704896540
transform 1 0 72488 0 1 45565
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2073
timestamp 1704896540
transform 1 0 72488 0 1 45837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2074
timestamp 1704896540
transform 1 0 71264 0 1 49781
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2075
timestamp 1704896540
transform 1 0 71264 0 1 49509
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2076
timestamp 1704896540
transform 1 0 71264 0 1 47877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2077
timestamp 1704896540
transform 1 0 72624 0 1 49781
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2078
timestamp 1704896540
transform 1 0 72488 0 1 45021
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2079
timestamp 1704896540
transform 1 0 72488 0 1 44749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2080
timestamp 1704896540
transform 1 0 72624 0 1 49509
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2081
timestamp 1704896540
transform 1 0 71400 0 1 45837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2082
timestamp 1704896540
transform 1 0 71672 0 1 45565
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2083
timestamp 1704896540
transform 1 0 71672 0 1 45837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2084
timestamp 1704896540
transform 1 0 71264 0 1 44749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2085
timestamp 1704896540
transform 1 0 71264 0 1 45021
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2086
timestamp 1704896540
transform 1 0 72216 0 1 47061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2087
timestamp 1704896540
transform 1 0 72216 0 1 47333
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2088
timestamp 1704896540
transform 1 0 73032 0 1 46245
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2089
timestamp 1704896540
transform 1 0 73032 0 1 45973
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2090
timestamp 1704896540
transform 1 0 71264 0 1 45429
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2091
timestamp 1704896540
transform 1 0 71264 0 1 45157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2092
timestamp 1704896540
transform 1 0 72896 0 1 45837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2093
timestamp 1704896540
transform 1 0 72896 0 1 45565
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2094
timestamp 1704896540
transform 1 0 72624 0 1 49101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2095
timestamp 1704896540
transform 1 0 72624 0 1 49373
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2096
timestamp 1704896540
transform 1 0 73032 0 1 45429
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2097
timestamp 1704896540
transform 1 0 73032 0 1 45157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2098
timestamp 1704896540
transform 1 0 73032 0 1 44749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2099
timestamp 1704896540
transform 1 0 73032 0 1 45021
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2100
timestamp 1704896540
transform 1 0 73032 0 1 48285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2101
timestamp 1704896540
transform 1 0 73032 0 1 48557
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2102
timestamp 1704896540
transform 1 0 72896 0 1 48693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2103
timestamp 1704896540
transform 1 0 72896 0 1 48965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2104
timestamp 1704896540
transform 1 0 71400 0 1 48693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2105
timestamp 1704896540
transform 1 0 71264 0 1 48285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2106
timestamp 1704896540
transform 1 0 71264 0 1 48557
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2107
timestamp 1704896540
transform 1 0 71400 0 1 45565
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2108
timestamp 1704896540
transform 1 0 71672 0 1 48285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2109
timestamp 1704896540
transform 1 0 72080 0 1 48149
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2110
timestamp 1704896540
transform 1 0 71672 0 1 48557
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2111
timestamp 1704896540
transform 1 0 71808 0 1 48965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2112
timestamp 1704896540
transform 1 0 71808 0 1 48693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2113
timestamp 1704896540
transform 1 0 70720 0 1 45157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2114
timestamp 1704896540
transform 1 0 71264 0 1 47333
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2115
timestamp 1704896540
transform 1 0 72080 0 1 47877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2116
timestamp 1704896540
transform 1 0 71808 0 1 47877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2117
timestamp 1704896540
transform 1 0 71808 0 1 48149
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2118
timestamp 1704896540
transform 1 0 71672 0 1 49373
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2119
timestamp 1704896540
transform 1 0 69360 0 1 45565
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2120
timestamp 1704896540
transform 1 0 72080 0 1 45565
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2121
timestamp 1704896540
transform 1 0 72488 0 1 46653
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2122
timestamp 1704896540
transform 1 0 71672 0 1 45021
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2123
timestamp 1704896540
transform 1 0 71672 0 1 44749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2124
timestamp 1704896540
transform 1 0 72216 0 1 48285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2125
timestamp 1704896540
transform 1 0 72216 0 1 48557
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2126
timestamp 1704896540
transform 1 0 72488 0 1 48965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2127
timestamp 1704896540
transform 1 0 72488 0 1 48693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2128
timestamp 1704896540
transform 1 0 71808 0 1 47333
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2129
timestamp 1704896540
transform 1 0 71808 0 1 47061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2130
timestamp 1704896540
transform 1 0 72488 0 1 46381
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2131
timestamp 1704896540
transform 1 0 73032 0 1 49781
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2132
timestamp 1704896540
transform 1 0 73032 0 1 49509
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2133
timestamp 1704896540
transform 1 0 73032 0 1 49101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2134
timestamp 1704896540
transform 1 0 73032 0 1 49373
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2135
timestamp 1704896540
transform 1 0 71264 0 1 47741
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2136
timestamp 1704896540
transform 1 0 72080 0 1 49509
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2137
timestamp 1704896540
transform 1 0 72080 0 1 49781
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2138
timestamp 1704896540
transform 1 0 71264 0 1 47469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2139
timestamp 1704896540
transform 1 0 71264 0 1 47061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2140
timestamp 1704896540
transform 1 0 72080 0 1 48693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2141
timestamp 1704896540
transform 1 0 72896 0 1 47061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2142
timestamp 1704896540
transform 1 0 72896 0 1 46789
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2143
timestamp 1704896540
transform 1 0 72896 0 1 46381
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2144
timestamp 1704896540
transform 1 0 72896 0 1 46653
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2145
timestamp 1704896540
transform 1 0 71672 0 1 49781
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2146
timestamp 1704896540
transform 1 0 71672 0 1 49509
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2147
timestamp 1704896540
transform 1 0 72896 0 1 49917
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2148
timestamp 1704896540
transform 1 0 71672 0 1 49101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2149
timestamp 1704896540
transform 1 0 72080 0 1 48965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2150
timestamp 1704896540
transform 1 0 71400 0 1 48965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2151
timestamp 1704896540
transform 1 0 71264 0 1 52501
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2152
timestamp 1704896540
transform 1 0 72624 0 1 52229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2153
timestamp 1704896540
transform 1 0 72624 0 1 52501
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2154
timestamp 1704896540
transform 1 0 72488 0 1 51277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2155
timestamp 1704896540
transform 1 0 72488 0 1 51005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2156
timestamp 1704896540
transform 1 0 73032 0 1 52909
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2157
timestamp 1704896540
transform 1 0 73032 0 1 52637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2158
timestamp 1704896540
transform 1 0 72896 0 1 53045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2159
timestamp 1704896540
transform 1 0 72896 0 1 53317
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2160
timestamp 1704896540
transform 1 0 72896 0 1 52501
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2161
timestamp 1704896540
transform 1 0 72896 0 1 52229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2162
timestamp 1704896540
transform 1 0 73032 0 1 53453
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2163
timestamp 1704896540
transform 1 0 73032 0 1 53725
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2164
timestamp 1704896540
transform 1 0 73032 0 1 54133
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2165
timestamp 1704896540
transform 1 0 73032 0 1 53861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2166
timestamp 1704896540
transform 1 0 72352 0 1 50325
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2167
timestamp 1704896540
transform 1 0 72352 0 1 50597
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2168
timestamp 1704896540
transform 1 0 72352 0 1 55221
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2169
timestamp 1704896540
transform 1 0 72896 0 1 50733
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2170
timestamp 1704896540
transform 1 0 72896 0 1 51005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2171
timestamp 1704896540
transform 1 0 72352 0 1 54949
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2172
timestamp 1704896540
transform 1 0 72216 0 1 55221
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2173
timestamp 1704896540
transform 1 0 72216 0 1 54949
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2174
timestamp 1704896540
transform 1 0 72352 0 1 53317
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2175
timestamp 1704896540
transform 1 0 72896 0 1 54269
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2176
timestamp 1704896540
transform 1 0 72896 0 1 54541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2177
timestamp 1704896540
transform 1 0 73032 0 1 54949
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2178
timestamp 1704896540
transform 1 0 73032 0 1 54677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2179
timestamp 1704896540
transform 1 0 72488 0 1 51685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2180
timestamp 1704896540
transform 1 0 72352 0 1 51413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2181
timestamp 1704896540
transform 1 0 72352 0 1 53045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2182
timestamp 1704896540
transform 1 0 72216 0 1 52637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2183
timestamp 1704896540
transform 1 0 72216 0 1 52909
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2184
timestamp 1704896540
transform 1 0 72080 0 1 53317
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2185
timestamp 1704896540
transform 1 0 72352 0 1 54269
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2186
timestamp 1704896540
transform 1 0 72352 0 1 54541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2187
timestamp 1704896540
transform 1 0 72080 0 1 53045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2188
timestamp 1704896540
transform 1 0 73032 0 1 50597
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2189
timestamp 1704896540
transform 1 0 73032 0 1 50325
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2190
timestamp 1704896540
transform 1 0 71264 0 1 52229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2191
timestamp 1704896540
transform 1 0 71400 0 1 53725
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2192
timestamp 1704896540
transform 1 0 71400 0 1 53453
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2193
timestamp 1704896540
transform 1 0 71400 0 1 53045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2194
timestamp 1704896540
transform 1 0 71400 0 1 53317
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2195
timestamp 1704896540
transform 1 0 71400 0 1 55357
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2196
timestamp 1704896540
transform 1 0 71400 0 1 55629
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2197
timestamp 1704896540
transform 1 0 72352 0 1 52093
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2198
timestamp 1704896540
transform 1 0 72352 0 1 51821
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2199
timestamp 1704896540
transform 1 0 71400 0 1 53861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2200
timestamp 1704896540
transform 1 0 71400 0 1 54133
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2201
timestamp 1704896540
transform 1 0 71400 0 1 51005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2202
timestamp 1704896540
transform 1 0 72080 0 1 53725
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2203
timestamp 1704896540
transform 1 0 71672 0 1 51005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2204
timestamp 1704896540
transform 1 0 71672 0 1 51277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2205
timestamp 1704896540
transform 1 0 72080 0 1 53453
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2206
timestamp 1704896540
transform 1 0 72080 0 1 52501
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2207
timestamp 1704896540
transform 1 0 72080 0 1 52229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2208
timestamp 1704896540
transform 1 0 71400 0 1 51277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2209
timestamp 1704896540
transform 1 0 71264 0 1 52093
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2210
timestamp 1704896540
transform 1 0 71264 0 1 51821
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2211
timestamp 1704896540
transform 1 0 71672 0 1 52637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2212
timestamp 1704896540
transform 1 0 71672 0 1 52909
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2213
timestamp 1704896540
transform 1 0 71672 0 1 52501
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2214
timestamp 1704896540
transform 1 0 71672 0 1 52229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2215
timestamp 1704896540
transform 1 0 71264 0 1 51413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2216
timestamp 1704896540
transform 1 0 71264 0 1 51685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2217
timestamp 1704896540
transform 1 0 71264 0 1 52909
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2218
timestamp 1704896540
transform 1 0 71672 0 1 51413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2219
timestamp 1704896540
transform 1 0 71672 0 1 51685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2220
timestamp 1704896540
transform 1 0 71672 0 1 52093
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2221
timestamp 1704896540
transform 1 0 71672 0 1 51821
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2222
timestamp 1704896540
transform 1 0 71808 0 1 53861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2223
timestamp 1704896540
transform 1 0 71808 0 1 54133
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2224
timestamp 1704896540
transform 1 0 71808 0 1 55629
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2225
timestamp 1704896540
transform 1 0 71808 0 1 55357
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2226
timestamp 1704896540
transform 1 0 71672 0 1 53725
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2227
timestamp 1704896540
transform 1 0 71672 0 1 53453
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2228
timestamp 1704896540
transform 1 0 71672 0 1 53045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2229
timestamp 1704896540
transform 1 0 71672 0 1 53317
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2230
timestamp 1704896540
transform 1 0 71264 0 1 52637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2231
timestamp 1704896540
transform 1 0 72896 0 1 50189
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2232
timestamp 1704896540
transform 1 0 72216 0 1 57261
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2233
timestamp 1704896540
transform 1 0 72216 0 1 56989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2234
timestamp 1704896540
transform 1 0 72352 0 1 58485
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2235
timestamp 1704896540
transform 1 0 72352 0 1 58213
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2236
timestamp 1704896540
transform 1 0 72488 0 1 56581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2237
timestamp 1704896540
transform 1 0 72080 0 1 61205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2238
timestamp 1704896540
transform 1 0 71400 0 1 56173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2239
timestamp 1704896540
transform 1 0 71400 0 1 56445
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2240
timestamp 1704896540
transform 1 0 72080 0 1 60933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2241
timestamp 1704896540
transform 1 0 73032 0 1 56989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2242
timestamp 1704896540
transform 1 0 73032 0 1 57261
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2243
timestamp 1704896540
transform 1 0 72896 0 1 58893
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2244
timestamp 1704896540
transform 1 0 72896 0 1 58621
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2245
timestamp 1704896540
transform 1 0 71264 0 1 59573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2246
timestamp 1704896540
transform 1 0 71264 0 1 59301
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2247
timestamp 1704896540
transform 1 0 71400 0 1 61205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2248
timestamp 1704896540
transform 1 0 71400 0 1 60933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2249
timestamp 1704896540
transform 1 0 72080 0 1 59709
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2250
timestamp 1704896540
transform 1 0 72080 0 1 59981
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2251
timestamp 1704896540
transform 1 0 72080 0 1 58213
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2252
timestamp 1704896540
transform 1 0 72080 0 1 58485
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2253
timestamp 1704896540
transform 1 0 73032 0 1 58485
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2254
timestamp 1704896540
transform 1 0 73032 0 1 58213
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2255
timestamp 1704896540
transform 1 0 71264 0 1 57261
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2256
timestamp 1704896540
transform 1 0 71264 0 1 56989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2257
timestamp 1704896540
transform 1 0 72624 0 1 55765
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2258
timestamp 1704896540
transform 1 0 72624 0 1 56037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2259
timestamp 1704896540
transform 1 0 73032 0 1 60389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2260
timestamp 1704896540
transform 1 0 73032 0 1 60117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2261
timestamp 1704896540
transform 1 0 71264 0 1 56581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2262
timestamp 1704896540
transform 1 0 71264 0 1 56853
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2263
timestamp 1704896540
transform 1 0 71264 0 1 57805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2264
timestamp 1704896540
transform 1 0 71264 0 1 58077
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2265
timestamp 1704896540
transform 1 0 72352 0 1 56445
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2266
timestamp 1704896540
transform 1 0 72352 0 1 56173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2267
timestamp 1704896540
transform 1 0 73032 0 1 60933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2268
timestamp 1704896540
transform 1 0 73032 0 1 61205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2269
timestamp 1704896540
transform 1 0 72896 0 1 57397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2270
timestamp 1704896540
transform 1 0 72896 0 1 57669
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2271
timestamp 1704896540
transform 1 0 72896 0 1 58077
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2272
timestamp 1704896540
transform 1 0 72896 0 1 57805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2273
timestamp 1704896540
transform 1 0 72624 0 1 60933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2274
timestamp 1704896540
transform 1 0 72624 0 1 61205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2275
timestamp 1704896540
transform 1 0 71400 0 1 59709
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2276
timestamp 1704896540
transform 1 0 71400 0 1 59981
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2277
timestamp 1704896540
transform 1 0 71400 0 1 57397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2278
timestamp 1704896540
transform 1 0 72896 0 1 56853
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2279
timestamp 1704896540
transform 1 0 72896 0 1 56581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2280
timestamp 1704896540
transform 1 0 72896 0 1 56173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2281
timestamp 1704896540
transform 1 0 72896 0 1 56445
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2282
timestamp 1704896540
transform 1 0 72896 0 1 59709
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2283
timestamp 1704896540
transform 1 0 72896 0 1 59437
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2284
timestamp 1704896540
transform 1 0 71672 0 1 59709
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2285
timestamp 1704896540
transform 1 0 71672 0 1 59981
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2286
timestamp 1704896540
transform 1 0 71808 0 1 57669
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2287
timestamp 1704896540
transform 1 0 71808 0 1 57397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2288
timestamp 1704896540
transform 1 0 71400 0 1 57669
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2289
timestamp 1704896540
transform 1 0 71264 0 1 60797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2290
timestamp 1704896540
transform 1 0 71808 0 1 57261
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2291
timestamp 1704896540
transform 1 0 71808 0 1 56989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2292
timestamp 1704896540
transform 1 0 71264 0 1 60525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2293
timestamp 1704896540
transform 1 0 71264 0 1 60117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2294
timestamp 1704896540
transform 1 0 71808 0 1 60933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2295
timestamp 1704896540
transform 1 0 71808 0 1 61205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2296
timestamp 1704896540
transform 1 0 71264 0 1 60389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2297
timestamp 1704896540
transform 1 0 72352 0 1 58893
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2298
timestamp 1704896540
transform 1 0 71808 0 1 57805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2299
timestamp 1704896540
transform 1 0 71808 0 1 58077
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2300
timestamp 1704896540
transform 1 0 71808 0 1 59573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2301
timestamp 1704896540
transform 1 0 71808 0 1 59301
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2302
timestamp 1704896540
transform 1 0 71672 0 1 60797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2303
timestamp 1704896540
transform 1 0 71672 0 1 60525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2304
timestamp 1704896540
transform 1 0 71672 0 1 60117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2305
timestamp 1704896540
transform 1 0 71672 0 1 60389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2306
timestamp 1704896540
transform 1 0 72352 0 1 59165
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2307
timestamp 1704896540
transform 1 0 72216 0 1 60117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2308
timestamp 1704896540
transform 1 0 71672 0 1 55765
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2309
timestamp 1704896540
transform 1 0 71672 0 1 56037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2310
timestamp 1704896540
transform 1 0 72216 0 1 60389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2311
timestamp 1704896540
transform 1 0 72352 0 1 57669
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2312
timestamp 1704896540
transform 1 0 72352 0 1 57397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2313
timestamp 1704896540
transform 1 0 72080 0 1 56853
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2314
timestamp 1704896540
transform 1 0 71672 0 1 56853
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2315
timestamp 1704896540
transform 1 0 71672 0 1 56581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2316
timestamp 1704896540
transform 1 0 71672 0 1 56173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2317
timestamp 1704896540
transform 1 0 71672 0 1 56445
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2318
timestamp 1704896540
transform 1 0 72080 0 1 56581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2319
timestamp 1704896540
transform 1 0 72624 0 1 60117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2320
timestamp 1704896540
transform 1 0 72624 0 1 60389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2321
timestamp 1704896540
transform 1 0 71264 0 1 56037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2322
timestamp 1704896540
transform 1 0 71264 0 1 55765
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2323
timestamp 1704896540
transform 1 0 72488 0 1 56853
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2324
timestamp 1704896540
transform 1 0 71400 0 1 62429
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2325
timestamp 1704896540
transform 1 0 71400 0 1 62157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2326
timestamp 1704896540
transform 1 0 72352 0 1 65693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2327
timestamp 1704896540
transform 1 0 73032 0 1 63381
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2328
timestamp 1704896540
transform 1 0 73032 0 1 63653
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2329
timestamp 1704896540
transform 1 0 73032 0 1 65965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2330
timestamp 1704896540
transform 1 0 73032 0 1 65693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2331
timestamp 1704896540
transform 1 0 72896 0 1 65557
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2332
timestamp 1704896540
transform 1 0 72896 0 1 65285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2333
timestamp 1704896540
transform 1 0 73032 0 1 65149
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2334
timestamp 1704896540
transform 1 0 73032 0 1 64877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2335
timestamp 1704896540
transform 1 0 72896 0 1 62565
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2336
timestamp 1704896540
transform 1 0 72896 0 1 62837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2337
timestamp 1704896540
transform 1 0 72896 0 1 63245
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2338
timestamp 1704896540
transform 1 0 72896 0 1 62973
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2339
timestamp 1704896540
transform 1 0 72896 0 1 62429
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2340
timestamp 1704896540
transform 1 0 72896 0 1 62157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2341
timestamp 1704896540
transform 1 0 72896 0 1 61749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2342
timestamp 1704896540
transform 1 0 72896 0 1 62021
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2343
timestamp 1704896540
transform 1 0 73032 0 1 61613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2344
timestamp 1704896540
transform 1 0 73032 0 1 61341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2345
timestamp 1704896540
transform 1 0 72896 0 1 66509
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2346
timestamp 1704896540
transform 1 0 72896 0 1 66101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2347
timestamp 1704896540
transform 1 0 72896 0 1 66373
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2348
timestamp 1704896540
transform 1 0 72896 0 1 64333
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2349
timestamp 1704896540
transform 1 0 72896 0 1 64061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2350
timestamp 1704896540
transform 1 0 71672 0 1 64061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2351
timestamp 1704896540
transform 1 0 71672 0 1 64333
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2352
timestamp 1704896540
transform 1 0 71672 0 1 61749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2353
timestamp 1704896540
transform 1 0 71672 0 1 62021
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2354
timestamp 1704896540
transform 1 0 71808 0 1 61613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2355
timestamp 1704896540
transform 1 0 71808 0 1 61341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2356
timestamp 1704896540
transform 1 0 71672 0 1 62157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2357
timestamp 1704896540
transform 1 0 71672 0 1 62429
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2358
timestamp 1704896540
transform 1 0 71808 0 1 66373
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2359
timestamp 1704896540
transform 1 0 71808 0 1 66101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2360
timestamp 1704896540
transform 1 0 71672 0 1 65693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2361
timestamp 1704896540
transform 1 0 71672 0 1 65965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2362
timestamp 1704896540
transform 1 0 71672 0 1 63925
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2363
timestamp 1704896540
transform 1 0 71672 0 1 63653
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2364
timestamp 1704896540
transform 1 0 71672 0 1 64469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2365
timestamp 1704896540
transform 1 0 71672 0 1 64741
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2366
timestamp 1704896540
transform 1 0 71672 0 1 65557
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2367
timestamp 1704896540
transform 1 0 71672 0 1 65285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2368
timestamp 1704896540
transform 1 0 71808 0 1 64877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2369
timestamp 1704896540
transform 1 0 71808 0 1 65149
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2370
timestamp 1704896540
transform 1 0 72352 0 1 65965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2371
timestamp 1704896540
transform 1 0 72216 0 1 65965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2372
timestamp 1704896540
transform 1 0 72216 0 1 65693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2373
timestamp 1704896540
transform 1 0 72080 0 1 62973
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2374
timestamp 1704896540
transform 1 0 72080 0 1 63245
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2375
timestamp 1704896540
transform 1 0 72352 0 1 65149
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2376
timestamp 1704896540
transform 1 0 72352 0 1 64877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2377
timestamp 1704896540
transform 1 0 72216 0 1 64741
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2378
timestamp 1704896540
transform 1 0 72216 0 1 64469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2379
timestamp 1704896540
transform 1 0 72352 0 1 63925
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2380
timestamp 1704896540
transform 1 0 72352 0 1 63653
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2381
timestamp 1704896540
transform 1 0 72080 0 1 63653
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2382
timestamp 1704896540
transform 1 0 72080 0 1 63925
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2383
timestamp 1704896540
transform 1 0 72080 0 1 65557
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2384
timestamp 1704896540
transform 1 0 72080 0 1 65285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2385
timestamp 1704896540
transform 1 0 71264 0 1 61613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2386
timestamp 1704896540
transform 1 0 71400 0 1 62021
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2387
timestamp 1704896540
transform 1 0 71400 0 1 61749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2388
timestamp 1704896540
transform 1 0 71264 0 1 61341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2389
timestamp 1704896540
transform 1 0 72352 0 1 61341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2390
timestamp 1704896540
transform 1 0 72352 0 1 61613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2391
timestamp 1704896540
transform 1 0 72352 0 1 62021
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2392
timestamp 1704896540
transform 1 0 72352 0 1 61749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2393
timestamp 1704896540
transform 1 0 72216 0 1 61341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2394
timestamp 1704896540
transform 1 0 72216 0 1 61613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2395
timestamp 1704896540
transform 1 0 72080 0 1 61749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2396
timestamp 1704896540
transform 1 0 72080 0 1 62021
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2397
timestamp 1704896540
transform 1 0 71264 0 1 64741
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2398
timestamp 1704896540
transform 1 0 71264 0 1 64469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2399
timestamp 1704896540
transform 1 0 71400 0 1 64333
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2400
timestamp 1704896540
transform 1 0 71400 0 1 64061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2401
timestamp 1704896540
transform 1 0 71264 0 1 65693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2402
timestamp 1704896540
transform 1 0 71264 0 1 65965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2403
timestamp 1704896540
transform 1 0 71264 0 1 63925
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2404
timestamp 1704896540
transform 1 0 71264 0 1 63653
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2405
timestamp 1704896540
transform 1 0 72080 0 1 66645
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2406
timestamp 1704896540
transform 1 0 72080 0 1 66237
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2407
timestamp 1704896540
transform 1 0 71400 0 1 66101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2408
timestamp 1704896540
transform 1 0 71400 0 1 66373
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2409
timestamp 1704896540
transform 1 0 71400 0 1 64877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2410
timestamp 1704896540
transform 1 0 71400 0 1 65149
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2411
timestamp 1704896540
transform 1 0 71400 0 1 65557
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2412
timestamp 1704896540
transform 1 0 71400 0 1 65285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2413
timestamp 1704896540
transform 1 0 72488 0 1 62429
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2414
timestamp 1704896540
transform 1 0 72488 0 1 62157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2415
timestamp 1704896540
transform 1 0 72488 0 1 64061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2416
timestamp 1704896540
transform 1 0 72488 0 1 64333
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2417
timestamp 1704896540
transform 1 0 72624 0 1 64741
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2418
timestamp 1704896540
transform 1 0 72624 0 1 64469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2419
timestamp 1704896540
transform 1 0 72488 0 1 65557
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2420
timestamp 1704896540
transform 1 0 72488 0 1 65285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2421
timestamp 1704896540
transform 1 0 89760 0 1 59165
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2422
timestamp 1704896540
transform 1 0 89760 0 1 57397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2423
timestamp 1704896540
transform 1 0 89760 0 1 55765
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2424
timestamp 1704896540
transform 1 0 89760 0 1 60933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2425
timestamp 1704896540
transform 1 0 90440 0 1 64469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2426
timestamp 1704896540
transform 1 0 87720 0 1 64605
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2427
timestamp 1704896540
transform 1 0 87720 0 1 61885
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2428
timestamp 1704896540
transform 1 0 87584 0 1 64469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2429
timestamp 1704896540
transform 1 0 88459 0 1 62425
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2430
timestamp 1704896540
transform 1 0 89760 0 1 62565
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2431
timestamp 1704896540
transform 1 0 89760 0 1 64197
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2432
timestamp 1704896540
transform 1 0 89760 0 1 65829
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2433
timestamp 1704896540
transform 1 0 89080 0 1 62565
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2434
timestamp 1704896540
transform 1 0 89080 0 1 63109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2435
timestamp 1704896540
transform 1 0 66368 0 1 50461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2436
timestamp 1704896540
transform 1 0 66504 0 1 63517
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2437
timestamp 1704896540
transform 1 0 66504 0 1 63789
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2438
timestamp 1704896540
transform 1 0 66504 0 1 55085
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2439
timestamp 1704896540
transform 1 0 66504 0 1 54813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2440
timestamp 1704896540
transform 1 0 66504 0 1 54405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2441
timestamp 1704896540
transform 1 0 66504 0 1 54677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2442
timestamp 1704896540
transform 1 0 66504 0 1 50325
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2443
timestamp 1704896540
transform 1 0 66504 0 1 58621
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2444
timestamp 1704896540
transform 1 0 66368 0 1 59573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2445
timestamp 1704896540
transform 1 0 66368 0 1 59845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2446
timestamp 1704896540
transform 1 0 66504 0 1 58349
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2447
timestamp 1704896540
transform 1 0 66368 0 1 63381
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2448
timestamp 1704896540
transform 1 0 66504 0 1 65829
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2449
timestamp 1704896540
transform 1 0 66504 0 1 66101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2450
timestamp 1704896540
transform 1 0 66504 0 1 46381
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2451
timestamp 1704896540
transform 1 0 66504 0 1 46109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2452
timestamp 1704896540
transform 1 0 66504 0 1 66645
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2453
timestamp 1704896540
transform 1 0 66368 0 1 63109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2454
timestamp 1704896540
transform 1 0 66368 0 1 62701
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2455
timestamp 1704896540
transform 1 0 66368 0 1 62973
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2456
timestamp 1704896540
transform 1 0 66504 0 1 62701
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2457
timestamp 1704896540
transform 1 0 66504 0 1 62429
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2458
timestamp 1704896540
transform 1 0 66504 0 1 50733
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2459
timestamp 1704896540
transform 1 0 66368 0 1 51141
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2460
timestamp 1704896540
transform 1 0 66368 0 1 50869
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2461
timestamp 1704896540
transform 1 0 66368 0 1 46517
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2462
timestamp 1704896540
transform 1 0 66368 0 1 46789
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2463
timestamp 1704896540
transform 1 0 66368 0 1 59029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2464
timestamp 1704896540
transform 1 0 66368 0 1 58757
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2465
timestamp 1704896540
transform 1 0 66504 0 1 59165
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2466
timestamp 1704896540
transform 1 0 66504 0 1 59573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2467
timestamp 1704896540
transform 1 0 66368 0 1 50733
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2468
timestamp 1704896540
transform 1 0 58888 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2469
timestamp 1704896540
transform 1 0 63920 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2470
timestamp 1704896540
transform 1 0 63920 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2471
timestamp 1704896540
transform 1 0 63104 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2472
timestamp 1704896540
transform 1 0 66504 0 1 67869
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2473
timestamp 1704896540
transform 1 0 66504 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2474
timestamp 1704896540
transform 1 0 66504 0 1 70453
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2475
timestamp 1704896540
transform 1 0 66504 0 1 70045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2476
timestamp 1704896540
transform 1 0 66368 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2477
timestamp 1704896540
transform 1 0 66368 0 1 68549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2478
timestamp 1704896540
transform 1 0 66504 0 1 66917
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2479
timestamp 1704896540
transform 1 0 66504 0 1 67325
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2480
timestamp 1704896540
transform 1 0 66504 0 1 67053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2481
timestamp 1704896540
transform 1 0 66776 0 1 71133
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2482
timestamp 1704896540
transform 1 0 66776 0 1 73309
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2483
timestamp 1704896540
transform 1 0 60928 0 1 73581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2484
timestamp 1704896540
transform 1 0 60928 0 1 76029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2485
timestamp 1704896540
transform 1 0 60792 0 1 76029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2486
timestamp 1704896540
transform 1 0 60928 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2487
timestamp 1704896540
transform 1 0 63104 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2488
timestamp 1704896540
transform 1 0 62696 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2489
timestamp 1704896540
transform 1 0 62696 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2490
timestamp 1704896540
transform 1 0 58208 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2491
timestamp 1704896540
transform 1 0 58208 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2492
timestamp 1704896540
transform 1 0 62016 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2493
timestamp 1704896540
transform 1 0 62016 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2494
timestamp 1704896540
transform 1 0 61472 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2495
timestamp 1704896540
transform 1 0 61472 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2496
timestamp 1704896540
transform 1 0 57664 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2497
timestamp 1704896540
transform 1 0 57664 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2498
timestamp 1704896540
transform 1 0 61472 0 1 71949
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2499
timestamp 1704896540
transform 1 0 61472 0 1 76573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2500
timestamp 1704896540
transform 1 0 60928 0 1 77525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2501
timestamp 1704896540
transform 1 0 60928 0 1 76845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2502
timestamp 1704896540
transform 1 0 60656 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2503
timestamp 1704896540
transform 1 0 60656 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2504
timestamp 1704896540
transform 1 0 56984 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2505
timestamp 1704896540
transform 1 0 56984 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2506
timestamp 1704896540
transform 1 0 67728 0 1 70997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2507
timestamp 1704896540
transform 1 0 67728 0 1 71269
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2508
timestamp 1704896540
transform 1 0 65688 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2509
timestamp 1704896540
transform 1 0 65688 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2510
timestamp 1704896540
transform 1 0 65144 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2511
timestamp 1704896540
transform 1 0 65144 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2512
timestamp 1704896540
transform 1 0 64464 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2513
timestamp 1704896540
transform 1 0 64464 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2514
timestamp 1704896540
transform 1 0 58888 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2515
timestamp 1704896540
transform 1 0 56168 0 1 76029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2516
timestamp 1704896540
transform 1 0 56032 0 1 76029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2517
timestamp 1704896540
transform 1 0 56032 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2518
timestamp 1704896540
transform 1 0 51000 0 1 73581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2519
timestamp 1704896540
transform 1 0 51000 0 1 76029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2520
timestamp 1704896540
transform 1 0 50864 0 1 76029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2521
timestamp 1704896540
transform 1 0 50864 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2522
timestamp 1704896540
transform 1 0 46104 0 1 73581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2523
timestamp 1704896540
transform 1 0 46104 0 1 76029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2524
timestamp 1704896540
transform 1 0 45968 0 1 76029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2525
timestamp 1704896540
transform 1 0 45968 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2526
timestamp 1704896540
transform 1 0 50184 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2527
timestamp 1704896540
transform 1 0 49368 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2528
timestamp 1704896540
transform 1 0 49368 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2529
timestamp 1704896540
transform 1 0 45696 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2530
timestamp 1704896540
transform 1 0 45696 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2531
timestamp 1704896540
transform 1 0 48960 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2532
timestamp 1704896540
transform 1 0 48960 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2533
timestamp 1704896540
transform 1 0 56440 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2534
timestamp 1704896540
transform 1 0 56440 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2535
timestamp 1704896540
transform 1 0 55896 0 1 77525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2536
timestamp 1704896540
transform 1 0 55896 0 1 76845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2537
timestamp 1704896540
transform 1 0 47736 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2538
timestamp 1704896540
transform 1 0 47736 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2539
timestamp 1704896540
transform 1 0 55760 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2540
timestamp 1704896540
transform 1 0 55760 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2541
timestamp 1704896540
transform 1 0 55352 0 1 76573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2542
timestamp 1704896540
transform 1 0 55352 0 1 71949
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2543
timestamp 1704896540
transform 1 0 45696 0 1 76573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2544
timestamp 1704896540
transform 1 0 45696 0 1 71949
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2545
timestamp 1704896540
transform 1 0 54128 0 1 71269
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2546
timestamp 1704896540
transform 1 0 54128 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2547
timestamp 1704896540
transform 1 0 52632 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2548
timestamp 1704896540
transform 1 0 52632 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2549
timestamp 1704896540
transform 1 0 46920 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2550
timestamp 1704896540
transform 1 0 46920 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2551
timestamp 1704896540
transform 1 0 51952 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2552
timestamp 1704896540
transform 1 0 51952 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2553
timestamp 1704896540
transform 1 0 51408 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2554
timestamp 1704896540
transform 1 0 51408 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2555
timestamp 1704896540
transform 1 0 50728 0 1 77525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2556
timestamp 1704896540
transform 1 0 50728 0 1 76845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2557
timestamp 1704896540
transform 1 0 45832 0 1 77525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2558
timestamp 1704896540
transform 1 0 45832 0 1 76845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2559
timestamp 1704896540
transform 1 0 50728 0 1 76573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2560
timestamp 1704896540
transform 1 0 50728 0 1 71949
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2561
timestamp 1704896540
transform 1 0 50184 0 1 71813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2562
timestamp 1704896540
transform 1 0 56168 0 1 73581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2563
timestamp 1704896540
transform 1 0 55624 0 1 77933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2564
timestamp 1704896540
transform 1 0 50456 0 1 77933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2565
timestamp 1704896540
transform 1 0 45560 0 1 77933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2566
timestamp 1704896540
transform 1 0 55896 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2567
timestamp 1704896540
transform 1 0 55896 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2568
timestamp 1704896540
transform 1 0 54264 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2569
timestamp 1704896540
transform 1 0 54264 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2570
timestamp 1704896540
transform 1 0 52496 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2571
timestamp 1704896540
transform 1 0 52496 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2572
timestamp 1704896540
transform 1 0 50864 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2573
timestamp 1704896540
transform 1 0 50864 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2574
timestamp 1704896540
transform 1 0 49096 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2575
timestamp 1704896540
transform 1 0 49096 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2576
timestamp 1704896540
transform 1 0 47328 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2577
timestamp 1704896540
transform 1 0 47328 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2578
timestamp 1704896540
transform 1 0 45832 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2579
timestamp 1704896540
transform 1 0 45832 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2580
timestamp 1704896540
transform 1 0 60656 0 1 77933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2581
timestamp 1704896540
transform 1 0 57392 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2582
timestamp 1704896540
transform 1 0 57392 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2583
timestamp 1704896540
transform 1 0 67592 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2584
timestamp 1704896540
transform 1 0 67592 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2585
timestamp 1704896540
transform 1 0 65960 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2586
timestamp 1704896540
transform 1 0 65960 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2587
timestamp 1704896540
transform 1 0 64328 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2588
timestamp 1704896540
transform 1 0 64328 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2589
timestamp 1704896540
transform 1 0 62560 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2590
timestamp 1704896540
transform 1 0 62560 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2591
timestamp 1704896540
transform 1 0 60928 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2592
timestamp 1704896540
transform 1 0 60928 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2593
timestamp 1704896540
transform 1 0 59296 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2594
timestamp 1704896540
transform 1 0 59296 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2595
timestamp 1704896540
transform 1 0 89760 0 1 67733
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2596
timestamp 1704896540
transform 1 0 90440 0 1 70181
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2597
timestamp 1704896540
transform 1 0 87720 0 1 67325
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2598
timestamp 1704896540
transform 1 0 89760 0 1 69365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2599
timestamp 1704896540
transform 1 0 89080 0 1 69229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2600
timestamp 1704896540
transform 1 0 89080 0 1 68957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2601
timestamp 1704896540
transform 1 0 89080 0 1 71677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2602
timestamp 1704896540
transform 1 0 89760 0 1 70861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2603
timestamp 1704896540
transform 1 0 79560 0 1 73173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2604
timestamp 1704896540
transform 1 0 79560 0 1 76029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2605
timestamp 1704896540
transform 1 0 79560 0 1 75757
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2606
timestamp 1704896540
transform 1 0 90440 0 1 73173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2607
timestamp 1704896540
transform 1 0 88459 0 1 72660
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2608
timestamp 1704896540
transform 1 0 89760 0 1 75893
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2609
timestamp 1704896540
transform 1 0 89760 0 1 77525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2610
timestamp 1704896540
transform 1 0 89760 0 1 74397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2611
timestamp 1704896540
transform 1 0 89760 0 1 72493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2612
timestamp 1704896540
transform 1 0 89080 0 1 72493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2613
timestamp 1704896540
transform 1 0 72760 0 1 70997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2614
timestamp 1704896540
transform 1 0 71400 0 1 70453
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2615
timestamp 1704896540
transform 1 0 71400 0 1 70861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2616
timestamp 1704896540
transform 1 0 79288 0 1 77389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2617
timestamp 1704896540
transform 1 0 72896 0 1 74805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2618
timestamp 1704896540
transform 1 0 79288 0 1 74397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2619
timestamp 1704896540
transform 1 0 79288 0 1 71677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2620
timestamp 1704896540
transform 1 0 72896 0 1 77525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2621
timestamp 1704896540
transform 1 0 71128 0 1 70453
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2622
timestamp 1704896540
transform 1 0 71128 0 1 70861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2623
timestamp 1704896540
transform 1 0 72624 0 1 69637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2624
timestamp 1704896540
transform 1 0 79288 0 1 77253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2625
timestamp 1704896540
transform 1 0 79288 0 1 76165
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2626
timestamp 1704896540
transform 1 0 72624 0 1 69909
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2627
timestamp 1704896540
transform 1 0 74120 0 1 76165
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2628
timestamp 1704896540
transform 1 0 72624 0 1 67189
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2629
timestamp 1704896540
transform 1 0 72624 0 1 66917
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2630
timestamp 1704896540
transform 1 0 72488 0 1 68413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2631
timestamp 1704896540
transform 1 0 72488 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2632
timestamp 1704896540
transform 1 0 74120 0 1 73173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2633
timestamp 1704896540
transform 1 0 74120 0 1 70453
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2634
timestamp 1704896540
transform 1 0 73032 0 1 70045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2635
timestamp 1704896540
transform 1 0 73032 0 1 70317
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2636
timestamp 1704896540
transform 1 0 73032 0 1 69093
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2637
timestamp 1704896540
transform 1 0 73032 0 1 68821
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2638
timestamp 1704896540
transform 1 0 72896 0 1 69909
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2639
timestamp 1704896540
transform 1 0 72896 0 1 69637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2640
timestamp 1704896540
transform 1 0 72896 0 1 69229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2641
timestamp 1704896540
transform 1 0 72896 0 1 69501
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2642
timestamp 1704896540
transform 1 0 72896 0 1 67597
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2643
timestamp 1704896540
transform 1 0 72896 0 1 67325
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2644
timestamp 1704896540
transform 1 0 72896 0 1 66917
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2645
timestamp 1704896540
transform 1 0 72896 0 1 67189
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2646
timestamp 1704896540
transform 1 0 72624 0 1 73445
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2647
timestamp 1704896540
transform 1 0 72624 0 1 76029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2648
timestamp 1704896540
transform 1 0 71808 0 1 69637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2649
timestamp 1704896540
transform 1 0 71808 0 1 69909
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2650
timestamp 1704896540
transform 1 0 71672 0 1 67869
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2651
timestamp 1704896540
transform 1 0 71672 0 1 67597
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2652
timestamp 1704896540
transform 1 0 71672 0 1 68821
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2653
timestamp 1704896540
transform 1 0 71672 0 1 69093
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2654
timestamp 1704896540
transform 1 0 71672 0 1 69501
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2655
timestamp 1704896540
transform 1 0 71672 0 1 69229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2656
timestamp 1704896540
transform 1 0 71808 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2657
timestamp 1704896540
transform 1 0 71808 0 1 68413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2658
timestamp 1704896540
transform 1 0 71808 0 1 68005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2659
timestamp 1704896540
transform 1 0 71808 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2660
timestamp 1704896540
transform 1 0 71672 0 1 70045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2661
timestamp 1704896540
transform 1 0 71672 0 1 70317
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2662
timestamp 1704896540
transform 1 0 72352 0 1 68821
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2663
timestamp 1704896540
transform 1 0 72352 0 1 69093
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2664
timestamp 1704896540
transform 1 0 72216 0 1 69501
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2665
timestamp 1704896540
transform 1 0 72216 0 1 69229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2666
timestamp 1704896540
transform 1 0 72080 0 1 66917
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2667
timestamp 1704896540
transform 1 0 72080 0 1 67189
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2668
timestamp 1704896540
transform 1 0 72352 0 1 70317
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2669
timestamp 1704896540
transform 1 0 72352 0 1 70045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2670
timestamp 1704896540
transform 1 0 72216 0 1 70317
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2671
timestamp 1704896540
transform 1 0 72216 0 1 70045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2672
timestamp 1704896540
transform 1 0 72080 0 1 68413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2673
timestamp 1704896540
transform 1 0 72080 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2674
timestamp 1704896540
transform 1 0 72352 0 1 67597
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2675
timestamp 1704896540
transform 1 0 72352 0 1 67869
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2676
timestamp 1704896540
transform 1 0 71264 0 1 70317
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2677
timestamp 1704896540
transform 1 0 71264 0 1 70045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2678
timestamp 1704896540
transform 1 0 71264 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2679
timestamp 1704896540
transform 1 0 71264 0 1 68005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2680
timestamp 1704896540
transform 1 0 71264 0 1 67597
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2681
timestamp 1704896540
transform 1 0 71264 0 1 67869
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2682
timestamp 1704896540
transform 1 0 71400 0 1 69229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2683
timestamp 1704896540
transform 1 0 71400 0 1 69501
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2684
timestamp 1704896540
transform 1 0 71400 0 1 69909
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2685
timestamp 1704896540
transform 1 0 71400 0 1 69637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2686
timestamp 1704896540
transform 1 0 71264 0 1 69093
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2687
timestamp 1704896540
transform 1 0 71264 0 1 68821
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2688
timestamp 1704896540
transform 1 0 71400 0 1 68413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2689
timestamp 1704896540
transform 1 0 79288 0 1 75757
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2690
timestamp 1704896540
transform 1 0 79288 0 1 74805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2691
timestamp 1704896540
transform 1 0 74256 0 1 77661
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2692
timestamp 1704896540
transform 1 0 71400 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2693
timestamp 1704896540
transform 1 0 72760 0 1 74669
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2694
timestamp 1704896540
transform 1 0 74120 0 1 83237
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2695
timestamp 1704896540
transform 1 0 74256 0 1 80245
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2696
timestamp 1704896540
transform 1 0 74256 0 1 83101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2697
timestamp 1704896540
transform 1 0 79288 0 1 80109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2698
timestamp 1704896540
transform 1 0 74256 0 1 80381
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2699
timestamp 1704896540
transform 1 0 74392 0 1 81877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2700
timestamp 1704896540
transform 1 0 74120 0 1 81741
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2701
timestamp 1704896540
transform 1 0 74120 0 1 79021
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2702
timestamp 1704896540
transform 1 0 74120 0 1 78885
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2703
timestamp 1704896540
transform 1 0 72624 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2704
timestamp 1704896540
transform 1 0 72624 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2705
timestamp 1704896540
transform 1 0 70856 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2706
timestamp 1704896540
transform 1 0 70856 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2707
timestamp 1704896540
transform 1 0 69360 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2708
timestamp 1704896540
transform 1 0 69360 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2709
timestamp 1704896540
transform 1 0 74392 0 1 84597
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2710
timestamp 1704896540
transform 1 0 73984 0 1 88677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2711
timestamp 1704896540
transform 1 0 73984 0 1 86909
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2712
timestamp 1704896540
transform 1 0 74256 0 1 84733
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2713
timestamp 1704896540
transform 1 0 74256 0 1 86773
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2714
timestamp 1704896540
transform 1 0 77656 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2715
timestamp 1704896540
transform 1 0 77656 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2716
timestamp 1704896540
transform 1 0 76024 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2717
timestamp 1704896540
transform 1 0 76024 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2718
timestamp 1704896540
transform 1 0 76296 0 1 85413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2719
timestamp 1704896540
transform 1 0 76296 0 1 87317
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2720
timestamp 1704896540
transform 1 0 74256 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2721
timestamp 1704896540
transform 1 0 74256 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2722
timestamp 1704896540
transform 1 0 74120 0 1 85277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2723
timestamp 1704896540
transform 1 0 74528 0 1 86229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2724
timestamp 1704896540
transform 1 0 75616 0 1 86229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2725
timestamp 1704896540
transform 1 0 76704 0 1 86229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2726
timestamp 1704896540
transform 1 0 90440 0 1 80109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2727
timestamp 1704896540
transform 1 0 89760 0 1 79293
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2728
timestamp 1704896540
transform 1 0 89760 0 1 80925
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2729
timestamp 1704896540
transform 1 0 89760 0 1 82693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2730
timestamp 1704896540
transform 1 0 89080 0 1 79293
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2731
timestamp 1704896540
transform 1 0 89080 0 1 78749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2732
timestamp 1704896540
transform 1 0 87992 0 1 79157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2733
timestamp 1704896540
transform 1 0 87992 0 1 79429
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2734
timestamp 1704896540
transform 1 0 79560 0 1 78613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2735
timestamp 1704896540
transform 1 0 84320 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2736
timestamp 1704896540
transform 1 0 84320 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2737
timestamp 1704896540
transform 1 0 82552 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2738
timestamp 1704896540
transform 1 0 82552 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2739
timestamp 1704896540
transform 1 0 81056 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2740
timestamp 1704896540
transform 1 0 81056 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2741
timestamp 1704896540
transform 1 0 89760 0 1 85957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2742
timestamp 1704896540
transform 1 0 89760 0 1 84325
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2743
timestamp 1704896540
transform 1 0 87856 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2744
timestamp 1704896540
transform 1 0 87856 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2745
timestamp 1704896540
transform 1 0 86088 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2746
timestamp 1704896540
transform 1 0 86088 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2747
timestamp 1704896540
transform 1 0 79424 0 1 77253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2748
timestamp 1704896540
transform 1 0 79424 0 1 74533
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2749
timestamp 1704896540
transform 1 0 79424 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2750
timestamp 1704896540
transform 1 0 79424 0 1 87589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2751
timestamp 1704896540
transform 1 0 72896 0 1 66781
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2752
timestamp 1704896540
transform 1 0 72896 0 1 44613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2753
timestamp 1704896540
transform 1 0 71808 0 1 44613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2754
timestamp 1704896540
transform 1 0 19176 0 1 44613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2755
timestamp 1704896540
transform 1 0 17816 0 1 44613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2756
timestamp 1704896540
transform 1 0 72352 0 1 44613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2757
timestamp 1704896540
transform 1 0 72080 0 1 44613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2758
timestamp 1704896540
transform 1 0 71400 0 1 44613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2759
timestamp 1704896540
transform 1 0 19584 0 1 44613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_33_2760
timestamp 1704896540
transform 1 0 18632 0 1 44613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_38  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_38_0
timestamp 1704896540
transform 1 0 89148 0 1 1672
box 0 0 192 192
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_38  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_38_1
timestamp 1704896540
transform 1 0 1650 0 1 1672
box 0 0 192 192
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_38  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_38_2
timestamp 1704896540
transform 1 0 1650 0 1 87400
box 0 0 192 192
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_38  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_38_3
timestamp 1704896540
transform 1 0 89148 0 1 87400
box 0 0 192 192
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_0
timestamp 1704896540
transform 1 0 90712 0 1 277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_1
timestamp 1704896540
transform 1 0 90032 0 1 957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_2
timestamp 1704896540
transform 1 0 90576 0 1 413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_3
timestamp 1704896540
transform 1 0 90440 0 1 277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_4
timestamp 1704896540
transform 1 0 90440 0 1 413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_5
timestamp 1704896540
transform 1 0 90440 0 1 549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_6
timestamp 1704896540
transform 1 0 90576 0 1 277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_7
timestamp 1704896540
transform 1 0 90712 0 1 549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_8
timestamp 1704896540
transform 1 0 90712 0 1 413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_9
timestamp 1704896540
transform 1 0 89760 0 1 1093
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_10
timestamp 1704896540
transform 1 0 90576 0 1 549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_11
timestamp 1704896540
transform 1 0 89896 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_12
timestamp 1704896540
transform 1 0 90032 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_13
timestamp 1704896540
transform 1 0 89760 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_14
timestamp 1704896540
transform 1 0 89896 0 1 957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_15
timestamp 1704896540
transform 1 0 89896 0 1 1093
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_16
timestamp 1704896540
transform 1 0 89760 0 1 957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_17
timestamp 1704896540
transform 1 0 90032 0 1 1093
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_18
timestamp 1704896540
transform 1 0 544 0 1 549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_19
timestamp 1704896540
transform 1 0 1088 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_20
timestamp 1704896540
transform 1 0 952 0 1 957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_21
timestamp 1704896540
transform 1 0 1224 0 1 957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_22
timestamp 1704896540
transform 1 0 1224 0 1 1093
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_23
timestamp 1704896540
transform 1 0 1088 0 1 957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_24
timestamp 1704896540
transform 1 0 272 0 1 549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_25
timestamp 1704896540
transform 1 0 272 0 1 413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_26
timestamp 1704896540
transform 1 0 408 0 1 549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_27
timestamp 1704896540
transform 1 0 544 0 1 277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_28
timestamp 1704896540
transform 1 0 408 0 1 413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_29
timestamp 1704896540
transform 1 0 1224 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_30
timestamp 1704896540
transform 1 0 952 0 1 1093
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_31
timestamp 1704896540
transform 1 0 272 0 1 277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_32
timestamp 1704896540
transform 1 0 952 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_33
timestamp 1704896540
transform 1 0 1088 0 1 1093
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_34
timestamp 1704896540
transform 1 0 544 0 1 413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_35
timestamp 1704896540
transform 1 0 408 0 1 277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_36
timestamp 1704896540
transform 1 0 952 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_37
timestamp 1704896540
transform 1 0 1224 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_38
timestamp 1704896540
transform 1 0 1224 0 1 88133
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_39
timestamp 1704896540
transform 1 0 1088 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_40
timestamp 1704896540
transform 1 0 952 0 1 88269
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_41
timestamp 1704896540
transform 1 0 1088 0 1 88133
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_42
timestamp 1704896540
transform 1 0 1224 0 1 88269
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_43
timestamp 1704896540
transform 1 0 952 0 1 88133
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_44
timestamp 1704896540
transform 1 0 1088 0 1 88269
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_45
timestamp 1704896540
transform 1 0 408 0 1 88813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_46
timestamp 1704896540
transform 1 0 544 0 1 88677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_47
timestamp 1704896540
transform 1 0 408 0 1 88949
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_48
timestamp 1704896540
transform 1 0 272 0 1 88677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_49
timestamp 1704896540
transform 1 0 408 0 1 88677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_50
timestamp 1704896540
transform 1 0 544 0 1 88813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_51
timestamp 1704896540
transform 1 0 272 0 1 88949
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_52
timestamp 1704896540
transform 1 0 272 0 1 88813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_53
timestamp 1704896540
transform 1 0 544 0 1 88949
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_54
timestamp 1704896540
transform 1 0 90576 0 1 88813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_55
timestamp 1704896540
transform 1 0 90440 0 1 88949
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_56
timestamp 1704896540
transform 1 0 90712 0 1 88813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_57
timestamp 1704896540
transform 1 0 90712 0 1 88949
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_58
timestamp 1704896540
transform 1 0 90440 0 1 88813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_59
timestamp 1704896540
transform 1 0 90576 0 1 88677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_60
timestamp 1704896540
transform 1 0 90712 0 1 88677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_61
timestamp 1704896540
transform 1 0 90576 0 1 88949
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_62
timestamp 1704896540
transform 1 0 90440 0 1 88677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_63
timestamp 1704896540
transform 1 0 89760 0 1 88133
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_64
timestamp 1704896540
transform 1 0 89896 0 1 88269
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_65
timestamp 1704896540
transform 1 0 90032 0 1 88269
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_66
timestamp 1704896540
transform 1 0 89760 0 1 88269
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_67
timestamp 1704896540
transform 1 0 89896 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_68
timestamp 1704896540
transform 1 0 89896 0 1 88133
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_69
timestamp 1704896540
transform 1 0 89760 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_70
timestamp 1704896540
transform 1 0 90032 0 1 88133
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_39_71
timestamp 1704896540
transform 1 0 90032 0 1 87997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_control_logic_r  sky130_sram_1kbyte_1rw1r_8x1024_8_control_logic_r_0
timestamp 1704896540
transform -1 0 88454 0 -1 80171
box -75 -49 9082 18431
use sky130_sram_1kbyte_1rw1r_8x1024_8_control_logic_rw  sky130_sram_1kbyte_1rw1r_8x1024_8_control_logic_rw_0
timestamp 1704896540
transform 1 0 2536 0 1 7987
box -75 -49 9166 18431
use sky130_sram_1kbyte_1rw1r_8x1024_8_cr_3  sky130_sram_1kbyte_1rw1r_8x1024_8_cr_3_0
timestamp 1704896540
transform 1 0 11870 0 1 6294
box 2083 -3207 4613 3549
use sky130_sram_1kbyte_1rw1r_8x1024_8_cr_4  sky130_sram_1kbyte_1rw1r_8x1024_8_cr_4_0
timestamp 1704896540
transform 1 0 11870 0 1 6294
box 5544 -3230 48961 4461
use sky130_sram_1kbyte_1rw1r_8x1024_8_cr_5  sky130_sram_1kbyte_1rw1r_8x1024_8_cr_5_0
timestamp 1704896540
transform 1 0 11870 0 1 6294
box 61683 74849 64083 79883
use sky130_sram_1kbyte_1rw1r_8x1024_8_data_dff  sky130_sram_1kbyte_1rw1r_8x1024_8_data_dff_0
timestamp 1704896540
transform 1 0 17542 0 1 2440
box -36 -49 9380 1467
use sky130_sram_1kbyte_1rw1r_8x1024_8_row_addr_dff  sky130_sram_1kbyte_1rw1r_8x1024_8_row_addr_dff_0
timestamp 1704896540
transform -1 0 80540 0 -1 20213
box -36 -49 1204 9951
use sky130_sram_1kbyte_1rw1r_8x1024_8_row_addr_dff  sky130_sram_1kbyte_1rw1r_8x1024_8_row_addr_dff_1
timestamp 1704896540
transform 1 0 10534 0 1 28113
box -36 -49 1204 9951
use sky130_sram_1kbyte_1rw1r_8x1024_8_wmask_dff  sky130_sram_1kbyte_1rw1r_8x1024_8_wmask_dff_0
timestamp 1704896540
transform 1 0 16374 0 1 2440
box -36 -49 1204 1467
<< labels >>
rlabel metal3 s 0 8568 212 8644 4 csb0
port 29 nsew default input
rlabel metal3 s 0 10200 212 10276 4 web0
port 31 nsew default input
rlabel metal3 s 0 8296 212 8372 4 clk0
port 32 nsew default input
rlabel metal3 s 0 28560 212 28636 4 addr0[3]
port 15 nsew default input
rlabel metal3 s 0 30192 212 30268 4 addr0[4]
port 14 nsew default input
rlabel metal3 s 0 31552 212 31628 4 addr0[5]
port 13 nsew default input
rlabel metal3 s 0 33184 212 33260 4 addr0[6]
port 12 nsew default input
rlabel metal3 s 0 34272 212 34348 4 addr0[7]
port 11 nsew default input
rlabel metal3 s 0 35904 212 35980 4 addr0[8]
port 10 nsew default input
rlabel metal3 s 0 36992 212 37068 4 addr0[9]
port 9 nsew default input
rlabel metal3 s 90848 79696 91060 79772 4 csb1
port 30 nsew default input
rlabel metal3 s 90848 79152 91060 79228 4 clk1
port 33 nsew default input
rlabel metal3 s 90848 19720 91060 19796 4 addr1[3]
port 25 nsew default input
rlabel metal3 s 90848 17952 91060 18028 4 addr1[4]
port 24 nsew default input
rlabel metal3 s 90848 16864 91060 16940 4 addr1[5]
port 23 nsew default input
rlabel metal3 s 90848 15096 91060 15172 4 addr1[6]
port 22 nsew default input
rlabel metal3 s 90848 14008 91060 14084 4 addr1[7]
port 21 nsew default input
rlabel metal3 s 90848 12376 91060 12452 4 addr1[8]
port 20 nsew default input
rlabel metal3 s 90848 11016 91060 11092 4 addr1[9]
port 19 nsew default input
rlabel metal3 s 952 87992 90108 88340 4 vccd1
port 51 nsew power bidirectional abutment
rlabel metal3 s 952 952 90108 1300 4 vccd1
port 51 nsew power bidirectional abutment
rlabel metal3 s 272 272 90788 620 4 vssd1
port 52 nsew ground bidirectional abutment
rlabel metal3 s 272 88672 90788 89020 4 vssd1
port 52 nsew ground bidirectional abutment
rlabel metal4 s 17680 0 17756 212 4 din0[0]
port 8 nsew default input
rlabel metal4 s 18904 0 18980 212 4 din0[1]
port 7 nsew default input
rlabel metal4 s 19992 0 20068 212 4 din0[2]
port 6 nsew default input
rlabel metal4 s 21080 0 21156 212 4 din0[3]
port 5 nsew default input
rlabel metal4 s 22304 0 22380 212 4 din0[4]
port 4 nsew default input
rlabel metal4 s 23392 0 23468 212 4 din0[5]
port 3 nsew default input
rlabel metal4 s 24752 0 24828 212 4 din0[6]
port 2 nsew default input
rlabel metal4 s 25704 0 25780 212 4 din0[7]
port 1 nsew default input
rlabel metal4 s 25296 0 25372 212 4 dout0[0]
port 42 nsew default output
rlabel metal4 s 30464 0 30540 212 4 dout0[1]
port 41 nsew default output
rlabel metal4 s 35496 0 35572 212 4 dout0[2]
port 40 nsew default output
rlabel metal4 s 40528 0 40604 212 4 dout0[3]
port 39 nsew default output
rlabel metal4 s 45560 0 45636 212 4 dout0[4]
port 38 nsew default output
rlabel metal4 s 50456 0 50532 212 4 dout0[5]
port 37 nsew default output
rlabel metal4 s 55488 0 55564 212 4 dout0[6]
port 36 nsew default output
rlabel metal4 s 60520 0 60596 212 4 dout0[7]
port 35 nsew default output
rlabel metal4 s 12920 0 12996 212 4 addr0[0]
port 18 nsew default input
rlabel metal4 s 14280 0 14356 212 4 addr0[1]
port 17 nsew default input
rlabel metal4 s 15368 0 15444 212 4 addr0[2]
port 16 nsew default input
rlabel metal4 s 16456 0 16532 212 4 wmask0[0]
port 34 nsew default input
rlabel metal4 s 25568 89080 25644 89292 4 dout1[0]
port 50 nsew default output
rlabel metal4 s 30600 89080 30676 89292 4 dout1[1]
port 49 nsew default output
rlabel metal4 s 35632 89080 35708 89292 4 dout1[2]
port 48 nsew default output
rlabel metal4 s 40664 89080 40740 89292 4 dout1[3]
port 47 nsew default output
rlabel metal4 s 45560 89080 45636 89292 4 dout1[4]
port 46 nsew default output
rlabel metal4 s 50456 89080 50532 89292 4 dout1[5]
port 45 nsew default output
rlabel metal4 s 55624 89080 55700 89292 4 dout1[6]
port 44 nsew default output
rlabel metal4 s 60656 89080 60732 89292 4 dout1[7]
port 43 nsew default output
rlabel metal4 s 76704 89080 76780 89292 4 addr1[0]
port 28 nsew default input
rlabel metal4 s 75616 89080 75692 89292 4 addr1[1]
port 27 nsew default input
rlabel metal4 s 74528 89080 74604 89292 4 addr1[2]
port 26 nsew default input
rlabel metal4 s 89760 952 90108 88340 4 vccd1
port 51 nsew power bidirectional abutment
rlabel metal4 s 952 952 1300 88340 4 vccd1
port 51 nsew power bidirectional abutment
rlabel metal4 s 272 272 620 89020 4 vssd1
port 52 nsew ground bidirectional abutment
rlabel metal4 s 90440 272 90788 89020 4 vssd1
port 52 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 91060 89292
string GDS_END 9277678
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_8x1024_8.gds
string GDS_START 7724596
string LEFclass BLOCK
string LEFsymmetry X Y R90
<< end >>
