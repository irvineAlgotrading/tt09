magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -119 -66 239 1066
<< mvpmos >>
rect 0 0 120 1000
<< mvpdiff >>
rect -50 0 0 1000
rect 120 0 170 1000
<< poly >>
rect 0 1000 120 1026
rect 0 -26 120 0
<< locali >>
rect -45 -4 -11 946
rect 131 -4 165 946
use hvDFL1sd_CDNS_52468879185112  hvDFL1sd_CDNS_52468879185112_0
timestamp 1704896540
transform -1 0 0 0 1 0
box -36 -36 89 1036
use hvDFL1sd_CDNS_52468879185112  hvDFL1sd_CDNS_52468879185112_1
timestamp 1704896540
transform 1 0 120 0 1 0
box -36 -36 89 1036
<< labels >>
flabel comment s -28 471 -28 471 0 FreeSans 300 0 0 0 S
flabel comment s 148 471 148 471 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 87728044
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 87727026
<< end >>
