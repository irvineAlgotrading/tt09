magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< pwell >>
rect -26 -26 82 1426
<< ndiff >>
rect 0 1338 56 1400
rect 0 1304 11 1338
rect 45 1304 56 1338
rect 0 1270 56 1304
rect 0 1236 11 1270
rect 45 1236 56 1270
rect 0 1202 56 1236
rect 0 1168 11 1202
rect 45 1168 56 1202
rect 0 1134 56 1168
rect 0 1100 11 1134
rect 45 1100 56 1134
rect 0 1066 56 1100
rect 0 1032 11 1066
rect 45 1032 56 1066
rect 0 998 56 1032
rect 0 964 11 998
rect 45 964 56 998
rect 0 930 56 964
rect 0 896 11 930
rect 45 896 56 930
rect 0 862 56 896
rect 0 828 11 862
rect 45 828 56 862
rect 0 794 56 828
rect 0 760 11 794
rect 45 760 56 794
rect 0 726 56 760
rect 0 692 11 726
rect 45 692 56 726
rect 0 658 56 692
rect 0 624 11 658
rect 45 624 56 658
rect 0 590 56 624
rect 0 556 11 590
rect 45 556 56 590
rect 0 522 56 556
rect 0 488 11 522
rect 45 488 56 522
rect 0 454 56 488
rect 0 420 11 454
rect 45 420 56 454
rect 0 386 56 420
rect 0 352 11 386
rect 45 352 56 386
rect 0 318 56 352
rect 0 284 11 318
rect 45 284 56 318
rect 0 250 56 284
rect 0 216 11 250
rect 45 216 56 250
rect 0 182 56 216
rect 0 148 11 182
rect 45 148 56 182
rect 0 114 56 148
rect 0 80 11 114
rect 45 80 56 114
rect 0 46 56 80
rect 0 12 11 46
rect 45 12 56 46
rect 0 0 56 12
<< ndiffc >>
rect 11 1304 45 1338
rect 11 1236 45 1270
rect 11 1168 45 1202
rect 11 1100 45 1134
rect 11 1032 45 1066
rect 11 964 45 998
rect 11 896 45 930
rect 11 828 45 862
rect 11 760 45 794
rect 11 692 45 726
rect 11 624 45 658
rect 11 556 45 590
rect 11 488 45 522
rect 11 420 45 454
rect 11 352 45 386
rect 11 284 45 318
rect 11 216 45 250
rect 11 148 45 182
rect 11 80 45 114
rect 11 12 45 46
<< locali >>
rect 11 1338 45 1354
rect 11 1270 45 1304
rect 11 1202 45 1236
rect 11 1134 45 1168
rect 11 1066 45 1100
rect 11 998 45 1032
rect 11 930 45 964
rect 11 862 45 896
rect 11 794 45 828
rect 11 726 45 760
rect 11 658 45 692
rect 11 590 45 624
rect 11 522 45 556
rect 11 454 45 488
rect 11 386 45 420
rect 11 318 45 352
rect 11 250 45 284
rect 11 182 45 216
rect 11 114 45 148
rect 11 46 45 80
rect 11 -4 45 12
<< properties >>
string GDS_END 34505992
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 34504516
<< end >>
