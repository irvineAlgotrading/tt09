magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< mvnsubdiff >>
rect 1526 2050 1600 2084
<< locali >>
rect 1526 2050 1600 2084
rect 458 947 496 981
rect 530 947 568 981
rect 424 928 602 947
rect 2251 947 2289 981
rect 2323 947 2361 981
rect 2395 947 2433 981
rect 1703 867 1741 901
rect 1775 867 1813 901
rect 2217 894 2467 947
rect 956 669 990 820
rect 956 597 990 635
rect 1132 669 1166 820
rect 1132 597 1166 635
rect 1308 669 1342 820
rect 1308 597 1342 635
rect 1444 669 1478 820
rect 1669 786 1847 867
rect 1444 597 1478 635
rect 2474 669 2508 820
rect 2474 597 2508 635
rect 2610 669 2644 820
rect 2610 597 2644 635
<< viali >>
rect 424 947 458 981
rect 496 947 530 981
rect 568 947 602 981
rect 2217 947 2251 981
rect 2289 947 2323 981
rect 2361 947 2395 981
rect 2433 947 2467 981
rect 1669 867 1703 901
rect 1741 867 1775 901
rect 1813 867 1847 901
rect 956 635 990 669
rect 956 563 990 597
rect 1132 635 1166 669
rect 1132 563 1166 597
rect 1308 635 1342 669
rect 1308 563 1342 597
rect 1444 635 1478 669
rect 1444 563 1478 597
rect 2474 635 2508 669
rect 2474 563 2508 597
rect 2610 635 2644 669
rect 2610 563 2644 597
<< metal1 >>
rect 636 1686 670 1720
rect 2100 1686 2134 1720
rect 2884 1228 2896 1430
rect 412 981 2479 987
rect 412 947 424 981
rect 458 947 496 981
rect 530 947 568 981
rect 602 947 2217 981
rect 2251 947 2289 981
rect 2323 947 2361 981
rect 2395 947 2433 981
rect 2467 947 2479 981
rect 412 941 2479 947
rect 1657 901 1859 907
rect 1657 867 1669 901
rect 1703 867 1741 901
rect 1775 867 1813 901
rect 1847 867 1859 901
rect 1657 861 1859 867
rect 944 669 2656 675
rect 944 635 956 669
rect 990 635 1132 669
rect 1166 635 1308 669
rect 1342 635 1444 669
rect 1478 635 2474 669
rect 2508 635 2610 669
rect 2644 635 2656 669
rect 944 597 2656 635
rect 944 563 956 597
rect 990 563 1132 597
rect 1166 563 1308 597
rect 1342 563 1444 597
rect 1478 563 2474 597
rect 2508 563 2610 597
rect 2644 563 2656 597
rect 944 557 2656 563
rect 1546 30 1592 217
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_0
timestamp 1704896540
transform 1 0 2610 0 -1 669
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_1
timestamp 1704896540
transform 1 0 2474 0 -1 669
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_2
timestamp 1704896540
transform 1 0 1444 0 -1 669
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_3
timestamp 1704896540
transform 1 0 1308 0 -1 669
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_4
timestamp 1704896540
transform 1 0 1132 0 -1 669
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_5
timestamp 1704896540
transform 1 0 956 0 -1 669
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1704896540
transform -1 0 602 0 1 947
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_1
timestamp 1704896540
transform -1 0 1847 0 1 867
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_0
timestamp 1704896540
transform 1 0 2217 0 1 947
box 0 0 1 1
use sky130_fd_io__sio_pupredrvr_reg  sky130_fd_io__sio_pupredrvr_reg_0
timestamp 1704896540
transform 1 0 0 0 1 10
box -108 0 1620 2140
use sky130_fd_io__sio_pupredrvr_reg_slow  sky130_fd_io__sio_pupredrvr_reg_slow_0
timestamp 1704896540
transform 1 0 1518 0 1 10
box -8 0 1378 2140
<< labels >>
flabel metal1 s 1741 867 1775 901 0 FreeSans 200 0 0 0 slow_h_n
port 2 nsew
flabel metal1 s 2884 1228 2896 1430 7 FreeSans 200 0 0 0 vcc_io
port 3 nsew
flabel metal1 s 2066 941 2111 987 0 FreeSans 200 0 0 0 drvhi_h
port 4 nsew
flabel metal1 s 2066 596 2111 635 0 FreeSans 200 0 0 0 puen_h
port 5 nsew
flabel metal1 s 636 1686 670 1720 7 FreeSans 200 0 0 0 pu_h_n<5>
port 6 nsew
flabel metal1 s 2100 1686 2134 1720 7 FreeSans 200 0 0 0 pu_h_n<4>
port 1 nsew
flabel metal1 s 1546 30 1571 217 7 FreeSans 200 0 0 0 vgnd_io
port 7 nsew
flabel metal1 s 1571 30 1592 217 3 FreeSans 200 0 0 0 vgnd_io
port 7 nsew
<< properties >>
string GDS_END 88144788
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 88142148
<< end >>
