magic
tech sky130A
magscale 1 2
timestamp 1704896540
use sky130_fd_pr__dfl1sd2__example_5595914180869  sky130_fd_pr__dfl1sd2__example_5595914180869_0
timestamp 1704896540
transform 1 0 120 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_5595914180869  sky130_fd_pr__dfl1sd2__example_5595914180869_1
timestamp 1704896540
transform 1 0 296 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_5595914180869  sky130_fd_pr__dfl1sd2__example_5595914180869_2
timestamp 1704896540
transform 1 0 472 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_5595914180869  sky130_fd_pr__dfl1sd2__example_5595914180869_3
timestamp 1704896540
transform 1 0 648 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_5595914180869  sky130_fd_pr__dfl1sd2__example_5595914180869_4
timestamp 1704896540
transform 1 0 824 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_5595914180869  sky130_fd_pr__dfl1sd2__example_5595914180869_5
timestamp 1704896540
transform 1 0 1000 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_5595914180868  sky130_fd_pr__dfl1sd__example_5595914180868_0
timestamp 1704896540
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_5595914180868  sky130_fd_pr__dfl1sd__example_5595914180868_1
timestamp 1704896540
transform 1 0 1176 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 21788310
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 21784304
<< end >>
