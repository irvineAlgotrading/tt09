magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect 4276 1557 5361 1725
rect 4282 1021 5361 1557
<< pwell >>
rect 4363 700 5279 916
rect 4316 614 5321 700
<< mvnmos >>
rect 4442 750 4562 890
rect 4618 750 4738 890
rect 4904 750 5024 890
rect 5080 750 5200 890
<< mvpmos >>
rect 4442 1356 4562 1556
rect 4618 1356 4738 1556
rect 4904 1356 5024 1556
rect 5080 1356 5200 1556
rect 4442 1088 4562 1288
rect 4618 1088 4738 1288
rect 4904 1088 5024 1288
rect 5080 1088 5200 1288
<< mvndiff >>
rect 4389 878 4442 890
rect 4389 844 4397 878
rect 4431 844 4442 878
rect 4389 810 4442 844
rect 4389 776 4397 810
rect 4431 776 4442 810
rect 4389 750 4442 776
rect 4562 878 4618 890
rect 4562 844 4573 878
rect 4607 844 4618 878
rect 4562 810 4618 844
rect 4562 776 4573 810
rect 4607 776 4618 810
rect 4562 750 4618 776
rect 4738 878 4791 890
rect 4738 844 4749 878
rect 4783 844 4791 878
rect 4738 810 4791 844
rect 4738 776 4749 810
rect 4783 776 4791 810
rect 4738 750 4791 776
rect 4851 878 4904 890
rect 4851 844 4859 878
rect 4893 844 4904 878
rect 4851 810 4904 844
rect 4851 776 4859 810
rect 4893 776 4904 810
rect 4851 750 4904 776
rect 5024 750 5080 890
rect 5200 878 5253 890
rect 5200 844 5211 878
rect 5245 844 5253 878
rect 5200 810 5253 844
rect 5200 776 5211 810
rect 5245 776 5253 810
rect 5200 750 5253 776
<< mvpdiff >>
rect 4389 1538 4442 1556
rect 4389 1504 4397 1538
rect 4431 1504 4442 1538
rect 4389 1470 4442 1504
rect 4389 1436 4397 1470
rect 4431 1436 4442 1470
rect 4389 1402 4442 1436
rect 4389 1368 4397 1402
rect 4431 1368 4442 1402
rect 4389 1356 4442 1368
rect 4562 1538 4618 1556
rect 4562 1504 4573 1538
rect 4607 1504 4618 1538
rect 4562 1470 4618 1504
rect 4562 1436 4573 1470
rect 4607 1436 4618 1470
rect 4562 1402 4618 1436
rect 4562 1368 4573 1402
rect 4607 1368 4618 1402
rect 4562 1356 4618 1368
rect 4738 1538 4791 1556
rect 4738 1504 4749 1538
rect 4783 1504 4791 1538
rect 4738 1470 4791 1504
rect 4738 1436 4749 1470
rect 4783 1436 4791 1470
rect 4738 1402 4791 1436
rect 4738 1368 4749 1402
rect 4783 1368 4791 1402
rect 4738 1356 4791 1368
rect 4851 1538 4904 1556
rect 4851 1504 4859 1538
rect 4893 1504 4904 1538
rect 4851 1470 4904 1504
rect 4851 1436 4859 1470
rect 4893 1436 4904 1470
rect 4851 1402 4904 1436
rect 4851 1368 4859 1402
rect 4893 1368 4904 1402
rect 4851 1356 4904 1368
rect 5024 1538 5080 1556
rect 5024 1504 5035 1538
rect 5069 1504 5080 1538
rect 5024 1470 5080 1504
rect 5024 1436 5035 1470
rect 5069 1436 5080 1470
rect 5024 1402 5080 1436
rect 5024 1368 5035 1402
rect 5069 1368 5080 1402
rect 5024 1356 5080 1368
rect 5200 1538 5253 1556
rect 5200 1504 5211 1538
rect 5245 1504 5253 1538
rect 5200 1470 5253 1504
rect 5200 1436 5211 1470
rect 5245 1436 5253 1470
rect 5200 1402 5253 1436
rect 5200 1368 5211 1402
rect 5245 1368 5253 1402
rect 5200 1356 5253 1368
rect 4389 1276 4442 1288
rect 4389 1242 4397 1276
rect 4431 1242 4442 1276
rect 4389 1208 4442 1242
rect 4389 1174 4397 1208
rect 4431 1174 4442 1208
rect 4389 1140 4442 1174
rect 4389 1106 4397 1140
rect 4431 1106 4442 1140
rect 4389 1088 4442 1106
rect 4562 1276 4618 1288
rect 4562 1242 4573 1276
rect 4607 1242 4618 1276
rect 4562 1208 4618 1242
rect 4562 1174 4573 1208
rect 4607 1174 4618 1208
rect 4562 1140 4618 1174
rect 4562 1106 4573 1140
rect 4607 1106 4618 1140
rect 4562 1088 4618 1106
rect 4738 1276 4791 1288
rect 4738 1242 4749 1276
rect 4783 1242 4791 1276
rect 4738 1208 4791 1242
rect 4738 1174 4749 1208
rect 4783 1174 4791 1208
rect 4738 1140 4791 1174
rect 4738 1106 4749 1140
rect 4783 1106 4791 1140
rect 4738 1088 4791 1106
rect 4851 1276 4904 1288
rect 4851 1242 4859 1276
rect 4893 1242 4904 1276
rect 4851 1208 4904 1242
rect 4851 1174 4859 1208
rect 4893 1174 4904 1208
rect 4851 1140 4904 1174
rect 4851 1106 4859 1140
rect 4893 1106 4904 1140
rect 4851 1088 4904 1106
rect 5024 1276 5080 1288
rect 5024 1242 5035 1276
rect 5069 1242 5080 1276
rect 5024 1208 5080 1242
rect 5024 1174 5035 1208
rect 5069 1174 5080 1208
rect 5024 1140 5080 1174
rect 5024 1106 5035 1140
rect 5069 1106 5080 1140
rect 5024 1088 5080 1106
rect 5200 1276 5253 1288
rect 5200 1242 5211 1276
rect 5245 1242 5253 1276
rect 5200 1208 5253 1242
rect 5200 1174 5211 1208
rect 5245 1174 5253 1208
rect 5200 1140 5253 1174
rect 5200 1106 5211 1140
rect 5245 1106 5253 1140
rect 5200 1088 5253 1106
<< mvndiffc >>
rect 4397 844 4431 878
rect 4397 776 4431 810
rect 4573 844 4607 878
rect 4573 776 4607 810
rect 4749 844 4783 878
rect 4749 776 4783 810
rect 4859 844 4893 878
rect 4859 776 4893 810
rect 5211 844 5245 878
rect 5211 776 5245 810
<< mvpdiffc >>
rect 4397 1504 4431 1538
rect 4397 1436 4431 1470
rect 4397 1368 4431 1402
rect 4573 1504 4607 1538
rect 4573 1436 4607 1470
rect 4573 1368 4607 1402
rect 4749 1504 4783 1538
rect 4749 1436 4783 1470
rect 4749 1368 4783 1402
rect 4859 1504 4893 1538
rect 4859 1436 4893 1470
rect 4859 1368 4893 1402
rect 5035 1504 5069 1538
rect 5035 1436 5069 1470
rect 5035 1368 5069 1402
rect 5211 1504 5245 1538
rect 5211 1436 5245 1470
rect 5211 1368 5245 1402
rect 4397 1242 4431 1276
rect 4397 1174 4431 1208
rect 4397 1106 4431 1140
rect 4573 1242 4607 1276
rect 4573 1174 4607 1208
rect 4573 1106 4607 1140
rect 4749 1242 4783 1276
rect 4749 1174 4783 1208
rect 4749 1106 4783 1140
rect 4859 1242 4893 1276
rect 4859 1174 4893 1208
rect 4859 1106 4893 1140
rect 5035 1242 5069 1276
rect 5035 1174 5069 1208
rect 5035 1106 5069 1140
rect 5211 1242 5245 1276
rect 5211 1174 5245 1208
rect 5211 1106 5245 1140
<< mvpsubdiff >>
rect 4342 640 4366 674
rect 4400 640 4439 674
rect 4473 640 4512 674
rect 4546 640 4585 674
rect 4619 640 4658 674
rect 4692 640 4731 674
rect 4765 640 4804 674
rect 4838 640 4877 674
rect 4911 640 4949 674
rect 4983 640 5021 674
rect 5055 640 5093 674
rect 5127 640 5165 674
rect 5199 640 5237 674
rect 5271 640 5295 674
<< mvnsubdiff >>
rect 4343 1624 4377 1658
rect 4411 1624 4445 1658
rect 4479 1624 4513 1658
rect 4547 1624 4581 1658
rect 4615 1624 4649 1658
rect 4683 1624 4717 1658
rect 4751 1624 4785 1658
rect 4819 1624 4853 1658
rect 4887 1624 4921 1658
rect 4955 1624 4989 1658
rect 5023 1624 5057 1658
rect 5091 1624 5125 1658
rect 5159 1624 5193 1658
rect 5227 1624 5294 1658
<< mvpsubdiffcont >>
rect 4366 640 4400 674
rect 4439 640 4473 674
rect 4512 640 4546 674
rect 4585 640 4619 674
rect 4658 640 4692 674
rect 4731 640 4765 674
rect 4804 640 4838 674
rect 4877 640 4911 674
rect 4949 640 4983 674
rect 5021 640 5055 674
rect 5093 640 5127 674
rect 5165 640 5199 674
rect 5237 640 5271 674
<< mvnsubdiffcont >>
rect 4377 1624 4411 1658
rect 4445 1624 4479 1658
rect 4513 1624 4547 1658
rect 4581 1624 4615 1658
rect 4649 1624 4683 1658
rect 4717 1624 4751 1658
rect 4785 1624 4819 1658
rect 4853 1624 4887 1658
rect 4921 1624 4955 1658
rect 4989 1624 5023 1658
rect 5057 1624 5091 1658
rect 5125 1624 5159 1658
rect 5193 1624 5227 1658
<< poly >>
rect 4442 1556 4562 1582
rect 4618 1556 4738 1582
rect 4904 1556 5024 1582
rect 5080 1556 5200 1582
rect 4442 1288 4562 1356
rect 4618 1288 4738 1356
rect 4904 1288 5024 1356
rect 5080 1288 5200 1356
rect 4442 1040 4562 1088
rect 4442 1006 4484 1040
rect 4518 1006 4562 1040
rect 4442 972 4562 1006
rect 4442 938 4484 972
rect 4518 938 4562 972
rect 4442 890 4562 938
rect 4618 1040 4738 1088
rect 4618 1006 4662 1040
rect 4696 1006 4738 1040
rect 4618 972 4738 1006
rect 4618 938 4662 972
rect 4696 938 4738 972
rect 4618 890 4738 938
rect 4904 1040 5024 1088
rect 4904 1006 4949 1040
rect 4983 1006 5024 1040
rect 4904 972 5024 1006
rect 4904 938 4949 972
rect 4983 938 5024 972
rect 4904 890 5024 938
rect 5080 1040 5200 1088
rect 5080 1006 5120 1040
rect 5154 1006 5200 1040
rect 5080 972 5200 1006
rect 5080 938 5120 972
rect 5154 938 5200 972
rect 5080 890 5200 938
rect 4442 724 4562 750
rect 4618 724 4738 750
rect 4904 724 5024 750
rect 5080 724 5200 750
<< polycont >>
rect 4484 1006 4518 1040
rect 4484 938 4518 972
rect 4662 1006 4696 1040
rect 4662 938 4696 972
rect 4949 1006 4983 1040
rect 4949 938 4983 972
rect 5120 1006 5154 1040
rect 5120 938 5154 972
<< locali >>
rect 4343 1624 4356 1658
rect 4411 1624 4431 1658
rect 4479 1624 4506 1658
rect 4547 1624 4581 1658
rect 4615 1624 4649 1658
rect 4690 1624 4717 1658
rect 4764 1624 4785 1658
rect 4838 1624 4853 1658
rect 4912 1624 4921 1658
rect 4986 1624 4989 1658
rect 5023 1624 5026 1658
rect 5091 1624 5100 1658
rect 5159 1624 5174 1658
rect 5227 1624 5248 1658
rect 5282 1624 5294 1658
rect 4397 1538 4431 1556
rect 4397 1470 4431 1504
rect 4397 1402 4431 1436
rect 4397 1276 4431 1368
rect 4397 1208 4431 1242
rect 4397 1140 4431 1169
rect 4397 1056 4431 1096
rect 4573 1538 4607 1550
rect 4573 1470 4607 1478
rect 4573 1402 4607 1436
rect 4573 1276 4607 1368
rect 4573 1208 4607 1242
rect 4573 1140 4607 1174
rect 4573 1090 4607 1106
rect 4749 1538 4783 1556
rect 4749 1470 4783 1504
rect 4749 1425 4783 1436
rect 4749 1353 4783 1368
rect 4749 1276 4783 1319
rect 4749 1208 4783 1242
rect 4749 1140 4783 1174
rect 4397 982 4431 1022
rect 4397 878 4431 948
rect 4468 1006 4484 1040
rect 4468 972 4534 1006
rect 4468 938 4484 972
rect 4518 968 4534 972
rect 4646 1006 4662 1040
rect 4699 1010 4712 1040
rect 4696 1006 4712 1010
rect 4646 972 4712 1006
rect 4646 938 4662 972
rect 4699 938 4712 972
rect 4397 810 4431 844
rect 4397 760 4431 776
rect 4573 878 4607 894
rect 4573 833 4607 844
rect 4573 761 4607 776
rect 4749 878 4783 1106
rect 4859 1538 4893 1550
rect 4859 1470 4893 1478
rect 4859 1402 4893 1436
rect 4859 1276 4893 1368
rect 4859 1208 4893 1242
rect 4859 1140 4893 1174
rect 4859 1090 4893 1106
rect 5035 1538 5069 1556
rect 5035 1470 5069 1504
rect 5035 1402 5069 1436
rect 5035 1276 5069 1368
rect 5035 1208 5069 1242
rect 5035 1140 5069 1174
rect 4933 1013 4939 1040
rect 4933 1006 4949 1013
rect 4983 1006 4999 1040
rect 4933 975 4999 1006
rect 4933 941 4939 975
rect 4973 972 4999 975
rect 4933 938 4949 941
rect 4983 938 4999 972
rect 5035 991 5069 1106
rect 5211 1538 5245 1550
rect 5211 1470 5245 1478
rect 5211 1402 5245 1436
rect 5211 1276 5245 1368
rect 5211 1208 5245 1242
rect 5211 1140 5245 1174
rect 5211 1090 5245 1106
rect 5035 919 5069 957
rect 5104 1006 5120 1040
rect 5154 1006 5170 1010
rect 5104 972 5170 1006
rect 5104 938 5120 972
rect 4749 810 4783 844
rect 4749 760 4783 776
rect 4859 878 4893 894
rect 5035 867 5069 885
rect 4893 844 5069 867
rect 4859 833 5069 844
rect 5211 878 5245 894
rect 5211 833 5245 844
rect 4859 810 4898 833
rect 4893 776 4898 810
rect 4859 760 4898 776
rect 5211 761 5245 776
rect 4342 640 4354 674
rect 4400 640 4429 674
rect 4473 640 4504 674
rect 4546 640 4579 674
rect 4619 640 4654 674
rect 4692 640 4729 674
rect 4765 640 4804 674
rect 4838 640 4877 674
rect 4913 640 4949 674
rect 4987 640 5021 674
rect 5061 640 5093 674
rect 5135 640 5165 674
rect 5209 640 5237 674
rect 5283 640 5295 674
<< viali >>
rect 4356 1624 4377 1658
rect 4377 1624 4390 1658
rect 4431 1624 4445 1658
rect 4445 1624 4465 1658
rect 4506 1624 4513 1658
rect 4513 1624 4540 1658
rect 4581 1624 4615 1658
rect 4656 1624 4683 1658
rect 4683 1624 4690 1658
rect 4730 1624 4751 1658
rect 4751 1624 4764 1658
rect 4804 1624 4819 1658
rect 4819 1624 4838 1658
rect 4878 1624 4887 1658
rect 4887 1624 4912 1658
rect 4952 1624 4955 1658
rect 4955 1624 4986 1658
rect 5026 1624 5057 1658
rect 5057 1624 5060 1658
rect 5100 1624 5125 1658
rect 5125 1624 5134 1658
rect 5174 1624 5193 1658
rect 5193 1624 5208 1658
rect 5248 1624 5282 1658
rect 4397 1242 4431 1276
rect 4397 1174 4431 1203
rect 4397 1169 4431 1174
rect 4397 1106 4431 1130
rect 4397 1096 4431 1106
rect 4573 1550 4607 1584
rect 4573 1504 4607 1512
rect 4573 1478 4607 1504
rect 4749 1402 4783 1425
rect 4749 1391 4783 1402
rect 4749 1319 4783 1353
rect 4397 1022 4431 1056
rect 4665 1040 4699 1044
rect 4397 948 4431 982
rect 4500 1006 4518 1040
rect 4518 1006 4534 1040
rect 4500 938 4518 968
rect 4518 938 4534 968
rect 4665 1010 4696 1040
rect 4696 1010 4699 1040
rect 4665 938 4696 972
rect 4696 938 4699 972
rect 4500 934 4534 938
rect 4573 810 4607 833
rect 4573 799 4607 810
rect 4573 727 4607 761
rect 4859 1550 4893 1584
rect 4859 1504 4893 1512
rect 4859 1478 4893 1504
rect 4939 1040 4973 1047
rect 4939 1013 4949 1040
rect 4949 1013 4973 1040
rect 4939 972 4973 975
rect 4939 941 4949 972
rect 4949 941 4973 972
rect 5211 1550 5245 1584
rect 5211 1504 5245 1512
rect 5211 1478 5245 1504
rect 5136 1040 5170 1044
rect 5035 957 5069 991
rect 5136 1010 5154 1040
rect 5154 1010 5170 1040
rect 5136 938 5154 972
rect 5154 938 5170 972
rect 5035 885 5069 919
rect 5211 810 5245 833
rect 5211 799 5245 810
rect 5211 727 5245 761
rect 4354 640 4366 674
rect 4366 640 4388 674
rect 4429 640 4439 674
rect 4439 640 4463 674
rect 4504 640 4512 674
rect 4512 640 4538 674
rect 4579 640 4585 674
rect 4585 640 4613 674
rect 4654 640 4658 674
rect 4658 640 4688 674
rect 4729 640 4731 674
rect 4731 640 4763 674
rect 4804 640 4838 674
rect 4879 640 4911 674
rect 4911 640 4913 674
rect 4953 640 4983 674
rect 4983 640 4987 674
rect 5027 640 5055 674
rect 5055 640 5061 674
rect 5101 640 5127 674
rect 5127 640 5135 674
rect 5175 640 5199 674
rect 5199 640 5209 674
rect 5249 640 5271 674
rect 5271 640 5283 674
<< metal1 >>
rect 8293 4271 8345 4277
rect 8293 4207 8345 4219
rect -92 4149 -86 4201
rect -34 4149 -22 4201
rect 30 4149 4234 4201
tri 4148 4121 4176 4149 ne
rect 4176 4121 4234 4149
rect 109 4069 583 4121
rect 635 4069 647 4121
rect 699 4069 3455 4121
rect 3507 4069 3519 4121
rect 3571 4069 3859 4121
rect 3911 4069 3926 4121
rect 3978 4069 3984 4121
tri 4176 4115 4182 4121 ne
rect 1412 3954 1612 3960
rect 1464 3902 1486 3954
rect 1538 3902 1560 3954
rect 1412 3885 1612 3902
rect 1464 3833 1486 3885
rect 1538 3833 1560 3885
rect 1412 3816 1612 3833
rect 1464 3764 1486 3816
rect 1538 3764 1560 3816
rect 2374 3793 2717 3928
rect 1412 3758 1612 3764
rect 3996 3758 4154 3960
rect 3836 3724 3964 3730
rect 3888 3672 3912 3724
rect 3836 3658 3964 3672
rect 3888 3606 3912 3658
rect 3836 3600 3964 3606
rect 4182 3718 4234 4121
rect 4182 3654 4234 3666
rect 653 3468 705 3474
rect 3449 3468 3501 3474
rect 194 3376 294 3406
rect 653 3398 705 3416
rect 1783 3409 1923 3438
rect 2146 3408 2248 3435
rect 653 3340 705 3346
rect 3449 3398 3501 3416
rect 3811 3370 3951 3404
rect 3449 3340 3501 3346
rect 1576 3085 1700 3118
rect 2381 3083 2512 3118
rect 1112 2961 1312 2962
rect 1112 2909 1118 2961
rect 1170 2909 1186 2961
rect 1238 2909 1254 2961
rect 1306 2909 1312 2961
rect 1112 2889 1312 2909
rect 1112 2837 1118 2889
rect 1170 2837 1186 2889
rect 1238 2837 1254 2889
rect 1306 2837 1312 2889
rect 1112 2817 1312 2837
rect 1112 2765 1118 2817
rect 1170 2765 1186 2817
rect 1238 2765 1254 2817
rect 1306 2765 1312 2817
rect 1112 2764 1312 2765
tri 76 2729 110 2763 ne
rect 110 2668 162 2763
tri 162 2729 196 2763 nw
tri 3958 2729 3992 2763 ne
rect 3992 2668 4044 2763
tri 4044 2729 4078 2763 nw
rect -92 2522 -40 2528
rect -92 2458 -40 2470
tri -40 2446 -6 2480 sw
tri 278 2446 310 2478 se
rect 310 2458 356 2552
rect 310 2446 344 2458
tri 344 2446 356 2458 nw
rect 3798 2458 3844 2552
tri 4180 2478 4182 2480 se
rect 4182 2478 4234 3602
tri 3798 2446 3810 2458 ne
rect 3810 2446 3844 2458
tri 3844 2446 3876 2478 sw
tri 4148 2446 4180 2478 se
rect 4180 2446 4234 2478
rect -40 2406 298 2446
rect -92 2400 298 2406
tri 298 2400 344 2446 nw
tri 3810 2412 3844 2446 ne
rect 3844 2412 4234 2446
tri 3844 2400 3856 2412 ne
rect 3856 2400 4234 2412
tri 4148 2366 4182 2400 ne
rect 2983 2120 3355 2238
tri 4148 1720 4182 1754 se
rect 4182 1720 4234 2400
rect -92 1714 298 1720
rect -40 1674 298 1714
rect -40 1662 -22 1674
rect -92 1658 -22 1662
tri -22 1658 -6 1674 nw
tri 278 1658 294 1674 ne
rect 294 1662 298 1674
tri 298 1662 356 1720 sw
rect 294 1658 356 1662
rect -92 1650 -40 1658
tri -40 1640 -22 1658 nw
tri 294 1654 298 1658 ne
rect 298 1654 356 1658
tri 298 1642 310 1654 ne
rect -92 1592 -40 1598
rect 310 1568 356 1654
tri 3798 1662 3856 1720 se
rect 3856 1674 4234 1720
rect 3856 1662 3864 1674
tri 3864 1662 3876 1674 nw
tri 4148 1662 4160 1674 ne
rect 4160 1662 4234 1674
rect 3798 1658 3860 1662
tri 3860 1658 3864 1662 nw
tri 4160 1658 4164 1662 ne
rect 4164 1658 4234 1662
rect 3798 1568 3844 1658
tri 3844 1642 3860 1658 nw
tri 4164 1642 4180 1658 ne
rect 4180 1642 4234 1658
tri 4180 1640 4182 1642 ne
tri 84 1319 110 1345 se
rect 110 1319 162 1406
tri 162 1319 188 1345 sw
tri 3966 1319 3992 1345 se
rect 3992 1319 4044 1406
tri 4044 1319 4070 1345 sw
tri 76 1311 84 1319 se
rect 84 1311 188 1319
tri 188 1311 196 1319 sw
tri 3958 1311 3966 1319 se
rect 3966 1311 4070 1319
tri 4070 1311 4078 1319 sw
rect 1112 1309 1312 1311
rect 1112 1257 1118 1309
rect 1170 1257 1186 1309
rect 1238 1257 1254 1309
rect 1306 1282 1312 1309
rect 3996 1305 4154 1311
rect 1306 1257 1349 1282
rect 1112 1237 1349 1257
rect 1112 1185 1118 1237
rect 1170 1185 1186 1237
rect 1238 1185 1254 1237
rect 1306 1185 1349 1237
rect 1112 1165 1349 1185
rect 1112 1113 1118 1165
rect 1170 1113 1186 1165
rect 1238 1113 1254 1165
rect 1306 1151 1349 1165
rect 4048 1253 4102 1305
rect 3996 1238 4154 1253
rect 4048 1186 4102 1238
rect 3996 1170 4154 1186
rect 1306 1113 1312 1151
rect 1112 1112 1312 1113
rect 4048 1118 4102 1170
rect 4182 1263 4234 1642
rect 4262 4069 4268 4121
rect 4320 4069 4332 4121
rect 4384 4069 4390 4121
rect 4262 1434 4314 4069
tri 4314 4035 4348 4069 nw
rect 8293 3718 8345 4155
rect 8519 4069 8525 4121
rect 8577 4069 8589 4121
rect 8641 4069 9765 4121
rect 9817 4069 9829 4121
rect 9881 4069 9887 4121
rect 8956 3954 9156 3960
rect 9008 3902 9030 3954
rect 9082 3902 9104 3954
rect 8956 3885 9156 3902
rect 9008 3833 9030 3885
rect 9082 3833 9104 3885
rect 8956 3816 9156 3833
rect 9008 3764 9030 3816
rect 9082 3764 9104 3816
rect 9256 3793 9599 3928
rect 8956 3758 9156 3764
rect 8293 3654 8345 3666
rect 8293 3596 8345 3602
rect 10222 3724 10350 3730
rect 10274 3672 10298 3724
rect 10222 3658 10350 3672
rect 10274 3606 10298 3658
rect 10222 3600 10350 3606
rect 9835 3468 9887 3474
rect 8546 3406 8681 3438
rect 9835 3398 9887 3416
rect 10195 3368 10313 3402
rect 9835 3340 9887 3346
rect 8777 3084 8880 3117
rect 10458 2956 10574 2962
rect 10510 2904 10522 2956
rect 10458 2889 10574 2904
rect 10510 2837 10522 2889
rect 10458 2821 10574 2837
rect 10510 2769 10522 2821
rect 10458 2763 10574 2769
tri 10344 2729 10378 2763 ne
rect 10378 2668 10430 2763
tri 10430 2729 10464 2763 nw
rect 10184 2412 10230 2520
rect 10378 2463 10430 2469
tri 10184 2366 10230 2412 ne
tri 10230 2387 10275 2432 sw
tri 10344 2387 10378 2421 se
rect 10378 2399 10430 2411
rect 10230 2366 10378 2387
tri 10230 2341 10255 2366 ne
rect 10255 2347 10378 2366
rect 10255 2341 10430 2347
rect 9332 2120 9704 2238
tri 10189 1681 10255 1747 se
rect 10255 1741 10430 1747
rect 10255 1701 10378 1741
tri 10255 1681 10275 1701 nw
tri 10344 1681 10364 1701 ne
rect 10364 1689 10378 1701
rect 10364 1681 10430 1689
tri 10184 1676 10189 1681 se
rect 10189 1676 10230 1681
rect 4342 1658 5294 1668
rect 4342 1624 4356 1658
rect 4390 1624 4431 1658
rect 4465 1624 4506 1658
rect 4540 1624 4581 1658
rect 4615 1624 4656 1658
rect 4690 1624 4730 1658
rect 4764 1624 4804 1658
rect 4838 1624 4878 1658
rect 4912 1624 4952 1658
rect 4986 1624 5026 1658
rect 5060 1624 5100 1658
rect 5134 1624 5174 1658
rect 5208 1624 5248 1658
rect 5282 1624 5294 1658
rect 4342 1584 5294 1624
rect 4342 1550 4573 1584
rect 4607 1550 4859 1584
rect 4893 1550 5211 1584
rect 5245 1550 5294 1584
rect 10184 1568 10230 1676
tri 10230 1656 10255 1681 nw
tri 10364 1667 10378 1681 ne
rect 10378 1677 10430 1681
rect 10378 1619 10430 1625
rect 4342 1512 5294 1550
rect 4342 1478 4573 1512
rect 4607 1478 4859 1512
rect 4893 1478 5211 1512
rect 5245 1478 5294 1512
rect 4342 1465 5294 1478
tri 4314 1434 4331 1451 sw
tri 4740 1434 4743 1437 se
rect 4743 1434 4789 1437
rect 4262 1429 4331 1434
tri 4262 1425 4266 1429 ne
rect 4266 1425 4331 1429
tri 4331 1425 4340 1434 sw
tri 4731 1425 4740 1434 se
rect 4740 1425 4789 1434
tri 4266 1391 4300 1425 ne
rect 4300 1412 4340 1425
tri 4340 1412 4353 1425 sw
tri 4718 1412 4731 1425 se
rect 4731 1412 4749 1425
rect 4300 1391 4749 1412
rect 4783 1391 4789 1425
tri 4300 1360 4331 1391 ne
rect 4331 1360 4789 1391
tri 4709 1353 4716 1360 ne
rect 4716 1353 4789 1360
tri 4716 1326 4743 1353 ne
rect 4743 1319 4749 1353
rect 4783 1319 4789 1353
rect 4743 1307 4789 1319
tri 10344 1311 10378 1345 se
rect 10378 1311 10430 1406
tri 10430 1311 10464 1345 sw
rect 10458 1305 10574 1311
rect 4182 1199 4234 1211
rect 4182 1141 4234 1147
rect 4388 1276 4440 1288
rect 4388 1263 4397 1276
rect 4431 1263 4440 1276
tri 4540 1214 4601 1275 se
rect 4601 1249 5101 1275
tri 5101 1249 5127 1275 sw
rect 4601 1229 5127 1249
rect 4601 1214 4606 1229
tri 4606 1214 4621 1229 nw
tri 5081 1214 5096 1229 ne
rect 5096 1214 5127 1229
rect 4388 1203 4440 1211
rect 4388 1199 4397 1203
rect 4431 1199 4440 1203
rect 3996 1112 4154 1118
rect 4388 1130 4440 1147
rect 4388 1096 4397 1130
rect 4431 1096 4440 1130
rect 4388 1056 4440 1096
rect 4388 1022 4397 1056
rect 4431 1022 4440 1056
rect 1589 956 1741 986
rect 2398 957 2565 992
rect 4388 982 4440 1022
rect 4388 948 4397 982
rect 4431 948 4440 982
rect 4388 936 4440 948
tri 4494 1168 4540 1214 se
rect 4494 1040 4540 1168
tri 4540 1148 4606 1214 nw
tri 5096 1183 5127 1214 ne
tri 5127 1197 5179 1249 sw
rect 4494 1006 4500 1040
rect 4534 1006 4540 1040
rect 4494 968 4540 1006
rect 4494 934 4500 968
rect 4534 934 4540 968
rect 4494 922 4540 934
rect 4659 1044 4705 1056
rect 4659 1010 4665 1044
rect 4699 1010 4705 1044
rect 4659 972 4705 1010
rect 4659 938 4665 972
rect 4699 938 4705 972
rect 4659 919 4705 938
rect 4933 1047 4979 1059
rect 4933 1013 4939 1047
rect 4973 1013 4979 1047
rect 5127 1044 5179 1197
rect 9221 1151 9409 1282
rect 10510 1253 10522 1305
rect 10458 1238 10574 1253
rect 10510 1186 10522 1238
rect 10458 1170 10574 1186
rect 10510 1118 10522 1170
rect 10458 1112 10574 1118
rect 5127 1014 5136 1044
rect 4933 975 4979 1013
rect 5130 1010 5136 1014
rect 5170 1014 5179 1044
rect 5170 1010 5176 1014
rect 4933 941 4939 975
rect 4973 941 4979 975
tri 4705 919 4721 935 sw
rect 4933 929 4979 941
rect 5029 991 5075 1003
rect 5029 957 5035 991
rect 5069 957 5075 991
tri 5023 929 5029 935 se
rect 5029 929 5075 957
tri 5013 919 5023 929 se
rect 5023 919 5075 929
rect 5130 972 5176 1010
rect 5130 938 5136 972
rect 5170 938 5176 972
rect 8782 960 8946 989
rect 5130 926 5176 938
rect 4659 901 4721 919
tri 4721 901 4739 919 sw
tri 4995 901 5013 919 se
rect 5013 901 5035 919
rect 4659 885 5035 901
rect 5069 885 5075 919
rect 4659 873 5075 885
rect 4342 844 5295 845
rect 4342 792 4348 844
rect 4400 792 4433 844
rect 4485 792 4518 844
rect 4570 833 4603 844
rect 4655 833 5295 844
rect 4570 799 4573 833
rect 4655 799 5211 833
rect 5245 799 5295 833
rect 4570 792 4603 799
rect 4655 792 5295 799
rect 4342 761 5295 792
rect 4342 740 4573 761
rect 4607 740 5211 761
rect 653 728 705 734
rect 225 667 347 704
rect 653 658 705 676
rect 3449 728 3501 734
rect 1839 641 1973 673
rect 2221 638 2363 664
rect 3449 658 3501 676
rect 3779 673 3893 702
rect 4342 688 4348 740
rect 4400 688 4433 740
rect 4485 688 4518 740
rect 4570 727 4573 740
rect 4655 727 5211 740
rect 5245 727 5295 761
rect 4570 688 4603 727
rect 4655 688 5295 727
rect 4342 674 5295 688
rect 653 600 705 606
rect 4342 640 4354 674
rect 4388 640 4429 674
rect 4463 640 4504 674
rect 4538 640 4579 674
rect 4613 640 4654 674
rect 4688 640 4729 674
rect 4763 640 4804 674
rect 4838 640 4879 674
rect 4913 640 4953 674
rect 4987 640 5027 674
rect 5061 640 5101 674
rect 5135 640 5175 674
rect 5209 640 5249 674
rect 5283 640 5295 674
rect 9835 728 9887 734
rect 4342 630 5295 640
rect 8552 638 8662 669
rect 9835 658 9887 676
rect 10229 669 10306 701
rect 3449 600 3501 606
rect 9835 600 9887 606
rect 3836 468 3964 474
rect 3888 416 3912 468
rect 3836 402 3964 416
rect 3888 350 3912 402
rect 3836 344 3964 350
rect 10222 468 10350 474
rect 10274 416 10298 468
rect 10222 402 10350 416
rect 10274 350 10298 402
rect 10222 344 10350 350
rect 1412 310 1612 316
rect 1464 258 1486 310
rect 1538 258 1560 310
rect 1412 241 1612 258
rect 1464 189 1486 241
rect 1538 189 1560 241
rect 1412 172 1612 189
rect 1464 120 1486 172
rect 1538 120 1560 172
rect 1412 114 1612 120
rect 8956 310 9156 316
rect 9008 258 9030 310
rect 9082 258 9104 310
rect 8956 241 9156 258
rect 9008 189 9030 241
rect 9082 189 9104 241
rect 8956 172 9156 189
rect 9008 120 9030 172
rect 9082 120 9104 172
rect 8956 114 9156 120
<< via1 >>
rect 8293 4219 8345 4271
rect -86 4149 -34 4201
rect -22 4149 30 4201
rect 8293 4155 8345 4207
rect 583 4069 635 4121
rect 647 4069 699 4121
rect 3455 4069 3507 4121
rect 3519 4069 3571 4121
rect 3859 4069 3911 4121
rect 3926 4069 3978 4121
rect 1412 3902 1464 3954
rect 1486 3902 1538 3954
rect 1560 3902 1612 3954
rect 1412 3833 1464 3885
rect 1486 3833 1538 3885
rect 1560 3833 1612 3885
rect 1412 3764 1464 3816
rect 1486 3764 1538 3816
rect 1560 3764 1612 3816
rect 3836 3672 3888 3724
rect 3912 3672 3964 3724
rect 3836 3606 3888 3658
rect 3912 3606 3964 3658
rect 4182 3666 4234 3718
rect 4182 3602 4234 3654
rect 653 3416 705 3468
rect 3449 3416 3501 3468
rect 653 3346 705 3398
rect 3449 3346 3501 3398
rect 1118 2909 1170 2961
rect 1186 2909 1238 2961
rect 1254 2909 1306 2961
rect 1118 2837 1170 2889
rect 1186 2837 1238 2889
rect 1254 2837 1306 2889
rect 1118 2765 1170 2817
rect 1186 2765 1238 2817
rect 1254 2765 1306 2817
rect -92 2470 -40 2522
rect -92 2406 -40 2458
rect -92 1662 -40 1714
rect -92 1598 -40 1650
rect 1118 1257 1170 1309
rect 1186 1257 1238 1309
rect 1254 1257 1306 1309
rect 1118 1185 1170 1237
rect 1186 1185 1238 1237
rect 1254 1185 1306 1237
rect 1118 1113 1170 1165
rect 1186 1113 1238 1165
rect 1254 1113 1306 1165
rect 3996 1253 4048 1305
rect 4102 1253 4154 1305
rect 3996 1186 4048 1238
rect 4102 1186 4154 1238
rect 3996 1118 4048 1170
rect 4102 1118 4154 1170
rect 4268 4069 4320 4121
rect 4332 4069 4384 4121
rect 8525 4069 8577 4121
rect 8589 4069 8641 4121
rect 9765 4069 9817 4121
rect 9829 4069 9881 4121
rect 8956 3902 9008 3954
rect 9030 3902 9082 3954
rect 9104 3902 9156 3954
rect 8956 3833 9008 3885
rect 9030 3833 9082 3885
rect 9104 3833 9156 3885
rect 8956 3764 9008 3816
rect 9030 3764 9082 3816
rect 9104 3764 9156 3816
rect 8293 3666 8345 3718
rect 8293 3602 8345 3654
rect 10222 3672 10274 3724
rect 10298 3672 10350 3724
rect 10222 3606 10274 3658
rect 10298 3606 10350 3658
rect 9835 3416 9887 3468
rect 9835 3346 9887 3398
rect 10458 2904 10510 2956
rect 10522 2904 10574 2956
rect 10458 2837 10510 2889
rect 10522 2837 10574 2889
rect 10458 2769 10510 2821
rect 10522 2769 10574 2821
rect 10378 2411 10430 2463
rect 10378 2347 10430 2399
rect 10378 1689 10430 1741
rect 10378 1625 10430 1677
rect 4182 1211 4234 1263
rect 4182 1147 4234 1199
rect 4388 1242 4397 1263
rect 4397 1242 4431 1263
rect 4431 1242 4440 1263
rect 4388 1211 4440 1242
rect 4388 1169 4397 1199
rect 4397 1169 4431 1199
rect 4431 1169 4440 1199
rect 4388 1147 4440 1169
rect 10458 1253 10510 1305
rect 10522 1253 10574 1305
rect 10458 1186 10510 1238
rect 10522 1186 10574 1238
rect 10458 1118 10510 1170
rect 10522 1118 10574 1170
rect 4348 792 4400 844
rect 4433 792 4485 844
rect 4518 792 4570 844
rect 4603 833 4655 844
rect 4603 799 4607 833
rect 4607 799 4655 833
rect 4603 792 4655 799
rect 653 676 705 728
rect 3449 676 3501 728
rect 653 606 705 658
rect 4348 688 4400 740
rect 4433 688 4485 740
rect 4518 688 4570 740
rect 4603 727 4607 740
rect 4607 727 4655 740
rect 4603 688 4655 727
rect 3449 606 3501 658
rect 9835 676 9887 728
rect 9835 606 9887 658
rect 3836 416 3888 468
rect 3912 416 3964 468
rect 3836 350 3888 402
rect 3912 350 3964 402
rect 10222 416 10274 468
rect 10298 416 10350 468
rect 10222 350 10274 402
rect 10298 350 10350 402
rect 1412 258 1464 310
rect 1486 258 1538 310
rect 1560 258 1612 310
rect 1412 189 1464 241
rect 1486 189 1538 241
rect 1560 189 1612 241
rect 1412 120 1464 172
rect 1486 120 1538 172
rect 1560 120 1612 172
rect 8956 258 9008 310
rect 9030 258 9082 310
rect 9104 258 9156 310
rect 8956 189 9008 241
rect 9030 189 9082 241
rect 9104 189 9156 241
rect 8956 120 9008 172
rect 9030 120 9082 172
rect 9104 120 9156 172
<< metal2 >>
rect 8293 4271 8345 4277
rect 8293 4207 8345 4219
rect -92 4149 -86 4201
rect -34 4149 -22 4201
rect 30 4149 36 4201
tri 8345 4201 8379 4235 sw
rect 8345 4155 10430 4201
rect 8293 4149 10430 4155
rect -92 4121 -34 4149
tri -34 4121 -6 4149 nw
tri 10344 4121 10372 4149 ne
rect 10372 4121 10430 4149
rect -92 2522 -40 4121
tri -40 4115 -34 4121 nw
rect 577 4069 583 4121
rect 635 4069 647 4121
rect 699 4069 705 4121
tri 619 4035 653 4069 ne
rect -92 2458 -40 2470
rect -92 1714 -40 2406
rect -92 1650 -40 1662
rect -92 1592 -40 1598
rect 653 3468 705 4069
rect 3449 4069 3455 4121
rect 3507 4069 3519 4121
rect 3571 4069 3577 4121
rect 3853 4069 3859 4121
rect 3911 4069 3926 4121
rect 3978 4069 4268 4121
rect 4320 4069 4332 4121
rect 4384 4069 5268 4121
tri 5268 4069 5320 4121 sw
tri 8085 4069 8137 4121 se
rect 8137 4069 8525 4121
rect 8577 4069 8589 4121
rect 8641 4069 8647 4121
rect 9759 4069 9765 4121
rect 9817 4069 9829 4121
rect 9881 4069 9887 4121
tri 10372 4115 10378 4121 ne
rect 653 3398 705 3416
rect 653 728 705 3346
rect 1412 3954 1612 3960
rect 1464 3902 1486 3954
rect 1538 3902 1560 3954
rect 1412 3885 1612 3902
rect 1464 3833 1486 3885
rect 1538 3833 1560 3885
rect 1412 3816 1612 3833
rect 1464 3764 1486 3816
rect 1538 3764 1560 3816
rect 1112 2961 1312 2962
rect 1112 2909 1118 2961
rect 1170 2909 1186 2961
rect 1238 2909 1254 2961
rect 1306 2909 1312 2961
rect 1112 2889 1312 2909
rect 1112 2837 1118 2889
rect 1170 2837 1186 2889
rect 1238 2837 1254 2889
rect 1306 2837 1312 2889
rect 1112 2817 1312 2837
rect 1112 2765 1118 2817
rect 1170 2765 1186 2817
rect 1238 2765 1254 2817
rect 1306 2765 1312 2817
rect 1112 1309 1312 2765
rect 1112 1257 1118 1309
rect 1170 1257 1186 1309
rect 1238 1257 1254 1309
rect 1306 1257 1312 1309
rect 1112 1237 1312 1257
rect 1112 1185 1118 1237
rect 1170 1185 1186 1237
rect 1238 1185 1254 1237
rect 1306 1185 1312 1237
rect 1112 1165 1312 1185
rect 1112 1113 1118 1165
rect 1170 1113 1186 1165
rect 1238 1113 1254 1165
rect 1306 1113 1312 1165
rect 1112 1112 1312 1113
rect 653 658 705 676
rect 653 600 705 606
rect 1412 310 1612 3764
rect 3449 3468 3501 4069
tri 3501 4035 3535 4069 nw
tri 5246 4047 5268 4069 ne
rect 5268 4061 5320 4069
tri 5320 4061 5328 4069 sw
tri 8077 4061 8085 4069 se
rect 8085 4061 8151 4069
tri 8151 4061 8159 4069 nw
tri 9801 4061 9809 4069 ne
rect 9809 4061 9887 4069
rect 5268 4047 8099 4061
tri 5268 4035 5280 4047 ne
rect 5280 4035 8099 4047
tri 5280 4009 5306 4035 ne
rect 5306 4009 8099 4035
tri 8099 4009 8151 4061 nw
tri 9809 4035 9835 4061 ne
rect 8956 3954 9156 3960
rect 9008 3902 9030 3954
rect 9082 3902 9104 3954
rect 8956 3885 9156 3902
rect 9008 3833 9030 3885
rect 9082 3833 9104 3885
rect 8956 3816 9156 3833
rect 9008 3764 9030 3816
rect 9082 3764 9104 3816
rect 3836 3724 3964 3730
rect 3888 3672 3912 3724
rect 3836 3658 3964 3672
rect 3888 3606 3912 3658
rect 3836 3565 3964 3606
rect 4182 3718 8345 3724
rect 4234 3672 8293 3718
rect 4234 3666 4262 3672
tri 4262 3666 4268 3672 nw
tri 8259 3666 8265 3672 ne
rect 8265 3666 8293 3672
rect 4182 3658 4254 3666
tri 4254 3658 4262 3666 nw
tri 8265 3658 8273 3666 ne
rect 8273 3658 8345 3666
rect 4182 3654 4250 3658
tri 4250 3654 4254 3658 nw
tri 8273 3654 8277 3658 ne
rect 8277 3654 8345 3658
tri 4234 3638 4250 3654 nw
tri 8277 3638 8293 3654 ne
rect 4182 3596 4234 3602
rect 8293 3596 8345 3602
rect 3449 3398 3501 3416
rect 3449 728 3501 3346
rect 3836 1949 3964 2102
rect 3996 1305 4154 1311
rect 4048 1253 4102 1305
rect 3996 1238 4154 1253
rect 4048 1186 4102 1238
rect 3996 1170 4154 1186
rect 4048 1118 4102 1170
rect 4182 1263 4440 1269
rect 4234 1211 4388 1263
rect 4182 1199 4440 1211
rect 4234 1147 4388 1199
rect 4182 1141 4440 1147
rect 3996 846 4154 1118
tri 4154 846 4194 886 sw
rect 3996 844 4661 846
rect 3996 822 4348 844
tri 3996 792 4026 822 ne
rect 4026 792 4348 822
rect 4400 792 4433 844
rect 4485 792 4518 844
rect 4570 792 4603 844
rect 4655 792 4661 844
tri 4026 740 4078 792 ne
rect 4078 740 4661 792
tri 4078 688 4130 740 ne
rect 4130 688 4348 740
rect 4400 688 4433 740
rect 4485 688 4518 740
rect 4570 688 4603 740
rect 4655 688 4661 740
rect 3449 658 3501 676
rect 3449 600 3501 606
rect 3836 468 3964 509
rect 3888 416 3912 468
rect 3836 402 3964 416
rect 3888 350 3912 402
rect 3836 344 3964 350
rect 1464 258 1486 310
rect 1538 258 1560 310
rect 1412 241 1612 258
rect 1464 189 1486 241
rect 1538 189 1560 241
rect 1412 172 1612 189
rect 1464 120 1486 172
rect 1538 120 1560 172
rect 1412 114 1612 120
rect 8956 310 9156 3764
rect 9835 3468 9887 4061
rect 10222 3724 10350 3730
rect 10274 3672 10298 3724
rect 10222 3658 10350 3672
rect 10274 3606 10298 3658
rect 10222 3558 10350 3606
rect 9835 3398 9887 3416
rect 9835 728 9887 3346
rect 10378 2463 10430 4121
rect 10378 2399 10430 2411
rect 10222 1983 10350 2096
rect 10378 1741 10430 2347
rect 10378 1677 10430 1689
rect 10378 1619 10430 1625
rect 10458 2956 10574 2962
rect 10510 2904 10522 2956
rect 10458 2889 10574 2904
rect 10510 2837 10522 2889
rect 10458 2821 10574 2837
rect 10510 2769 10522 2821
rect 10458 1305 10574 2769
rect 10510 1253 10522 1305
rect 10458 1238 10574 1253
rect 10510 1186 10522 1238
rect 10458 1170 10574 1186
rect 10510 1118 10522 1170
rect 10458 1112 10574 1118
rect 9835 658 9887 676
rect 9835 600 9887 606
rect 10222 468 10350 508
rect 10274 416 10298 468
rect 10222 402 10350 416
rect 10274 350 10298 402
rect 10222 344 10350 350
rect 9008 258 9030 310
rect 9082 258 9104 310
rect 8956 241 9156 258
rect 9008 189 9030 241
rect 9082 189 9104 241
rect 8956 172 9156 189
rect 9008 120 9030 172
rect 9082 120 9104 172
rect 8956 114 9156 120
use sky130_fd_io__com_ctl_ls  sky130_fd_io__com_ctl_ls_0
timestamp 1704896540
transform -1 0 2077 0 1 -10
box -71 10 2077 2019
use sky130_fd_io__com_ctl_ls  sky130_fd_io__com_ctl_ls_1
timestamp 1704896540
transform -1 0 2077 0 -1 4084
box -71 10 2077 2019
use sky130_fd_io__com_ctl_ls  sky130_fd_io__com_ctl_ls_2
timestamp 1704896540
transform 1 0 2077 0 -1 4084
box -71 10 2077 2019
use sky130_fd_io__com_ctl_ls  sky130_fd_io__com_ctl_ls_3
timestamp 1704896540
transform 1 0 8463 0 -1 4084
box -71 10 2077 2019
use sky130_fd_io__com_ctl_ls  sky130_fd_io__com_ctl_ls_4
timestamp 1704896540
transform 1 0 2077 0 1 -10
box -71 10 2077 2019
use sky130_fd_io__com_ctl_ls  sky130_fd_io__com_ctl_ls_5
timestamp 1704896540
transform 1 0 8463 0 1 -10
box -71 10 2077 2019
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_0
timestamp 1704896540
transform -1 0 4681 0 1 606
box 107 226 240 873
use sky130_fd_io__hvsbt_inv_x1  sky130_fd_io__hvsbt_inv_x1_1
timestamp 1704896540
transform 1 0 4499 0 1 606
box 107 226 240 873
use sky130_fd_io__hvsbt_nand2  sky130_fd_io__hvsbt_nand2_0
timestamp 1704896540
transform -1 0 5319 0 1 606
box 107 226 460 873
<< labels >>
flabel metal1 s 2398 957 2565 992 3 FreeSans 200 0 0 0 vrefgen_en_h_n
port 1 nsew
flabel metal1 s 2221 638 2363 664 3 FreeSans 200 0 0 0 vrefgen_en_h
port 2 nsew
flabel metal1 s 1161 1151 1349 1282 3 FreeSans 200 0 0 0 vssd
port 3 nsew
flabel metal1 s 9221 1151 9409 1282 3 FreeSans 200 0 0 0 vssd
port 3 nsew
flabel metal1 s 9256 3793 9599 3928 3 FreeSans 200 0 0 0 vddio_q
port 4 nsew
flabel metal1 s 2374 3793 2717 3928 3 FreeSans 200 0 0 0 vddio_q
port 4 nsew
flabel metal1 s 9332 2120 9704 2238 3 FreeSans 200 0 0 0 vccd
port 5 nsew
flabel metal1 s 2983 2120 3355 2238 3 FreeSans 200 0 0 0 vccd
port 5 nsew
flabel metal1 s 4352 1488 4634 1623 3 FreeSans 200 0 0 0 vddio_q
port 4 nsew
flabel metal1 s 4935 957 4979 1043 3 FreeSans 200 0 0 0 hld_h_n
port 6 nsew
flabel metal1 s 4500 964 4529 1026 3 FreeSans 200 0 0 0 enable_h
port 7 nsew
flabel metal1 s 8777 3084 8880 3117 3 FreeSans 200 0 0 0 selb_h<1>
port 9 nsew
flabel metal1 s 8782 960 8946 989 3 FreeSans 200 0 0 0 selb_h<0>
port 20 nsew
flabel metal1 s 8546 3406 8681 3438 3 FreeSans 200 0 0 0 sel_h<1>
port 12 nsew
flabel metal1 s 2146 3408 2248 3435 3 FreeSans 200 0 0 0 sel_h<2>
port 10 nsew
flabel metal1 s 8552 638 8662 669 3 FreeSans 200 0 0 0 sel_h<0>
port 13 nsew
flabel metal1 s 3779 673 3893 702 3 FreeSans 200 0 0 0 vrefgen_en
port 22 nsew
flabel metal1 s 10229 669 10306 701 3 FreeSans 200 0 0 0 sel<0>
port 23 nsew
flabel metal1 s 194 3376 294 3406 3 FreeSans 200 0 0 0 sel<3>
port 17 nsew
flabel metal1 s 10195 3368 10313 3402 3 FreeSans 200 0 0 0 sel<1>
port 14 nsew
flabel metal1 s 3811 3370 3951 3404 3 FreeSans 200 0 0 0 sel<2>
port 16 nsew
flabel metal1 s 1576 3085 1700 3118 3 FreeSans 200 0 0 0 selb_h<3>
port 18 nsew
flabel metal1 s 1589 956 1741 986 3 FreeSans 200 0 0 0 selb_h<4>
port 19 nsew
flabel metal1 s 1839 641 1973 673 3 FreeSans 200 0 0 0 sel_h<4>
port 21 nsew
flabel metal1 s 1783 3409 1923 3438 3 FreeSans 200 0 0 0 sel_h<3>
port 11 nsew
flabel metal1 s 225 667 347 704 3 FreeSans 200 0 0 0 sel<4>
port 15 nsew
flabel metal1 s 2381 3083 2512 3118 3 FreeSans 200 0 0 0 selb_h<2>
port 8 nsew
<< properties >>
string GDS_END 25922622
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 25895538
string path 246.525 15.000 246.525 18.350 
<< end >>
