magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect 1005 1982 1501 2714
rect 1127 1892 1501 1982
<< pwell >>
rect 1028 102 1114 432
rect 1327 356 1461 444
<< nsubdiff >>
rect 1041 2593 1091 2642
rect 1041 2570 1049 2593
rect 1083 2570 1091 2593
<< mvpsubdiff >>
rect 1054 382 1088 406
rect 1054 284 1088 348
rect 1353 416 1435 418
rect 1353 382 1377 416
rect 1411 382 1435 416
rect 1054 186 1088 250
rect 1054 128 1088 152
<< mvnsubdiff >>
rect 1041 2559 1049 2570
rect 1083 2559 1091 2570
rect 1041 2525 1091 2559
rect 1041 2491 1049 2525
rect 1083 2491 1091 2525
rect 1041 2457 1091 2491
rect 1041 2423 1049 2457
rect 1083 2423 1091 2457
rect 1041 2389 1091 2423
rect 1041 2355 1049 2389
rect 1083 2355 1091 2389
rect 1041 2321 1091 2355
rect 1041 2287 1049 2321
rect 1083 2287 1091 2321
rect 1041 2253 1091 2287
rect 1041 2219 1049 2253
rect 1083 2219 1091 2253
rect 1041 2185 1091 2219
rect 1041 2151 1049 2185
rect 1083 2151 1091 2185
rect 1041 2054 1091 2151
<< nsubdiffcont >>
rect 1049 2570 1083 2593
<< mvpsubdiffcont >>
rect 1054 348 1088 382
rect 1377 382 1411 416
rect 1054 250 1088 284
rect 1054 152 1088 186
<< mvnsubdiffcont >>
rect 1049 2559 1083 2570
rect 1049 2491 1083 2525
rect 1049 2423 1083 2457
rect 1049 2355 1083 2389
rect 1049 2287 1083 2321
rect 1049 2219 1083 2253
rect 1049 2151 1083 2185
<< poly >>
rect 162 2730 886 2746
rect 162 2696 178 2730
rect 212 2696 252 2730
rect 286 2696 325 2730
rect 359 2696 398 2730
rect 432 2696 471 2730
rect 505 2696 544 2730
rect 578 2696 617 2730
rect 651 2696 690 2730
rect 724 2696 763 2730
rect 797 2696 836 2730
rect 870 2696 886 2730
rect 162 2680 886 2696
rect 1239 2730 1373 2746
rect 1239 2696 1255 2730
rect 1289 2696 1323 2730
rect 1357 2696 1373 2730
rect 1239 2680 1373 2696
rect 1246 2674 1366 2680
rect 1246 334 1342 2022
rect 1246 76 1366 82
rect 162 54 886 70
rect 162 20 178 54
rect 212 20 252 54
rect 286 20 325 54
rect 359 20 398 54
rect 432 20 471 54
rect 505 20 544 54
rect 578 20 617 54
rect 651 20 690 54
rect 724 20 763 54
rect 797 20 836 54
rect 870 20 886 54
rect 162 4 886 20
rect 1239 60 1373 76
rect 1239 26 1255 60
rect 1289 26 1323 60
rect 1357 26 1373 60
rect 1239 10 1373 26
<< polycont >>
rect 178 2696 212 2730
rect 252 2696 286 2730
rect 325 2696 359 2730
rect 398 2696 432 2730
rect 471 2696 505 2730
rect 544 2696 578 2730
rect 617 2696 651 2730
rect 690 2696 724 2730
rect 763 2696 797 2730
rect 836 2696 870 2730
rect 1255 2696 1289 2730
rect 1323 2696 1357 2730
rect 178 20 212 54
rect 252 20 286 54
rect 325 20 359 54
rect 398 20 432 54
rect 471 20 505 54
rect 544 20 578 54
rect 617 20 651 54
rect 690 20 724 54
rect 763 20 797 54
rect 836 20 870 54
rect 1255 26 1289 60
rect 1323 26 1357 60
<< locali >>
rect 162 2696 178 2730
rect 213 2696 252 2730
rect 287 2696 325 2730
rect 361 2696 398 2730
rect 435 2696 471 2730
rect 509 2696 544 2730
rect 582 2696 617 2730
rect 655 2696 690 2730
rect 728 2696 763 2730
rect 801 2696 836 2730
rect 874 2696 886 2730
rect 1041 2593 1091 2827
rect 1255 2730 1357 2746
rect 1289 2696 1323 2730
rect 1255 2680 1357 2696
rect 77 1606 191 2586
rect 111 1572 157 1606
rect 77 1534 191 1572
rect 111 1500 157 1534
rect 77 130 191 1500
rect 267 2552 313 2586
rect 233 2514 347 2552
rect 267 2480 313 2514
rect 233 2442 347 2480
rect 267 2408 313 2442
rect 233 2369 347 2408
rect 267 2335 313 2369
rect 233 130 347 2335
rect 389 1606 503 2586
rect 423 1572 469 1606
rect 389 1534 503 1572
rect 423 1500 469 1534
rect 389 130 503 1500
rect 579 2552 625 2586
rect 545 2514 659 2552
rect 579 2480 625 2514
rect 545 2442 659 2480
rect 579 2408 625 2442
rect 545 2369 659 2408
rect 579 2335 625 2369
rect 545 130 659 2335
rect 701 1606 815 2586
rect 735 1572 781 1606
rect 701 1534 815 1572
rect 735 1500 781 1534
rect 701 130 815 1500
rect 891 2552 937 2586
rect 857 2514 971 2552
rect 891 2480 937 2514
rect 857 2442 971 2480
rect 891 2408 937 2442
rect 857 2369 971 2408
rect 891 2335 937 2369
rect 857 130 971 2335
rect 1041 2559 1049 2593
rect 1083 2559 1091 2593
rect 1041 2525 1091 2559
rect 1041 2491 1049 2525
rect 1083 2491 1091 2525
rect 1041 2457 1091 2491
rect 1041 2423 1049 2457
rect 1083 2423 1091 2457
rect 1041 2389 1091 2423
rect 1041 2355 1049 2389
rect 1083 2355 1091 2389
rect 1041 2321 1091 2355
rect 1041 2287 1049 2321
rect 1083 2287 1091 2321
rect 1041 2253 1091 2287
rect 1041 2200 1049 2253
rect 1083 2200 1091 2253
rect 1041 2185 1091 2200
rect 1041 2128 1049 2185
rect 1083 2128 1091 2185
rect 1041 2089 1091 2128
rect 1041 2055 1049 2089
rect 1083 2055 1091 2089
rect 1041 2054 1091 2055
rect 1201 2575 1235 2613
rect 1049 2016 1083 2054
rect 1054 394 1088 406
rect 1054 322 1088 348
rect 1054 284 1088 288
rect 1054 249 1088 250
rect 1054 186 1088 215
rect 1054 128 1088 142
rect 1201 110 1235 2541
rect 1269 76 1343 2680
rect 1377 2234 1411 2246
rect 1377 2162 1411 2200
rect 1377 2090 1411 2128
rect 1377 2044 1411 2056
rect 1377 416 1411 432
rect 1377 248 1411 286
rect 1377 176 1411 214
rect 1377 130 1411 142
rect 1255 60 1357 76
rect 162 20 170 54
rect 212 20 245 54
rect 286 20 320 54
rect 359 20 395 54
rect 432 20 470 54
rect 505 20 544 54
rect 578 20 617 54
rect 652 20 690 54
rect 726 20 763 54
rect 800 20 836 54
rect 874 20 886 54
rect 1289 26 1323 60
rect 1285 20 1323 26
rect 1255 10 1357 20
<< viali >>
rect 179 2696 212 2730
rect 212 2696 213 2730
rect 253 2696 286 2730
rect 286 2696 287 2730
rect 327 2696 359 2730
rect 359 2696 361 2730
rect 401 2696 432 2730
rect 432 2696 435 2730
rect 475 2696 505 2730
rect 505 2696 509 2730
rect 548 2696 578 2730
rect 578 2696 582 2730
rect 621 2696 651 2730
rect 651 2696 655 2730
rect 694 2696 724 2730
rect 724 2696 728 2730
rect 767 2696 797 2730
rect 797 2696 801 2730
rect 840 2696 870 2730
rect 870 2696 874 2730
rect 77 1572 111 1606
rect 157 1572 191 1606
rect 77 1500 111 1534
rect 157 1500 191 1534
rect 233 2552 267 2586
rect 313 2552 347 2586
rect 233 2480 267 2514
rect 313 2480 347 2514
rect 233 2408 267 2442
rect 313 2408 347 2442
rect 233 2335 267 2369
rect 313 2335 347 2369
rect 389 1572 423 1606
rect 469 1572 503 1606
rect 389 1500 423 1534
rect 469 1500 503 1534
rect 545 2552 579 2586
rect 625 2552 659 2586
rect 545 2480 579 2514
rect 625 2480 659 2514
rect 545 2408 579 2442
rect 625 2408 659 2442
rect 545 2335 579 2369
rect 625 2335 659 2369
rect 701 1572 735 1606
rect 781 1572 815 1606
rect 701 1500 735 1534
rect 781 1500 815 1534
rect 857 2552 891 2586
rect 937 2552 971 2586
rect 857 2480 891 2514
rect 937 2480 971 2514
rect 857 2408 891 2442
rect 937 2408 971 2442
rect 857 2335 891 2369
rect 937 2335 971 2369
rect 1049 2219 1083 2234
rect 1049 2200 1083 2219
rect 1049 2151 1083 2162
rect 1049 2128 1083 2151
rect 1049 2055 1083 2089
rect 1201 2613 1235 2647
rect 1201 2541 1235 2575
rect 1049 1982 1083 2016
rect 1054 382 1088 394
rect 1054 360 1088 382
rect 1054 288 1088 322
rect 1054 215 1088 249
rect 1054 152 1088 176
rect 1054 142 1088 152
rect 1377 2200 1411 2234
rect 1377 2128 1411 2162
rect 1377 2056 1411 2090
rect 1377 382 1411 400
rect 1377 366 1411 382
rect 1377 286 1411 320
rect 1377 214 1411 248
rect 1377 142 1411 176
rect 170 20 178 54
rect 178 20 204 54
rect 245 20 252 54
rect 252 20 279 54
rect 320 20 325 54
rect 325 20 354 54
rect 395 20 398 54
rect 398 20 429 54
rect 470 20 471 54
rect 471 20 504 54
rect 544 20 578 54
rect 618 20 651 54
rect 651 20 652 54
rect 692 20 724 54
rect 724 20 726 54
rect 766 20 797 54
rect 797 20 800 54
rect 840 20 870 54
rect 870 20 874 54
rect 1251 26 1255 54
rect 1255 26 1285 54
rect 1323 26 1357 54
rect 1251 20 1285 26
rect 1323 20 1357 26
<< metal1 >>
rect 167 2730 1241 2736
rect 167 2696 179 2730
rect 213 2696 253 2730
rect 287 2696 327 2730
rect 361 2696 401 2730
rect 435 2696 475 2730
rect 509 2696 548 2730
rect 582 2696 621 2730
rect 655 2696 694 2730
rect 728 2696 767 2730
rect 801 2696 840 2730
rect 874 2696 1241 2730
rect 167 2690 1241 2696
tri 1133 2647 1176 2690 ne
rect 1176 2647 1241 2690
tri 1176 2628 1195 2647 ne
rect 1195 2613 1201 2647
rect 1235 2613 1241 2647
rect 227 2586 977 2598
rect 227 2552 233 2586
rect 267 2552 313 2586
rect 347 2552 545 2586
rect 579 2552 625 2586
rect 659 2552 857 2586
rect 891 2552 937 2586
rect 971 2552 977 2586
rect 227 2514 977 2552
rect 1195 2575 1241 2613
rect 1195 2541 1201 2575
rect 1235 2541 1241 2575
rect 1195 2529 1241 2541
rect 227 2480 233 2514
rect 267 2480 313 2514
rect 347 2480 545 2514
rect 579 2480 625 2514
rect 659 2480 857 2514
rect 891 2480 937 2514
rect 971 2480 977 2514
rect 227 2442 977 2480
rect 227 2408 233 2442
rect 267 2408 313 2442
rect 347 2408 545 2442
rect 579 2408 625 2442
rect 659 2408 857 2442
rect 891 2408 937 2442
rect 971 2408 977 2442
rect 227 2369 977 2408
rect 227 2335 233 2369
rect 267 2335 313 2369
rect 347 2335 545 2369
rect 579 2335 625 2369
rect 659 2335 857 2369
rect 891 2335 937 2369
rect 971 2335 977 2369
rect 227 2323 977 2335
rect 1041 2234 1423 2246
rect 1041 2200 1049 2234
rect 1083 2200 1377 2234
rect 1411 2200 1423 2234
rect 1041 2162 1423 2200
rect 1041 2128 1049 2162
rect 1083 2128 1377 2162
rect 1411 2128 1423 2162
rect 1041 2090 1423 2128
rect 1041 2089 1377 2090
rect 1041 2055 1049 2089
rect 1083 2056 1377 2089
rect 1411 2056 1423 2090
rect 1083 2055 1423 2056
rect 1041 2016 1423 2055
rect 1041 1982 1049 2016
rect 1083 1982 1423 2016
rect 1041 1970 1423 1982
rect 71 1606 821 1618
rect 71 1572 77 1606
rect 111 1572 157 1606
rect 191 1572 389 1606
rect 423 1572 469 1606
rect 503 1572 701 1606
rect 735 1572 781 1606
rect 815 1572 821 1606
rect 71 1534 821 1572
rect 71 1500 77 1534
rect 111 1500 157 1534
rect 191 1500 389 1534
rect 423 1500 469 1534
rect 503 1500 701 1534
rect 735 1500 781 1534
rect 815 1500 821 1534
rect 71 1488 821 1500
rect 1048 400 1423 406
rect 1048 394 1377 400
rect 1048 360 1054 394
rect 1088 366 1377 394
rect 1411 366 1423 400
rect 1088 360 1423 366
rect 1048 322 1423 360
rect 1048 288 1054 322
rect 1088 320 1423 322
rect 1088 288 1377 320
rect 1048 286 1377 288
rect 1411 286 1423 320
rect 1048 249 1423 286
rect 1048 215 1054 249
rect 1088 248 1423 249
rect 1088 215 1377 248
rect 1048 214 1377 215
rect 1411 214 1423 248
rect 1048 176 1423 214
rect 1048 142 1054 176
rect 1088 142 1377 176
rect 1411 142 1423 176
rect 1048 130 1423 142
rect 158 54 1369 60
rect 158 20 170 54
rect 204 20 245 54
rect 279 20 320 54
rect 354 20 395 54
rect 429 20 470 54
rect 504 20 544 54
rect 578 20 618 54
rect 652 20 692 54
rect 726 20 766 54
rect 800 20 840 54
rect 874 20 1251 54
rect 1285 20 1323 54
rect 1357 20 1369 54
rect 158 14 1369 20
use hvnTran_CDNS_52468879185404  hvnTran_CDNS_52468879185404_0
timestamp 1704896540
transform -1 0 1366 0 -1 308
box -79 -26 199 226
use hvpTran_CDNS_52468879185406  hvpTran_CDNS_52468879185406_0
timestamp 1704896540
transform -1 0 1366 0 1 2048
box -119 -66 239 666
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1704896540
transform 0 1 1377 -1 0 320
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_1
timestamp 1704896540
transform 0 1 1377 1 0 2056
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_0
timestamp 1704896540
transform -1 0 1411 0 -1 400
box 0 0 1 1
use nfet_CDNS_52468879185937  nfet_CDNS_52468879185937_0
timestamp 1704896540
transform 1 0 162 0 -1 396
box -79 -26 803 326
use pfet_CDNS_52468879185936  pfet_CDNS_52468879185936_0
timestamp 1704896540
transform 1 0 162 0 1 2048
box -119 -66 843 666
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_0
timestamp 1704896540
transform 1 0 1239 0 -1 2746
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_1
timestamp 1704896540
transform 1 0 1239 0 1 10
box 0 0 1 1
<< labels >>
flabel metal1 s 1047 2705 1047 2705 0 FreeSans 200 0 0 0 sel_b
flabel metal1 s 1118 221 1196 302 0 FreeSans 200 0 0 0 vgnd
port 1 nsew
flabel metal1 s 1129 2088 1245 2150 0 FreeSans 200 0 0 0 vcc_io
port 2 nsew
flabel metal1 s 401 2423 494 2514 0 FreeSans 200 0 0 0 out
port 3 nsew
flabel metal1 s 1023 14 1086 60 0 FreeSans 200 0 0 0 sel
port 4 nsew
flabel metal1 s 213 1516 375 1595 0 FreeSans 200 0 0 0 in
port 5 nsew
<< properties >>
string GDS_END 80606504
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 80594926
string path 26.650 66.075 26.650 51.325 
<< end >>
