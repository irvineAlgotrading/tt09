magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -38 261 1418 582
<< pwell >>
rect 1 21 1303 203
rect 30 -17 64 21
<< locali >>
rect 975 325 1025 425
rect 1143 325 1193 425
rect 1311 325 1352 483
rect 975 291 1352 325
rect 22 215 89 257
rect 207 215 538 257
rect 607 215 860 257
rect 1284 181 1352 291
rect 191 145 1352 181
rect 191 51 257 145
rect 359 51 425 145
rect 631 51 697 145
rect 799 51 865 145
rect 967 51 1033 145
rect 1135 51 1201 145
rect 1303 63 1352 145
<< obsli1 >>
rect 0 527 1380 561
rect 22 325 81 493
rect 115 359 165 527
rect 199 393 249 493
rect 283 427 333 527
rect 367 393 417 493
rect 451 427 501 527
rect 555 459 1277 493
rect 555 427 605 459
rect 723 427 773 459
rect 639 393 689 425
rect 807 393 857 425
rect 199 359 857 393
rect 891 359 941 459
rect 1059 359 1109 459
rect 1227 359 1277 459
rect 22 291 941 325
rect 123 181 157 291
rect 907 257 941 291
rect 907 215 1225 257
rect 22 147 157 181
rect 22 51 89 147
rect 123 17 157 111
rect 291 17 325 111
rect 459 17 597 111
rect 731 17 765 111
rect 899 17 933 111
rect 1067 17 1101 111
rect 1235 17 1269 111
rect 0 -17 1380 17
<< metal1 >>
rect 0 496 1380 592
rect 0 -48 1380 48
<< labels >>
rlabel locali s 207 215 538 257 6 A
port 1 nsew signal input
rlabel locali s 607 215 860 257 6 B
port 2 nsew signal input
rlabel locali s 22 215 89 257 6 C_N
port 3 nsew signal input
rlabel metal1 s 0 -48 1380 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 21 1303 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 1418 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 1380 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1303 63 1352 145 6 Y
port 8 nsew signal output
rlabel locali s 1135 51 1201 145 6 Y
port 8 nsew signal output
rlabel locali s 967 51 1033 145 6 Y
port 8 nsew signal output
rlabel locali s 799 51 865 145 6 Y
port 8 nsew signal output
rlabel locali s 631 51 697 145 6 Y
port 8 nsew signal output
rlabel locali s 359 51 425 145 6 Y
port 8 nsew signal output
rlabel locali s 191 51 257 145 6 Y
port 8 nsew signal output
rlabel locali s 191 145 1352 181 6 Y
port 8 nsew signal output
rlabel locali s 1284 181 1352 291 6 Y
port 8 nsew signal output
rlabel locali s 975 291 1352 325 6 Y
port 8 nsew signal output
rlabel locali s 1311 325 1352 483 6 Y
port 8 nsew signal output
rlabel locali s 1143 325 1193 425 6 Y
port 8 nsew signal output
rlabel locali s 975 325 1025 425 6 Y
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1380 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1123316
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1113216
<< end >>
