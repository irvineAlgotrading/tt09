magic
tech sky130B
magscale 1 2
timestamp 1704896540
use sky130_fd_pr__hvdfl1sd__example_55959141808122  sky130_fd_pr__hvdfl1sd__example_55959141808122_0
timestamp 1704896540
transform -1 0 -18 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd__example_55959141808452  sky130_fd_pr__hvdfm1sd__example_55959141808452_0
timestamp 1704896540
transform 1 0 100 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 22078598
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 22077480
<< end >>
