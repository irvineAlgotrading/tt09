magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< pwell >>
rect -76 -26 876 2026
<< mvnnmos >>
rect 0 0 800 2000
<< mvndiff >>
rect -50 0 0 2000
rect 800 0 850 2000
<< poly >>
rect 0 2000 800 2026
rect 0 -26 800 0
<< locali >>
rect -45 -4 -11 1966
rect 811 -4 845 1966
use DFL1sd_CDNS_52468879185709  DFL1sd_CDNS_52468879185709_0
timestamp 1704896540
transform 1 0 800 0 1 0
box -26 -26 79 2026
use hvDFL1sd_CDNS_52468879185990  hvDFL1sd_CDNS_52468879185990_0
timestamp 1704896540
transform -1 0 0 0 1 0
box -26 -26 79 2026
<< labels >>
flabel comment s -28 981 -28 981 0 FreeSans 300 0 0 0 S
flabel comment s 828 981 828 981 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 96486774
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 96485822
<< end >>
