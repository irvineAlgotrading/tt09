magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect 37 3488 661 4329
<< pwell >>
rect -28 1922 1320 2008
rect -28 100 58 1922
rect 1234 100 1320 1922
rect -28 14 1320 100
<< mvpsubdiff >>
rect -2 1948 104 1982
rect 138 1948 172 1982
rect 206 1948 240 1982
rect 274 1948 308 1982
rect 342 1948 376 1982
rect 410 1948 444 1982
rect 478 1948 512 1982
rect 546 1948 580 1982
rect 614 1948 648 1982
rect 682 1948 716 1982
rect 750 1948 784 1982
rect 818 1948 852 1982
rect 886 1948 920 1982
rect 954 1948 988 1982
rect 1022 1948 1056 1982
rect 1090 1948 1124 1982
rect 1158 1948 1192 1982
rect 1226 1948 1294 1982
rect -2 1914 32 1948
rect 1260 1910 1294 1948
rect -2 1846 32 1880
rect 1260 1842 1294 1876
rect -2 1778 32 1812
rect -2 1710 32 1744
rect -2 1642 32 1676
rect -2 1574 32 1608
rect -2 1506 32 1540
rect -2 1438 32 1472
rect -2 1370 32 1404
rect -2 1302 32 1336
rect -2 1234 32 1268
rect -2 1166 32 1200
rect -2 1098 32 1132
rect -2 1030 32 1064
rect -2 962 32 996
rect -2 894 32 928
rect -2 826 32 860
rect 1260 1774 1294 1808
rect 1260 1706 1294 1740
rect 1260 1638 1294 1672
rect 1260 1570 1294 1604
rect 1260 1502 1294 1536
rect 1260 1434 1294 1468
rect 1260 1366 1294 1400
rect 1260 1298 1294 1332
rect 1260 1230 1294 1264
rect 1260 1162 1294 1196
rect 1260 1094 1294 1128
rect 1260 1026 1294 1060
rect 1260 958 1294 992
rect 1260 890 1294 924
rect -2 758 32 792
rect 1260 822 1294 856
rect -2 690 32 724
rect -2 622 32 656
rect -2 554 32 588
rect -2 486 32 520
rect 1260 754 1294 788
rect 1260 686 1294 720
rect 1260 618 1294 652
rect 1260 550 1294 584
rect 1260 482 1294 516
rect -2 418 32 452
rect 1260 414 1294 448
rect -2 350 32 384
rect -2 282 32 316
rect -2 214 32 248
rect -2 74 32 180
rect 1260 346 1294 380
rect 1260 278 1294 312
rect 1260 210 1294 244
rect 1260 142 1294 176
rect 1260 74 1294 108
rect -2 40 66 74
rect 100 40 134 74
rect 168 40 202 74
rect 236 40 270 74
rect 304 40 338 74
rect 372 40 406 74
rect 440 40 474 74
rect 508 40 542 74
rect 576 40 610 74
rect 644 40 678 74
rect 712 40 746 74
rect 780 40 814 74
rect 848 40 882 74
rect 916 40 950 74
rect 984 40 1018 74
rect 1052 40 1086 74
rect 1120 40 1154 74
rect 1188 40 1294 74
<< mvnsubdiff >>
rect 104 4228 138 4262
rect 172 4228 206 4262
rect 240 4228 274 4262
rect 308 4228 342 4262
rect 376 4228 410 4262
rect 444 4228 478 4262
rect 512 4228 594 4262
<< mvpsubdiffcont >>
rect 104 1948 138 1982
rect 172 1948 206 1982
rect 240 1948 274 1982
rect 308 1948 342 1982
rect 376 1948 410 1982
rect 444 1948 478 1982
rect 512 1948 546 1982
rect 580 1948 614 1982
rect 648 1948 682 1982
rect 716 1948 750 1982
rect 784 1948 818 1982
rect 852 1948 886 1982
rect 920 1948 954 1982
rect 988 1948 1022 1982
rect 1056 1948 1090 1982
rect 1124 1948 1158 1982
rect 1192 1948 1226 1982
rect -2 1880 32 1914
rect -2 1812 32 1846
rect 1260 1876 1294 1910
rect -2 1744 32 1778
rect -2 1676 32 1710
rect -2 1608 32 1642
rect -2 1540 32 1574
rect -2 1472 32 1506
rect -2 1404 32 1438
rect -2 1336 32 1370
rect -2 1268 32 1302
rect -2 1200 32 1234
rect -2 1132 32 1166
rect -2 1064 32 1098
rect -2 996 32 1030
rect -2 928 32 962
rect -2 860 32 894
rect 1260 1808 1294 1842
rect 1260 1740 1294 1774
rect 1260 1672 1294 1706
rect 1260 1604 1294 1638
rect 1260 1536 1294 1570
rect 1260 1468 1294 1502
rect 1260 1400 1294 1434
rect 1260 1332 1294 1366
rect 1260 1264 1294 1298
rect 1260 1196 1294 1230
rect 1260 1128 1294 1162
rect 1260 1060 1294 1094
rect 1260 992 1294 1026
rect 1260 924 1294 958
rect 1260 856 1294 890
rect -2 792 32 826
rect 1260 788 1294 822
rect -2 724 32 758
rect -2 656 32 690
rect -2 588 32 622
rect -2 520 32 554
rect -2 452 32 486
rect 1260 720 1294 754
rect 1260 652 1294 686
rect 1260 584 1294 618
rect 1260 516 1294 550
rect -2 384 32 418
rect 1260 448 1294 482
rect -2 316 32 350
rect -2 248 32 282
rect -2 180 32 214
rect 1260 380 1294 414
rect 1260 312 1294 346
rect 1260 244 1294 278
rect 1260 176 1294 210
rect 1260 108 1294 142
rect 66 40 100 74
rect 134 40 168 74
rect 202 40 236 74
rect 270 40 304 74
rect 338 40 372 74
rect 406 40 440 74
rect 474 40 508 74
rect 542 40 576 74
rect 610 40 644 74
rect 678 40 712 74
rect 746 40 780 74
rect 814 40 848 74
rect 882 40 916 74
rect 950 40 984 74
rect 1018 40 1052 74
rect 1086 40 1120 74
rect 1154 40 1188 74
<< mvnsubdiffcont >>
rect 138 4228 172 4262
rect 206 4228 240 4262
rect 274 4228 308 4262
rect 342 4228 376 4262
rect 410 4228 444 4262
rect 478 4228 512 4262
<< poly >>
rect 122 3956 256 3972
rect 122 3922 138 3956
rect 172 3922 206 3956
rect 240 3922 256 3956
rect 122 3906 256 3922
rect 156 3786 290 3802
rect 156 3752 172 3786
rect 206 3752 240 3786
rect 274 3752 290 3786
rect 156 3736 290 3752
rect 203 1872 609 1888
rect 203 1838 219 1872
rect 253 1838 287 1872
rect 321 1838 355 1872
rect 389 1838 423 1872
rect 457 1838 491 1872
rect 525 1838 559 1872
rect 593 1838 609 1872
rect 203 1822 609 1838
rect 651 1872 785 1888
rect 651 1838 667 1872
rect 701 1838 735 1872
rect 769 1838 785 1872
rect 651 1822 785 1838
rect 203 836 1091 852
rect 203 802 219 836
rect 253 802 287 836
rect 321 802 355 836
rect 389 802 423 836
rect 457 802 491 836
rect 525 802 559 836
rect 593 802 627 836
rect 661 802 696 836
rect 730 802 765 836
rect 799 802 834 836
rect 868 802 903 836
rect 937 802 972 836
rect 1006 802 1041 836
rect 1075 802 1091 836
rect 203 786 1091 802
rect 203 442 491 458
rect 203 408 219 442
rect 253 408 293 442
rect 327 408 367 442
rect 401 408 441 442
rect 475 408 491 442
rect 203 392 491 408
rect 547 442 835 458
rect 547 408 563 442
rect 597 408 637 442
rect 671 408 711 442
rect 745 408 785 442
rect 819 408 835 442
rect 547 392 835 408
<< polycont >>
rect 138 3922 172 3956
rect 206 3922 240 3956
rect 172 3752 206 3786
rect 240 3752 274 3786
rect 219 1838 253 1872
rect 287 1838 321 1872
rect 355 1838 389 1872
rect 423 1838 457 1872
rect 491 1838 525 1872
rect 559 1838 593 1872
rect 667 1838 701 1872
rect 735 1838 769 1872
rect 219 802 253 836
rect 287 802 321 836
rect 355 802 389 836
rect 423 802 457 836
rect 491 802 525 836
rect 559 802 593 836
rect 627 802 661 836
rect 696 802 730 836
rect 765 802 799 836
rect 834 802 868 836
rect 903 802 937 836
rect 972 802 1006 836
rect 1041 802 1075 836
rect 219 408 253 442
rect 293 408 327 442
rect 367 408 401 442
rect 441 408 475 442
rect 563 408 597 442
rect 637 408 671 442
rect 711 408 745 442
rect 785 408 819 442
<< locali >>
rect 172 4228 178 4262
rect 240 4228 252 4262
rect 308 4228 326 4262
rect 376 4228 400 4262
rect 444 4228 474 4262
rect 512 4228 548 4262
rect 582 4228 594 4262
rect 111 4050 145 4088
rect 267 4050 301 4088
rect 149 3956 187 3957
rect 172 3923 187 3956
rect 122 3922 138 3923
rect 172 3922 206 3923
rect 240 3922 256 3956
rect 156 3752 172 3786
rect 227 3752 240 3786
rect 111 3620 145 3658
rect 267 3600 301 3638
rect -8 1982 1300 1988
rect -8 1948 70 1982
rect 138 1948 142 1982
rect 206 1948 215 1982
rect 274 1948 288 1982
rect 342 1948 361 1982
rect 410 1948 444 1982
rect 505 1948 512 1982
rect 546 1948 550 1982
rect 614 1948 629 1982
rect 682 1948 708 1982
rect 750 1948 784 1982
rect 822 1948 852 1982
rect 902 1948 920 1982
rect 982 1948 988 1982
rect 1022 1948 1028 1982
rect 1090 1948 1108 1982
rect 1158 1948 1188 1982
rect 1226 1948 1300 1982
rect -8 1942 1300 1948
rect -8 1914 38 1942
rect -8 1876 -2 1914
rect 32 1876 38 1914
rect -8 1846 38 1876
rect 1254 1910 1300 1942
rect 1254 1875 1260 1910
rect 1294 1875 1300 1910
rect -8 1802 -2 1846
rect 32 1802 38 1846
rect 203 1838 219 1872
rect 272 1838 287 1872
rect 351 1838 355 1872
rect 389 1838 397 1872
rect 457 1838 477 1872
rect 525 1838 557 1872
rect 593 1838 609 1872
rect 651 1838 667 1872
rect 701 1838 735 1872
rect 773 1838 785 1872
rect 1254 1842 1300 1875
rect -8 1778 38 1802
rect -8 1728 -2 1778
rect 32 1728 38 1778
rect -8 1710 38 1728
rect 1254 1802 1260 1842
rect 1294 1802 1300 1842
rect 1254 1774 1300 1802
rect 1254 1729 1260 1774
rect 1294 1729 1300 1774
rect -8 1654 -2 1710
rect 32 1654 38 1710
rect -8 1642 38 1654
rect -8 1580 -2 1642
rect 32 1580 38 1642
rect -8 1574 38 1580
rect -8 1472 -2 1574
rect 32 1472 38 1574
rect -8 1466 38 1472
rect -8 1404 -2 1466
rect 32 1404 38 1466
rect -8 1392 38 1404
rect -8 1336 -2 1392
rect 32 1336 38 1392
rect -8 1318 38 1336
rect -8 1268 -2 1318
rect 32 1268 38 1318
rect -8 1244 38 1268
rect -8 1200 -2 1244
rect 32 1200 38 1244
rect -8 1170 38 1200
rect 158 1635 192 1682
rect 158 1554 192 1601
rect 158 1473 192 1520
rect 158 1392 192 1439
rect 158 1312 192 1358
rect 158 1232 192 1278
rect 334 1635 368 1682
rect 334 1554 368 1601
rect 334 1473 368 1520
rect 334 1392 368 1439
rect 334 1312 368 1358
rect 334 1232 368 1278
rect 444 1635 478 1682
rect 444 1554 478 1601
rect 444 1473 478 1520
rect 444 1392 478 1439
rect 444 1312 478 1358
rect 444 1232 478 1278
rect 620 1635 654 1682
rect 620 1554 654 1601
rect 620 1473 654 1520
rect 620 1392 654 1439
rect 620 1312 654 1358
rect 620 1232 654 1278
rect 796 1635 830 1682
rect 796 1554 830 1601
rect 796 1473 830 1520
rect 796 1392 830 1439
rect 796 1312 830 1358
rect 796 1232 830 1278
rect 1254 1706 1300 1729
rect 1254 1656 1260 1706
rect 1294 1656 1300 1706
rect 1254 1638 1300 1656
rect 1254 1583 1260 1638
rect 1294 1583 1300 1638
rect 1254 1570 1300 1583
rect 1254 1510 1260 1570
rect 1294 1510 1300 1570
rect 1254 1502 1300 1510
rect 1254 1437 1260 1502
rect 1294 1437 1300 1502
rect 1254 1434 1300 1437
rect 1254 1400 1260 1434
rect 1294 1400 1300 1434
rect 1254 1398 1300 1400
rect 1254 1332 1260 1398
rect 1294 1332 1300 1398
rect 1254 1324 1300 1332
rect 1254 1264 1260 1324
rect 1294 1264 1300 1324
rect 1254 1250 1300 1264
rect -8 1132 -2 1170
rect 32 1132 38 1170
rect -8 1098 38 1132
rect -8 1062 -2 1098
rect 32 1062 38 1098
rect 1254 1196 1260 1250
rect 1294 1196 1300 1250
rect 1254 1176 1300 1196
rect 1254 1128 1260 1176
rect 1294 1128 1300 1176
rect 1254 1102 1300 1128
rect -8 1030 38 1062
rect -8 989 -2 1030
rect 32 989 38 1030
rect -8 962 38 989
rect 158 1010 192 1048
rect 630 1010 664 1048
rect -8 916 -2 962
rect 32 916 38 962
rect -8 894 38 916
rect 1102 1010 1136 1048
rect 394 930 428 968
rect 1254 1060 1260 1102
rect 1294 1060 1300 1102
rect 1254 1028 1300 1060
rect 1254 992 1260 1028
rect 1294 992 1300 1028
rect 866 930 900 968
rect 1254 958 1300 992
rect 1254 920 1260 958
rect 1294 920 1300 958
rect -8 843 -2 894
rect 32 843 38 894
rect -8 826 38 843
rect 1254 890 1300 920
rect 1254 846 1260 890
rect 1294 846 1300 890
rect -8 770 -2 826
rect 32 770 38 826
rect 203 802 219 836
rect 253 802 276 836
rect 321 802 355 836
rect 389 802 423 836
rect 468 802 491 836
rect 547 802 559 836
rect 626 802 627 836
rect 661 802 671 836
rect 730 802 751 836
rect 799 802 831 836
rect 868 802 903 836
rect 945 802 972 836
rect 1025 802 1041 836
rect 1075 802 1091 836
rect 1254 822 1300 846
rect -8 758 38 770
rect -8 697 -2 758
rect 32 697 38 758
rect 1254 772 1260 822
rect 1294 772 1300 822
rect 1254 754 1300 772
rect -8 690 38 697
rect -8 624 -2 690
rect 32 624 38 690
rect 394 680 428 718
rect -8 622 38 624
rect -8 588 -2 622
rect 32 588 38 622
rect -8 585 38 588
rect -8 520 -2 585
rect 32 520 38 585
rect 866 680 900 718
rect 158 600 192 638
rect 1254 698 1260 754
rect 1294 698 1300 754
rect 1254 686 1300 698
rect 630 600 664 638
rect 1254 660 1260 686
rect 1102 600 1136 638
rect 1294 660 1300 686
rect 1260 618 1294 652
rect -8 512 38 520
rect -8 452 -2 512
rect 32 452 38 512
rect -8 439 38 452
rect 1260 550 1294 584
rect 1260 482 1294 516
rect -8 384 -2 439
rect 32 384 38 439
rect 203 408 219 442
rect 286 408 293 442
rect 327 408 328 442
rect 362 408 367 442
rect 401 408 404 442
rect 438 408 441 442
rect 475 408 491 442
rect 547 408 563 442
rect 616 408 637 442
rect 692 408 711 442
rect 768 408 785 442
rect 819 408 835 442
rect 1260 414 1294 448
rect -8 366 38 384
rect -8 316 -2 366
rect 32 316 38 366
rect 1254 380 1260 389
rect 1294 380 1300 389
rect -8 293 38 316
rect -8 248 -2 293
rect 32 248 38 293
rect 244 283 278 321
rect -8 220 38 248
rect -8 180 -2 220
rect 32 180 38 220
rect -8 147 38 180
rect 416 283 450 321
rect 158 190 192 228
rect 588 283 622 321
rect 330 190 364 228
rect 760 283 794 321
rect 502 190 536 228
rect 1254 351 1300 380
rect 1254 312 1260 351
rect 1294 312 1300 351
rect 1254 278 1300 312
rect 674 190 708 228
rect 846 190 880 228
rect 1254 215 1260 278
rect 1294 215 1300 278
rect 1254 210 1300 215
rect 1254 176 1260 210
rect 1294 176 1300 210
rect -8 113 -2 147
rect 32 113 38 147
rect -8 80 38 113
rect 1254 146 1300 176
rect 1254 108 1260 146
rect 1294 108 1300 146
rect 1254 80 1300 108
rect -8 74 1300 80
rect -8 40 66 74
rect 104 40 134 74
rect 179 40 202 74
rect 254 40 270 74
rect 329 40 338 74
rect 404 40 406 74
rect 440 40 445 74
rect 508 40 520 74
rect 576 40 594 74
rect 644 40 668 74
rect 712 40 742 74
rect 780 40 814 74
rect 850 40 882 74
rect 924 40 950 74
rect 998 40 1018 74
rect 1072 40 1086 74
rect 1146 40 1154 74
rect 1220 40 1300 74
rect -8 34 1300 40
<< viali >>
rect 104 4228 138 4262
rect 178 4228 206 4262
rect 206 4228 212 4262
rect 252 4228 274 4262
rect 274 4228 286 4262
rect 326 4228 342 4262
rect 342 4228 360 4262
rect 400 4228 410 4262
rect 410 4228 434 4262
rect 474 4228 478 4262
rect 478 4228 508 4262
rect 548 4228 582 4262
rect 111 4088 145 4122
rect 111 4016 145 4050
rect 267 4088 301 4122
rect 267 4016 301 4050
rect 115 3956 149 3957
rect 187 3956 221 3957
rect 115 3923 138 3956
rect 138 3923 149 3956
rect 187 3923 206 3956
rect 206 3923 221 3956
rect 193 3752 206 3786
rect 206 3752 227 3786
rect 265 3752 274 3786
rect 274 3752 299 3786
rect 111 3658 145 3692
rect 111 3586 145 3620
rect 267 3638 301 3672
rect 267 3566 301 3600
rect 70 1948 104 1982
rect 142 1948 172 1982
rect 172 1948 176 1982
rect 215 1948 240 1982
rect 240 1948 249 1982
rect 288 1948 308 1982
rect 308 1948 322 1982
rect 361 1948 376 1982
rect 376 1948 395 1982
rect 471 1948 478 1982
rect 478 1948 505 1982
rect 550 1948 580 1982
rect 580 1948 584 1982
rect 629 1948 648 1982
rect 648 1948 663 1982
rect 708 1948 716 1982
rect 716 1948 742 1982
rect 788 1948 818 1982
rect 818 1948 822 1982
rect 868 1948 886 1982
rect 886 1948 902 1982
rect 948 1948 954 1982
rect 954 1948 982 1982
rect 1028 1948 1056 1982
rect 1056 1948 1062 1982
rect 1108 1948 1124 1982
rect 1124 1948 1142 1982
rect 1188 1948 1192 1982
rect 1192 1948 1222 1982
rect -2 1880 32 1910
rect -2 1876 32 1880
rect 1260 1876 1294 1909
rect 1260 1875 1294 1876
rect -2 1812 32 1836
rect -2 1802 32 1812
rect 238 1838 253 1872
rect 253 1838 272 1872
rect 317 1838 321 1872
rect 321 1838 351 1872
rect 397 1838 423 1872
rect 423 1838 431 1872
rect 477 1838 491 1872
rect 491 1838 511 1872
rect 557 1838 559 1872
rect 559 1838 591 1872
rect 667 1838 701 1872
rect 739 1838 769 1872
rect 769 1838 773 1872
rect -2 1744 32 1762
rect -2 1728 32 1744
rect 1260 1808 1294 1836
rect 1260 1802 1294 1808
rect 1260 1740 1294 1763
rect 1260 1729 1294 1740
rect -2 1676 32 1688
rect -2 1654 32 1676
rect -2 1608 32 1614
rect -2 1580 32 1608
rect -2 1506 32 1540
rect -2 1438 32 1466
rect -2 1432 32 1438
rect -2 1370 32 1392
rect -2 1358 32 1370
rect -2 1302 32 1318
rect -2 1284 32 1302
rect -2 1234 32 1244
rect -2 1210 32 1234
rect 158 1682 192 1716
rect 158 1601 192 1635
rect 158 1520 192 1554
rect 158 1439 192 1473
rect 158 1358 192 1392
rect 158 1278 192 1312
rect 158 1198 192 1232
rect 334 1682 368 1716
rect 334 1601 368 1635
rect 334 1520 368 1554
rect 334 1439 368 1473
rect 334 1358 368 1392
rect 334 1278 368 1312
rect 334 1198 368 1232
rect 444 1682 478 1716
rect 444 1601 478 1635
rect 444 1520 478 1554
rect 444 1439 478 1473
rect 444 1358 478 1392
rect 444 1278 478 1312
rect 444 1198 478 1232
rect 620 1682 654 1716
rect 620 1601 654 1635
rect 620 1520 654 1554
rect 620 1439 654 1473
rect 620 1358 654 1392
rect 620 1278 654 1312
rect 620 1198 654 1232
rect 796 1682 830 1716
rect 796 1601 830 1635
rect 796 1520 830 1554
rect 796 1439 830 1473
rect 796 1358 830 1392
rect 796 1278 830 1312
rect 796 1198 830 1232
rect 1260 1672 1294 1690
rect 1260 1656 1294 1672
rect 1260 1604 1294 1617
rect 1260 1583 1294 1604
rect 1260 1536 1294 1544
rect 1260 1510 1294 1536
rect 1260 1468 1294 1471
rect 1260 1437 1294 1468
rect 1260 1366 1294 1398
rect 1260 1364 1294 1366
rect 1260 1298 1294 1324
rect 1260 1290 1294 1298
rect -2 1166 32 1170
rect -2 1136 32 1166
rect -2 1064 32 1096
rect -2 1062 32 1064
rect 1260 1230 1294 1250
rect 1260 1216 1294 1230
rect 1260 1162 1294 1176
rect 1260 1142 1294 1162
rect -2 996 32 1023
rect -2 989 32 996
rect 158 1048 192 1082
rect 158 976 192 1010
rect 630 1048 664 1082
rect -2 928 32 950
rect -2 916 32 928
rect 394 968 428 1002
rect 630 976 664 1010
rect 1102 1048 1136 1082
rect 394 896 428 930
rect 866 968 900 1002
rect 1102 976 1136 1010
rect 1260 1094 1294 1102
rect 1260 1068 1294 1094
rect 1260 1026 1294 1028
rect 1260 994 1294 1026
rect 866 896 900 930
rect 1260 924 1294 954
rect 1260 920 1294 924
rect -2 860 32 877
rect -2 843 32 860
rect 1260 856 1294 880
rect 1260 846 1294 856
rect -2 792 32 804
rect -2 770 32 792
rect 276 802 287 836
rect 287 802 310 836
rect 355 802 389 836
rect 434 802 457 836
rect 457 802 468 836
rect 513 802 525 836
rect 525 802 547 836
rect 592 802 593 836
rect 593 802 626 836
rect 671 802 696 836
rect 696 802 705 836
rect 751 802 765 836
rect 765 802 785 836
rect 831 802 834 836
rect 834 802 865 836
rect 911 802 937 836
rect 937 802 945 836
rect 991 802 1006 836
rect 1006 802 1025 836
rect -2 724 32 731
rect -2 697 32 724
rect 1260 788 1294 806
rect 1260 772 1294 788
rect -2 656 32 658
rect -2 624 32 656
rect 394 718 428 752
rect -2 554 32 585
rect -2 551 32 554
rect 158 638 192 672
rect 394 646 428 680
rect 866 718 900 752
rect 158 566 192 600
rect 630 638 664 672
rect 866 646 900 680
rect 1260 720 1294 732
rect 1260 698 1294 720
rect 630 566 664 600
rect 1102 638 1136 672
rect 1102 566 1136 600
rect -2 486 32 512
rect -2 478 32 486
rect -2 418 32 439
rect -2 405 32 418
rect 252 408 253 442
rect 253 408 286 442
rect 328 408 362 442
rect 404 408 438 442
rect 582 408 597 442
rect 597 408 616 442
rect 658 408 671 442
rect 671 408 692 442
rect 734 408 745 442
rect 745 408 768 442
rect -2 350 32 366
rect -2 332 32 350
rect -2 282 32 293
rect -2 259 32 282
rect 244 321 278 355
rect -2 214 32 220
rect -2 186 32 214
rect 158 228 192 262
rect 244 249 278 283
rect 416 321 450 355
rect 158 156 192 190
rect 330 228 364 262
rect 416 249 450 283
rect 588 321 622 355
rect 330 156 364 190
rect 502 228 536 262
rect 588 249 622 283
rect 760 321 794 355
rect 502 156 536 190
rect 674 228 708 262
rect 760 249 794 283
rect 1260 346 1294 351
rect 1260 317 1294 346
rect 674 156 708 190
rect 846 228 880 262
rect 846 156 880 190
rect 1260 244 1294 249
rect 1260 215 1294 244
rect -2 113 32 147
rect 1260 142 1294 146
rect 1260 112 1294 142
rect 70 40 100 74
rect 100 40 104 74
rect 145 40 168 74
rect 168 40 179 74
rect 220 40 236 74
rect 236 40 254 74
rect 295 40 304 74
rect 304 40 329 74
rect 370 40 372 74
rect 372 40 404 74
rect 445 40 474 74
rect 474 40 479 74
rect 520 40 542 74
rect 542 40 554 74
rect 594 40 610 74
rect 610 40 628 74
rect 668 40 678 74
rect 678 40 702 74
rect 742 40 746 74
rect 746 40 776 74
rect 816 40 848 74
rect 848 40 850 74
rect 890 40 916 74
rect 916 40 924 74
rect 964 40 984 74
rect 984 40 998 74
rect 1038 40 1052 74
rect 1052 40 1072 74
rect 1112 40 1120 74
rect 1120 40 1146 74
rect 1186 40 1188 74
rect 1188 40 1220 74
<< metal1 >>
rect 91 4262 594 4268
rect 91 4228 104 4262
rect 138 4228 178 4262
rect 212 4228 252 4262
rect 286 4228 326 4262
rect 360 4228 400 4262
rect 434 4228 474 4262
rect 508 4228 548 4262
rect 582 4228 594 4262
rect 91 4222 594 4228
rect 91 4122 151 4222
tri 151 4188 185 4222 nw
rect 91 4088 111 4122
rect 145 4088 151 4122
rect 91 4050 151 4088
rect 91 4016 111 4050
rect 145 4016 151 4050
rect 91 4004 151 4016
rect 261 4122 313 4134
rect 261 4088 267 4122
rect 301 4088 313 4122
rect 261 4050 313 4088
rect 261 4016 267 4050
rect 301 4016 313 4050
rect 101 3957 233 3963
rect 101 3923 115 3957
rect 149 3923 187 3957
rect 221 3923 233 3957
rect 101 3917 233 3923
rect 101 3695 153 3917
tri 153 3883 187 3917 nw
rect 261 3868 313 4016
tri 227 3792 261 3826 se
rect 261 3804 313 3816
rect 181 3786 261 3792
rect 181 3752 193 3786
rect 227 3752 261 3786
rect 181 3746 313 3752
rect 101 3631 153 3643
rect 101 3573 153 3579
rect 261 3672 307 3684
rect 261 3638 267 3672
rect 301 3638 307 3672
rect 261 3600 307 3638
rect 261 3566 267 3600
rect 301 3566 307 3600
tri 227 3369 261 3403 se
rect 261 3369 307 3566
tri 307 3369 341 3403 sw
rect 121 3169 687 3369
rect 116 2938 267 2990
rect 319 2938 360 2990
rect 412 2938 1037 2990
rect 101 2858 107 2910
rect 159 2858 171 2910
rect 223 2858 1037 2910
rect 116 2824 1037 2830
rect 116 2772 824 2824
rect 876 2772 1037 2824
rect 116 2756 1037 2772
rect 116 2704 824 2756
rect 876 2704 1037 2756
rect 116 2688 1037 2704
rect 116 2636 824 2688
rect 876 2636 1037 2688
rect 116 2630 1037 2636
rect 116 2538 674 2590
rect 726 2538 738 2590
rect 790 2538 1037 2590
rect 116 2458 211 2510
rect 263 2458 275 2510
rect 327 2458 1037 2510
rect -8 1982 1300 1988
rect -8 1948 70 1982
rect 104 1948 142 1982
rect 176 1948 215 1982
rect 249 1948 288 1982
rect 322 1948 361 1982
rect 395 1948 471 1982
rect 505 1948 550 1982
rect 584 1948 629 1982
rect 663 1948 708 1982
rect 742 1948 788 1982
rect 822 1948 868 1982
rect 902 1948 948 1982
rect 982 1948 1028 1982
rect 1062 1948 1108 1982
rect 1142 1948 1188 1982
rect 1222 1948 1300 1982
rect -8 1942 1300 1948
rect -8 1910 39 1942
rect -8 1876 -2 1910
rect 32 1909 39 1910
tri 39 1909 72 1942 nw
tri 1220 1909 1253 1942 ne
rect 1253 1909 1300 1942
rect 32 1876 38 1909
tri 38 1908 39 1909 nw
tri 1253 1908 1254 1909 ne
rect -8 1836 38 1876
rect -8 1802 -2 1836
rect 32 1802 38 1836
rect 205 1829 211 1881
rect 263 1872 275 1881
rect 327 1872 603 1881
rect 272 1838 275 1872
rect 351 1838 397 1872
rect 431 1838 477 1872
rect 511 1838 557 1872
rect 591 1838 603 1872
rect 263 1829 275 1838
rect 327 1829 603 1838
rect 655 1829 663 1881
rect 715 1829 727 1881
rect 779 1829 785 1881
rect 1254 1875 1260 1909
rect 1294 1875 1300 1909
rect 1254 1836 1300 1875
rect -8 1762 38 1802
rect -8 1728 -2 1762
rect 32 1728 38 1762
rect 1254 1802 1260 1836
rect 1294 1802 1300 1836
rect 1254 1763 1300 1802
rect 1254 1729 1260 1763
rect 1294 1729 1300 1763
rect -8 1688 38 1728
rect -8 1654 -2 1688
rect 32 1654 38 1688
rect -8 1614 38 1654
rect -8 1580 -2 1614
rect 32 1580 38 1614
rect -8 1540 38 1580
rect -8 1506 -2 1540
rect 32 1506 38 1540
rect -8 1466 38 1506
rect -8 1432 -2 1466
rect 32 1432 38 1466
rect -8 1392 38 1432
rect -8 1358 -2 1392
rect 32 1358 38 1392
rect -8 1318 38 1358
rect -8 1284 -2 1318
rect 32 1284 38 1318
rect -8 1244 38 1284
rect -8 1210 -2 1244
rect 32 1210 38 1244
rect -8 1170 38 1210
rect 149 1716 201 1728
rect 149 1682 158 1716
rect 192 1682 201 1716
rect 149 1635 201 1682
rect 149 1601 158 1635
rect 192 1601 201 1635
rect 149 1554 201 1601
rect 149 1520 158 1554
rect 192 1520 201 1554
rect 149 1473 201 1520
rect 149 1439 158 1473
rect 192 1439 201 1473
rect 149 1392 201 1439
rect 149 1358 158 1392
rect 192 1358 201 1392
rect 149 1312 201 1358
rect 149 1308 158 1312
rect 192 1308 201 1312
rect 149 1244 201 1256
rect 149 1186 201 1192
rect 321 1716 374 1728
rect 321 1682 334 1716
rect 368 1682 374 1716
rect 321 1635 374 1682
rect 321 1601 334 1635
rect 368 1601 374 1635
rect 321 1557 374 1601
rect 373 1505 374 1557
rect 321 1493 374 1505
rect 373 1441 374 1493
rect 321 1439 334 1441
rect 368 1439 374 1441
rect 321 1392 374 1439
rect 321 1358 334 1392
rect 368 1358 374 1392
rect 321 1312 374 1358
rect 321 1278 334 1312
rect 368 1278 374 1312
rect 321 1232 374 1278
rect 321 1198 334 1232
rect 368 1198 374 1232
rect 321 1186 374 1198
rect 435 1716 487 1728
rect 435 1682 444 1716
rect 478 1682 487 1716
rect 435 1635 487 1682
rect 435 1601 444 1635
rect 478 1601 487 1635
rect 435 1554 487 1601
rect 435 1520 444 1554
rect 478 1520 487 1554
rect 435 1473 487 1520
rect 435 1439 444 1473
rect 478 1439 487 1473
rect 435 1392 487 1439
rect 435 1358 444 1392
rect 478 1358 487 1392
rect 435 1312 487 1358
rect 435 1308 444 1312
rect 478 1308 487 1312
rect 435 1244 487 1256
rect 435 1186 487 1192
rect 611 1716 663 1728
rect 611 1682 620 1716
rect 654 1682 663 1716
rect 611 1635 663 1682
rect 611 1601 620 1635
rect 654 1601 663 1635
rect 611 1600 663 1601
rect 611 1536 620 1548
rect 654 1536 663 1548
rect 611 1473 663 1484
rect 611 1439 620 1473
rect 654 1439 663 1473
rect 611 1392 663 1439
rect 611 1358 620 1392
rect 654 1358 663 1392
rect 611 1312 663 1358
rect 611 1278 620 1312
rect 654 1278 663 1312
rect 611 1232 663 1278
rect 611 1198 620 1232
rect 654 1198 663 1232
rect 611 1186 663 1198
rect 790 1716 836 1728
rect 790 1682 796 1716
rect 830 1682 836 1716
rect 790 1635 836 1682
rect 790 1601 796 1635
rect 830 1601 836 1635
rect 790 1554 836 1601
rect 790 1520 796 1554
rect 830 1520 836 1554
rect 790 1473 836 1520
rect 790 1439 796 1473
rect 830 1439 836 1473
rect 1254 1690 1300 1729
rect 1254 1656 1260 1690
rect 1294 1656 1300 1690
rect 1254 1617 1300 1656
rect 1254 1583 1260 1617
rect 1294 1583 1300 1617
rect 1254 1544 1300 1583
rect 1254 1510 1260 1544
rect 1294 1510 1300 1544
rect 1254 1471 1300 1510
rect 790 1437 836 1439
tri 836 1437 866 1467 sw
tri 1224 1437 1254 1467 se
rect 1254 1437 1260 1471
rect 1294 1437 1300 1471
rect 790 1433 866 1437
tri 866 1433 870 1437 sw
tri 1220 1433 1224 1437 se
rect 1224 1433 1300 1437
rect 790 1398 1300 1433
rect 790 1392 1260 1398
rect 790 1358 796 1392
rect 830 1364 1260 1392
rect 1294 1364 1300 1398
rect 830 1358 1300 1364
rect 790 1324 1300 1358
rect 790 1312 1260 1324
rect 790 1278 796 1312
rect 830 1290 1260 1312
rect 1294 1290 1300 1324
rect 830 1278 1300 1290
rect 790 1250 1300 1278
rect 790 1232 1260 1250
rect 790 1198 796 1232
rect 830 1216 1260 1232
rect 1294 1216 1300 1250
rect 830 1198 1300 1216
rect 790 1186 1300 1198
tri 1220 1176 1230 1186 ne
rect 1230 1176 1300 1186
rect -8 1136 -2 1170
rect 32 1136 38 1170
tri 1230 1152 1254 1176 ne
rect -8 1096 38 1136
rect -8 1062 -2 1096
rect 32 1062 38 1096
rect 1254 1142 1260 1176
rect 1294 1142 1300 1176
rect 1254 1102 1300 1142
rect -8 1023 38 1062
rect -8 989 -2 1023
rect 32 989 38 1023
rect -8 950 38 989
rect 152 1082 441 1094
rect 152 1048 158 1082
rect 192 1048 441 1082
rect 152 1042 441 1048
rect 493 1042 505 1094
rect 557 1082 1142 1094
rect 557 1048 630 1082
rect 664 1048 1102 1082
rect 1136 1048 1142 1082
rect 557 1042 1142 1048
rect 152 1028 218 1042
tri 218 1028 232 1042 nw
tri 590 1028 604 1042 ne
rect 604 1028 690 1042
tri 690 1028 704 1042 nw
tri 1062 1028 1076 1042 ne
rect 1076 1028 1142 1042
rect 152 1010 200 1028
tri 200 1010 218 1028 nw
tri 604 1014 618 1028 ne
rect 618 1014 672 1028
rect 152 976 158 1010
rect 192 976 198 1010
tri 198 1008 200 1010 nw
rect 152 964 198 976
rect 388 1002 434 1014
tri 618 1010 622 1014 ne
rect 622 1010 672 1014
tri 672 1010 690 1028 nw
tri 1076 1014 1090 1028 ne
rect 1090 1014 1142 1028
tri 622 1008 624 1010 ne
rect 388 968 394 1002
rect 428 968 434 1002
rect 624 976 630 1010
rect 664 976 670 1010
tri 670 1008 672 1010 nw
tri 434 968 436 970 sw
rect -8 916 -2 950
rect 32 916 38 950
rect -8 877 38 916
rect 388 954 436 968
tri 436 954 450 968 sw
rect 624 964 670 976
rect 860 1002 906 1014
tri 1090 1010 1094 1014 ne
rect 1094 1010 1142 1014
tri 1094 1008 1096 1010 ne
tri 858 968 860 970 se
rect 860 968 866 1002
rect 900 968 906 1002
tri 854 964 858 968 se
rect 858 964 906 968
rect 1096 976 1102 1010
rect 1136 976 1142 1010
rect 1096 964 1142 976
rect 1254 1068 1260 1102
rect 1294 1068 1300 1102
rect 1254 1028 1300 1068
rect 1254 994 1260 1028
rect 1294 994 1300 1028
tri 844 954 854 964 se
rect 854 954 906 964
rect 388 936 450 954
tri 450 936 468 954 sw
tri 826 936 844 954 se
rect 844 936 906 954
rect 388 930 512 936
rect 388 896 394 930
rect 428 896 512 930
rect 388 884 512 896
rect 564 884 576 936
rect 628 930 906 936
rect 628 896 866 930
rect 900 896 906 930
rect 628 884 906 896
rect 1254 954 1300 994
rect 1254 920 1260 954
rect 1294 920 1300 954
rect -8 843 -2 877
rect 32 843 38 877
rect 1254 880 1300 920
rect -8 804 38 843
rect -8 770 -2 804
rect 32 770 38 804
rect 264 836 672 847
rect 264 802 276 836
rect 310 802 355 836
rect 389 802 434 836
rect 468 802 513 836
rect 547 802 592 836
rect 626 802 671 836
rect 264 795 672 802
rect 724 795 736 847
rect 788 836 1037 847
rect 788 802 831 836
rect 865 802 911 836
rect 945 802 991 836
rect 1025 802 1037 836
rect 788 795 1037 802
rect 1254 846 1260 880
rect 1294 846 1300 880
rect 1254 806 1300 846
rect -8 731 38 770
rect 1254 772 1260 806
rect 1294 772 1300 806
rect -8 697 -2 731
rect 32 697 38 731
rect 314 712 320 764
rect 372 712 384 764
rect 436 752 906 764
rect 436 718 866 752
rect 900 718 906 752
rect 436 712 906 718
tri 354 698 368 712 ne
rect 368 698 454 712
tri 454 698 468 712 nw
tri 826 698 840 712 ne
rect 840 698 906 712
rect -8 658 38 697
tri 368 684 382 698 ne
rect 382 684 436 698
rect -8 624 -2 658
rect 32 624 38 658
rect -8 585 38 624
rect -8 551 -2 585
rect 32 551 38 585
rect 152 672 198 684
tri 382 680 386 684 ne
rect 386 680 436 684
tri 436 680 454 698 nw
tri 840 684 854 698 ne
rect 854 684 906 698
rect 1254 732 1300 772
rect 1254 698 1260 732
rect 1294 698 1300 732
tri 386 678 388 680 ne
rect 152 638 158 672
rect 192 638 198 672
rect 388 646 394 680
rect 428 646 434 680
tri 434 678 436 680 nw
tri 198 638 200 640 sw
rect 152 606 200 638
tri 200 606 232 638 sw
rect 388 634 434 646
rect 624 672 670 684
tri 854 680 858 684 ne
rect 858 680 906 684
tri 858 678 860 680 ne
tri 622 638 624 640 se
rect 624 638 630 672
rect 664 638 670 672
rect 860 646 866 680
rect 900 646 906 680
tri 670 638 672 640 sw
tri 618 634 622 638 se
rect 622 634 672 638
tri 590 606 618 634 se
rect 618 606 672 634
tri 672 606 704 638 sw
rect 860 634 906 646
rect 1096 672 1142 684
tri 1094 638 1096 640 se
rect 1096 638 1102 672
rect 1136 638 1142 672
rect 1254 660 1300 698
tri 1090 634 1094 638 se
rect 1094 634 1142 638
tri 1062 606 1090 634 se
rect 1090 606 1142 634
rect 152 554 158 606
rect 210 554 222 606
rect 274 600 1142 606
rect 274 566 630 600
rect 664 566 1102 600
rect 1136 566 1142 600
rect 274 554 1142 566
rect -8 512 38 551
rect -8 478 -2 512
rect 32 478 38 512
rect -8 439 38 478
tri 462 458 520 516 se
rect 520 484 906 516
tri 520 458 546 484 nw
tri 452 448 462 458 se
rect 462 448 504 458
rect -8 405 -2 439
rect 32 405 38 439
rect -8 366 38 405
rect 240 442 504 448
tri 504 442 520 458 nw
rect 570 442 780 448
rect 240 408 252 442
rect 286 408 328 442
rect 362 408 404 442
rect 438 408 470 442
tri 470 408 504 442 nw
rect 570 408 582 442
rect 616 408 658 442
rect 692 408 734 442
rect 768 408 780 442
rect 240 402 464 408
tri 464 402 470 408 nw
rect 570 402 780 408
rect -8 332 -2 366
rect 32 332 38 366
rect -8 293 38 332
rect -8 259 -2 293
rect 32 259 38 293
rect 238 315 244 367
rect 296 315 308 367
rect 360 355 456 367
rect 360 321 416 355
rect 450 321 456 355
rect 360 315 456 321
rect 238 283 286 315
tri 286 283 318 315 nw
tri 376 283 408 315 ne
rect 408 283 456 315
rect -8 228 38 259
rect 152 262 198 274
tri 38 228 46 236 sw
tri 144 228 152 236 se
rect 152 228 158 262
rect 192 228 198 262
rect 238 249 244 283
rect 278 249 284 283
tri 284 281 286 283 nw
tri 408 281 410 283 ne
rect 238 237 284 249
rect 324 262 370 274
tri 198 228 206 236 sw
tri 316 228 324 236 se
rect 324 228 330 262
rect 364 228 370 262
rect 410 249 416 283
rect 450 249 456 283
rect 582 315 588 367
rect 640 315 652 367
rect 704 355 800 367
rect 704 321 760 355
rect 794 321 800 355
rect 704 315 800 321
rect 582 283 630 315
tri 630 283 662 315 nw
tri 720 283 752 315 ne
rect 752 283 800 315
rect 410 237 456 249
rect 496 262 542 274
tri 370 228 378 236 sw
tri 488 228 496 236 se
rect 496 228 502 262
rect 536 228 542 262
rect 582 249 588 283
rect 622 249 628 283
tri 628 281 630 283 nw
tri 752 281 754 283 ne
rect 582 237 628 249
rect 668 262 714 274
tri 542 228 550 236 sw
tri 660 228 668 236 se
rect 668 228 674 262
rect 708 228 714 262
rect 754 249 760 283
rect 794 249 800 283
rect 1254 351 1300 389
rect 1254 317 1260 351
rect 1294 317 1300 351
rect 754 237 800 249
rect 840 262 886 274
tri 714 228 722 236 sw
tri 832 228 840 236 se
rect 840 228 846 262
rect 880 228 886 262
rect 1254 249 1300 317
rect -8 220 46 228
rect -8 186 -2 220
rect 32 215 46 220
tri 46 215 59 228 sw
tri 131 215 144 228 se
rect 144 215 206 228
tri 206 215 219 228 sw
tri 303 215 316 228 se
rect 316 215 378 228
tri 378 215 391 228 sw
tri 475 215 488 228 se
rect 488 215 550 228
tri 550 215 563 228 sw
tri 647 215 660 228 se
rect 660 215 722 228
tri 722 215 735 228 sw
tri 819 215 832 228 se
rect 832 215 886 228
tri 886 215 907 236 sw
tri 1233 215 1254 236 se
rect 1254 215 1260 249
rect 1294 215 1300 249
rect 32 202 59 215
tri 59 202 72 215 sw
tri 118 202 131 215 se
rect 131 202 219 215
tri 219 202 232 215 sw
tri 290 202 303 215 se
rect 303 202 391 215
tri 391 202 404 215 sw
tri 462 202 475 215 se
rect 475 202 563 215
tri 563 202 576 215 sw
tri 634 202 647 215 se
rect 647 202 735 215
tri 735 202 748 215 sw
tri 806 202 819 215 se
rect 819 202 907 215
tri 907 202 920 215 sw
tri 1220 202 1233 215 se
rect 1233 202 1300 215
rect 32 190 1300 202
rect 32 186 158 190
rect -8 156 158 186
rect 192 156 330 190
rect 364 156 502 190
rect 536 156 674 190
rect 708 156 846 190
rect 880 156 1300 190
rect -8 147 1300 156
rect -8 113 -2 147
rect 32 146 1300 147
rect 32 113 1260 146
rect -8 112 1260 113
rect 1294 112 1300 146
rect -8 74 1300 112
rect -8 40 70 74
rect 104 40 145 74
rect 179 40 220 74
rect 254 40 295 74
rect 329 40 370 74
rect 404 40 445 74
rect 479 40 520 74
rect 554 40 594 74
rect 628 40 668 74
rect 702 40 742 74
rect 776 40 816 74
rect 850 40 890 74
rect 924 40 964 74
rect 998 40 1038 74
rect 1072 40 1112 74
rect 1146 40 1186 74
rect 1220 40 1300 74
rect -8 34 1300 40
<< via1 >>
rect 261 3816 313 3868
rect 261 3786 313 3804
rect 261 3752 265 3786
rect 265 3752 299 3786
rect 299 3752 313 3786
rect 101 3692 153 3695
rect 101 3658 111 3692
rect 111 3658 145 3692
rect 145 3658 153 3692
rect 101 3643 153 3658
rect 101 3620 153 3631
rect 101 3586 111 3620
rect 111 3586 145 3620
rect 145 3586 153 3620
rect 101 3579 153 3586
rect 267 2938 319 2990
rect 360 2938 412 2990
rect 107 2858 159 2910
rect 171 2858 223 2910
rect 824 2772 876 2824
rect 824 2704 876 2756
rect 824 2636 876 2688
rect 674 2538 726 2590
rect 738 2538 790 2590
rect 211 2458 263 2510
rect 275 2458 327 2510
rect 211 1872 263 1881
rect 275 1872 327 1881
rect 211 1838 238 1872
rect 238 1838 263 1872
rect 275 1838 317 1872
rect 317 1838 327 1872
rect 211 1829 263 1838
rect 275 1829 327 1838
rect 663 1872 715 1881
rect 663 1838 667 1872
rect 667 1838 701 1872
rect 701 1838 715 1872
rect 663 1829 715 1838
rect 727 1872 779 1881
rect 727 1838 739 1872
rect 739 1838 773 1872
rect 773 1838 779 1872
rect 727 1829 779 1838
rect 149 1278 158 1308
rect 158 1278 192 1308
rect 192 1278 201 1308
rect 149 1256 201 1278
rect 149 1232 201 1244
rect 149 1198 158 1232
rect 158 1198 192 1232
rect 192 1198 201 1232
rect 149 1192 201 1198
rect 321 1554 373 1557
rect 321 1520 334 1554
rect 334 1520 368 1554
rect 368 1520 373 1554
rect 321 1505 373 1520
rect 321 1473 373 1493
rect 321 1441 334 1473
rect 334 1441 368 1473
rect 368 1441 373 1473
rect 435 1278 444 1308
rect 444 1278 478 1308
rect 478 1278 487 1308
rect 435 1256 487 1278
rect 435 1232 487 1244
rect 435 1198 444 1232
rect 444 1198 478 1232
rect 478 1198 487 1232
rect 435 1192 487 1198
rect 611 1554 663 1600
rect 611 1548 620 1554
rect 620 1548 654 1554
rect 654 1548 663 1554
rect 611 1520 620 1536
rect 620 1520 654 1536
rect 654 1520 663 1536
rect 611 1484 663 1520
rect 441 1042 493 1094
rect 505 1042 557 1094
rect 512 884 564 936
rect 576 884 628 936
rect 672 836 724 847
rect 672 802 705 836
rect 705 802 724 836
rect 672 795 724 802
rect 736 836 788 847
rect 736 802 751 836
rect 751 802 785 836
rect 785 802 788 836
rect 736 795 788 802
rect 320 712 372 764
rect 384 752 436 764
rect 384 718 394 752
rect 394 718 428 752
rect 428 718 436 752
rect 384 712 436 718
rect 158 600 210 606
rect 158 566 192 600
rect 192 566 210 600
rect 158 554 210 566
rect 222 554 274 606
rect 244 355 296 367
rect 244 321 278 355
rect 278 321 296 355
rect 244 315 296 321
rect 308 315 360 367
rect 588 355 640 367
rect 588 321 622 355
rect 622 321 640 355
rect 588 315 640 321
rect 652 315 704 367
<< metal2 >>
rect 261 3868 313 3874
rect 261 3804 313 3816
rect 101 3695 153 3701
rect 101 3631 153 3643
rect 101 2938 153 3579
rect 261 2990 313 3752
tri 313 2990 347 3024 sw
tri 153 2938 159 2944 sw
rect 261 2938 267 2990
rect 319 2938 360 2990
rect 412 2938 418 2990
rect 101 2910 159 2938
tri 159 2910 187 2938 sw
tri 332 2910 360 2938 ne
rect 360 2910 418 2938
rect 101 2858 107 2910
rect 159 2858 171 2910
rect 223 2858 229 2910
tri 360 2904 366 2910 ne
rect 101 1769 153 2858
tri 153 2824 187 2858 nw
rect 205 2458 211 2510
rect 263 2458 275 2510
rect 327 2458 333 2510
rect 205 1881 257 2458
tri 257 2424 291 2458 nw
rect 366 1929 418 2910
rect 824 2824 876 2830
rect 824 2756 876 2772
rect 824 2688 876 2704
rect 668 2538 674 2590
rect 726 2538 738 2590
rect 790 2538 796 2590
tri 418 1929 420 1931 sw
tri 257 1881 291 1915 sw
rect 366 1902 420 1929
tri 366 1881 387 1902 ne
rect 387 1881 420 1902
tri 420 1881 468 1929 sw
tri 657 1881 668 1892 se
rect 668 1881 720 2538
tri 720 2504 754 2538 nw
tri 720 1881 754 1915 sw
rect 205 1829 211 1881
rect 263 1829 275 1881
rect 327 1829 333 1881
tri 387 1848 420 1881 ne
rect 420 1848 468 1881
tri 468 1848 501 1881 sw
tri 420 1829 439 1848 ne
rect 439 1829 501 1848
tri 501 1829 520 1848 sw
rect 657 1829 663 1881
rect 715 1829 727 1881
rect 779 1829 785 1881
tri 439 1791 477 1829 ne
rect 477 1791 520 1829
tri 101 1717 153 1769 ne
tri 153 1719 225 1791 sw
tri 477 1767 501 1791 ne
rect 501 1767 520 1791
tri 520 1767 582 1829 sw
tri 794 1773 824 1803 se
rect 824 1781 876 2636
rect 824 1773 868 1781
tri 868 1773 876 1781 nw
tri 788 1767 794 1773 se
tri 501 1719 549 1767 ne
rect 549 1719 582 1767
rect 153 1717 225 1719
tri 153 1645 225 1717 ne
tri 225 1645 299 1719 sw
tri 549 1686 582 1719 ne
tri 582 1686 663 1767 sw
tri 582 1657 611 1686 ne
tri 225 1600 270 1645 ne
rect 270 1600 299 1645
tri 299 1600 344 1645 sw
rect 611 1600 663 1686
tri 270 1571 299 1600 ne
rect 299 1571 344 1600
tri 344 1571 373 1600 sw
tri 299 1557 313 1571 ne
rect 313 1557 373 1571
tri 313 1549 321 1557 ne
rect 321 1493 373 1505
rect 611 1536 663 1548
rect 611 1478 663 1484
tri 742 1721 788 1767 se
rect 788 1721 794 1767
rect 321 1435 373 1441
rect 149 1308 201 1314
rect 149 1244 201 1256
rect 149 606 201 1192
rect 435 1308 487 1314
rect 435 1244 487 1256
rect 435 1094 487 1192
tri 487 1094 521 1128 sw
rect 435 1042 441 1094
rect 493 1042 505 1094
rect 557 1042 563 1094
rect 506 884 512 936
rect 564 884 576 936
rect 628 884 634 936
tri 548 850 582 884 ne
rect 314 712 320 764
rect 372 712 384 764
rect 436 712 442 764
tri 201 606 235 640 sw
rect 149 554 158 606
rect 210 554 222 606
rect 274 554 280 606
tri 287 367 314 394 se
rect 314 367 366 712
tri 366 678 400 712 nw
rect 238 315 244 367
rect 296 315 308 367
rect 360 315 366 367
rect 582 367 634 884
tri 708 847 742 881 se
rect 742 847 794 1721
tri 794 1699 868 1773 nw
rect 666 795 672 847
rect 724 795 736 847
rect 788 795 794 847
tri 634 367 661 394 sw
rect 582 315 588 367
rect 640 315 652 367
rect 704 315 710 367
use nfet_CDNS_5595914180818  nfet_CDNS_5595914180818_0
timestamp 1704896540
transform 1 0 665 0 1 1190
box -79 -32 199 632
use nfet_CDNS_5595914180818  nfet_CDNS_5595914180818_1
timestamp 1704896540
transform 1 0 489 0 1 1190
box -79 -32 199 632
use nfet_CDNS_5595914180818  nfet_CDNS_5595914180818_2
timestamp 1704896540
transform 1 0 203 0 1 1190
box -79 -32 199 632
use nfet_CDNS_5595914180820  nfet_CDNS_5595914180820_0
timestamp 1704896540
transform -1 0 1091 0 1 884
box -79 -32 967 232
use nfet_CDNS_5595914180820  nfet_CDNS_5595914180820_1
timestamp 1704896540
transform -1 0 1091 0 1 554
box -79 -32 967 232
use nfet_CDNS_5595914180821  nfet_CDNS_5595914180821_0
timestamp 1704896540
transform -1 0 491 0 1 160
box -79 -32 367 232
use nfet_CDNS_5595914180821  nfet_CDNS_5595914180821_1
timestamp 1704896540
transform -1 0 835 0 1 160
box -79 -32 367 232
use pfet_CDNS_5595914180822  pfet_CDNS_5595914180822_0
timestamp 1704896540
transform 1 0 156 0 1 4004
box -119 -66 219 216
use pfet_CDNS_5595914180822  pfet_CDNS_5595914180822_1
timestamp 1704896540
transform 1 0 156 0 1 3554
box -119 -66 219 216
<< labels >>
flabel metal1 s 146 2644 301 2738 3 FreeSans 200 0 0 0 vpwr_lv
port 2 nsew
flabel metal1 s 135 4234 228 4259 3 FreeSans 200 0 0 0 vpwr_hv
port 3 nsew
flabel metal1 s 144 2870 225 2900 3 FreeSans 200 0 0 0 fbk_n
port 4 nsew
flabel metal1 s 144 2947 244 2980 3 FreeSans 200 0 0 0 fbk
port 5 nsew
flabel metal1 s 146 2547 237 2581 3 FreeSans 200 0 0 0 reset
port 6 nsew
flabel metal1 s 143 2464 207 2501 3 FreeSans 200 0 0 0 hold
port 7 nsew
flabel metal1 s 637 412 732 437 3 FreeSans 200 0 0 0 switch_lv_n
port 8 nsew
flabel metal1 s 278 413 393 440 3 FreeSans 200 0 0 0 switch_lv
port 9 nsew
flabel metal1 s 133 67 301 127 3 FreeSans 200 0 0 0 vgnd
port 1 nsew
<< properties >>
string GDS_END 694224
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 653874
<< end >>
