magic
tech sky130A
timestamp 1704896540
<< metal1 >>
rect 0 0 3 122
rect 189 0 192 122
<< via1 >>
rect 3 0 189 122
<< metal2 >>
rect 0 0 3 122
rect 189 0 192 122
<< properties >>
string GDS_END 88155338
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 88153670
<< end >>
