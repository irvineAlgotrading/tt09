magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect 675 6574 2933 7988
rect 675 6464 2563 6574
rect 725 5278 1465 6064
rect 635 2182 1229 4878
rect 665 122 1189 1782
<< pwell >>
rect 467 7143 553 8102
rect 27 6816 545 6902
rect -433 4602 -288 4771
rect 27 4602 113 6816
rect -433 4516 113 4602
rect -433 4314 72 4516
rect -433 3521 -288 4314
rect -419 3507 -288 3521
rect -406 725 -288 3507
rect 459 2288 545 6816
rect 2993 7882 3917 7968
rect 2993 6680 3079 7882
rect 3831 6680 3917 7882
rect 2993 6594 3917 6680
rect 135 1744 545 2288
rect -400 348 -288 725
rect -400 198 72 348
rect 459 198 545 1744
rect -400 112 545 198
<< pdiff >>
rect 925 5928 1051 5940
rect 925 5894 1005 5928
rect 1039 5894 1051 5928
rect 925 5886 1051 5894
rect 1129 5928 1255 5940
rect 1129 5894 1209 5928
rect 1243 5894 1255 5928
rect 1129 5886 1255 5894
rect 925 5448 1051 5456
rect 925 5414 1005 5448
rect 1039 5414 1051 5448
rect 925 5402 1051 5414
rect 1129 5448 1255 5456
rect 1129 5414 1209 5448
rect 1243 5414 1255 5448
rect 1129 5402 1255 5414
<< mvndiff >>
rect -240 4450 -156 4458
rect -240 4416 -228 4450
rect -194 4416 -156 4450
rect -240 4382 -156 4416
rect -38 4450 46 4458
rect -38 4416 0 4450
rect 34 4416 46 4450
rect -38 4382 46 4416
rect -240 4348 -228 4382
rect -194 4352 -156 4382
rect -194 4348 -182 4352
rect -240 4340 -182 4348
rect -12 4348 0 4382
rect 34 4348 46 4382
rect -12 4340 46 4348
rect -240 314 46 322
rect -240 280 -109 314
rect -75 280 46 314
rect -240 264 46 280
<< ndiffc >>
rect -228 4348 -194 4382
rect 0 4348 34 4382
<< pdiffc >>
rect 1005 5894 1039 5928
rect 1209 5894 1243 5928
rect 1005 5414 1039 5448
rect 1209 5414 1243 5448
<< mvndiffc >>
rect -228 4416 -194 4450
rect 0 4416 34 4450
rect -109 280 -75 314
<< psubdiff >>
rect 493 8052 527 8076
rect 493 7983 527 8018
rect 493 7914 527 7949
rect 493 7845 527 7880
rect 493 7776 527 7811
rect 493 7707 527 7742
rect 493 7638 527 7673
rect 493 7569 527 7604
rect 493 7500 527 7535
rect 493 7431 527 7466
rect 493 7363 527 7397
rect 493 7295 527 7329
rect 493 7227 527 7261
rect 493 7169 527 7193
rect 161 2110 185 2144
rect 219 2110 254 2144
rect 288 2110 323 2144
rect 357 2110 392 2144
rect 426 2110 461 2144
rect 495 2110 519 2144
rect 161 2076 519 2110
rect 161 2042 185 2076
rect 219 2042 254 2076
rect 288 2042 323 2076
rect 357 2042 392 2076
rect 426 2042 461 2076
rect 495 2042 519 2076
rect 161 2008 519 2042
rect 161 1974 185 2008
rect 219 1974 254 2008
rect 288 1974 323 2008
rect 357 1974 392 2008
rect 426 1974 461 2008
rect 495 1974 519 2008
rect 161 1940 519 1974
rect 161 1906 185 1940
rect 219 1906 254 1940
rect 288 1906 323 1940
rect 357 1906 392 1940
rect 426 1906 461 1940
rect 495 1906 519 1940
rect 161 1872 519 1906
rect 161 1838 185 1872
rect 219 1838 254 1872
rect 288 1838 323 1872
rect 357 1838 392 1872
rect 426 1838 461 1872
rect 495 1838 519 1872
rect 161 1804 519 1838
rect 161 1770 185 1804
rect 219 1770 254 1804
rect 288 1770 323 1804
rect 357 1770 392 1804
rect 426 1770 461 1804
rect 495 1770 519 1804
rect 485 1694 519 1770
rect 485 1622 519 1660
rect 485 1378 519 1588
rect 485 1306 519 1344
rect 485 1127 519 1272
rect 485 928 519 1093
rect 485 856 519 894
rect 485 784 519 822
rect 485 712 519 750
rect 485 640 519 678
rect 485 568 519 606
rect 485 496 519 534
rect 485 424 519 462
rect 485 352 519 390
rect 485 280 519 318
rect 485 172 519 246
rect 150 138 231 172
rect 265 138 303 172
rect 337 138 375 172
rect 409 138 447 172
rect 481 138 519 172
<< nsubdiff >>
rect 761 6004 891 6028
rect 795 5994 891 6004
rect 925 5994 968 6028
rect 1002 5994 1045 6028
rect 1079 5994 1122 6028
rect 1156 5994 1199 6028
rect 1233 5994 1276 6028
rect 1310 5994 1429 6028
rect 761 5935 795 5970
rect 761 5866 795 5901
rect 1395 5926 1429 5960
rect 761 5797 795 5832
rect 761 5728 795 5763
rect 761 5659 795 5694
rect 761 5590 795 5625
rect 761 5521 795 5556
rect 761 5452 795 5487
rect 1395 5858 1429 5892
rect 1395 5790 1429 5824
rect 1395 5722 1429 5756
rect 1395 5654 1429 5688
rect 1395 5586 1429 5620
rect 1395 5518 1429 5552
rect 761 5382 795 5418
rect 1395 5450 1429 5484
rect 761 5314 867 5348
rect 901 5314 937 5348
rect 971 5314 1007 5348
rect 1041 5314 1077 5348
rect 1111 5314 1148 5348
rect 1182 5314 1219 5348
rect 1253 5314 1290 5348
rect 1324 5314 1361 5348
rect 1395 5314 1429 5416
rect 701 1712 725 1746
rect 759 1712 797 1746
rect 831 1712 869 1746
rect 903 1712 940 1746
rect 974 1712 1011 1746
rect 1045 1712 1153 1746
rect 701 1581 735 1712
rect 701 1523 735 1547
rect 1119 1641 1153 1678
rect 1119 1570 1153 1607
rect 1119 1499 1153 1536
rect 1119 1428 1153 1465
rect 701 1303 735 1406
rect 701 1104 735 1269
rect 1119 1357 1153 1394
rect 1119 1286 1153 1323
rect 1119 1215 1153 1252
rect 1119 1144 1153 1181
rect 1119 1073 1153 1110
rect 701 920 735 1070
rect 701 851 735 886
rect 1119 1002 1153 1039
rect 1119 931 1153 968
rect 1119 860 1153 897
rect 701 782 735 817
rect 701 713 735 748
rect 701 644 735 679
rect 701 575 735 610
rect 701 506 735 541
rect 701 436 735 472
rect 701 366 735 402
rect 701 296 735 332
rect 1119 789 1153 826
rect 1119 718 1153 755
rect 1119 648 1153 684
rect 1119 578 1153 614
rect 1119 508 1153 544
rect 1119 438 1153 474
rect 1119 368 1153 404
rect 701 226 735 262
rect 1119 298 1153 334
rect 701 158 805 192
rect 839 158 875 192
rect 909 158 945 192
rect 979 158 1015 192
rect 1049 158 1085 192
rect 1119 158 1153 264
<< mvpsubdiff >>
rect 53 6852 123 6876
rect 87 6842 123 6852
rect 157 6842 203 6876
rect 237 6842 282 6876
rect 316 6842 361 6876
rect 395 6842 519 6876
rect 53 6782 87 6818
rect 53 6712 87 6748
rect 485 6773 519 6808
rect 53 6642 87 6678
rect 53 6572 87 6608
rect 53 6502 87 6538
rect 53 6432 87 6468
rect 485 6704 519 6739
rect 485 6635 519 6670
rect 485 6566 519 6601
rect 485 6497 519 6532
rect 3019 7908 3143 7942
rect 3177 7908 3211 7942
rect 3245 7908 3279 7942
rect 3313 7908 3347 7942
rect 3381 7908 3415 7942
rect 3449 7908 3483 7942
rect 3517 7908 3551 7942
rect 3585 7908 3619 7942
rect 3653 7908 3687 7942
rect 3721 7908 3755 7942
rect 3789 7908 3823 7942
rect 3019 7840 3053 7874
rect 3019 7772 3053 7806
rect 3857 7844 3891 7942
rect 3019 7704 3053 7738
rect 3019 7636 3053 7670
rect 3019 7568 3053 7602
rect 3019 7500 3053 7534
rect 3019 7432 3053 7466
rect 3019 7364 3053 7398
rect 3019 7296 3053 7330
rect 3019 7228 3053 7262
rect 3019 7160 3053 7194
rect 3857 7776 3891 7810
rect 3857 7708 3891 7742
rect 3857 7640 3891 7674
rect 3857 7572 3891 7606
rect 3857 7504 3891 7538
rect 3857 7436 3891 7470
rect 3857 7368 3891 7402
rect 3857 7300 3891 7334
rect 3857 7232 3891 7266
rect 3857 7164 3891 7198
rect 3019 7092 3053 7126
rect 3857 7096 3891 7130
rect 3019 7024 3053 7058
rect 3019 6956 3053 6990
rect 3019 6888 3053 6922
rect 3019 6820 3053 6854
rect 3019 6752 3053 6786
rect 3857 7028 3891 7062
rect 3857 6960 3891 6994
rect 3857 6892 3891 6926
rect 3857 6824 3891 6858
rect 3019 6620 3053 6718
rect 3857 6756 3891 6790
rect 3857 6688 3891 6722
rect 3087 6620 3121 6654
rect 3155 6620 3189 6654
rect 3223 6620 3257 6654
rect 3291 6620 3325 6654
rect 3359 6620 3393 6654
rect 3427 6620 3461 6654
rect 3495 6620 3529 6654
rect 3563 6620 3597 6654
rect 3631 6620 3665 6654
rect 3699 6620 3733 6654
rect 3767 6620 3891 6654
rect 53 6362 87 6398
rect 53 6292 87 6328
rect 485 6428 519 6463
rect 485 6359 519 6394
rect 53 6222 87 6258
rect 53 6152 87 6188
rect 485 6290 519 6325
rect 485 6221 519 6256
rect 485 6152 519 6187
rect 53 6082 87 6118
rect 485 6083 519 6118
rect 53 6012 87 6048
rect 53 5942 87 5978
rect 53 5872 87 5908
rect 53 5802 87 5838
rect 53 5732 87 5768
rect 53 5662 87 5698
rect 53 5592 87 5628
rect 53 5522 87 5558
rect 53 5452 87 5488
rect 53 5382 87 5418
rect 485 6014 519 6049
rect 485 5945 519 5980
rect 485 5876 519 5911
rect 485 5807 519 5842
rect 485 5738 519 5773
rect 485 5669 519 5704
rect 485 5600 519 5635
rect 485 5531 519 5566
rect 485 5462 519 5497
rect 485 5393 519 5428
rect 53 5312 87 5348
rect 485 5324 519 5359
rect 53 5242 87 5278
rect 53 5172 87 5208
rect 53 5102 87 5138
rect 53 5032 87 5068
rect 53 4962 87 4998
rect 485 5255 519 5290
rect 485 5186 519 5221
rect 485 5117 519 5152
rect 485 5048 519 5083
rect 485 4979 519 5014
rect 53 4892 87 4928
rect 485 4910 519 4945
rect 53 4822 87 4858
rect 53 4752 87 4788
rect -407 4576 -314 4745
rect 53 4681 87 4718
rect 53 4610 87 4647
rect -407 4542 -264 4576
rect -230 4542 -193 4576
rect -159 4542 -123 4576
rect -89 4542 -53 4576
rect -19 4542 87 4576
rect -407 3547 -314 4542
rect 485 4841 519 4876
rect 485 4772 519 4807
rect 485 4703 519 4738
rect 485 4634 519 4669
rect 485 4565 519 4600
rect 485 4496 519 4531
rect -393 3533 -314 3547
rect -380 3493 -314 3533
rect -380 3459 -348 3493
rect -380 3423 -314 3459
rect -380 3389 -348 3423
rect -380 3353 -314 3389
rect -380 3319 -348 3353
rect -380 3283 -314 3319
rect -380 3249 -348 3283
rect -380 3213 -314 3249
rect -380 3179 -348 3213
rect -380 3143 -314 3179
rect -380 3109 -348 3143
rect -380 3073 -314 3109
rect -380 3039 -348 3073
rect -380 3003 -314 3039
rect -380 2969 -348 3003
rect -380 2933 -314 2969
rect -380 2899 -348 2933
rect -380 2863 -314 2899
rect -380 2829 -348 2863
rect -380 2793 -314 2829
rect -380 2759 -348 2793
rect -380 2723 -314 2759
rect -380 2689 -348 2723
rect -380 2653 -314 2689
rect -380 2619 -348 2653
rect -380 2583 -314 2619
rect -380 2549 -348 2583
rect -380 2513 -314 2549
rect -380 2479 -348 2513
rect -380 2443 -314 2479
rect -380 2409 -348 2443
rect -380 2373 -314 2409
rect -380 2339 -348 2373
rect -380 2303 -314 2339
rect -380 2269 -348 2303
rect -380 2233 -314 2269
rect -380 2199 -348 2233
rect -380 2163 -314 2199
rect -380 2129 -348 2163
rect -380 2093 -314 2129
rect -380 2059 -348 2093
rect -380 2023 -314 2059
rect -380 1989 -348 2023
rect -380 1953 -314 1989
rect -380 1919 -348 1953
rect -380 1883 -314 1919
rect -380 1849 -348 1883
rect -380 1813 -314 1849
rect -380 1779 -348 1813
rect -380 1743 -314 1779
rect -380 1709 -348 1743
rect -380 1673 -314 1709
rect -380 1639 -348 1673
rect -380 1603 -314 1639
rect -380 1569 -348 1603
rect -380 1533 -314 1569
rect -380 1499 -348 1533
rect -380 1463 -314 1499
rect -380 1429 -348 1463
rect -380 1393 -314 1429
rect -380 1359 -348 1393
rect -380 1323 -314 1359
rect -380 1289 -348 1323
rect -380 1253 -314 1289
rect -380 1219 -348 1253
rect -380 1184 -314 1219
rect -380 1150 -348 1184
rect -380 1115 -314 1150
rect -380 1081 -348 1115
rect -380 1046 -314 1081
rect -380 1012 -348 1046
rect -380 751 -314 1012
rect -374 172 -314 751
rect 485 4427 519 4462
rect 485 4358 519 4393
rect 485 4289 519 4324
rect 485 4220 519 4255
rect 485 4151 519 4186
rect 485 4082 519 4117
rect 485 4013 519 4048
rect 485 3944 519 3979
rect 485 3875 519 3910
rect 485 3806 519 3841
rect 485 3737 519 3772
rect 485 3668 519 3703
rect 485 3599 519 3634
rect 485 3530 519 3565
rect 485 3461 519 3496
rect 485 3392 519 3427
rect 485 3323 519 3358
rect 485 3254 519 3289
rect 485 3185 519 3220
rect 485 3116 519 3151
rect 485 3047 519 3082
rect 485 2978 519 3013
rect 485 2909 519 2944
rect 485 2840 519 2875
rect 485 2772 519 2806
rect 485 2704 519 2738
rect 485 2636 519 2670
rect 485 2568 519 2602
rect 485 2500 519 2534
rect 485 2432 519 2466
rect 485 2364 519 2398
rect 161 2228 185 2262
rect 219 2228 273 2262
rect 307 2228 362 2262
rect 396 2228 451 2262
rect 485 2228 519 2330
rect -374 138 -280 172
rect -246 138 -210 172
rect -176 138 -140 172
rect -106 138 -70 172
rect -36 138 1 172
rect 35 138 59 172
<< mvnsubdiff >>
rect 741 7888 765 7922
rect 799 7888 836 7922
rect 870 7888 907 7922
rect 941 7888 977 7922
rect 1011 7888 1047 7922
rect 1081 7888 1117 7922
rect 1151 7888 1187 7922
rect 1221 7888 1257 7922
rect 1291 7888 1327 7922
rect 1361 7888 1397 7922
rect 1431 7888 1467 7922
rect 1501 7888 1537 7922
rect 1571 7888 1607 7922
rect 1641 7888 1677 7922
rect 1711 7888 1747 7922
rect 1781 7888 1817 7922
rect 1851 7888 1887 7922
rect 1921 7888 1957 7922
rect 1991 7888 2027 7922
rect 2061 7888 2097 7922
rect 2131 7888 2167 7922
rect 2201 7888 2237 7922
rect 2271 7888 2307 7922
rect 2341 7888 2377 7922
rect 2411 7888 2447 7922
rect 2481 7888 2517 7922
rect 2551 7888 2587 7922
rect 2621 7888 2657 7922
rect 2691 7888 2727 7922
rect 2761 7888 2867 7922
rect 741 7792 775 7888
rect 2833 7818 2867 7854
rect 741 7722 775 7758
rect 741 7652 775 7688
rect 741 7582 775 7618
rect 741 7512 775 7548
rect 741 7442 775 7478
rect 741 7372 775 7408
rect 741 7302 775 7338
rect 741 7232 775 7268
rect 741 7162 775 7198
rect 2833 7748 2867 7784
rect 2833 7678 2867 7714
rect 2833 7608 2867 7644
rect 2833 7538 2867 7574
rect 2833 7468 2867 7504
rect 2833 7399 2867 7434
rect 2833 7330 2867 7365
rect 2833 7261 2867 7296
rect 2833 7192 2867 7227
rect 741 7092 775 7128
rect 2833 7123 2867 7158
rect 741 7022 775 7058
rect 741 6952 775 6988
rect 741 6882 775 6918
rect 741 6811 775 6848
rect 741 6740 775 6777
rect 741 6669 775 6706
rect 2833 7054 2867 7089
rect 2833 6985 2867 7020
rect 2833 6916 2867 6951
rect 2833 6847 2867 6882
rect 2833 6778 2867 6813
rect 741 6598 775 6635
rect 1573 6640 1679 6674
rect 1713 6640 1749 6674
rect 1783 6640 1819 6674
rect 1853 6640 1889 6674
rect 1923 6640 1959 6674
rect 1993 6640 2029 6674
rect 2063 6640 2099 6674
rect 2133 6640 2169 6674
rect 2203 6640 2239 6674
rect 2273 6640 2309 6674
rect 2343 6640 2379 6674
rect 2413 6640 2449 6674
rect 2483 6640 2519 6674
rect 2553 6640 2589 6674
rect 2623 6640 2659 6674
rect 2693 6640 2729 6674
rect 2763 6640 2799 6674
rect 2833 6640 2867 6744
rect 741 6530 845 6564
rect 879 6530 914 6564
rect 948 6530 983 6564
rect 1017 6530 1052 6564
rect 1086 6530 1121 6564
rect 1155 6530 1190 6564
rect 1224 6530 1259 6564
rect 1293 6530 1329 6564
rect 1363 6530 1399 6564
rect 1433 6530 1469 6564
rect 1503 6530 1539 6564
rect 1573 6530 1607 6640
rect 701 4788 831 4812
rect 735 4778 831 4788
rect 865 4778 912 4812
rect 946 4778 993 4812
rect 1027 4778 1153 4812
rect 701 4720 735 4754
rect 701 4652 735 4686
rect 1119 4709 1153 4744
rect 701 4584 735 4618
rect 701 4516 735 4550
rect 1119 4640 1153 4675
rect 1119 4571 1153 4606
rect 701 4448 735 4482
rect 1119 4502 1153 4537
rect 701 4380 735 4414
rect 701 4312 735 4346
rect 1119 4433 1153 4468
rect 1119 4364 1153 4399
rect 701 4244 735 4278
rect 701 4176 735 4210
rect 701 4108 735 4142
rect 1119 4295 1153 4330
rect 1119 4226 1153 4261
rect 1119 4157 1153 4192
rect 701 4040 735 4074
rect 701 3972 735 4006
rect 701 3903 735 3938
rect 1119 4088 1153 4123
rect 1119 4019 1153 4054
rect 1119 3950 1153 3985
rect 701 3834 735 3869
rect 1119 3881 1153 3916
rect 701 3765 735 3800
rect 701 3696 735 3731
rect 701 3627 735 3662
rect 1119 3812 1153 3847
rect 1119 3744 1153 3778
rect 1119 3676 1153 3710
rect 701 3558 735 3593
rect 701 3489 735 3524
rect 1119 3608 1153 3642
rect 1119 3540 1153 3574
rect 1119 3472 1153 3506
rect 701 3420 735 3455
rect 701 3351 735 3386
rect 701 3282 735 3317
rect 1119 3404 1153 3438
rect 1119 3336 1153 3370
rect 1119 3268 1153 3302
rect 701 3213 735 3248
rect 701 3144 735 3179
rect 701 3075 735 3110
rect 701 3006 735 3041
rect 1119 3200 1153 3234
rect 1119 3132 1153 3166
rect 1119 3064 1153 3098
rect 701 2937 735 2972
rect 701 2868 735 2903
rect 1119 2996 1153 3030
rect 1119 2928 1153 2962
rect 1119 2860 1153 2894
rect 701 2799 735 2834
rect 701 2730 735 2765
rect 701 2661 735 2696
rect 1119 2792 1153 2826
rect 1119 2724 1153 2758
rect 1119 2656 1153 2690
rect 701 2592 735 2627
rect 701 2523 735 2558
rect 701 2454 735 2489
rect 701 2385 735 2420
rect 1119 2588 1153 2622
rect 1119 2520 1153 2554
rect 1119 2452 1153 2486
rect 701 2316 735 2351
rect 1119 2384 1153 2418
rect 701 2248 805 2282
rect 839 2248 875 2282
rect 909 2248 945 2282
rect 979 2248 1015 2282
rect 1049 2248 1085 2282
rect 1119 2248 1153 2350
<< psubdiffcont >>
rect 493 8018 527 8052
rect 493 7949 527 7983
rect 493 7880 527 7914
rect 493 7811 527 7845
rect 493 7742 527 7776
rect 493 7673 527 7707
rect 493 7604 527 7638
rect 493 7535 527 7569
rect 493 7466 527 7500
rect 493 7397 527 7431
rect 493 7329 527 7363
rect 493 7261 527 7295
rect 493 7193 527 7227
rect 185 2110 219 2144
rect 254 2110 288 2144
rect 323 2110 357 2144
rect 392 2110 426 2144
rect 461 2110 495 2144
rect 185 2042 219 2076
rect 254 2042 288 2076
rect 323 2042 357 2076
rect 392 2042 426 2076
rect 461 2042 495 2076
rect 185 1974 219 2008
rect 254 1974 288 2008
rect 323 1974 357 2008
rect 392 1974 426 2008
rect 461 1974 495 2008
rect 185 1906 219 1940
rect 254 1906 288 1940
rect 323 1906 357 1940
rect 392 1906 426 1940
rect 461 1906 495 1940
rect 185 1838 219 1872
rect 254 1838 288 1872
rect 323 1838 357 1872
rect 392 1838 426 1872
rect 461 1838 495 1872
rect 185 1770 219 1804
rect 254 1770 288 1804
rect 323 1770 357 1804
rect 392 1770 426 1804
rect 461 1770 495 1804
rect 485 1660 519 1694
rect 485 1588 519 1622
rect 485 1344 519 1378
rect 485 1272 519 1306
rect 485 1093 519 1127
rect 485 894 519 928
rect 485 822 519 856
rect 485 750 519 784
rect 485 678 519 712
rect 485 606 519 640
rect 485 534 519 568
rect 485 462 519 496
rect 485 390 519 424
rect 485 318 519 352
rect 485 246 519 280
rect 231 138 265 172
rect 303 138 337 172
rect 375 138 409 172
rect 447 138 481 172
<< nsubdiffcont >>
rect 761 5970 795 6004
rect 891 5994 925 6028
rect 968 5994 1002 6028
rect 1045 5994 1079 6028
rect 1122 5994 1156 6028
rect 1199 5994 1233 6028
rect 1276 5994 1310 6028
rect 1395 5960 1429 5994
rect 761 5901 795 5935
rect 1395 5892 1429 5926
rect 761 5832 795 5866
rect 761 5763 795 5797
rect 761 5694 795 5728
rect 761 5625 795 5659
rect 761 5556 795 5590
rect 761 5487 795 5521
rect 1395 5824 1429 5858
rect 1395 5756 1429 5790
rect 1395 5688 1429 5722
rect 1395 5620 1429 5654
rect 1395 5552 1429 5586
rect 1395 5484 1429 5518
rect 761 5418 795 5452
rect 1395 5416 1429 5450
rect 761 5348 795 5382
rect 867 5314 901 5348
rect 937 5314 971 5348
rect 1007 5314 1041 5348
rect 1077 5314 1111 5348
rect 1148 5314 1182 5348
rect 1219 5314 1253 5348
rect 1290 5314 1324 5348
rect 1361 5314 1395 5348
rect 725 1712 759 1746
rect 797 1712 831 1746
rect 869 1712 903 1746
rect 940 1712 974 1746
rect 1011 1712 1045 1746
rect 1119 1678 1153 1712
rect 701 1547 735 1581
rect 1119 1607 1153 1641
rect 1119 1536 1153 1570
rect 1119 1465 1153 1499
rect 1119 1394 1153 1428
rect 701 1269 735 1303
rect 1119 1323 1153 1357
rect 1119 1252 1153 1286
rect 701 1070 735 1104
rect 1119 1181 1153 1215
rect 1119 1110 1153 1144
rect 701 886 735 920
rect 1119 1039 1153 1073
rect 1119 968 1153 1002
rect 1119 897 1153 931
rect 701 817 735 851
rect 1119 826 1153 860
rect 701 748 735 782
rect 701 679 735 713
rect 701 610 735 644
rect 701 541 735 575
rect 701 472 735 506
rect 701 402 735 436
rect 701 332 735 366
rect 1119 755 1153 789
rect 1119 684 1153 718
rect 1119 614 1153 648
rect 1119 544 1153 578
rect 1119 474 1153 508
rect 1119 404 1153 438
rect 1119 334 1153 368
rect 701 262 735 296
rect 701 192 735 226
rect 1119 264 1153 298
rect 805 158 839 192
rect 875 158 909 192
rect 945 158 979 192
rect 1015 158 1049 192
rect 1085 158 1119 192
<< mvpsubdiffcont >>
rect 53 6818 87 6852
rect 123 6842 157 6876
rect 203 6842 237 6876
rect 282 6842 316 6876
rect 361 6842 395 6876
rect 53 6748 87 6782
rect 485 6808 519 6842
rect 485 6739 519 6773
rect 53 6678 87 6712
rect 53 6608 87 6642
rect 53 6538 87 6572
rect 53 6468 87 6502
rect 485 6670 519 6704
rect 485 6601 519 6635
rect 485 6532 519 6566
rect 3143 7908 3177 7942
rect 3211 7908 3245 7942
rect 3279 7908 3313 7942
rect 3347 7908 3381 7942
rect 3415 7908 3449 7942
rect 3483 7908 3517 7942
rect 3551 7908 3585 7942
rect 3619 7908 3653 7942
rect 3687 7908 3721 7942
rect 3755 7908 3789 7942
rect 3823 7908 3857 7942
rect 3019 7874 3053 7908
rect 3019 7806 3053 7840
rect 3857 7810 3891 7844
rect 3019 7738 3053 7772
rect 3019 7670 3053 7704
rect 3019 7602 3053 7636
rect 3019 7534 3053 7568
rect 3019 7466 3053 7500
rect 3019 7398 3053 7432
rect 3019 7330 3053 7364
rect 3019 7262 3053 7296
rect 3019 7194 3053 7228
rect 3019 7126 3053 7160
rect 3857 7742 3891 7776
rect 3857 7674 3891 7708
rect 3857 7606 3891 7640
rect 3857 7538 3891 7572
rect 3857 7470 3891 7504
rect 3857 7402 3891 7436
rect 3857 7334 3891 7368
rect 3857 7266 3891 7300
rect 3857 7198 3891 7232
rect 3019 7058 3053 7092
rect 3857 7130 3891 7164
rect 3019 6990 3053 7024
rect 3019 6922 3053 6956
rect 3019 6854 3053 6888
rect 3019 6786 3053 6820
rect 3857 7062 3891 7096
rect 3857 6994 3891 7028
rect 3857 6926 3891 6960
rect 3857 6858 3891 6892
rect 3857 6790 3891 6824
rect 3019 6718 3053 6752
rect 3857 6722 3891 6756
rect 3857 6654 3891 6688
rect 3053 6620 3087 6654
rect 3121 6620 3155 6654
rect 3189 6620 3223 6654
rect 3257 6620 3291 6654
rect 3325 6620 3359 6654
rect 3393 6620 3427 6654
rect 3461 6620 3495 6654
rect 3529 6620 3563 6654
rect 3597 6620 3631 6654
rect 3665 6620 3699 6654
rect 3733 6620 3767 6654
rect 485 6463 519 6497
rect 53 6398 87 6432
rect 53 6328 87 6362
rect 485 6394 519 6428
rect 485 6325 519 6359
rect 53 6258 87 6292
rect 53 6188 87 6222
rect 53 6118 87 6152
rect 485 6256 519 6290
rect 485 6187 519 6221
rect 53 6048 87 6082
rect 485 6118 519 6152
rect 53 5978 87 6012
rect 53 5908 87 5942
rect 53 5838 87 5872
rect 53 5768 87 5802
rect 53 5698 87 5732
rect 53 5628 87 5662
rect 53 5558 87 5592
rect 53 5488 87 5522
rect 53 5418 87 5452
rect 53 5348 87 5382
rect 485 6049 519 6083
rect 485 5980 519 6014
rect 485 5911 519 5945
rect 485 5842 519 5876
rect 485 5773 519 5807
rect 485 5704 519 5738
rect 485 5635 519 5669
rect 485 5566 519 5600
rect 485 5497 519 5531
rect 485 5428 519 5462
rect 485 5359 519 5393
rect 53 5278 87 5312
rect 53 5208 87 5242
rect 53 5138 87 5172
rect 53 5068 87 5102
rect 53 4998 87 5032
rect 53 4928 87 4962
rect 485 5290 519 5324
rect 485 5221 519 5255
rect 485 5152 519 5186
rect 485 5083 519 5117
rect 485 5014 519 5048
rect 485 4945 519 4979
rect 53 4858 87 4892
rect 53 4788 87 4822
rect 53 4718 87 4752
rect 53 4647 87 4681
rect 53 4576 87 4610
rect -264 4542 -230 4576
rect -193 4542 -159 4576
rect -123 4542 -89 4576
rect -53 4542 -19 4576
rect 485 4876 519 4910
rect 485 4807 519 4841
rect 485 4738 519 4772
rect 485 4669 519 4703
rect 485 4600 519 4634
rect 485 4531 519 4565
rect 485 4462 519 4496
rect -348 3459 -314 3493
rect -348 3389 -314 3423
rect -348 3319 -314 3353
rect -348 3249 -314 3283
rect -348 3179 -314 3213
rect -348 3109 -314 3143
rect -348 3039 -314 3073
rect -348 2969 -314 3003
rect -348 2899 -314 2933
rect -348 2829 -314 2863
rect -348 2759 -314 2793
rect -348 2689 -314 2723
rect -348 2619 -314 2653
rect -348 2549 -314 2583
rect -348 2479 -314 2513
rect -348 2409 -314 2443
rect -348 2339 -314 2373
rect -348 2269 -314 2303
rect -348 2199 -314 2233
rect -348 2129 -314 2163
rect -348 2059 -314 2093
rect -348 1989 -314 2023
rect -348 1919 -314 1953
rect -348 1849 -314 1883
rect -348 1779 -314 1813
rect -348 1709 -314 1743
rect -348 1639 -314 1673
rect -348 1569 -314 1603
rect -348 1499 -314 1533
rect -348 1429 -314 1463
rect -348 1359 -314 1393
rect -348 1289 -314 1323
rect -348 1219 -314 1253
rect -348 1150 -314 1184
rect -348 1081 -314 1115
rect -348 1012 -314 1046
rect 485 4393 519 4427
rect 485 4324 519 4358
rect 485 4255 519 4289
rect 485 4186 519 4220
rect 485 4117 519 4151
rect 485 4048 519 4082
rect 485 3979 519 4013
rect 485 3910 519 3944
rect 485 3841 519 3875
rect 485 3772 519 3806
rect 485 3703 519 3737
rect 485 3634 519 3668
rect 485 3565 519 3599
rect 485 3496 519 3530
rect 485 3427 519 3461
rect 485 3358 519 3392
rect 485 3289 519 3323
rect 485 3220 519 3254
rect 485 3151 519 3185
rect 485 3082 519 3116
rect 485 3013 519 3047
rect 485 2944 519 2978
rect 485 2875 519 2909
rect 485 2806 519 2840
rect 485 2738 519 2772
rect 485 2670 519 2704
rect 485 2602 519 2636
rect 485 2534 519 2568
rect 485 2466 519 2500
rect 485 2398 519 2432
rect 485 2330 519 2364
rect 185 2228 219 2262
rect 273 2228 307 2262
rect 362 2228 396 2262
rect 451 2228 485 2262
rect -280 138 -246 172
rect -210 138 -176 172
rect -140 138 -106 172
rect -70 138 -36 172
rect 1 138 35 172
<< mvnsubdiffcont >>
rect 765 7888 799 7922
rect 836 7888 870 7922
rect 907 7888 941 7922
rect 977 7888 1011 7922
rect 1047 7888 1081 7922
rect 1117 7888 1151 7922
rect 1187 7888 1221 7922
rect 1257 7888 1291 7922
rect 1327 7888 1361 7922
rect 1397 7888 1431 7922
rect 1467 7888 1501 7922
rect 1537 7888 1571 7922
rect 1607 7888 1641 7922
rect 1677 7888 1711 7922
rect 1747 7888 1781 7922
rect 1817 7888 1851 7922
rect 1887 7888 1921 7922
rect 1957 7888 1991 7922
rect 2027 7888 2061 7922
rect 2097 7888 2131 7922
rect 2167 7888 2201 7922
rect 2237 7888 2271 7922
rect 2307 7888 2341 7922
rect 2377 7888 2411 7922
rect 2447 7888 2481 7922
rect 2517 7888 2551 7922
rect 2587 7888 2621 7922
rect 2657 7888 2691 7922
rect 2727 7888 2761 7922
rect 741 7758 775 7792
rect 2833 7854 2867 7888
rect 2833 7784 2867 7818
rect 741 7688 775 7722
rect 741 7618 775 7652
rect 741 7548 775 7582
rect 741 7478 775 7512
rect 741 7408 775 7442
rect 741 7338 775 7372
rect 741 7268 775 7302
rect 741 7198 775 7232
rect 741 7128 775 7162
rect 2833 7714 2867 7748
rect 2833 7644 2867 7678
rect 2833 7574 2867 7608
rect 2833 7504 2867 7538
rect 2833 7434 2867 7468
rect 2833 7365 2867 7399
rect 2833 7296 2867 7330
rect 2833 7227 2867 7261
rect 2833 7158 2867 7192
rect 741 7058 775 7092
rect 2833 7089 2867 7123
rect 741 6988 775 7022
rect 741 6918 775 6952
rect 741 6848 775 6882
rect 741 6777 775 6811
rect 741 6706 775 6740
rect 2833 7020 2867 7054
rect 2833 6951 2867 6985
rect 2833 6882 2867 6916
rect 2833 6813 2867 6847
rect 2833 6744 2867 6778
rect 741 6635 775 6669
rect 741 6564 775 6598
rect 1679 6640 1713 6674
rect 1749 6640 1783 6674
rect 1819 6640 1853 6674
rect 1889 6640 1923 6674
rect 1959 6640 1993 6674
rect 2029 6640 2063 6674
rect 2099 6640 2133 6674
rect 2169 6640 2203 6674
rect 2239 6640 2273 6674
rect 2309 6640 2343 6674
rect 2379 6640 2413 6674
rect 2449 6640 2483 6674
rect 2519 6640 2553 6674
rect 2589 6640 2623 6674
rect 2659 6640 2693 6674
rect 2729 6640 2763 6674
rect 2799 6640 2833 6674
rect 845 6530 879 6564
rect 914 6530 948 6564
rect 983 6530 1017 6564
rect 1052 6530 1086 6564
rect 1121 6530 1155 6564
rect 1190 6530 1224 6564
rect 1259 6530 1293 6564
rect 1329 6530 1363 6564
rect 1399 6530 1433 6564
rect 1469 6530 1503 6564
rect 1539 6530 1573 6564
rect 701 4754 735 4788
rect 831 4778 865 4812
rect 912 4778 946 4812
rect 993 4778 1027 4812
rect 701 4686 735 4720
rect 1119 4744 1153 4778
rect 1119 4675 1153 4709
rect 701 4618 735 4652
rect 701 4550 735 4584
rect 701 4482 735 4516
rect 1119 4606 1153 4640
rect 1119 4537 1153 4571
rect 1119 4468 1153 4502
rect 701 4414 735 4448
rect 701 4346 735 4380
rect 1119 4399 1153 4433
rect 1119 4330 1153 4364
rect 701 4278 735 4312
rect 701 4210 735 4244
rect 701 4142 735 4176
rect 701 4074 735 4108
rect 1119 4261 1153 4295
rect 1119 4192 1153 4226
rect 1119 4123 1153 4157
rect 701 4006 735 4040
rect 701 3938 735 3972
rect 701 3869 735 3903
rect 1119 4054 1153 4088
rect 1119 3985 1153 4019
rect 1119 3916 1153 3950
rect 701 3800 735 3834
rect 1119 3847 1153 3881
rect 701 3731 735 3765
rect 701 3662 735 3696
rect 1119 3778 1153 3812
rect 1119 3710 1153 3744
rect 1119 3642 1153 3676
rect 701 3593 735 3627
rect 701 3524 735 3558
rect 701 3455 735 3489
rect 1119 3574 1153 3608
rect 1119 3506 1153 3540
rect 701 3386 735 3420
rect 701 3317 735 3351
rect 701 3248 735 3282
rect 1119 3438 1153 3472
rect 1119 3370 1153 3404
rect 1119 3302 1153 3336
rect 701 3179 735 3213
rect 1119 3234 1153 3268
rect 701 3110 735 3144
rect 701 3041 735 3075
rect 1119 3166 1153 3200
rect 1119 3098 1153 3132
rect 1119 3030 1153 3064
rect 701 2972 735 3006
rect 701 2903 735 2937
rect 701 2834 735 2868
rect 1119 2962 1153 2996
rect 1119 2894 1153 2928
rect 701 2765 735 2799
rect 701 2696 735 2730
rect 701 2627 735 2661
rect 1119 2826 1153 2860
rect 1119 2758 1153 2792
rect 1119 2690 1153 2724
rect 701 2558 735 2592
rect 1119 2622 1153 2656
rect 701 2489 735 2523
rect 701 2420 735 2454
rect 1119 2554 1153 2588
rect 1119 2486 1153 2520
rect 1119 2418 1153 2452
rect 701 2351 735 2385
rect 701 2282 735 2316
rect 1119 2350 1153 2384
rect 805 2248 839 2282
rect 875 2248 909 2282
rect 945 2248 979 2282
rect 1015 2248 1049 2282
rect 1085 2248 1119 2282
<< poly >>
rect 1161 7765 1253 7781
rect 1161 7731 1203 7765
rect 1237 7731 1253 7765
rect 1161 7670 1253 7731
rect 1161 7636 1203 7670
rect 1237 7636 1253 7670
rect 1161 7575 1253 7636
rect 1161 7541 1203 7575
rect 1237 7541 1253 7575
rect 1161 7525 1253 7541
rect 1999 7765 2077 7781
rect 1999 7731 2021 7765
rect 2055 7731 2077 7765
rect 1999 7692 2077 7731
rect 1999 7658 2021 7692
rect 2055 7658 2077 7692
rect 1999 7619 2077 7658
rect 1999 7585 2021 7619
rect 2055 7585 2077 7619
rect 1999 7546 2077 7585
rect 1999 7512 2021 7546
rect 2055 7512 2077 7546
rect 1999 7473 2077 7512
rect 1161 7453 1253 7469
rect 1161 7419 1203 7453
rect 1237 7419 1253 7453
rect 1161 7358 1253 7419
rect 1161 7324 1203 7358
rect 1237 7324 1253 7358
rect 1161 7263 1253 7324
rect 1161 7229 1203 7263
rect 1237 7229 1253 7263
rect 1161 7213 1253 7229
rect 1999 7439 2021 7473
rect 2055 7439 2077 7473
rect 1999 7400 2077 7439
rect 1999 7366 2021 7400
rect 2055 7366 2077 7400
rect 1999 7327 2077 7366
rect 1999 7293 2021 7327
rect 2055 7293 2077 7327
rect 1999 7255 2077 7293
rect 1999 7221 2021 7255
rect 2055 7221 2077 7255
rect 1999 7183 2077 7221
rect 1999 7149 2021 7183
rect 2055 7149 2077 7183
rect 1999 7133 2077 7149
rect 2729 7765 2801 7781
rect 2729 7731 2751 7765
rect 2785 7731 2801 7765
rect 2729 7692 2801 7731
rect 2729 7658 2751 7692
rect 2785 7658 2801 7692
rect 2729 7619 2801 7658
rect 2729 7585 2751 7619
rect 2785 7585 2801 7619
rect 2729 7546 2801 7585
rect 2729 7512 2751 7546
rect 2785 7512 2801 7546
rect 2729 7473 2801 7512
rect 2729 7439 2751 7473
rect 2785 7439 2801 7473
rect 2729 7400 2801 7439
rect 2729 7366 2751 7400
rect 2785 7366 2801 7400
rect 2729 7327 2801 7366
rect 2729 7293 2751 7327
rect 2785 7293 2801 7327
rect 2729 7255 2801 7293
rect 2729 7221 2751 7255
rect 2785 7221 2801 7255
rect 2729 7183 2801 7221
rect 2729 7149 2751 7183
rect 2785 7149 2801 7183
rect 2729 7133 2801 7149
rect 1999 7061 2077 7077
rect 1061 7031 1133 7047
rect 1061 6997 1083 7031
rect 1117 6997 1133 7031
rect 1061 6937 1133 6997
rect 1061 6903 1083 6937
rect 1117 6903 1133 6937
rect 1061 6887 1133 6903
rect 1999 7027 2021 7061
rect 2055 7027 2077 7061
rect 1999 6984 2077 7027
rect 1999 6950 2021 6984
rect 2055 6950 2077 6984
rect 1999 6907 2077 6950
rect 387 6699 453 6715
rect 387 6665 403 6699
rect 437 6665 453 6699
rect 387 6604 453 6665
rect 387 6570 403 6604
rect 437 6570 453 6604
rect 387 6509 453 6570
rect 387 6475 403 6509
rect 437 6475 453 6509
rect 387 6459 453 6475
rect 1999 6873 2021 6907
rect 2055 6873 2077 6907
rect 1999 6831 2077 6873
rect 1061 6815 1198 6831
rect 1061 6781 1148 6815
rect 1182 6781 1198 6815
rect 1999 6797 2021 6831
rect 2055 6797 2077 6831
rect 1999 6781 2077 6797
rect 2729 7061 2801 7077
rect 2729 7027 2751 7061
rect 2785 7027 2801 7061
rect 2729 6984 2801 7027
rect 2729 6950 2751 6984
rect 2785 6950 2801 6984
rect 2729 6907 2801 6950
rect 2729 6873 2751 6907
rect 2785 6873 2801 6907
rect 2729 6831 2801 6873
rect 2729 6797 2751 6831
rect 2785 6797 2801 6831
rect 2729 6781 2801 6797
rect 1061 6721 1198 6781
rect 1061 6687 1148 6721
rect 1182 6687 1198 6721
rect 1061 6671 1198 6687
rect 3085 7765 3157 7781
rect 3085 7731 3101 7765
rect 3135 7731 3157 7765
rect 3085 7693 3157 7731
rect 3085 7659 3101 7693
rect 3135 7659 3157 7693
rect 3085 7621 3157 7659
rect 3085 7587 3101 7621
rect 3135 7587 3157 7621
rect 3085 7548 3157 7587
rect 3085 7514 3101 7548
rect 3135 7514 3157 7548
rect 3085 7475 3157 7514
rect 3085 7441 3101 7475
rect 3135 7441 3157 7475
rect 3085 7402 3157 7441
rect 3085 7368 3101 7402
rect 3135 7368 3157 7402
rect 3085 7329 3157 7368
rect 3085 7295 3101 7329
rect 3135 7295 3157 7329
rect 3085 7256 3157 7295
rect 3085 7222 3101 7256
rect 3135 7222 3157 7256
rect 3085 7183 3157 7222
rect 3085 7149 3101 7183
rect 3135 7149 3157 7183
rect 3085 7133 3157 7149
rect 3085 7061 3157 7077
rect 3085 7027 3101 7061
rect 3135 7027 3157 7061
rect 3085 6984 3157 7027
rect 3085 6950 3101 6984
rect 3135 6950 3157 6984
rect 3085 6907 3157 6950
rect 3085 6873 3101 6907
rect 3135 6873 3157 6907
rect 3085 6831 3157 6873
rect 3085 6797 3101 6831
rect 3135 6797 3157 6831
rect 3085 6781 3157 6797
rect 387 6277 453 6293
rect 387 6243 403 6277
rect 437 6243 453 6277
rect 387 6183 453 6243
rect 387 6149 403 6183
rect 437 6149 453 6183
rect 387 6133 453 6149
rect 387 6061 453 6077
rect 387 6027 403 6061
rect 437 6027 453 6061
rect 387 5967 453 6027
rect 387 5933 403 5967
rect 437 5933 453 5967
rect 387 5735 453 5933
rect 387 5701 403 5735
rect 437 5701 453 5735
rect 387 5657 453 5701
rect 387 5623 403 5657
rect 437 5623 453 5657
rect 387 5579 453 5623
rect 387 5545 403 5579
rect 437 5545 453 5579
rect 387 5502 453 5545
rect 387 5468 403 5502
rect 437 5468 453 5502
rect 387 5425 453 5468
rect 387 5391 403 5425
rect 437 5391 453 5425
rect 387 5375 453 5391
rect 387 5303 453 5319
rect 387 5269 403 5303
rect 437 5269 453 5303
rect 387 5225 453 5269
rect 387 5191 403 5225
rect 437 5191 453 5225
rect 387 5147 453 5191
rect 387 5113 403 5147
rect 437 5113 453 5147
rect 387 5070 453 5113
rect 387 5036 403 5070
rect 437 5036 453 5070
rect 387 4993 453 5036
rect 387 4959 403 4993
rect 437 4959 453 4993
rect 387 4943 453 4959
rect 827 5855 899 5871
rect 827 5821 843 5855
rect 877 5821 899 5855
rect 827 5772 899 5821
rect 827 5738 843 5772
rect 877 5738 899 5772
rect 827 5689 899 5738
rect 827 5655 843 5689
rect 877 5655 899 5689
rect 827 5605 899 5655
rect 827 5571 843 5605
rect 877 5571 899 5605
rect 827 5521 899 5571
rect 827 5487 843 5521
rect 877 5487 899 5521
rect 827 5471 899 5487
rect 1265 5855 1363 5871
rect 1265 5821 1313 5855
rect 1347 5821 1363 5855
rect 1265 5771 1363 5821
rect 1265 5737 1313 5771
rect 1347 5737 1363 5771
rect 1265 5687 1363 5737
rect 1265 5653 1313 5687
rect 1347 5653 1363 5687
rect 1265 5604 1363 5653
rect 1265 5570 1313 5604
rect 1347 5570 1363 5604
rect 1265 5521 1363 5570
rect 1265 5487 1313 5521
rect 1347 5487 1363 5521
rect 1265 5471 1363 5487
rect 387 4871 453 4887
rect 387 4837 403 4871
rect 437 4837 453 4871
rect 387 4793 453 4837
rect 387 4759 403 4793
rect 437 4759 453 4793
rect 387 4715 453 4759
rect 387 4681 403 4715
rect 437 4681 453 4715
rect 387 4638 453 4681
rect 387 4604 403 4638
rect 437 4604 453 4638
rect 387 4561 453 4604
rect 387 4527 403 4561
rect 437 4527 453 4561
rect 387 4511 453 4527
rect 387 4439 453 4455
rect 387 4405 403 4439
rect 437 4405 453 4439
rect 387 4371 453 4405
rect 387 4337 403 4371
rect 437 4337 453 4371
rect -130 4321 -64 4337
rect 387 4321 453 4337
rect -130 4287 -114 4321
rect -80 4287 -64 4321
rect -130 4252 -64 4287
rect -130 4218 -114 4252
rect -80 4218 -64 4252
rect -130 4183 -64 4218
rect -130 4149 -114 4183
rect -80 4149 -64 4183
rect -130 4114 -64 4149
rect -130 4080 -114 4114
rect -80 4080 -64 4114
rect -130 4045 -64 4080
rect -130 4011 -114 4045
rect -80 4011 -64 4045
rect -130 3976 -64 4011
rect -130 3942 -114 3976
rect -80 3942 -64 3976
rect 387 4073 453 4089
rect 387 4039 403 4073
rect 437 4039 453 4073
rect 387 3996 453 4039
rect 387 3962 403 3996
rect 437 3962 453 3996
rect 387 3946 453 3962
rect -130 3907 -64 3942
rect -130 3873 -114 3907
rect -80 3873 -64 3907
rect -130 3838 -64 3873
rect -130 3804 -114 3838
rect -80 3804 -64 3838
rect -130 3769 -64 3804
rect -130 3735 -114 3769
rect -80 3735 -64 3769
rect -130 3700 -64 3735
rect -130 3666 -114 3700
rect -80 3666 -64 3700
rect -130 3631 -64 3666
rect 387 3817 453 3833
rect 387 3783 403 3817
rect 437 3783 453 3817
rect 387 3706 453 3783
rect 387 3672 403 3706
rect 437 3672 453 3706
rect 387 3656 453 3672
rect -130 3597 -114 3631
rect -80 3597 -64 3631
rect -130 3562 -64 3597
rect -130 3528 -114 3562
rect -80 3528 -64 3562
rect -130 3493 -64 3528
rect -130 3459 -114 3493
rect -80 3459 -64 3493
rect -130 3424 -64 3459
rect -130 3390 -114 3424
rect -80 3390 -64 3424
rect -130 3355 -64 3390
rect -130 3321 -114 3355
rect -80 3321 -64 3355
rect -130 3286 -64 3321
rect -130 3252 -114 3286
rect -80 3252 -64 3286
rect 387 3451 453 3467
rect 387 3417 403 3451
rect 437 3417 453 3451
rect 387 3317 453 3417
rect 387 3283 403 3317
rect 437 3283 453 3317
rect 387 3267 453 3283
rect -130 3217 -64 3252
rect -130 3183 -114 3217
rect -80 3183 -64 3217
rect -130 3148 -64 3183
rect -130 3114 -114 3148
rect -80 3114 -64 3148
rect -130 3079 -64 3114
rect -130 3045 -114 3079
rect -80 3045 -64 3079
rect -130 3010 -64 3045
rect 387 3195 453 3211
rect 387 3161 403 3195
rect 437 3161 453 3195
rect 387 3084 453 3161
rect 387 3050 403 3084
rect 437 3050 453 3084
rect 387 3034 453 3050
rect -130 2976 -114 3010
rect -80 2976 -64 3010
rect -130 2941 -64 2976
rect -130 2907 -114 2941
rect -80 2907 -64 2941
rect -130 2872 -64 2907
rect -130 2838 -114 2872
rect -80 2838 -64 2872
rect -130 2803 -64 2838
rect -130 2769 -114 2803
rect -80 2769 -64 2803
rect -130 2734 -64 2769
rect -130 2700 -114 2734
rect -80 2700 -64 2734
rect -130 2665 -64 2700
rect -130 2631 -114 2665
rect -80 2631 -64 2665
rect 387 2829 453 2845
rect 387 2795 403 2829
rect 437 2795 453 2829
rect 387 2695 453 2795
rect 387 2661 403 2695
rect 437 2661 453 2695
rect 387 2645 453 2661
rect -130 2596 -64 2631
rect -130 2562 -114 2596
rect -80 2562 -64 2596
rect -130 2527 -64 2562
rect -130 2493 -114 2527
rect -80 2493 -64 2527
rect -130 2458 -64 2493
rect -130 2424 -114 2458
rect -80 2424 -64 2458
rect -130 2389 -64 2424
rect 387 2573 453 2589
rect 387 2539 403 2573
rect 437 2539 453 2573
rect 387 2439 453 2539
rect 387 2405 403 2439
rect 437 2405 453 2439
rect 387 2389 453 2405
rect -130 2355 -114 2389
rect -80 2355 -64 2389
rect -130 2320 -64 2355
rect -130 2286 -114 2320
rect -80 2286 -64 2320
rect -130 2251 -64 2286
rect -130 2217 -114 2251
rect -80 2217 -64 2251
rect 767 4655 839 4671
rect 767 4621 783 4655
rect 817 4621 839 4655
rect 767 4561 839 4621
rect 767 4527 783 4561
rect 817 4527 839 4561
rect 767 4511 839 4527
rect 767 4439 839 4455
rect 767 4405 783 4439
rect 817 4405 839 4439
rect 767 4371 839 4405
rect 767 4337 783 4371
rect 817 4337 839 4371
rect 767 4321 839 4337
rect 767 4073 839 4089
rect 767 4039 783 4073
rect 817 4039 839 4073
rect 767 3939 839 4039
rect 767 3905 783 3939
rect 817 3905 839 3939
rect 767 3889 839 3905
rect 767 3817 839 3833
rect 767 3783 783 3817
rect 817 3783 839 3817
rect 767 3706 839 3783
rect 767 3672 783 3706
rect 817 3672 839 3706
rect 767 3656 839 3672
rect 833 3633 839 3656
rect 767 3451 839 3467
rect 767 3417 783 3451
rect 817 3417 839 3451
rect 767 3317 839 3417
rect 767 3283 783 3317
rect 817 3283 839 3317
rect 767 3267 839 3283
rect 767 3195 839 3211
rect 767 3161 783 3195
rect 817 3161 839 3195
rect 767 3084 839 3161
rect 767 3050 783 3084
rect 817 3050 839 3084
rect 767 3034 839 3050
rect 833 3011 839 3034
rect 767 2829 839 2845
rect 767 2795 783 2829
rect 817 2795 839 2829
rect 767 2695 839 2795
rect 767 2661 783 2695
rect 817 2661 839 2695
rect 767 2645 839 2661
rect 767 2573 839 2589
rect 767 2539 783 2573
rect 817 2539 839 2573
rect 767 2439 839 2539
rect 767 2405 783 2439
rect 817 2405 839 2439
rect 767 2389 839 2405
rect -130 2182 -64 2217
rect -130 2148 -114 2182
rect -80 2148 -64 2182
rect -130 2113 -64 2148
rect -130 2079 -114 2113
rect -80 2079 -64 2113
rect -130 2044 -64 2079
rect -130 2010 -114 2044
rect -80 2010 -64 2044
rect -130 1975 -64 2010
rect -130 1941 -114 1975
rect -80 1941 -64 1975
rect -130 1906 -64 1941
rect -130 1872 -114 1906
rect -80 1872 -64 1906
rect -130 1838 -64 1872
rect -130 1804 -114 1838
rect -80 1804 -64 1838
rect -130 1770 -64 1804
rect -130 1736 -114 1770
rect -80 1736 -64 1770
rect -130 1702 -64 1736
rect -130 1668 -114 1702
rect -80 1668 -64 1702
rect -130 1634 -64 1668
rect -130 1600 -114 1634
rect -80 1600 -64 1634
rect -130 1566 -64 1600
rect -130 1532 -114 1566
rect -80 1532 -64 1566
rect 387 1677 453 1693
rect 387 1643 403 1677
rect 437 1643 453 1677
rect 387 1609 453 1643
rect 387 1575 403 1609
rect 437 1575 453 1609
rect 387 1559 453 1575
rect -130 1498 -64 1532
rect -130 1464 -114 1498
rect -80 1464 -64 1498
rect -130 1430 -64 1464
rect -130 1396 -114 1430
rect -80 1396 -64 1430
rect -130 1362 -64 1396
rect 387 1487 453 1503
rect 387 1453 403 1487
rect 437 1453 453 1487
rect 387 1419 453 1453
rect 387 1385 403 1419
rect 437 1385 453 1419
rect 387 1369 453 1385
rect 767 1662 839 1678
rect 767 1628 783 1662
rect 817 1628 839 1662
rect 767 1594 839 1628
rect 767 1560 783 1594
rect 817 1560 839 1594
rect 767 1544 839 1560
rect 699 1485 839 1501
rect 699 1451 715 1485
rect 749 1451 783 1485
rect 817 1451 839 1485
rect 699 1435 839 1451
rect -130 1328 -114 1362
rect -80 1328 -64 1362
rect -130 1294 -64 1328
rect -130 1260 -114 1294
rect -80 1260 -64 1294
rect -130 1226 -64 1260
rect -130 1192 -114 1226
rect -80 1192 -64 1226
rect -130 1158 -64 1192
rect 387 1311 453 1327
rect 387 1277 403 1311
rect 437 1277 453 1311
rect 387 1227 453 1277
rect 387 1193 403 1227
rect 437 1193 453 1227
rect 387 1177 453 1193
rect -130 1124 -114 1158
rect -80 1124 -64 1158
rect -130 1090 -64 1124
rect -130 1056 -114 1090
rect -80 1056 -64 1090
rect -130 1022 -64 1056
rect -130 988 -114 1022
rect -80 988 -64 1022
rect -130 954 -64 988
rect -130 920 -114 954
rect -80 920 -64 954
rect -130 886 -64 920
rect -130 852 -114 886
rect -80 852 -64 886
rect -130 818 -64 852
rect 387 1055 453 1071
rect 387 1021 403 1055
rect 437 1021 453 1055
rect 387 978 453 1021
rect 387 944 403 978
rect 437 944 453 978
rect 387 901 453 944
rect 387 867 403 901
rect 437 867 453 901
rect 387 851 453 867
rect -130 784 -114 818
rect -80 784 -64 818
rect -130 750 -64 784
rect -130 716 -114 750
rect -80 716 -64 750
rect -130 682 -64 716
rect -130 648 -114 682
rect -80 648 -64 682
rect -130 614 -64 648
rect -130 580 -114 614
rect -80 580 -64 614
rect -130 546 -64 580
rect -130 512 -114 546
rect -80 512 -64 546
rect -130 478 -64 512
rect -130 444 -114 478
rect -80 444 -64 478
rect -130 410 -64 444
rect -130 376 -114 410
rect -80 376 -64 410
rect -130 337 -64 376
rect 387 779 453 795
rect 387 745 403 779
rect 437 745 453 779
rect 387 707 453 745
rect 387 673 403 707
rect 437 673 453 707
rect 387 635 453 673
rect 387 601 403 635
rect 437 601 453 635
rect 387 563 453 601
rect 387 529 403 563
rect 437 529 453 563
rect 387 491 453 529
rect 387 457 403 491
rect 437 457 453 491
rect 387 420 453 457
rect 387 386 403 420
rect 437 386 453 420
rect 387 349 453 386
rect 387 315 403 349
rect 437 315 453 349
rect 387 299 453 315
rect 767 1377 839 1393
rect 767 1343 783 1377
rect 817 1343 839 1377
rect 767 1287 839 1343
rect 767 1253 783 1287
rect 817 1253 839 1287
rect 767 1237 839 1253
rect 767 1055 839 1071
rect 767 1021 783 1055
rect 817 1021 839 1055
rect 767 978 839 1021
rect 767 944 783 978
rect 817 944 839 978
rect 767 901 839 944
rect 767 867 783 901
rect 817 867 839 901
rect 767 851 839 867
rect 767 779 839 795
rect 767 745 783 779
rect 817 745 839 779
rect 767 707 839 745
rect 767 673 783 707
rect 817 673 839 707
rect 767 635 839 673
rect 767 601 783 635
rect 817 601 839 635
rect 767 563 839 601
rect 767 529 783 563
rect 817 529 839 563
rect 767 491 839 529
rect 767 457 783 491
rect 817 457 839 491
rect 767 420 839 457
rect 767 386 783 420
rect 817 386 839 420
rect 767 349 839 386
rect 767 315 783 349
rect 817 315 839 349
rect 767 299 839 315
<< polycont >>
rect 1203 7731 1237 7765
rect 1203 7636 1237 7670
rect 1203 7541 1237 7575
rect 2021 7731 2055 7765
rect 2021 7658 2055 7692
rect 2021 7585 2055 7619
rect 2021 7512 2055 7546
rect 1203 7419 1237 7453
rect 1203 7324 1237 7358
rect 1203 7229 1237 7263
rect 2021 7439 2055 7473
rect 2021 7366 2055 7400
rect 2021 7293 2055 7327
rect 2021 7221 2055 7255
rect 2021 7149 2055 7183
rect 2751 7731 2785 7765
rect 2751 7658 2785 7692
rect 2751 7585 2785 7619
rect 2751 7512 2785 7546
rect 2751 7439 2785 7473
rect 2751 7366 2785 7400
rect 2751 7293 2785 7327
rect 2751 7221 2785 7255
rect 2751 7149 2785 7183
rect 1083 6997 1117 7031
rect 1083 6903 1117 6937
rect 2021 7027 2055 7061
rect 2021 6950 2055 6984
rect 403 6665 437 6699
rect 403 6570 437 6604
rect 403 6475 437 6509
rect 2021 6873 2055 6907
rect 1148 6781 1182 6815
rect 2021 6797 2055 6831
rect 2751 7027 2785 7061
rect 2751 6950 2785 6984
rect 2751 6873 2785 6907
rect 2751 6797 2785 6831
rect 1148 6687 1182 6721
rect 3101 7731 3135 7765
rect 3101 7659 3135 7693
rect 3101 7587 3135 7621
rect 3101 7514 3135 7548
rect 3101 7441 3135 7475
rect 3101 7368 3135 7402
rect 3101 7295 3135 7329
rect 3101 7222 3135 7256
rect 3101 7149 3135 7183
rect 3101 7027 3135 7061
rect 3101 6950 3135 6984
rect 3101 6873 3135 6907
rect 3101 6797 3135 6831
rect 403 6243 437 6277
rect 403 6149 437 6183
rect 403 6027 437 6061
rect 403 5933 437 5967
rect 403 5701 437 5735
rect 403 5623 437 5657
rect 403 5545 437 5579
rect 403 5468 437 5502
rect 403 5391 437 5425
rect 403 5269 437 5303
rect 403 5191 437 5225
rect 403 5113 437 5147
rect 403 5036 437 5070
rect 403 4959 437 4993
rect 843 5821 877 5855
rect 843 5738 877 5772
rect 843 5655 877 5689
rect 843 5571 877 5605
rect 843 5487 877 5521
rect 1313 5821 1347 5855
rect 1313 5737 1347 5771
rect 1313 5653 1347 5687
rect 1313 5570 1347 5604
rect 1313 5487 1347 5521
rect 403 4837 437 4871
rect 403 4759 437 4793
rect 403 4681 437 4715
rect 403 4604 437 4638
rect 403 4527 437 4561
rect 403 4405 437 4439
rect 403 4337 437 4371
rect -114 4287 -80 4321
rect -114 4218 -80 4252
rect -114 4149 -80 4183
rect -114 4080 -80 4114
rect -114 4011 -80 4045
rect -114 3942 -80 3976
rect 403 4039 437 4073
rect 403 3962 437 3996
rect -114 3873 -80 3907
rect -114 3804 -80 3838
rect -114 3735 -80 3769
rect -114 3666 -80 3700
rect 403 3783 437 3817
rect 403 3672 437 3706
rect -114 3597 -80 3631
rect -114 3528 -80 3562
rect -114 3459 -80 3493
rect -114 3390 -80 3424
rect -114 3321 -80 3355
rect -114 3252 -80 3286
rect 403 3417 437 3451
rect 403 3283 437 3317
rect -114 3183 -80 3217
rect -114 3114 -80 3148
rect -114 3045 -80 3079
rect 403 3161 437 3195
rect 403 3050 437 3084
rect -114 2976 -80 3010
rect -114 2907 -80 2941
rect -114 2838 -80 2872
rect -114 2769 -80 2803
rect -114 2700 -80 2734
rect -114 2631 -80 2665
rect 403 2795 437 2829
rect 403 2661 437 2695
rect -114 2562 -80 2596
rect -114 2493 -80 2527
rect -114 2424 -80 2458
rect 403 2539 437 2573
rect 403 2405 437 2439
rect -114 2355 -80 2389
rect -114 2286 -80 2320
rect -114 2217 -80 2251
rect 783 4621 817 4655
rect 783 4527 817 4561
rect 783 4405 817 4439
rect 783 4337 817 4371
rect 783 4039 817 4073
rect 783 3905 817 3939
rect 783 3783 817 3817
rect 783 3672 817 3706
rect 783 3417 817 3451
rect 783 3283 817 3317
rect 783 3161 817 3195
rect 783 3050 817 3084
rect 783 2795 817 2829
rect 783 2661 817 2695
rect 783 2539 817 2573
rect 783 2405 817 2439
rect -114 2148 -80 2182
rect -114 2079 -80 2113
rect -114 2010 -80 2044
rect -114 1941 -80 1975
rect -114 1872 -80 1906
rect -114 1804 -80 1838
rect -114 1736 -80 1770
rect -114 1668 -80 1702
rect -114 1600 -80 1634
rect -114 1532 -80 1566
rect 403 1643 437 1677
rect 403 1575 437 1609
rect -114 1464 -80 1498
rect -114 1396 -80 1430
rect 403 1453 437 1487
rect 403 1385 437 1419
rect 783 1628 817 1662
rect 783 1560 817 1594
rect 715 1451 749 1485
rect 783 1451 817 1485
rect -114 1328 -80 1362
rect -114 1260 -80 1294
rect -114 1192 -80 1226
rect 403 1277 437 1311
rect 403 1193 437 1227
rect -114 1124 -80 1158
rect -114 1056 -80 1090
rect -114 988 -80 1022
rect -114 920 -80 954
rect -114 852 -80 886
rect 403 1021 437 1055
rect 403 944 437 978
rect 403 867 437 901
rect -114 784 -80 818
rect -114 716 -80 750
rect -114 648 -80 682
rect -114 580 -80 614
rect -114 512 -80 546
rect -114 444 -80 478
rect -114 376 -80 410
rect 403 745 437 779
rect 403 673 437 707
rect 403 601 437 635
rect 403 529 437 563
rect 403 457 437 491
rect 403 386 437 420
rect 403 315 437 349
rect 783 1343 817 1377
rect 783 1253 817 1287
rect 783 1021 817 1055
rect 783 944 817 978
rect 783 867 817 901
rect 783 745 817 779
rect 783 673 817 707
rect 783 601 817 635
rect 783 529 817 563
rect 783 457 817 491
rect 783 386 817 420
rect 783 315 817 349
<< locali >>
rect 493 8052 527 8056
rect 493 7983 527 8018
rect 493 7914 527 7941
rect 493 7845 527 7880
rect 493 7776 527 7811
rect 493 7707 527 7742
rect 493 7638 527 7673
rect 493 7569 527 7604
rect 493 7500 527 7535
rect 493 7431 527 7450
rect 493 7363 527 7378
rect 493 7295 527 7329
rect 493 7227 527 7261
rect 493 7169 527 7193
rect 741 7888 765 7922
rect 799 7888 836 7922
rect 885 7888 907 7922
rect 957 7888 977 7922
rect 1029 7888 1047 7922
rect 1101 7888 1117 7922
rect 1173 7888 1187 7922
rect 1245 7888 1257 7922
rect 1317 7888 1327 7922
rect 1389 7888 1397 7922
rect 1461 7888 1467 7922
rect 1533 7888 1537 7922
rect 1605 7888 1607 7922
rect 1641 7888 1643 7922
rect 1711 7888 1715 7922
rect 1781 7888 1787 7922
rect 1851 7888 1859 7922
rect 1921 7888 1931 7922
rect 1991 7888 2003 7922
rect 2061 7888 2075 7922
rect 2131 7888 2147 7922
rect 2201 7888 2219 7922
rect 2271 7888 2291 7922
rect 2341 7888 2363 7922
rect 2411 7888 2435 7922
rect 2481 7888 2507 7922
rect 2551 7888 2579 7922
rect 2621 7888 2651 7922
rect 2691 7888 2723 7922
rect 2761 7888 2795 7922
rect 2829 7888 2867 7922
rect 741 7884 775 7888
rect 741 7809 775 7850
rect 1101 7792 1169 7826
rect 741 7734 775 7758
rect 741 7660 775 7688
rect 741 7586 775 7618
rect 741 7512 775 7548
rect 1135 7514 1169 7792
rect 2833 7818 2867 7854
rect 1203 7765 1237 7781
rect 2021 7765 2055 7781
rect 2751 7765 2785 7781
rect 1237 7710 1276 7744
rect 2055 7710 2094 7744
rect 2705 7710 2744 7744
rect 2778 7710 2785 7731
rect 1203 7670 1237 7710
rect 1203 7575 1237 7636
rect 1203 7525 1237 7541
rect 2021 7692 2055 7710
rect 2021 7619 2055 7658
rect 2021 7546 2055 7585
rect 1101 7480 1169 7514
rect 741 7442 775 7478
rect 741 7372 775 7404
rect 741 7302 775 7338
rect 741 7232 775 7244
rect 1135 7202 1169 7480
rect 2021 7473 2055 7512
rect 1203 7453 1237 7469
rect 1203 7375 1237 7419
rect 2021 7400 2055 7439
rect 1237 7341 1276 7375
rect 1203 7263 1237 7324
rect 1203 7213 1237 7229
rect 2021 7327 2055 7366
rect 2021 7255 2055 7293
rect 741 7162 775 7198
rect 1101 7168 1169 7202
rect 2021 7183 2055 7221
rect 2021 7133 2055 7149
rect 2751 7692 2785 7710
rect 2751 7619 2785 7658
rect 2751 7546 2785 7585
rect 2751 7473 2785 7512
rect 2751 7400 2785 7439
rect 2751 7327 2785 7366
rect 2751 7255 2785 7293
rect 2751 7183 2785 7221
rect 2751 7133 2785 7149
rect 2833 7748 2867 7771
rect 2833 7678 2867 7695
rect 2833 7608 2867 7619
rect 2833 7538 2867 7574
rect 2833 7468 2867 7504
rect 3019 7908 3057 7942
rect 3091 7908 3133 7942
rect 3177 7908 3209 7942
rect 3245 7908 3279 7942
rect 3319 7908 3347 7942
rect 3395 7908 3415 7942
rect 3471 7908 3483 7942
rect 3547 7908 3551 7942
rect 3585 7908 3589 7942
rect 3653 7908 3665 7942
rect 3721 7908 3741 7942
rect 3789 7908 3823 7942
rect 3019 7840 3053 7874
rect 3857 7904 3891 7942
rect 3857 7844 3891 7870
rect 3019 7772 3053 7773
rect 3019 7722 3053 7738
rect 3019 7637 3053 7670
rect 3019 7568 3053 7602
rect 3019 7500 3053 7534
rect 2833 7399 2867 7434
rect 2975 7432 3013 7466
rect 3047 7432 3053 7466
rect 2833 7330 2867 7365
rect 2833 7295 2867 7296
rect 2833 7202 2867 7227
rect 741 7092 775 7128
rect 2833 7123 2867 7158
rect 741 7022 775 7058
rect 2021 7061 2055 7077
rect 741 6952 775 6988
rect 741 6882 775 6910
rect 53 6852 123 6876
rect 87 6842 123 6852
rect 157 6842 189 6876
rect 237 6842 275 6876
rect 316 6842 361 6876
rect 395 6842 447 6876
rect 481 6842 519 6876
rect 53 6782 87 6804
rect 53 6712 87 6729
rect 485 6773 519 6808
rect 53 6642 87 6678
rect 53 6607 87 6608
rect 53 6572 87 6573
rect 53 6527 87 6538
rect 53 6447 87 6468
rect 403 6713 437 6715
rect 403 6641 437 6665
rect 403 6604 437 6607
rect 403 6509 437 6570
rect 403 6459 437 6475
rect 485 6704 519 6739
rect 485 6635 519 6670
rect 485 6566 519 6601
rect 485 6497 519 6532
rect 741 6811 775 6828
rect 741 6740 775 6777
rect 741 6669 775 6706
rect 1067 7031 1117 7047
rect 1067 6997 1083 7031
rect 1067 6937 1117 6997
rect 1067 6903 1083 6937
rect 1067 6887 1117 6903
rect 2021 7020 2055 7027
rect 2751 7061 2785 7065
rect 2751 7026 2785 7027
rect 2055 6986 2094 7020
rect 2021 6984 2055 6986
rect 2021 6907 2055 6950
rect 1067 6660 1101 6887
rect 1148 6815 1182 6835
rect 2021 6831 2055 6873
rect 2021 6781 2055 6797
rect 2751 6984 2785 6992
rect 2751 6907 2785 6950
rect 2751 6831 2785 6873
rect 2751 6781 2785 6797
rect 2833 7054 2867 7074
rect 2833 6985 2867 7020
rect 2833 6916 2867 6951
rect 2833 6866 2867 6882
rect 1148 6721 1182 6763
rect 1148 6671 1182 6687
rect 2833 6778 2867 6813
rect 741 6598 775 6635
rect 1033 6626 1101 6660
rect 1573 6640 1679 6674
rect 1713 6640 1749 6674
rect 1783 6640 1819 6674
rect 1853 6640 1889 6674
rect 1923 6640 1959 6674
rect 1993 6640 2029 6674
rect 2063 6640 2099 6674
rect 2133 6640 2169 6674
rect 2203 6640 2239 6674
rect 2273 6640 2309 6674
rect 2343 6640 2379 6674
rect 2413 6640 2449 6674
rect 2483 6640 2519 6674
rect 2553 6640 2589 6674
rect 2623 6640 2659 6674
rect 2693 6640 2729 6674
rect 2763 6640 2799 6674
rect 2833 6640 2867 6739
rect 1573 6637 2867 6640
rect 1573 6603 1612 6637
rect 1646 6603 1688 6637
rect 1722 6603 1764 6637
rect 1798 6603 1840 6637
rect 1874 6603 1916 6637
rect 1950 6603 1992 6637
rect 2026 6603 2068 6637
rect 2102 6603 2144 6637
rect 2178 6603 2220 6637
rect 2254 6603 2296 6637
rect 2330 6603 2372 6637
rect 2406 6603 2448 6637
rect 2482 6603 2525 6637
rect 2559 6603 2602 6637
rect 2636 6603 2679 6637
rect 2713 6603 2756 6637
rect 2790 6603 2833 6637
rect 3019 7364 3053 7398
rect 3019 7296 3053 7330
rect 3019 7228 3053 7261
rect 3019 7160 3053 7177
rect 3101 7765 3135 7781
rect 3101 7693 3135 7731
rect 3101 7621 3135 7659
rect 3101 7551 3135 7587
rect 3857 7776 3891 7794
rect 3857 7708 3891 7718
rect 3857 7640 3891 7642
rect 3857 7600 3891 7606
rect 3101 7548 3111 7551
rect 3145 7517 3184 7551
rect 3857 7524 3891 7538
rect 3101 7475 3135 7514
rect 3101 7402 3135 7441
rect 3101 7329 3135 7368
rect 3101 7256 3135 7295
rect 3101 7183 3135 7222
rect 3101 7133 3135 7149
rect 3857 7448 3891 7470
rect 3857 7373 3891 7402
rect 3857 7300 3891 7334
rect 3857 7232 3891 7264
rect 3857 7164 3891 7189
rect 3857 7096 3891 7114
rect 3019 7024 3053 7058
rect 3019 6956 3053 6990
rect 3019 6888 3053 6922
rect 3019 6820 3053 6832
rect 3019 6773 3053 6786
rect 3101 7061 3135 7077
rect 3101 7020 3135 7027
rect 3857 7028 3891 7039
rect 3135 6986 3174 7020
rect 3101 6984 3135 6986
rect 3101 6907 3135 6950
rect 3101 6831 3135 6873
rect 3101 6781 3135 6797
rect 3857 6960 3891 6964
rect 3857 6923 3891 6926
rect 3857 6848 3891 6858
rect 3019 6637 3053 6718
rect 3857 6773 3891 6790
rect 3857 6688 3891 6722
rect 3087 6637 3121 6654
rect 3155 6637 3189 6654
rect 3223 6637 3257 6654
rect 3019 6620 3036 6637
rect 3087 6620 3109 6637
rect 3155 6620 3182 6637
rect 3223 6620 3255 6637
rect 3291 6620 3325 6654
rect 3359 6637 3393 6654
rect 3427 6637 3461 6654
rect 3495 6637 3529 6654
rect 3563 6637 3597 6654
rect 3631 6637 3665 6654
rect 3699 6637 3733 6654
rect 3767 6637 3891 6654
rect 3362 6620 3393 6637
rect 3435 6620 3461 6637
rect 3508 6620 3529 6637
rect 3581 6620 3597 6637
rect 3654 6620 3665 6637
rect 3727 6620 3733 6637
rect 3070 6603 3109 6620
rect 3143 6603 3182 6620
rect 3216 6603 3255 6620
rect 3289 6603 3328 6620
rect 3362 6603 3401 6620
rect 3435 6603 3474 6620
rect 3508 6603 3547 6620
rect 3581 6603 3620 6620
rect 3654 6603 3693 6620
rect 3727 6603 3766 6620
rect 3800 6603 3840 6637
rect 3874 6620 3891 6637
rect 1573 6564 1607 6603
rect 741 6530 769 6564
rect 803 6530 843 6564
rect 879 6530 914 6564
rect 950 6530 983 6564
rect 1023 6530 1052 6564
rect 1096 6530 1121 6564
rect 1169 6530 1190 6564
rect 1242 6530 1259 6564
rect 1315 6530 1329 6564
rect 1388 6530 1399 6564
rect 1461 6530 1469 6564
rect 1534 6530 1539 6564
rect 741 6523 1607 6530
rect 53 6368 87 6398
rect 53 6292 87 6328
rect 485 6428 519 6463
rect 485 6359 519 6394
rect 53 6222 87 6255
rect 53 6152 87 6176
rect 403 6281 437 6293
rect 403 6209 437 6243
rect 403 6133 437 6149
rect 485 6290 519 6325
rect 485 6221 519 6256
rect 485 6155 519 6187
rect 53 6082 87 6097
rect 485 6083 519 6118
rect 403 6061 437 6077
rect 53 6012 87 6018
rect 343 6011 381 6045
rect 415 6011 437 6027
rect 53 5942 87 5978
rect 403 5967 437 6011
rect 403 5917 437 5933
rect 485 6014 519 6049
rect 485 5945 519 5980
rect 53 5900 87 5908
rect 53 5822 87 5838
rect 53 5744 87 5768
rect 485 5876 519 5911
rect 485 5826 519 5842
rect 53 5667 87 5698
rect 53 5592 87 5628
rect 53 5522 87 5556
rect 53 5452 87 5479
rect 53 5382 87 5402
rect 403 5735 437 5751
rect 403 5657 437 5701
rect 403 5579 437 5623
rect 403 5502 437 5545
rect 403 5425 437 5468
rect 403 5375 437 5391
rect 485 5749 519 5773
rect 485 5671 519 5704
rect 485 5600 519 5635
rect 485 5531 519 5566
rect 485 5462 519 5465
rect 485 5414 519 5428
rect 53 5312 87 5325
rect 485 5329 519 5359
rect 53 5242 87 5248
rect 53 5172 87 5208
rect 403 5303 437 5319
rect 403 5225 437 5269
rect 53 5102 87 5138
rect 263 5114 301 5148
rect 403 5147 437 5191
rect 403 5074 437 5113
rect 53 5032 87 5068
rect 365 5040 403 5074
rect 53 4962 87 4998
rect 403 4993 437 5036
rect 403 4943 437 4959
rect 485 5255 519 5290
rect 761 6004 816 6028
rect 795 5994 816 6004
rect 850 5994 891 6028
rect 927 5994 968 6028
rect 1004 5994 1045 6028
rect 1081 5994 1122 6028
rect 1158 5994 1199 6028
rect 1235 5994 1276 6028
rect 1311 5994 1429 6028
rect 795 5970 812 5994
rect 761 5952 812 5970
rect 761 5935 795 5952
rect 761 5866 795 5901
rect 921 5919 1005 5928
rect 921 5885 933 5919
rect 967 5885 1005 5919
rect 1039 5885 1059 5928
rect 921 5882 1059 5885
rect 1125 5919 1209 5928
rect 1125 5885 1137 5919
rect 1171 5885 1209 5919
rect 1243 5885 1263 5928
rect 1125 5882 1263 5885
rect 1395 5926 1429 5956
rect 761 5797 795 5832
rect 761 5741 795 5763
rect 761 5660 795 5694
rect 761 5590 795 5625
rect 761 5521 795 5556
rect 761 5452 795 5487
rect 843 5855 877 5871
rect 843 5772 877 5821
rect 843 5689 877 5738
rect 843 5605 877 5655
rect 1309 5855 1347 5871
rect 1309 5821 1313 5855
rect 1309 5771 1347 5821
rect 1309 5737 1313 5771
rect 1309 5687 1347 5737
rect 1309 5653 1313 5687
rect 1309 5604 1347 5653
rect 1125 5580 1263 5586
rect 843 5546 854 5571
rect 888 5546 926 5580
rect 1125 5546 1137 5580
rect 1171 5546 1209 5580
rect 1243 5546 1263 5580
rect 843 5521 877 5546
rect 843 5471 877 5487
rect 761 5382 795 5418
rect 921 5469 1059 5476
rect 921 5435 933 5469
rect 967 5435 1005 5469
rect 921 5414 1005 5435
rect 1039 5414 1059 5469
rect 1125 5448 1263 5546
rect 1125 5414 1209 5448
rect 1243 5414 1263 5448
rect 1309 5570 1313 5604
rect 1309 5521 1347 5570
rect 1309 5509 1313 5521
rect 1343 5475 1347 5487
rect 1309 5437 1347 5475
rect 1343 5403 1347 5437
rect 1395 5858 1429 5876
rect 1395 5790 1429 5796
rect 1395 5751 1429 5756
rect 1395 5672 1429 5688
rect 1395 5593 1429 5620
rect 1395 5518 1429 5552
rect 1395 5450 1429 5480
rect 761 5314 867 5348
rect 901 5314 937 5348
rect 971 5314 1007 5348
rect 1041 5314 1077 5348
rect 1111 5314 1148 5348
rect 1182 5314 1219 5348
rect 1253 5314 1290 5348
rect 1324 5314 1361 5348
rect 1395 5314 1429 5401
rect 761 5311 1429 5314
rect 795 5277 835 5311
rect 869 5277 909 5311
rect 943 5277 983 5311
rect 1017 5277 1057 5311
rect 1091 5277 1132 5311
rect 1166 5277 1207 5311
rect 1241 5277 1282 5311
rect 1316 5277 1357 5311
rect 1391 5277 1429 5311
rect 485 5186 519 5209
rect 485 5117 519 5152
rect 485 5048 519 5083
rect 485 4979 519 5014
rect 53 4892 87 4897
rect 485 4910 519 4945
rect 53 4822 87 4825
rect 53 4752 87 4788
rect -396 4576 -314 4745
rect 53 4681 87 4718
rect 53 4610 87 4647
rect 403 4880 437 4887
rect 403 4808 437 4837
rect 403 4715 437 4759
rect 403 4642 437 4681
rect 365 4608 403 4642
rect -396 4542 -264 4576
rect -230 4542 -193 4576
rect -159 4542 -123 4576
rect -89 4542 -53 4576
rect -19 4542 87 4576
rect 403 4561 437 4604
rect -396 4006 -314 4542
rect 191 4512 255 4546
rect 157 4507 289 4512
rect 403 4511 437 4527
rect 485 4841 519 4876
rect 485 4772 519 4807
rect 485 4703 519 4738
rect 485 4634 519 4669
rect 485 4565 519 4600
rect 157 4500 359 4507
rect 289 4473 359 4500
rect 485 4496 519 4523
rect -244 4450 -194 4454
rect -244 4416 -228 4450
rect -194 4416 -160 4420
rect -244 4382 -160 4416
rect -244 4348 -194 4382
rect -26 4416 0 4420
rect 34 4416 50 4450
rect 403 4439 437 4455
rect -26 4382 50 4416
rect 8 4348 50 4382
rect 157 4372 168 4406
rect 202 4372 240 4406
rect 274 4372 275 4406
rect -396 3972 -348 4006
rect -396 3864 -314 3972
rect -396 3830 -348 3864
rect -396 3493 -314 3830
rect -396 3459 -348 3493
rect -396 3423 -314 3459
rect -396 3364 -348 3423
rect -396 3353 -314 3364
rect -396 3319 -348 3353
rect -396 3305 -314 3319
rect -396 3249 -348 3305
rect -396 3213 -314 3249
rect -396 3178 -348 3213
rect -396 3143 -314 3178
rect -396 3084 -348 3143
rect -396 3073 -314 3084
rect -396 3039 -348 3073
rect -396 3003 -314 3039
rect -396 2969 -348 3003
rect -396 2933 -314 2969
rect -396 2899 -348 2933
rect -396 2863 -314 2899
rect -396 2829 -348 2863
rect -396 2814 -314 2829
rect -396 2759 -348 2814
rect -396 2737 -314 2759
rect -396 2689 -348 2737
rect -396 2653 -314 2689
rect -396 2619 -348 2653
rect -396 2583 -314 2619
rect -396 2549 -348 2583
rect -396 2513 -314 2549
rect -396 2479 -348 2513
rect -396 2443 -314 2479
rect -396 2409 -348 2443
rect -396 2373 -314 2409
rect -396 2339 -348 2373
rect -396 2303 -314 2339
rect -396 2269 -348 2303
rect -396 2233 -314 2269
rect -396 2199 -348 2233
rect -396 2163 -314 2199
rect -396 2129 -348 2163
rect -396 2093 -314 2129
rect -396 2059 -348 2093
rect -396 2023 -314 2059
rect -396 1989 -348 2023
rect -396 1953 -314 1989
rect -396 1919 -348 1953
rect -396 1895 -314 1919
rect -396 1849 -348 1895
rect -396 1819 -314 1849
rect -396 1779 -348 1819
rect -396 1743 -314 1779
rect -396 1708 -348 1743
rect -396 1673 -314 1708
rect -396 1631 -348 1673
rect -396 1603 -314 1631
rect -396 1569 -348 1603
rect -396 1533 -314 1569
rect -396 1499 -348 1533
rect -396 1495 -314 1499
rect -396 1429 -348 1495
rect -396 1415 -314 1429
rect -396 1359 -348 1415
rect -396 1323 -314 1359
rect -396 1289 -348 1323
rect -396 1253 -314 1289
rect -396 1219 -348 1253
rect -396 1184 -314 1219
rect -396 1150 -348 1184
rect -396 1115 -314 1150
rect -396 1065 -348 1115
rect -396 1046 -314 1065
rect -396 984 -348 1046
rect -396 384 -314 984
rect -396 350 -348 384
rect -114 4325 -80 4337
rect -114 4253 -80 4287
rect 157 4244 275 4372
rect 354 4405 403 4427
rect 354 4393 437 4405
rect 320 4371 437 4393
rect 320 4355 403 4371
rect 354 4337 403 4355
rect 354 4321 437 4337
rect 485 4427 519 4462
rect 485 4358 519 4393
rect 485 4289 519 4314
rect 403 4286 437 4287
rect -114 4183 -80 4218
rect -114 4114 -80 4149
rect 403 4214 437 4252
rect 230 4100 294 4134
rect -114 4045 -80 4080
rect -114 3976 -80 4011
rect 403 4073 437 4180
rect 403 3996 437 4039
rect 403 3946 437 3962
rect 485 4220 519 4255
rect 485 4151 519 4186
rect 485 4082 519 4117
rect 485 4046 519 4048
rect 485 3960 519 3979
rect -114 3907 -80 3942
rect -114 3838 -80 3873
rect 485 3875 519 3910
rect -114 3769 -80 3804
rect -114 3700 -80 3735
rect -114 3631 -80 3666
rect 403 3735 437 3783
rect 403 3656 437 3672
rect 485 3806 519 3840
rect 485 3737 519 3754
rect 485 3702 519 3703
rect -114 3562 -80 3597
rect 359 3588 437 3622
rect -114 3493 -80 3528
rect -114 3424 -80 3459
rect -114 3355 -80 3390
rect -114 3286 -80 3321
rect 403 3451 437 3588
rect 403 3317 437 3417
rect 403 3267 437 3283
rect 485 3599 519 3634
rect 485 3530 519 3565
rect 485 3461 519 3496
rect 485 3420 519 3427
rect 485 3335 519 3358
rect -114 3217 -80 3252
rect 485 3254 519 3289
rect -114 3148 -80 3183
rect -114 3079 -80 3114
rect -114 3010 -80 3045
rect 403 3113 437 3161
rect 403 3034 437 3050
rect 485 3185 519 3216
rect 485 3116 519 3131
rect 485 3080 519 3082
rect -114 2941 -80 2976
rect 359 2966 437 3000
rect -114 2872 -80 2907
rect -114 2803 -80 2838
rect -114 2734 -80 2769
rect -114 2665 -80 2700
rect 403 2829 437 2966
rect 403 2695 437 2795
rect 403 2645 437 2661
rect 485 2978 519 3013
rect 485 2909 519 2944
rect 485 2840 519 2875
rect 485 2795 519 2806
rect 485 2711 519 2738
rect -114 2596 -80 2631
rect 485 2636 519 2670
rect -114 2527 -80 2562
rect -114 2458 -80 2493
rect -114 2389 -80 2424
rect 403 2491 437 2539
rect 403 2439 437 2457
rect 403 2389 437 2405
rect 485 2568 519 2593
rect 485 2500 519 2509
rect 485 2458 519 2466
rect -114 2320 -80 2355
rect -114 2251 -80 2286
rect 485 2364 519 2398
rect 485 2262 519 2330
rect 161 2228 185 2262
rect 219 2228 237 2262
rect 271 2228 273 2262
rect 307 2228 315 2262
rect 349 2228 362 2262
rect 428 2228 451 2262
rect 507 2228 519 2262
rect 701 4788 739 4812
rect 735 4778 739 4788
rect 773 4778 822 4812
rect 865 4778 905 4812
rect 946 4778 988 4812
rect 1027 4778 1153 4812
rect 701 4720 735 4754
rect 701 4652 735 4686
rect 1119 4709 1153 4740
rect 701 4584 735 4618
rect 701 4516 735 4550
rect 783 4655 817 4671
rect 817 4608 855 4642
rect 1119 4640 1153 4667
rect 783 4561 817 4608
rect 783 4511 817 4527
rect 1119 4571 1153 4595
rect 701 4448 735 4482
rect 1119 4502 1153 4523
rect 701 4380 735 4414
rect 701 4312 735 4346
rect 783 4439 817 4455
rect 1119 4433 1153 4451
rect 783 4389 803 4405
rect 837 4389 901 4423
rect 783 4371 817 4389
rect 783 4321 817 4337
rect 1119 4364 1153 4379
rect 1119 4295 1153 4307
rect 701 4244 735 4278
rect 701 4176 735 4210
rect 701 4108 735 4142
rect 701 4040 735 4074
rect 701 3972 735 4004
rect 701 3903 735 3922
rect 783 4286 817 4287
rect 783 4214 817 4252
rect 967 4210 1031 4244
rect 1119 4226 1153 4235
rect 783 4073 817 4180
rect 783 3939 817 4039
rect 783 3889 817 3905
rect 1119 4157 1153 4163
rect 1119 4088 1153 4091
rect 1119 4053 1153 4054
rect 1119 3981 1153 3985
rect 1119 3909 1153 3916
rect 701 3834 735 3840
rect 1119 3837 1153 3847
rect 701 3792 735 3800
rect 701 3711 735 3731
rect 701 3627 735 3662
rect 783 3735 817 3783
rect 783 3656 817 3672
rect 1119 3765 1153 3778
rect 1119 3693 1153 3710
rect 701 3558 735 3593
rect 701 3489 735 3524
rect 701 3423 735 3455
rect 701 3351 735 3386
rect 701 3282 735 3306
rect 783 3588 867 3622
rect 1119 3621 1153 3642
rect 783 3451 817 3588
rect 783 3317 817 3417
rect 783 3267 817 3283
rect 1119 3549 1153 3574
rect 1119 3477 1153 3506
rect 1119 3405 1153 3438
rect 1119 3336 1153 3370
rect 1119 3268 1153 3299
rect 701 3213 735 3223
rect 701 3173 735 3179
rect 701 3089 735 3110
rect 701 3006 735 3041
rect 783 3113 817 3161
rect 783 3034 817 3050
rect 1119 3200 1153 3227
rect 1119 3132 1153 3155
rect 1119 3064 1153 3083
rect 701 2937 735 2972
rect 701 2868 735 2903
rect 701 2801 735 2834
rect 701 2730 735 2765
rect 701 2661 735 2685
rect 783 2966 863 3000
rect 897 2966 937 3000
rect 971 2966 1011 3000
rect 1119 2996 1153 3011
rect 783 2829 817 2966
rect 1119 2928 1153 2939
rect 897 2856 937 2890
rect 971 2856 1011 2890
rect 1119 2860 1153 2867
rect 783 2695 817 2795
rect 783 2645 817 2661
rect 1119 2792 1153 2795
rect 1119 2724 1153 2758
rect 1119 2656 1153 2690
rect 701 2592 735 2603
rect 909 2600 962 2634
rect 996 2600 1048 2634
rect 701 2555 735 2558
rect 701 2473 735 2489
rect 701 2385 735 2420
rect 783 2573 817 2589
rect 783 2518 817 2539
rect 1119 2588 1153 2622
rect 1119 2520 1153 2554
rect 783 2484 799 2518
rect 833 2484 897 2518
rect 783 2439 817 2484
rect 783 2389 817 2405
rect 1119 2452 1153 2478
rect 1119 2384 1153 2390
rect 701 2316 735 2351
rect 863 2362 1069 2378
rect 897 2328 937 2362
rect 971 2328 1011 2362
rect 1045 2328 1069 2362
rect 701 2248 749 2282
rect 783 2248 805 2282
rect 866 2248 875 2282
rect 909 2248 915 2282
rect 979 2248 998 2282
rect 1049 2248 1081 2282
rect 1119 2248 1153 2350
rect -114 2182 -80 2217
rect -114 2113 -80 2148
rect -114 2044 -80 2079
rect -114 1975 -80 2010
rect -114 1906 -80 1941
rect -114 1838 -80 1872
rect -114 1770 -80 1804
rect 161 2110 185 2144
rect 219 2136 254 2144
rect 288 2136 323 2144
rect 219 2110 237 2136
rect 288 2110 315 2136
rect 357 2110 392 2144
rect 426 2136 461 2144
rect 495 2136 519 2144
rect 428 2110 461 2136
rect 161 2102 237 2110
rect 271 2102 315 2110
rect 349 2102 394 2110
rect 428 2102 473 2110
rect 507 2102 519 2136
rect 161 2076 519 2102
rect 161 2042 185 2076
rect 219 2042 254 2076
rect 288 2042 323 2076
rect 357 2042 392 2076
rect 426 2042 461 2076
rect 495 2042 519 2076
rect 161 2008 519 2042
rect 161 1974 185 2008
rect 219 1974 254 2008
rect 288 1974 323 2008
rect 357 1974 392 2008
rect 426 1974 461 2008
rect 495 1974 519 2008
rect 161 1940 519 1974
rect 161 1906 185 1940
rect 219 1906 254 1940
rect 288 1906 323 1940
rect 357 1906 392 1940
rect 426 1906 461 1940
rect 495 1906 519 1940
rect 161 1872 519 1906
rect 161 1867 185 1872
rect 219 1867 254 1872
rect 161 1833 173 1867
rect 219 1838 248 1867
rect 288 1838 323 1872
rect 357 1838 392 1872
rect 426 1867 461 1872
rect 495 1867 519 1872
rect 432 1838 461 1867
rect 207 1833 248 1838
rect 282 1833 323 1838
rect 357 1833 398 1838
rect 432 1833 473 1838
rect 507 1833 519 1867
rect 161 1804 519 1833
rect 161 1795 185 1804
rect 219 1795 254 1804
rect 161 1770 173 1795
rect 219 1770 248 1795
rect 288 1770 323 1804
rect 357 1770 392 1804
rect 426 1795 461 1804
rect 495 1795 519 1804
rect 432 1770 461 1795
rect 162 1761 173 1770
rect 207 1761 248 1770
rect 282 1761 323 1770
rect 357 1761 398 1770
rect 432 1761 473 1770
rect 507 1761 519 1795
rect -114 1702 -80 1736
rect -114 1634 -80 1668
rect -114 1566 -80 1600
rect 403 1637 437 1643
rect 403 1559 437 1575
rect 485 1694 519 1761
rect 485 1622 519 1660
rect -114 1498 -80 1532
rect 280 1515 318 1549
rect 485 1535 519 1588
rect 614 1740 713 1774
rect 747 1746 795 1774
rect 829 1746 877 1774
rect 911 1746 959 1774
rect 993 1746 1041 1774
rect 759 1740 795 1746
rect 614 1712 725 1740
rect 759 1712 797 1740
rect 831 1712 869 1746
rect 911 1740 940 1746
rect 993 1740 1011 1746
rect 1075 1740 1205 1774
rect 903 1712 940 1740
rect 974 1712 1011 1740
rect 1045 1736 1205 1740
rect 1045 1712 1171 1736
rect 614 1605 676 1712
rect 1153 1702 1171 1712
rect 1153 1678 1205 1702
rect 710 1644 711 1678
rect 745 1644 783 1678
rect 614 1581 735 1605
rect 614 1547 701 1581
rect 614 1523 735 1547
rect 783 1594 817 1628
rect 783 1544 817 1560
rect 1119 1652 1205 1678
rect 1119 1641 1171 1652
rect 1153 1618 1171 1641
rect 1153 1607 1205 1618
rect 1119 1570 1205 1607
rect 1153 1568 1205 1570
rect 1153 1536 1171 1568
rect 1119 1534 1171 1536
rect -114 1430 -80 1464
rect -114 1362 -80 1396
rect 403 1487 437 1503
rect 1119 1499 1205 1534
rect 437 1475 715 1485
rect 437 1453 543 1475
rect 403 1441 543 1453
rect 577 1441 615 1475
rect 649 1451 715 1475
rect 749 1451 783 1485
rect 817 1451 833 1485
rect 649 1441 833 1451
rect 403 1440 833 1441
rect 1153 1484 1205 1499
rect 1153 1465 1171 1484
rect 1119 1450 1171 1465
rect 403 1419 437 1440
rect 1119 1428 1205 1450
rect 403 1369 437 1385
rect 485 1392 519 1394
rect 485 1378 488 1392
rect -114 1294 -80 1328
rect 522 1358 560 1392
rect 701 1372 704 1394
rect 1153 1400 1205 1428
rect 1153 1394 1171 1400
rect 783 1377 817 1393
rect 157 1292 241 1298
rect 275 1292 313 1326
rect 403 1311 437 1327
rect 347 1292 359 1298
rect -114 1226 -80 1260
rect 403 1227 437 1277
rect 485 1306 519 1344
rect 485 1245 519 1272
rect 701 1303 735 1372
rect 701 1245 735 1269
rect 783 1287 817 1343
rect 1119 1366 1171 1394
rect 1119 1357 1205 1366
rect 867 1292 879 1298
rect 913 1292 951 1326
rect 985 1292 1023 1326
rect 1153 1323 1205 1357
rect 1119 1317 1205 1323
rect 1057 1292 1069 1298
rect 191 1192 229 1226
rect 263 1192 301 1226
rect 783 1211 817 1253
rect 1119 1286 1171 1317
rect 1153 1283 1171 1286
rect 1153 1252 1205 1283
rect 1119 1234 1205 1252
rect -114 1158 -80 1192
rect 403 1177 405 1193
rect 439 1177 477 1211
rect 511 1177 817 1211
rect 901 1197 939 1231
rect 973 1197 1011 1231
rect 1045 1197 1069 1231
rect 1119 1215 1171 1234
rect 1153 1200 1171 1215
rect 1119 1144 1153 1181
rect -114 1090 -80 1124
rect 485 1127 519 1143
rect 157 1098 359 1116
rect 157 1064 169 1098
rect 203 1064 241 1098
rect 275 1064 359 1098
rect -114 1022 -80 1056
rect -114 954 -80 988
rect -114 886 -80 920
rect -114 818 -80 852
rect 403 1055 437 1071
rect 485 1046 519 1089
rect 701 1104 735 1143
rect 701 1046 735 1056
rect 783 1055 817 1071
rect 911 1064 949 1098
rect 983 1064 1021 1098
rect 1055 1064 1069 1098
rect 1119 1092 1153 1110
rect 1119 1073 1171 1092
rect 403 1012 437 1021
rect 783 1012 817 1021
rect 403 978 539 1012
rect 573 978 611 1012
rect 645 978 817 1012
rect 403 901 437 944
rect 403 851 437 867
rect 485 928 519 944
rect 485 856 519 894
rect -114 750 -80 784
rect -114 682 -80 716
rect -114 614 -80 648
rect -114 546 -80 580
rect -114 478 -80 512
rect -114 410 -80 444
rect -114 360 -80 376
rect 403 787 437 795
rect 403 708 437 745
rect 403 635 437 673
rect 403 563 437 596
rect 403 491 437 518
rect 403 420 437 457
rect -396 244 -314 350
rect 403 349 437 386
rect -178 292 -172 326
rect -138 314 -100 326
rect -138 292 -109 314
rect -66 292 -28 326
rect 403 299 437 315
rect 485 784 519 818
rect 485 712 519 738
rect 485 640 519 658
rect 485 568 519 578
rect 485 533 519 534
rect 485 496 519 499
rect 485 454 519 462
rect 485 375 519 390
rect 485 296 519 318
rect -244 280 -109 292
rect -75 280 50 292
rect -244 274 50 280
rect -396 210 -348 244
rect -396 172 -314 210
rect 485 172 519 246
rect -427 138 -386 172
rect -352 138 -311 172
rect -246 138 -236 172
rect -176 138 -161 172
rect -106 138 -85 172
rect -36 138 -9 172
rect 35 138 67 172
rect 101 138 143 172
rect 177 138 219 172
rect 265 138 295 172
rect 337 138 371 172
rect 409 138 447 172
rect 481 138 519 172
rect 701 920 735 944
rect 701 858 735 886
rect 783 901 817 944
rect 783 851 817 867
rect 1153 1058 1171 1073
rect 1153 1039 1205 1058
rect 1119 1014 1205 1039
rect 1119 1002 1171 1014
rect 1153 980 1171 1002
rect 1153 968 1205 980
rect 1119 936 1205 968
rect 1119 931 1171 936
rect 1153 902 1171 931
rect 1153 897 1205 902
rect 1119 860 1205 897
rect 701 786 735 817
rect 1153 858 1205 860
rect 1153 826 1171 858
rect 1119 824 1171 826
rect 701 713 735 748
rect 701 644 735 679
rect 701 604 735 610
rect 701 529 735 541
rect 701 454 735 472
rect 701 380 735 402
rect 701 306 735 332
rect 783 779 817 795
rect 783 707 817 745
rect 783 635 817 662
rect 783 563 817 575
rect 783 522 817 529
rect 783 436 817 457
rect 783 350 817 386
rect 783 299 817 315
rect 1119 789 1205 824
rect 1153 780 1205 789
rect 1153 755 1171 780
rect 1119 746 1171 755
rect 1119 718 1205 746
rect 1153 702 1205 718
rect 1153 684 1171 702
rect 1119 668 1171 684
rect 1119 648 1205 668
rect 1153 624 1205 648
rect 1153 614 1171 624
rect 1119 590 1171 614
rect 1119 578 1205 590
rect 1153 546 1205 578
rect 1153 544 1171 546
rect 1119 512 1171 544
rect 1119 508 1205 512
rect 1153 474 1205 508
rect 1119 467 1205 474
rect 1119 438 1171 467
rect 1153 433 1171 438
rect 1153 404 1205 433
rect 1119 388 1205 404
rect 1119 368 1171 388
rect 1153 354 1171 368
rect 1153 334 1205 354
rect 1119 309 1205 334
rect 701 226 735 262
rect 1119 298 1171 309
rect 1153 275 1171 298
rect 1153 264 1205 275
rect 1119 230 1205 264
rect 1119 196 1171 230
rect 701 158 739 192
rect 773 158 805 192
rect 851 158 875 192
rect 929 158 945 192
rect 1007 158 1015 192
rect 1049 158 1051 192
rect 1119 158 1205 196
<< viali >>
rect 493 8056 527 8090
rect 493 7949 527 7975
rect 493 7941 527 7949
rect 493 7466 527 7484
rect 493 7450 527 7466
rect 493 7397 527 7412
rect 493 7378 527 7397
rect 851 7888 870 7922
rect 870 7888 885 7922
rect 923 7888 941 7922
rect 941 7888 957 7922
rect 995 7888 1011 7922
rect 1011 7888 1029 7922
rect 1067 7888 1081 7922
rect 1081 7888 1101 7922
rect 1139 7888 1151 7922
rect 1151 7888 1173 7922
rect 1211 7888 1221 7922
rect 1221 7888 1245 7922
rect 1283 7888 1291 7922
rect 1291 7888 1317 7922
rect 1355 7888 1361 7922
rect 1361 7888 1389 7922
rect 1427 7888 1431 7922
rect 1431 7888 1461 7922
rect 1499 7888 1501 7922
rect 1501 7888 1533 7922
rect 1571 7888 1605 7922
rect 1643 7888 1677 7922
rect 1715 7888 1747 7922
rect 1747 7888 1749 7922
rect 1787 7888 1817 7922
rect 1817 7888 1821 7922
rect 1859 7888 1887 7922
rect 1887 7888 1893 7922
rect 1931 7888 1957 7922
rect 1957 7888 1965 7922
rect 2003 7888 2027 7922
rect 2027 7888 2037 7922
rect 2075 7888 2097 7922
rect 2097 7888 2109 7922
rect 2147 7888 2167 7922
rect 2167 7888 2181 7922
rect 2219 7888 2237 7922
rect 2237 7888 2253 7922
rect 2291 7888 2307 7922
rect 2307 7888 2325 7922
rect 2363 7888 2377 7922
rect 2377 7888 2397 7922
rect 2435 7888 2447 7922
rect 2447 7888 2469 7922
rect 2507 7888 2517 7922
rect 2517 7888 2541 7922
rect 2579 7888 2587 7922
rect 2587 7888 2613 7922
rect 2651 7888 2657 7922
rect 2657 7888 2685 7922
rect 2723 7888 2727 7922
rect 2727 7888 2757 7922
rect 2795 7888 2829 7922
rect 741 7850 775 7884
rect 741 7792 775 7809
rect 741 7775 775 7792
rect 741 7722 775 7734
rect 741 7700 775 7722
rect 741 7652 775 7660
rect 741 7626 775 7652
rect 741 7582 775 7586
rect 741 7552 775 7582
rect 2833 7784 2867 7805
rect 1203 7731 1237 7744
rect 1203 7710 1237 7731
rect 1276 7710 1310 7744
rect 2021 7731 2055 7744
rect 2021 7710 2055 7731
rect 2094 7710 2128 7744
rect 2671 7710 2705 7744
rect 2744 7731 2751 7744
rect 2751 7731 2778 7744
rect 2744 7710 2778 7731
rect 741 7478 775 7512
rect 741 7408 775 7438
rect 741 7404 775 7408
rect 741 7268 775 7278
rect 741 7244 775 7268
rect 1203 7358 1237 7375
rect 1203 7341 1237 7358
rect 1276 7341 1310 7375
rect 2833 7771 2867 7784
rect 2833 7714 2867 7729
rect 2833 7695 2867 7714
rect 2833 7644 2867 7653
rect 2833 7619 2867 7644
rect 3057 7908 3091 7942
rect 3133 7908 3143 7942
rect 3143 7908 3167 7942
rect 3209 7908 3211 7942
rect 3211 7908 3243 7942
rect 3285 7908 3313 7942
rect 3313 7908 3319 7942
rect 3361 7908 3381 7942
rect 3381 7908 3395 7942
rect 3437 7908 3449 7942
rect 3449 7908 3471 7942
rect 3513 7908 3517 7942
rect 3517 7908 3547 7942
rect 3589 7908 3619 7942
rect 3619 7908 3623 7942
rect 3665 7908 3687 7942
rect 3687 7908 3699 7942
rect 3741 7908 3755 7942
rect 3755 7908 3775 7942
rect 3019 7806 3053 7807
rect 3019 7773 3053 7806
rect 3857 7870 3891 7904
rect 3857 7810 3891 7828
rect 3857 7794 3891 7810
rect 3019 7704 3053 7722
rect 3019 7688 3053 7704
rect 3019 7636 3053 7637
rect 3019 7603 3053 7636
rect 2941 7432 2975 7466
rect 3013 7432 3047 7466
rect 2833 7261 2867 7295
rect 2833 7192 2867 7202
rect 2833 7168 2867 7192
rect 741 6918 775 6944
rect 741 6910 775 6918
rect 189 6842 203 6876
rect 203 6842 223 6876
rect 275 6842 282 6876
rect 282 6842 309 6876
rect 361 6842 395 6876
rect 447 6842 481 6876
rect 53 6818 87 6838
rect 53 6804 87 6818
rect 53 6748 87 6763
rect 53 6729 87 6748
rect 53 6573 87 6607
rect 53 6502 87 6527
rect 53 6493 87 6502
rect 403 6699 437 6713
rect 403 6679 437 6699
rect 403 6607 437 6641
rect 741 6848 775 6862
rect 741 6828 775 6848
rect 2751 7065 2785 7099
rect 2021 6986 2055 7020
rect 2094 6986 2128 7020
rect 2751 6992 2785 7026
rect 1148 6835 1182 6869
rect 1148 6781 1182 6797
rect 2833 7089 2867 7108
rect 2833 7074 2867 7089
rect 2833 6847 2867 6866
rect 2833 6832 2867 6847
rect 1148 6763 1182 6781
rect 2833 6744 2867 6773
rect 2833 6739 2867 6744
rect 1612 6603 1646 6637
rect 1688 6603 1722 6637
rect 1764 6603 1798 6637
rect 1840 6603 1874 6637
rect 1916 6603 1950 6637
rect 1992 6603 2026 6637
rect 2068 6603 2102 6637
rect 2144 6603 2178 6637
rect 2220 6603 2254 6637
rect 2296 6603 2330 6637
rect 2372 6603 2406 6637
rect 2448 6603 2482 6637
rect 2525 6603 2559 6637
rect 2602 6603 2636 6637
rect 2679 6603 2713 6637
rect 2756 6603 2790 6637
rect 2833 6603 2867 6637
rect 3019 7262 3053 7295
rect 3019 7261 3053 7262
rect 3019 7194 3053 7211
rect 3019 7177 3053 7194
rect 3857 7742 3891 7752
rect 3857 7718 3891 7742
rect 3857 7674 3891 7676
rect 3857 7642 3891 7674
rect 3857 7572 3891 7600
rect 3857 7566 3891 7572
rect 3111 7548 3145 7551
rect 3111 7517 3135 7548
rect 3135 7517 3145 7548
rect 3184 7517 3218 7551
rect 3857 7504 3891 7524
rect 3857 7490 3891 7504
rect 3857 7436 3891 7448
rect 3857 7414 3891 7436
rect 3857 7368 3891 7373
rect 3857 7339 3891 7368
rect 3857 7266 3891 7298
rect 3857 7264 3891 7266
rect 3857 7198 3891 7223
rect 3857 7189 3891 7198
rect 3019 7092 3053 7126
rect 3857 7130 3891 7148
rect 3857 7114 3891 7130
rect 3019 6854 3053 6866
rect 3019 6832 3053 6854
rect 3857 7062 3891 7073
rect 3857 7039 3891 7062
rect 3101 6986 3135 7020
rect 3174 6986 3208 7020
rect 3857 6994 3891 6998
rect 3857 6964 3891 6994
rect 3857 6892 3891 6923
rect 3857 6889 3891 6892
rect 3857 6824 3891 6848
rect 3857 6814 3891 6824
rect 3019 6752 3053 6773
rect 3019 6739 3053 6752
rect 3857 6756 3891 6773
rect 3857 6739 3891 6756
rect 3036 6620 3053 6637
rect 3053 6620 3070 6637
rect 3109 6620 3121 6637
rect 3121 6620 3143 6637
rect 3182 6620 3189 6637
rect 3189 6620 3216 6637
rect 3255 6620 3257 6637
rect 3257 6620 3289 6637
rect 3328 6620 3359 6637
rect 3359 6620 3362 6637
rect 3401 6620 3427 6637
rect 3427 6620 3435 6637
rect 3474 6620 3495 6637
rect 3495 6620 3508 6637
rect 3547 6620 3563 6637
rect 3563 6620 3581 6637
rect 3620 6620 3631 6637
rect 3631 6620 3654 6637
rect 3693 6620 3699 6637
rect 3699 6620 3727 6637
rect 3766 6620 3767 6637
rect 3767 6620 3800 6637
rect 3036 6603 3070 6620
rect 3109 6603 3143 6620
rect 3182 6603 3216 6620
rect 3255 6603 3289 6620
rect 3328 6603 3362 6620
rect 3401 6603 3435 6620
rect 3474 6603 3508 6620
rect 3547 6603 3581 6620
rect 3620 6603 3654 6620
rect 3693 6603 3727 6620
rect 3766 6603 3800 6620
rect 3840 6603 3874 6637
rect 769 6530 803 6564
rect 843 6530 845 6564
rect 845 6530 877 6564
rect 916 6530 948 6564
rect 948 6530 950 6564
rect 989 6530 1017 6564
rect 1017 6530 1023 6564
rect 1062 6530 1086 6564
rect 1086 6530 1096 6564
rect 1135 6530 1155 6564
rect 1155 6530 1169 6564
rect 1208 6530 1224 6564
rect 1224 6530 1242 6564
rect 1281 6530 1293 6564
rect 1293 6530 1315 6564
rect 1354 6530 1363 6564
rect 1363 6530 1388 6564
rect 1427 6530 1433 6564
rect 1433 6530 1461 6564
rect 1500 6530 1503 6564
rect 1503 6530 1534 6564
rect 1573 6530 1607 6564
rect 53 6432 87 6447
rect 53 6413 87 6432
rect 53 6362 87 6368
rect 53 6334 87 6362
rect 53 6258 87 6289
rect 53 6255 87 6258
rect 53 6188 87 6210
rect 53 6176 87 6188
rect 403 6277 437 6281
rect 403 6247 437 6277
rect 403 6183 437 6209
rect 403 6175 437 6183
rect 485 6152 519 6155
rect 53 6118 87 6131
rect 53 6097 87 6118
rect 485 6121 519 6152
rect 53 6048 87 6052
rect 53 6018 87 6048
rect 309 6011 343 6045
rect 381 6027 403 6045
rect 403 6027 415 6045
rect 381 6011 415 6027
rect 53 5872 87 5900
rect 53 5866 87 5872
rect 53 5802 87 5822
rect 53 5788 87 5802
rect 485 5807 519 5826
rect 485 5792 519 5807
rect 53 5732 87 5744
rect 53 5710 87 5732
rect 53 5662 87 5667
rect 53 5633 87 5662
rect 53 5558 87 5590
rect 53 5556 87 5558
rect 53 5488 87 5513
rect 53 5479 87 5488
rect 53 5418 87 5436
rect 53 5402 87 5418
rect 485 5738 519 5749
rect 485 5715 519 5738
rect 485 5669 519 5671
rect 485 5637 519 5669
rect 485 5497 519 5499
rect 485 5465 519 5497
rect 485 5393 519 5414
rect 485 5380 519 5393
rect 53 5348 87 5359
rect 53 5325 87 5348
rect 485 5324 519 5329
rect 53 5278 87 5282
rect 53 5248 87 5278
rect 229 5114 263 5148
rect 301 5114 335 5148
rect 331 5040 365 5074
rect 403 5070 437 5074
rect 403 5040 437 5070
rect 485 5295 519 5324
rect 816 5994 850 6028
rect 893 5994 925 6028
rect 925 5994 927 6028
rect 970 5994 1002 6028
rect 1002 5994 1004 6028
rect 1047 5994 1079 6028
rect 1079 5994 1081 6028
rect 1124 5994 1156 6028
rect 1156 5994 1158 6028
rect 1201 5994 1233 6028
rect 1233 5994 1235 6028
rect 1277 5994 1310 6028
rect 1310 5994 1311 6028
rect 1395 5960 1429 5990
rect 1395 5956 1429 5960
rect 933 5885 967 5919
rect 1005 5894 1039 5919
rect 1005 5885 1039 5894
rect 1137 5885 1171 5919
rect 1209 5894 1243 5919
rect 1209 5885 1243 5894
rect 1395 5892 1429 5910
rect 1395 5876 1429 5892
rect 761 5728 795 5741
rect 761 5707 795 5728
rect 761 5659 795 5660
rect 761 5626 795 5659
rect 854 5571 877 5580
rect 877 5571 888 5580
rect 854 5546 888 5571
rect 926 5546 960 5580
rect 1137 5546 1171 5580
rect 1209 5546 1243 5580
rect 933 5435 967 5469
rect 1005 5448 1039 5469
rect 1005 5435 1039 5448
rect 1309 5487 1313 5509
rect 1313 5487 1343 5509
rect 1309 5475 1343 5487
rect 1309 5403 1343 5437
rect 1395 5824 1429 5830
rect 1395 5796 1429 5824
rect 1395 5722 1429 5751
rect 1395 5717 1429 5722
rect 1395 5654 1429 5672
rect 1395 5638 1429 5654
rect 1395 5586 1429 5593
rect 1395 5559 1429 5586
rect 1395 5484 1429 5514
rect 1395 5480 1429 5484
rect 1395 5416 1429 5435
rect 1395 5401 1429 5416
rect 761 5277 795 5311
rect 835 5277 869 5311
rect 909 5277 943 5311
rect 983 5277 1017 5311
rect 1057 5277 1091 5311
rect 1132 5277 1166 5311
rect 1207 5277 1241 5311
rect 1282 5277 1316 5311
rect 1357 5277 1391 5311
rect 485 5221 519 5243
rect 485 5209 519 5221
rect 53 4928 87 4931
rect 53 4897 87 4928
rect 53 4858 87 4859
rect 53 4825 87 4858
rect 403 4871 437 4880
rect 403 4846 437 4871
rect 403 4793 437 4808
rect 403 4774 437 4793
rect 331 4608 365 4642
rect 403 4638 437 4642
rect 403 4608 437 4638
rect 157 4512 191 4546
rect 255 4512 289 4546
rect 485 4531 519 4557
rect 485 4523 519 4531
rect -194 4420 -160 4454
rect -194 4348 -160 4382
rect -26 4450 8 4454
rect -26 4420 0 4450
rect 0 4420 8 4450
rect -26 4348 8 4382
rect 168 4372 202 4406
rect 240 4372 274 4406
rect -348 3972 -314 4006
rect -348 3830 -314 3864
rect -348 3389 -314 3398
rect -348 3364 -314 3389
rect -348 3283 -314 3305
rect -348 3271 -314 3283
rect -348 3179 -314 3212
rect -348 3178 -314 3179
rect -348 3109 -314 3118
rect -348 3084 -314 3109
rect -348 2793 -314 2814
rect -348 2780 -314 2793
rect -348 2723 -314 2737
rect -348 2703 -314 2723
rect -348 1883 -314 1895
rect -348 1861 -314 1883
rect -348 1813 -314 1819
rect -348 1785 -314 1813
rect -348 1709 -314 1742
rect -348 1708 -314 1709
rect -348 1639 -314 1665
rect -348 1631 -314 1639
rect -348 1463 -314 1495
rect -348 1461 -314 1463
rect -348 1393 -314 1415
rect -348 1381 -314 1393
rect -348 1081 -314 1099
rect -348 1065 -314 1081
rect -348 1012 -314 1018
rect -348 984 -314 1012
rect -348 350 -314 384
rect -114 4321 -80 4325
rect -114 4291 -80 4321
rect -114 4252 -80 4253
rect -114 4219 -80 4252
rect 320 4393 354 4427
rect 320 4321 354 4355
rect 485 4324 519 4348
rect 485 4314 519 4324
rect 403 4252 437 4286
rect 403 4180 437 4214
rect 196 4100 230 4134
rect 294 4100 328 4134
rect 485 4013 519 4046
rect 485 4012 519 4013
rect 485 3944 519 3960
rect 485 3926 519 3944
rect 485 3841 519 3874
rect 485 3840 519 3841
rect 403 3817 437 3833
rect 403 3799 437 3817
rect 403 3706 437 3735
rect 403 3701 437 3706
rect 485 3772 519 3788
rect 485 3754 519 3772
rect 485 3668 519 3702
rect 485 3392 519 3420
rect 485 3386 519 3392
rect 485 3323 519 3335
rect 485 3301 519 3323
rect 485 3220 519 3250
rect 485 3216 519 3220
rect 403 3195 437 3211
rect 403 3177 437 3195
rect 403 3084 437 3113
rect 403 3079 437 3084
rect 485 3151 519 3165
rect 485 3131 519 3151
rect 485 3047 519 3080
rect 485 3046 519 3047
rect 485 2772 519 2795
rect 485 2761 519 2772
rect 485 2704 519 2711
rect 485 2677 519 2704
rect 485 2602 519 2627
rect 485 2593 519 2602
rect 403 2573 437 2589
rect 403 2555 437 2573
rect 403 2457 437 2491
rect 485 2534 519 2543
rect 485 2509 519 2534
rect 485 2432 519 2458
rect 485 2424 519 2432
rect 237 2228 271 2262
rect 315 2228 349 2262
rect 394 2228 396 2262
rect 396 2228 428 2262
rect 473 2228 485 2262
rect 485 2228 507 2262
rect 739 4778 773 4812
rect 822 4778 831 4812
rect 831 4778 856 4812
rect 905 4778 912 4812
rect 912 4778 939 4812
rect 988 4778 993 4812
rect 993 4778 1022 4812
rect 1119 4744 1153 4774
rect 1119 4740 1153 4744
rect 1119 4675 1153 4701
rect 1119 4667 1153 4675
rect 783 4621 817 4642
rect 783 4608 817 4621
rect 855 4608 889 4642
rect 1119 4606 1153 4629
rect 1119 4595 1153 4606
rect 1119 4537 1153 4557
rect 1119 4523 1153 4537
rect 1119 4468 1153 4485
rect 1119 4451 1153 4468
rect 803 4405 817 4423
rect 817 4405 837 4423
rect 803 4389 837 4405
rect 901 4389 935 4423
rect 1119 4399 1153 4413
rect 1119 4379 1153 4399
rect 1119 4330 1153 4341
rect 1119 4307 1153 4330
rect 701 4006 735 4038
rect 701 4004 735 4006
rect 701 3938 735 3956
rect 701 3922 735 3938
rect 783 4252 817 4286
rect 1119 4261 1153 4269
rect 783 4180 817 4214
rect 933 4210 967 4244
rect 1031 4210 1065 4244
rect 1119 4235 1153 4261
rect 1119 4192 1153 4197
rect 1119 4163 1153 4192
rect 1119 4123 1153 4125
rect 1119 4091 1153 4123
rect 1119 4019 1153 4053
rect 1119 3950 1153 3981
rect 1119 3947 1153 3950
rect 701 3869 735 3874
rect 701 3840 735 3869
rect 1119 3881 1153 3909
rect 1119 3875 1153 3881
rect 701 3765 735 3792
rect 701 3758 735 3765
rect 701 3696 735 3711
rect 701 3677 735 3696
rect 783 3817 817 3833
rect 783 3799 817 3817
rect 783 3706 817 3735
rect 783 3701 817 3706
rect 1119 3812 1153 3837
rect 1119 3803 1153 3812
rect 1119 3744 1153 3765
rect 1119 3731 1153 3744
rect 1119 3676 1153 3693
rect 1119 3659 1153 3676
rect 701 3420 735 3423
rect 701 3389 735 3420
rect 701 3317 735 3340
rect 701 3306 735 3317
rect 1119 3608 1153 3621
rect 1119 3587 1153 3608
rect 1119 3540 1153 3549
rect 1119 3515 1153 3540
rect 1119 3472 1153 3477
rect 1119 3443 1153 3472
rect 1119 3404 1153 3405
rect 1119 3371 1153 3404
rect 1119 3302 1153 3333
rect 1119 3299 1153 3302
rect 701 3248 735 3257
rect 701 3223 735 3248
rect 1119 3234 1153 3261
rect 1119 3227 1153 3234
rect 701 3144 735 3173
rect 701 3139 735 3144
rect 701 3075 735 3089
rect 701 3055 735 3075
rect 783 3195 817 3211
rect 783 3177 817 3195
rect 783 3084 817 3113
rect 783 3079 817 3084
rect 1119 3166 1153 3189
rect 1119 3155 1153 3166
rect 1119 3098 1153 3117
rect 1119 3083 1153 3098
rect 1119 3030 1153 3045
rect 1119 3011 1153 3030
rect 701 2799 735 2801
rect 701 2767 735 2799
rect 701 2696 735 2719
rect 701 2685 735 2696
rect 863 2966 897 3000
rect 937 2966 971 3000
rect 1011 2966 1045 3000
rect 1119 2962 1153 2973
rect 1119 2939 1153 2962
rect 1119 2894 1153 2901
rect 863 2856 897 2890
rect 937 2856 971 2890
rect 1011 2856 1045 2890
rect 1119 2867 1153 2894
rect 1119 2826 1153 2829
rect 1119 2795 1153 2826
rect 701 2627 735 2637
rect 701 2603 735 2627
rect 875 2600 909 2634
rect 962 2600 996 2634
rect 1048 2600 1082 2634
rect 701 2523 735 2555
rect 701 2521 735 2523
rect 701 2454 735 2473
rect 701 2439 735 2454
rect 799 2484 833 2518
rect 897 2484 931 2518
rect 1119 2486 1153 2512
rect 1119 2478 1153 2486
rect 1119 2418 1153 2424
rect 1119 2390 1153 2418
rect 863 2328 897 2362
rect 937 2328 971 2362
rect 1011 2328 1045 2362
rect 749 2248 783 2282
rect 832 2248 839 2282
rect 839 2248 866 2282
rect 915 2248 945 2282
rect 945 2248 949 2282
rect 998 2248 1015 2282
rect 1015 2248 1032 2282
rect 1081 2248 1085 2282
rect 1085 2248 1115 2282
rect 237 2110 254 2136
rect 254 2110 271 2136
rect 315 2110 323 2136
rect 323 2110 349 2136
rect 394 2110 426 2136
rect 426 2110 428 2136
rect 473 2110 495 2136
rect 495 2110 507 2136
rect 237 2102 271 2110
rect 315 2102 349 2110
rect 394 2102 428 2110
rect 473 2102 507 2110
rect 173 1838 185 1867
rect 185 1838 207 1867
rect 248 1838 254 1867
rect 254 1838 282 1867
rect 323 1838 357 1867
rect 398 1838 426 1867
rect 426 1838 432 1867
rect 473 1838 495 1867
rect 495 1838 507 1867
rect 173 1833 207 1838
rect 248 1833 282 1838
rect 323 1833 357 1838
rect 398 1833 432 1838
rect 473 1833 507 1838
rect 173 1770 185 1795
rect 185 1770 207 1795
rect 248 1770 254 1795
rect 254 1770 282 1795
rect 323 1770 357 1795
rect 398 1770 426 1795
rect 426 1770 432 1795
rect 473 1770 495 1795
rect 495 1770 507 1795
rect 173 1761 207 1770
rect 248 1761 282 1770
rect 323 1761 357 1770
rect 398 1761 432 1770
rect 473 1761 507 1770
rect 403 1677 437 1709
rect 403 1675 437 1677
rect 403 1609 437 1637
rect 403 1603 437 1609
rect 246 1515 280 1549
rect 318 1515 352 1549
rect 713 1746 747 1774
rect 795 1746 829 1774
rect 877 1746 911 1774
rect 959 1746 993 1774
rect 1041 1746 1075 1774
rect 713 1740 725 1746
rect 725 1740 747 1746
rect 795 1740 797 1746
rect 797 1740 829 1746
rect 877 1740 903 1746
rect 903 1740 911 1746
rect 959 1740 974 1746
rect 974 1740 993 1746
rect 1041 1740 1045 1746
rect 1045 1740 1075 1746
rect 1171 1702 1205 1736
rect 711 1644 745 1678
rect 783 1662 817 1678
rect 783 1644 817 1662
rect 1171 1618 1205 1652
rect 1171 1534 1205 1568
rect 543 1441 577 1475
rect 615 1441 649 1475
rect 1171 1450 1205 1484
rect 488 1378 522 1392
rect 488 1358 519 1378
rect 519 1358 522 1378
rect 560 1358 594 1392
rect 704 1372 738 1406
rect 241 1292 275 1326
rect 313 1292 347 1326
rect 1171 1366 1205 1400
rect 879 1292 913 1326
rect 951 1292 985 1326
rect 1023 1292 1057 1326
rect 157 1192 191 1226
rect 229 1192 263 1226
rect 301 1192 335 1226
rect 1171 1283 1205 1317
rect 405 1193 437 1211
rect 437 1193 439 1211
rect 405 1177 439 1193
rect 477 1177 511 1211
rect 867 1197 901 1231
rect 939 1197 973 1231
rect 1011 1197 1045 1231
rect 1171 1200 1205 1234
rect 169 1064 203 1098
rect 241 1064 275 1098
rect 485 1093 519 1123
rect 485 1089 519 1093
rect 701 1070 735 1090
rect 701 1056 735 1070
rect 877 1064 911 1098
rect 949 1064 983 1098
rect 1021 1064 1055 1098
rect 539 978 573 1012
rect 611 978 645 1012
rect 485 822 519 852
rect 485 818 519 822
rect 403 779 437 787
rect 403 753 437 779
rect 403 707 437 708
rect 403 674 437 707
rect 403 601 437 630
rect 403 596 437 601
rect 403 529 437 552
rect 403 518 437 529
rect -172 292 -138 326
rect -100 314 -66 326
rect -100 292 -75 314
rect -75 292 -66 314
rect -28 292 6 326
rect 485 750 519 772
rect 485 738 519 750
rect 485 678 519 692
rect 485 658 519 678
rect 485 606 519 612
rect 485 578 519 606
rect 485 499 519 533
rect 485 424 519 454
rect 485 420 519 424
rect 485 352 519 375
rect 485 341 519 352
rect 485 280 519 296
rect -348 210 -314 244
rect 485 262 519 280
rect -461 138 -427 172
rect -386 138 -352 172
rect -311 138 -280 172
rect -280 138 -277 172
rect -236 138 -210 172
rect -210 138 -202 172
rect -161 138 -140 172
rect -140 138 -127 172
rect -85 138 -70 172
rect -70 138 -51 172
rect -9 138 1 172
rect 1 138 25 172
rect 67 138 101 172
rect 143 138 177 172
rect 219 138 231 172
rect 231 138 253 172
rect 295 138 303 172
rect 303 138 329 172
rect 371 138 375 172
rect 375 138 405 172
rect 447 138 481 172
rect 701 851 735 858
rect 1171 1058 1205 1092
rect 1171 980 1205 1014
rect 1171 902 1205 936
rect 701 824 735 851
rect 1171 824 1205 858
rect 701 782 735 786
rect 701 752 735 782
rect 701 575 735 604
rect 701 570 735 575
rect 701 506 735 529
rect 701 495 735 506
rect 701 436 735 454
rect 701 420 735 436
rect 701 366 735 380
rect 701 346 735 366
rect 701 296 735 306
rect 783 673 817 696
rect 783 662 817 673
rect 783 601 817 609
rect 783 575 817 601
rect 783 491 817 522
rect 783 488 817 491
rect 783 420 817 436
rect 783 402 817 420
rect 783 349 817 350
rect 783 316 817 349
rect 1171 746 1205 780
rect 1171 668 1205 702
rect 1171 590 1205 624
rect 1171 512 1205 546
rect 1171 433 1205 467
rect 1171 354 1205 388
rect 701 272 735 296
rect 1171 275 1205 309
rect 1171 196 1205 230
rect 739 158 773 192
rect 817 158 839 192
rect 839 158 851 192
rect 895 158 909 192
rect 909 158 929 192
rect 973 158 979 192
rect 979 158 1007 192
rect 1051 158 1085 192
<< metal1 >>
tri 647 8303 901 8557 se
rect 901 8505 1522 8557
rect 1574 8505 1592 8557
rect 1644 8505 1662 8557
rect 1714 8505 1732 8557
rect 1784 8505 1803 8557
rect 1855 8505 1861 8557
rect 901 8493 1861 8505
rect 901 8441 1522 8493
rect 1574 8441 1592 8493
rect 1644 8441 1662 8493
rect 1714 8441 1732 8493
rect 1784 8441 1803 8493
rect 1855 8441 1861 8493
tri 4817 8484 4883 8550 se
rect 4883 8504 5255 8550
tri 4883 8484 4903 8504 nw
rect 901 8429 1861 8441
rect 901 8377 1522 8429
rect 1574 8377 1592 8429
rect 1644 8377 1662 8429
rect 1714 8377 1732 8429
rect 1784 8377 1803 8429
rect 1855 8377 1861 8429
tri 4751 8418 4817 8484 se
tri 4817 8418 4883 8484 nw
tri 4710 8377 4751 8418 se
rect 901 8333 931 8377
tri 931 8333 975 8377 nw
tri 4685 8352 4710 8377 se
rect 4710 8352 4751 8377
tri 4751 8352 4817 8418 nw
tri 4666 8333 4685 8352 se
rect 4685 8333 4686 8352
tri 901 8303 931 8333 nw
tri 968 8303 998 8333 se
rect 998 8303 4686 8333
tri 601 8257 647 8303 se
rect 647 8267 865 8303
tri 865 8267 901 8303 nw
tri 932 8267 968 8303 se
rect 968 8287 4686 8303
tri 4686 8287 4751 8352 nw
rect 968 8267 998 8287
tri 998 8267 1018 8287 nw
rect 647 8257 799 8267
rect 344 8205 350 8257
rect 402 8205 420 8257
rect 472 8205 489 8257
rect 541 8205 553 8257
tri 462 8180 487 8205 ne
rect 487 8090 553 8205
rect 487 8056 493 8090
rect 527 8077 553 8090
rect 669 8201 799 8257
tri 799 8201 865 8267 nw
tri 866 8201 932 8267 se
tri 932 8201 998 8267 nw
rect 1516 8205 1522 8257
rect 1574 8205 1592 8257
rect 1644 8205 1662 8257
rect 1714 8205 1732 8257
rect 1784 8205 1803 8257
rect 1855 8205 2789 8257
rect 2841 8205 2859 8257
rect 2911 8205 2930 8257
rect 2982 8205 3001 8257
rect 3053 8205 3387 8257
rect 669 8135 733 8201
tri 733 8135 799 8201 nw
tri 800 8135 866 8201 se
tri 866 8135 932 8201 nw
rect 1516 8193 3387 8205
rect 1516 8141 1522 8193
rect 1574 8141 1592 8193
rect 1644 8141 1662 8193
rect 1714 8141 1732 8193
rect 1784 8141 1803 8193
rect 1855 8141 2789 8193
rect 2841 8141 2859 8193
rect 2911 8141 2930 8193
rect 2982 8141 3001 8193
rect 3053 8141 3387 8193
rect 669 8077 675 8135
tri 675 8077 733 8135 nw
tri 742 8077 800 8135 se
rect 527 8056 558 8077
tri 462 7987 487 8012 se
rect 487 7987 558 8056
tri 558 8052 583 8077 nw
tri 734 8069 742 8077 se
rect 742 8069 800 8077
tri 800 8069 866 8135 nw
rect 1516 8129 3387 8141
rect 1516 8077 1522 8129
rect 1574 8077 1592 8129
rect 1644 8077 1662 8129
rect 1714 8077 1732 8129
rect 1784 8077 1803 8129
rect 1855 8077 2789 8129
rect 2841 8077 2859 8129
rect 2911 8077 2930 8129
rect 2982 8077 3001 8129
rect 3053 8077 3387 8129
rect 3567 8205 4503 8257
rect 4555 8205 4568 8257
rect 4620 8205 4633 8257
rect 4685 8205 4698 8257
rect 4750 8205 4763 8257
rect 4815 8205 4829 8257
rect 4881 8205 4895 8257
rect 4947 8205 4961 8257
rect 5013 8205 5027 8257
rect 5079 8205 5093 8257
rect 5145 8205 5159 8257
rect 5211 8205 5217 8257
rect 3567 8193 5217 8205
rect 3567 8141 4503 8193
rect 4555 8141 4568 8193
rect 4620 8141 4633 8193
rect 4685 8141 4698 8193
rect 4750 8141 4763 8193
rect 4815 8141 4829 8193
rect 4881 8141 4895 8193
rect 4947 8141 4961 8193
rect 5013 8141 5027 8193
rect 5079 8141 5093 8193
rect 5145 8141 5159 8193
rect 5211 8141 5217 8193
rect 3567 8129 5217 8141
rect 3567 8077 4503 8129
rect 4555 8077 4568 8129
rect 4620 8077 4633 8129
rect 4685 8077 4698 8129
rect 4750 8077 4763 8129
rect 4815 8077 4829 8129
rect 4881 8077 4895 8129
rect 4947 8077 4961 8129
rect 5013 8077 5027 8129
rect 5079 8077 5093 8129
rect 5145 8077 5159 8129
rect 5211 8077 5217 8129
tri 717 8052 734 8069 se
tri 668 8003 717 8052 se
rect 717 8003 734 8052
tri 734 8003 800 8069 nw
rect 382 7935 388 7987
rect 440 7935 489 7987
rect 541 7935 547 7987
tri 547 7976 558 7987 nw
tri 641 7976 668 8003 se
rect 668 7976 677 8003
tri 611 7946 641 7976 se
rect 641 7946 677 7976
tri 677 7946 734 8003 nw
rect 611 7942 673 7946
tri 673 7942 677 7946 nw
rect 3007 7942 3445 7951
rect 3497 7942 3515 7951
rect 3567 7942 3897 7951
rect 487 7929 533 7935
tri 604 7744 611 7751 se
rect 611 7744 657 7942
tri 657 7926 673 7942 nw
tri 594 7734 604 7744 se
rect 604 7734 657 7744
tri 560 7700 594 7734 se
rect 594 7731 657 7734
rect 594 7700 626 7731
tri 626 7700 657 7731 nw
rect 735 7922 2010 7931
rect 2062 7922 2083 7931
rect 2135 7922 2156 7931
rect 2208 7922 2229 7931
rect 2281 7922 2302 7931
rect 2354 7922 2374 7931
rect 2426 7922 2446 7931
rect 2498 7922 2873 7931
rect 735 7888 851 7922
rect 885 7888 923 7922
rect 957 7888 995 7922
rect 1029 7888 1067 7922
rect 1101 7888 1139 7922
rect 1173 7888 1211 7922
rect 1245 7888 1283 7922
rect 1317 7888 1355 7922
rect 1389 7888 1427 7922
rect 1461 7888 1499 7922
rect 1533 7888 1571 7922
rect 1605 7888 1643 7922
rect 1677 7888 1715 7922
rect 1749 7888 1787 7922
rect 1821 7888 1859 7922
rect 1893 7888 1931 7922
rect 1965 7888 2003 7922
rect 2062 7888 2075 7922
rect 2135 7888 2147 7922
rect 2208 7888 2219 7922
rect 2281 7888 2291 7922
rect 2354 7888 2363 7922
rect 2426 7888 2435 7922
rect 2498 7888 2507 7922
rect 2541 7888 2579 7922
rect 2613 7888 2651 7922
rect 2685 7888 2723 7922
rect 2757 7888 2795 7922
rect 2829 7888 2873 7922
rect 735 7884 2010 7888
rect 735 7850 741 7884
rect 775 7879 2010 7884
rect 2062 7879 2083 7888
rect 2135 7879 2156 7888
rect 2208 7879 2229 7888
rect 2281 7879 2302 7888
rect 2354 7879 2374 7888
rect 2426 7879 2446 7888
rect 2498 7879 2873 7888
rect 775 7870 797 7879
tri 797 7870 806 7879 nw
tri 2802 7870 2811 7879 ne
rect 2811 7870 2873 7879
rect 775 7850 781 7870
tri 781 7854 797 7870 nw
tri 2811 7854 2827 7870 ne
rect 735 7809 781 7850
rect 735 7775 741 7809
rect 775 7775 781 7809
rect 1357 7784 1854 7836
rect 1906 7784 1918 7836
rect 1970 7784 2649 7836
rect 2827 7805 2873 7870
rect 735 7734 781 7775
rect 2827 7771 2833 7805
rect 2867 7771 2873 7805
rect 735 7700 741 7734
rect 775 7700 781 7734
rect 1191 7744 1602 7756
rect 1191 7710 1203 7744
rect 1237 7710 1276 7744
rect 1310 7710 1602 7744
rect 1191 7704 1602 7710
rect 1654 7704 1669 7756
rect 1721 7744 2790 7756
rect 1721 7710 2021 7744
rect 2055 7710 2094 7744
rect 2128 7710 2671 7744
rect 2705 7710 2744 7744
rect 2778 7710 2790 7744
rect 1721 7704 2790 7710
rect 2827 7729 2873 7771
tri 555 7695 560 7700 se
rect 560 7695 621 7700
tri 621 7695 626 7700 nw
rect 735 7695 781 7700
tri 781 7695 787 7701 sw
tri 2821 7695 2827 7701 se
rect 2827 7695 2833 7729
rect 2867 7695 2873 7729
tri 548 7688 555 7695 se
rect 555 7688 614 7695
tri 614 7688 621 7695 nw
rect 735 7688 787 7695
tri 787 7688 794 7695 sw
tri 2814 7688 2821 7695 se
rect 2821 7688 2873 7695
tri 545 7685 548 7688 se
rect 548 7685 611 7688
tri 611 7685 614 7688 nw
tri 536 7676 545 7685 se
rect 545 7676 602 7685
tri 602 7676 611 7685 nw
rect 735 7676 794 7688
tri 794 7676 806 7688 sw
tri 2802 7676 2814 7688 se
rect 2814 7676 2873 7688
tri 520 7660 536 7676 se
rect 536 7660 586 7676
tri 586 7660 602 7676 nw
rect 735 7660 2873 7676
tri 486 7626 520 7660 se
rect 520 7626 552 7660
tri 552 7626 586 7660 nw
rect 735 7626 741 7660
rect 775 7659 2873 7660
rect 775 7626 2010 7659
tri 479 7619 486 7626 se
rect 486 7619 545 7626
tri 545 7619 552 7626 nw
tri 463 7603 479 7619 se
rect 479 7603 529 7619
tri 529 7603 545 7619 nw
rect 735 7607 2010 7626
rect 2062 7607 2083 7659
rect 2135 7607 2156 7659
rect 2208 7607 2229 7659
rect 2281 7607 2302 7659
rect 2354 7607 2374 7659
rect 2426 7607 2446 7659
rect 2498 7653 2873 7659
rect 2498 7619 2833 7653
rect 2867 7619 2873 7653
rect 2498 7607 2873 7619
rect 3007 7912 3057 7942
rect 3091 7908 3133 7942
rect 3167 7908 3209 7942
rect 3243 7908 3285 7942
rect 3319 7908 3361 7942
rect 3395 7908 3437 7942
rect 3497 7908 3513 7942
rect 3567 7908 3589 7942
rect 3623 7908 3665 7942
rect 3699 7908 3741 7942
rect 3775 7908 3897 7942
rect 3059 7899 3445 7908
rect 3497 7899 3515 7908
rect 3567 7904 3897 7908
rect 3567 7899 3857 7904
tri 3059 7874 3084 7899 nw
tri 3826 7874 3851 7899 ne
rect 3007 7846 3059 7860
rect 3851 7870 3857 7899
rect 3891 7870 3897 7904
rect 3007 7780 3019 7794
rect 3053 7780 3059 7794
rect 3167 7786 3823 7836
tri 3732 7761 3757 7786 ne
rect 3007 7722 3059 7728
rect 3007 7714 3019 7722
rect 3053 7714 3059 7722
rect 3007 7649 3059 7662
rect 735 7603 802 7607
tri 802 7603 806 7607 nw
rect 3091 7607 3097 7659
rect 3149 7607 3161 7659
rect 3213 7607 3225 7659
rect 3277 7607 3289 7659
rect 3341 7607 3353 7659
rect 3405 7607 3729 7659
tri 460 7600 463 7603 se
rect 463 7600 526 7603
tri 526 7600 529 7603 nw
rect 735 7600 799 7603
tri 799 7600 802 7603 nw
tri 459 7599 460 7600 se
rect 460 7599 512 7600
rect 425 7586 512 7599
tri 512 7586 526 7600 nw
rect 735 7586 781 7600
rect 425 7553 479 7586
tri 479 7553 512 7586 nw
rect 735 7552 741 7586
rect 775 7552 781 7586
tri 781 7582 799 7600 nw
rect 3007 7591 3059 7597
rect 735 7512 781 7552
rect 344 7444 350 7496
rect 402 7444 428 7496
rect 480 7484 507 7496
rect 480 7450 493 7484
rect 480 7444 507 7450
rect 559 7444 565 7496
rect 344 7432 565 7444
rect 344 7380 350 7432
rect 402 7380 428 7432
rect 480 7412 507 7432
rect 480 7380 493 7412
rect 559 7380 565 7432
rect 735 7478 741 7512
rect 775 7478 781 7512
rect 1685 7511 1691 7563
rect 1743 7511 1758 7563
rect 1810 7551 3230 7563
rect 1810 7517 3111 7551
rect 3145 7517 3184 7551
rect 3218 7517 3230 7551
rect 1810 7511 3230 7517
tri 3742 7490 3757 7505 se
rect 3757 7490 3823 7786
tri 3735 7483 3742 7490 se
rect 3742 7483 3823 7490
rect 735 7438 781 7478
rect 735 7404 741 7438
rect 775 7404 781 7438
rect 1357 7431 1854 7483
rect 1906 7431 1918 7483
rect 1970 7431 2649 7483
tri 3732 7480 3735 7483 se
rect 3735 7480 3823 7483
rect 2929 7423 2937 7475
rect 2989 7423 3001 7475
rect 3053 7423 3059 7475
rect 3167 7434 3823 7480
tri 3732 7423 3743 7434 ne
rect 3743 7423 3823 7434
tri 3743 7414 3752 7423 ne
rect 3752 7414 3823 7423
tri 3752 7409 3757 7414 ne
rect 735 7392 781 7404
rect 344 7378 493 7380
rect 527 7378 565 7380
rect 344 7366 565 7378
rect 1191 7375 3607 7387
rect 612 7358 819 7364
rect 664 7318 819 7358
rect 1191 7341 1203 7375
rect 1237 7341 1276 7375
rect 1310 7341 3607 7375
rect 1191 7335 3607 7341
rect 3659 7335 3671 7387
rect 3723 7335 3729 7387
rect 664 7306 669 7318
rect 612 7298 669 7306
tri 669 7298 689 7318 nw
rect 612 7295 666 7298
tri 666 7295 669 7298 nw
rect 612 7291 664 7295
tri 664 7293 666 7295 nw
rect 612 7233 664 7239
rect 735 7278 781 7290
rect 735 7244 741 7278
rect 775 7244 781 7278
rect 1357 7255 2010 7307
rect 2062 7255 2083 7307
rect 2135 7255 2156 7307
rect 2208 7255 2229 7307
rect 2281 7255 2302 7307
rect 2354 7255 2374 7307
rect 2426 7255 2446 7307
rect 2498 7295 2873 7307
rect 2498 7261 2833 7295
rect 2867 7261 2873 7295
rect 2498 7255 2873 7261
rect 735 7211 781 7244
tri 2802 7230 2827 7255 ne
rect 692 7177 744 7183
rect 2561 7165 2567 7217
rect 2619 7165 2631 7217
rect 2683 7165 2791 7217
tri 2720 7148 2737 7165 ne
rect 2737 7148 2791 7165
tri 2737 7140 2745 7148 ne
tri 744 7126 747 7129 sw
rect 744 7125 747 7126
rect 692 7110 747 7125
tri -82 7065 -55 7092 se
rect -55 7065 544 7092
tri 544 7065 571 7092 sw
tri -108 7039 -82 7065 se
rect -82 7064 571 7065
rect -82 7039 -46 7064
tri -46 7039 -21 7064 nw
tri 512 7039 537 7064 ne
rect 537 7052 571 7064
tri 571 7052 584 7065 sw
rect 744 7108 747 7110
tri 747 7108 765 7126 sw
rect 744 7104 765 7108
tri 765 7104 769 7108 sw
rect 744 7058 1021 7104
rect 1357 7079 1854 7131
rect 1906 7079 1918 7131
rect 1970 7079 2649 7131
rect 2745 7099 2791 7148
rect 692 7052 1021 7058
rect 2745 7065 2751 7099
rect 2785 7065 2791 7099
rect 537 7039 584 7052
tri 2733 7039 2745 7051 se
rect 2745 7039 2791 7065
rect 2827 7202 2873 7255
rect 2827 7168 2833 7202
rect 2867 7168 2873 7202
rect 2827 7108 2873 7168
rect 2827 7074 2833 7108
rect 2867 7074 2873 7108
rect 3013 7295 3059 7307
rect 3013 7261 3019 7295
rect 3053 7261 3059 7295
rect 3013 7223 3059 7261
rect 3091 7255 3097 7307
rect 3149 7255 3174 7307
rect 3226 7255 3251 7307
rect 3303 7255 3328 7307
rect 3380 7255 3729 7307
tri 3059 7223 3078 7242 sw
rect 3013 7217 3078 7223
tri 3078 7217 3084 7223 sw
rect 3013 7211 3411 7217
rect 3013 7177 3019 7211
rect 3053 7177 3411 7211
rect 3013 7165 3411 7177
rect 3463 7165 3514 7217
rect 3566 7165 3572 7217
rect 3013 7148 3067 7165
tri 3067 7148 3084 7165 nw
tri 3752 7148 3757 7153 se
rect 3757 7148 3823 7414
rect 3013 7126 3059 7148
tri 3059 7140 3067 7148 nw
tri 3744 7140 3752 7148 se
rect 3752 7140 3823 7148
tri 3732 7128 3744 7140 se
rect 3744 7128 3823 7140
rect 3013 7092 3019 7126
rect 3053 7092 3059 7126
rect 3013 7080 3059 7092
rect 3167 7082 3823 7128
tri 3732 7080 3734 7082 ne
rect 3734 7080 3823 7082
rect 2827 7062 2873 7074
tri 3734 7073 3741 7080 ne
rect 3741 7073 3823 7080
tri 3741 7062 3752 7073 ne
rect 3752 7062 3823 7073
tri 3752 7057 3757 7062 ne
tri 2791 7039 2803 7051 sw
tri -117 7030 -108 7039 se
rect -108 7030 -55 7039
tri -55 7030 -46 7039 nw
tri 537 7032 544 7039 ne
rect 544 7032 584 7039
tri 544 7030 546 7032 ne
rect 546 7030 584 7032
tri -121 7026 -117 7030 se
rect -117 7026 -59 7030
tri -59 7026 -55 7030 nw
tri 546 7026 550 7030 ne
rect 550 7026 584 7030
tri 2720 7026 2733 7039 se
rect 2733 7026 2803 7039
tri 2803 7026 2816 7039 sw
tri -127 7020 -121 7026 se
rect -121 7020 -65 7026
tri -65 7020 -59 7026 nw
tri 550 7020 556 7026 ne
tri -138 7009 -127 7020 se
rect -127 7009 -99 7020
rect -138 6986 -99 7009
tri -99 6986 -65 7020 nw
tri -141 6838 -138 6841 se
rect -138 6838 -110 6986
tri -110 6975 -99 6986 nw
tri -175 6804 -141 6838 se
rect -141 6804 -110 6838
tri -182 6797 -175 6804 se
rect -175 6797 -110 6804
tri -202 6777 -182 6797 se
rect -182 6777 -110 6797
rect 44 6876 525 6882
rect 96 6842 189 6876
rect 223 6842 275 6876
rect 309 6842 361 6876
rect 395 6842 447 6876
rect 481 6842 525 6876
rect 96 6836 525 6842
rect 96 6828 113 6836
tri 113 6828 121 6836 nw
tri 454 6828 462 6836 ne
rect 462 6828 525 6836
rect 96 6824 99 6828
rect 44 6804 53 6824
rect 87 6814 99 6824
tri 99 6814 113 6828 nw
tri 462 6814 476 6828 ne
rect 476 6814 525 6828
rect 87 6804 96 6814
tri 96 6811 99 6814 nw
tri 476 6811 479 6814 ne
rect 479 6810 525 6814
rect 44 6775 96 6804
tri -1642 6713 -1630 6725 ne
rect -1630 6713 -1610 6725
rect 44 6717 96 6723
rect 145 6717 151 6769
rect 203 6717 220 6769
rect 272 6717 289 6769
rect 341 6717 347 6769
rect 556 6739 584 7026
rect 2009 7020 2751 7026
rect 2009 6986 2021 7020
rect 2055 6986 2094 7020
rect 2128 6992 2751 7020
rect 2785 7020 3220 7026
rect 2785 6992 3101 7020
rect 2128 6986 3101 6992
rect 3135 6986 3174 7020
rect 3208 6986 3220 7020
rect 2009 6980 3220 6986
rect 735 6944 781 6956
rect 735 6910 741 6944
rect 775 6910 781 6944
rect 612 6887 664 6893
rect 612 6820 664 6835
rect 735 6889 781 6910
rect 1516 6946 1568 6952
tri 781 6889 799 6907 sw
tri 1491 6889 1508 6906 ne
rect 1508 6894 1516 6906
rect 1919 6906 3729 6952
rect 1568 6894 1576 6906
rect 1508 6889 1576 6894
tri 1576 6889 1593 6906 nw
rect 735 6882 799 6889
tri 799 6882 806 6889 sw
tri 1508 6882 1515 6889 ne
rect 1515 6882 1568 6889
rect 735 6862 819 6882
tri 1515 6881 1516 6882 ne
rect 735 6828 741 6862
rect 775 6836 819 6862
rect 1142 6869 1188 6881
rect 775 6835 800 6836
tri 800 6835 801 6836 nw
rect 1142 6835 1148 6869
rect 1182 6835 1188 6869
rect 775 6832 797 6835
tri 797 6832 800 6835 nw
rect 775 6828 781 6832
rect 735 6816 781 6828
tri 781 6816 797 6832 nw
tri 664 6797 680 6813 sw
tri 1126 6797 1142 6813 se
rect 1142 6797 1188 6835
rect 1516 6879 1568 6882
tri 1568 6881 1576 6889 nw
rect 1516 6821 1568 6827
rect 2827 6866 2873 6878
rect 2827 6832 2833 6866
rect 2867 6832 2873 6866
rect 664 6788 680 6797
tri 680 6788 689 6797 sw
tri 1117 6788 1126 6797 se
rect 1126 6788 1148 6797
rect 664 6768 1148 6788
rect 612 6763 1148 6768
rect 1182 6763 1188 6797
rect 612 6762 1188 6763
tri 646 6751 657 6762 ne
rect 657 6751 1188 6762
tri 584 6739 594 6749 sw
tri 396 6713 397 6714 se
rect 397 6713 443 6725
tri -1630 6693 -1610 6713 ne
tri 376 6693 396 6713 se
rect 396 6693 403 6713
tri 372 6689 376 6693 se
rect 376 6689 403 6693
tri -29 6679 -19 6689 se
rect -19 6679 403 6689
rect 437 6679 443 6713
tri -67 6641 -29 6679 se
rect -29 6647 443 6679
rect -29 6641 -9 6647
tri -9 6641 -3 6647 nw
tri 372 6641 378 6647 ne
rect 378 6641 443 6647
tri -77 6631 -67 6641 se
rect -67 6631 -19 6641
tri -19 6631 -9 6641 nw
tri 378 6631 388 6641 ne
rect 388 6631 403 6641
tri -101 6607 -77 6631 se
rect -77 6607 -43 6631
tri -43 6607 -19 6631 nw
tri 388 6622 397 6631 ne
rect 44 6613 96 6619
tri -119 6589 -101 6607 se
rect -101 6589 -67 6607
rect -119 6471 -67 6589
tri -67 6583 -43 6607 nw
rect -119 6407 -67 6419
rect -119 6349 -67 6355
rect 397 6607 403 6631
rect 437 6607 443 6641
rect 397 6595 443 6607
rect 556 6723 594 6739
tri 594 6723 610 6739 sw
rect 1357 6727 1854 6779
rect 1906 6727 1918 6779
rect 1970 6727 2649 6779
rect 2827 6773 2873 6832
rect 2827 6739 2833 6773
rect 2867 6739 2873 6773
rect 2827 6727 2873 6739
rect 3013 6866 3163 6878
rect 3013 6832 3019 6866
rect 3053 6832 3163 6866
rect 3013 6826 3163 6832
rect 3215 6826 3233 6878
rect 3285 6826 3303 6878
rect 3355 6826 3373 6878
rect 3425 6826 3431 6878
rect 3013 6814 3146 6826
tri 3146 6814 3158 6826 nw
rect 3013 6773 3105 6814
tri 3105 6773 3146 6814 nw
tri 3732 6776 3757 6801 se
rect 3757 6776 3823 7062
rect 3013 6739 3019 6773
rect 3053 6739 3071 6773
tri 3071 6739 3105 6773 nw
rect 3013 6727 3059 6739
tri 3059 6727 3071 6739 nw
rect 3167 6730 3823 6776
rect 3851 7828 3897 7870
rect 3851 7794 3857 7828
rect 3891 7794 3897 7828
rect 3851 7752 3897 7794
rect 3851 7718 3857 7752
rect 3891 7718 3897 7752
rect 3851 7676 3897 7718
rect 3851 7642 3857 7676
rect 3891 7642 3897 7676
rect 3851 7600 3897 7642
rect 3851 7566 3857 7600
rect 3891 7566 3897 7600
rect 3851 7524 3897 7566
rect 3851 7490 3857 7524
rect 3891 7490 3897 7524
rect 3851 7448 3897 7490
rect 3851 7414 3857 7448
rect 3891 7414 3897 7448
rect 3851 7373 3897 7414
rect 3851 7339 3857 7373
rect 3891 7339 3897 7373
rect 3851 7298 3897 7339
rect 3851 7264 3857 7298
rect 3891 7264 3897 7298
rect 3851 7223 3897 7264
rect 3851 7189 3857 7223
rect 3891 7189 3897 7223
rect 3851 7148 3897 7189
rect 3851 7114 3857 7148
rect 3891 7114 3897 7148
rect 3851 7073 3897 7114
rect 3851 7039 3857 7073
rect 3891 7039 3897 7073
rect 3851 6998 3897 7039
rect 3851 6964 3857 6998
rect 3891 6964 3897 6998
rect 3851 6923 3897 6964
rect 3851 6889 3857 6923
rect 3891 6889 3897 6923
rect 3851 6848 3897 6889
rect 3851 6814 3857 6848
rect 3891 6814 3897 6848
rect 3851 6773 3897 6814
rect 3851 6739 3857 6773
rect 3891 6739 3897 6773
rect 3851 6727 3897 6739
rect 556 6719 1208 6723
rect 608 6699 1208 6719
tri 1208 6699 1232 6723 sw
rect 608 6694 4647 6699
tri 608 6669 633 6694 nw
tri 1197 6671 1220 6694 ne
rect 1220 6671 4647 6694
tri 4576 6669 4578 6671 ne
rect 4578 6669 4647 6671
rect 556 6652 608 6667
tri 4578 6666 4581 6669 ne
rect 4581 6666 4647 6669
rect 556 6582 608 6600
rect 701 6620 819 6666
tri 4581 6646 4601 6666 ne
rect 1573 6637 2010 6643
rect 2062 6637 2083 6643
rect 2135 6637 2156 6643
rect 2208 6637 2229 6643
rect 2281 6637 2302 6643
rect 2354 6637 2374 6643
rect 701 6603 737 6620
tri 737 6603 754 6620 nw
rect 1573 6603 1612 6637
rect 1646 6603 1688 6637
rect 1722 6603 1764 6637
rect 1798 6603 1840 6637
rect 1874 6603 1916 6637
rect 1950 6603 1992 6637
rect 2062 6603 2068 6637
rect 2135 6603 2144 6637
rect 2208 6603 2220 6637
rect 2281 6603 2296 6637
rect 2354 6603 2372 6637
tri 347 6564 356 6573 sw
rect 44 6544 96 6561
rect 145 6548 356 6564
tri 356 6548 372 6564 sw
rect 145 6542 664 6548
rect 145 6515 612 6542
rect 44 6475 96 6492
tri 587 6490 612 6515 ne
rect 612 6475 664 6490
rect 44 6413 53 6423
rect 87 6413 96 6423
rect 44 6406 96 6413
rect 145 6405 151 6457
rect 203 6405 220 6457
rect 272 6405 289 6457
rect 341 6405 347 6457
rect 612 6417 664 6423
tri 676 6354 701 6379 se
rect 701 6354 729 6603
tri 729 6595 737 6603 nw
tri 1548 6570 1573 6595 se
rect 1573 6591 2010 6603
rect 2062 6591 2083 6603
rect 2135 6591 2156 6603
rect 2208 6591 2229 6603
rect 2281 6591 2302 6603
rect 2354 6591 2374 6603
rect 2426 6591 2446 6643
rect 2498 6637 2880 6643
rect 2498 6603 2525 6637
rect 2559 6603 2602 6637
rect 2636 6603 2679 6637
rect 2713 6603 2756 6637
rect 2790 6603 2833 6637
rect 2867 6603 2880 6637
rect 2498 6591 2880 6603
rect 3013 6637 3163 6643
rect 3215 6637 3233 6643
rect 3285 6637 3303 6643
rect 3355 6637 3373 6643
rect 3425 6637 3897 6643
rect 3013 6603 3036 6637
rect 3070 6603 3109 6637
rect 3143 6603 3163 6637
rect 3216 6603 3233 6637
rect 3289 6603 3303 6637
rect 3362 6603 3373 6637
rect 3435 6603 3474 6637
rect 3508 6603 3547 6637
rect 3581 6603 3620 6637
rect 3654 6603 3693 6637
rect 3727 6603 3766 6637
rect 3800 6603 3840 6637
rect 3874 6603 3897 6637
rect 3013 6591 3163 6603
rect 3215 6591 3233 6603
rect 3285 6591 3303 6603
rect 3355 6591 3373 6603
rect 3425 6591 3897 6603
rect 1573 6570 1619 6591
rect 757 6564 1619 6570
tri 1619 6566 1644 6591 nw
rect 757 6530 769 6564
rect 803 6530 843 6564
rect 877 6530 916 6564
rect 950 6530 989 6564
rect 1023 6530 1062 6564
rect 1096 6530 1135 6564
rect 1169 6530 1208 6564
rect 1242 6530 1281 6564
rect 1315 6530 1354 6564
rect 1388 6530 1427 6564
rect 1461 6530 1500 6564
rect 1534 6530 1573 6564
rect 1607 6530 1619 6564
rect 757 6524 1619 6530
rect 1685 6511 1691 6563
rect 1743 6511 1758 6563
rect 1810 6511 4439 6563
rect 4491 6511 4503 6563
rect 4555 6511 4561 6563
rect 4601 6503 4647 6666
tri 1076 6433 1126 6483 se
rect 1126 6455 1683 6483
tri 1126 6433 1148 6455 nw
tri 1026 6383 1076 6433 se
tri 1076 6383 1126 6433 nw
rect 44 6337 53 6354
rect 87 6337 96 6354
rect 145 6321 729 6354
tri 976 6333 1026 6383 se
tri 1026 6333 1076 6383 nw
tri 347 6298 370 6321 nw
tri 676 6298 699 6321 ne
rect 699 6298 729 6321
tri 699 6296 701 6298 ne
rect 44 6268 53 6285
rect 87 6268 96 6285
rect 44 6210 96 6216
rect 44 6200 53 6210
rect 87 6200 96 6210
rect 397 6287 664 6293
rect 397 6281 612 6287
rect 397 6247 403 6281
rect 437 6260 612 6281
rect 437 6247 443 6260
rect 397 6209 443 6247
tri 443 6235 468 6260 nw
tri 587 6235 612 6260 ne
rect 397 6175 403 6209
rect 437 6175 443 6209
rect 397 6163 443 6175
rect 476 6216 528 6222
rect 44 6132 96 6148
rect 476 6155 528 6164
rect 612 6220 664 6235
rect 612 6162 664 6168
rect 44 6064 96 6080
rect 145 6079 151 6131
rect 203 6079 220 6131
rect 272 6079 289 6131
rect 341 6079 347 6131
rect 476 6121 485 6155
rect 519 6121 528 6155
rect 476 6105 528 6121
tri 662 6105 701 6144 se
rect 701 6126 729 6298
tri 926 6283 976 6333 se
tri 976 6283 1026 6333 nw
tri 876 6233 926 6283 se
tri 926 6233 976 6283 nw
tri 826 6183 876 6233 se
tri 876 6183 926 6233 nw
tri 776 6133 826 6183 se
tri 826 6133 876 6183 nw
tri 655 6098 662 6105 se
rect 662 6098 701 6105
tri 701 6098 729 6126 nw
tri 741 6098 776 6133 se
tri 636 6079 655 6098 se
rect 655 6079 676 6098
tri 609 6052 636 6079 se
rect 636 6073 676 6079
tri 676 6073 701 6098 nw
tri 726 6083 741 6098 se
rect 741 6083 776 6098
tri 776 6083 826 6133 nw
tri 716 6073 726 6083 se
rect 726 6073 730 6083
rect 636 6052 655 6073
tri 655 6052 676 6073 nw
tri 695 6052 716 6073 se
rect 716 6052 730 6073
tri 608 6051 609 6052 se
rect 609 6051 654 6052
tri 654 6051 655 6052 nw
tri 694 6051 695 6052 se
rect 695 6051 730 6052
rect 44 6006 96 6012
rect 297 6045 631 6051
rect 297 6011 309 6045
rect 343 6011 381 6045
rect 415 6028 631 6045
tri 631 6028 654 6051 nw
tri 676 6033 694 6051 se
rect 694 6037 730 6051
tri 730 6037 776 6083 nw
rect 694 6033 726 6037
tri 726 6033 730 6037 nw
tri 671 6028 676 6033 se
rect 676 6028 721 6033
tri 721 6028 726 6033 nw
rect 772 6028 1178 6037
rect 1230 6028 1270 6037
rect 415 6023 626 6028
tri 626 6023 631 6028 nw
tri 666 6023 671 6028 se
rect 671 6023 687 6028
rect 415 6011 608 6023
rect 297 6005 608 6011
tri 608 6005 626 6023 nw
tri 648 6005 666 6023 se
rect 666 6005 687 6023
tri 637 5994 648 6005 se
rect 648 5994 687 6005
tri 687 5994 721 6028 nw
rect 772 5994 816 6028
rect 850 5994 893 6028
rect 927 5994 970 6028
rect 1004 5994 1047 6028
rect 1081 5994 1124 6028
rect 1158 5994 1178 6028
rect 1235 5994 1270 6028
tri 633 5990 637 5994 se
rect 637 5990 683 5994
tri 683 5990 687 5994 nw
tri 626 5983 633 5990 se
rect 633 5983 676 5990
tri 676 5983 683 5990 nw
rect 772 5985 1178 5994
rect 1230 5985 1270 5994
rect 1322 5985 1363 6037
rect 1415 5990 1438 6037
tri 620 5977 626 5983 se
rect 626 5977 649 5983
rect -29 5956 649 5977
tri 649 5956 676 5983 nw
rect -29 5940 633 5956
tri 633 5940 649 5956 nw
rect 772 5940 818 5985
tri 818 5960 843 5985 nw
tri 1361 5960 1386 5985 ne
rect 1386 5956 1395 5985
rect 1429 5956 1438 5990
rect 1386 5944 1438 5956
rect 44 5906 96 5912
rect 347 5906 744 5912
rect 347 5866 692 5906
rect 44 5838 96 5854
tri 667 5841 692 5866 ne
rect 851 5873 857 5925
rect 909 5919 940 5925
rect 992 5919 1023 5925
rect 1075 5919 1255 5925
rect 909 5885 933 5919
rect 992 5885 1005 5919
rect 1075 5885 1137 5919
rect 1171 5885 1209 5919
rect 1243 5885 1255 5919
rect 909 5873 940 5885
rect 992 5873 1023 5885
rect 1075 5873 1255 5885
rect 1386 5877 1395 5892
rect 1429 5877 1438 5892
rect 692 5839 744 5854
rect 476 5832 528 5838
rect 44 5770 96 5786
rect 145 5753 151 5805
rect 203 5753 220 5805
rect 272 5753 289 5805
rect 341 5753 347 5805
rect 393 5778 445 5784
rect 44 5710 53 5718
rect 87 5710 96 5718
rect 44 5702 96 5710
rect 44 5634 53 5650
rect 87 5634 96 5650
rect 393 5711 445 5726
rect 393 5652 445 5659
rect 394 5650 444 5651
rect 393 5614 445 5650
rect 692 5781 744 5787
rect 1386 5810 1395 5825
rect 1429 5810 1438 5825
rect 476 5757 528 5780
rect 476 5683 528 5705
rect 476 5625 528 5631
rect 755 5741 801 5753
rect 755 5707 761 5741
rect 795 5707 801 5741
rect 755 5660 801 5707
rect 755 5626 761 5660
rect 795 5626 801 5660
rect 755 5614 801 5626
rect 1386 5751 1438 5758
rect 1386 5743 1395 5751
rect 1429 5743 1438 5751
rect 1386 5676 1438 5691
rect 394 5613 444 5614
tri 375 5593 393 5611 se
rect 393 5593 445 5612
tri 445 5593 463 5611 sw
rect 1386 5609 1438 5624
tri 368 5586 375 5593 se
rect 375 5586 463 5593
tri 463 5586 470 5593 sw
rect 44 5566 53 5582
rect 87 5566 96 5582
rect 347 5580 1255 5586
rect 347 5546 854 5580
rect 888 5546 926 5580
rect 960 5546 1137 5580
rect 1171 5546 1209 5580
rect 1243 5546 1255 5580
rect 347 5540 1255 5546
rect 1386 5542 1438 5557
rect 44 5513 96 5514
rect 44 5498 53 5513
rect 87 5498 96 5513
rect 44 5436 96 5446
rect 44 5430 53 5436
rect 87 5430 96 5436
rect 44 5362 96 5378
rect 476 5505 528 5511
rect 1303 5509 1349 5521
rect 1303 5475 1309 5509
rect 1343 5475 1349 5509
rect 476 5421 528 5453
rect 921 5469 1051 5475
rect 921 5435 933 5469
rect 967 5435 1005 5469
rect 1039 5435 1051 5469
tri 908 5403 921 5416 se
rect 921 5403 1051 5435
rect 1303 5437 1349 5475
tri 1051 5403 1064 5416 sw
tri 1290 5403 1303 5416 se
rect 1303 5403 1309 5437
rect 1343 5403 1349 5437
tri 906 5401 908 5403 se
rect 908 5401 1064 5403
tri 1064 5401 1066 5403 sw
tri 1288 5401 1290 5403 se
rect 1290 5401 1349 5403
tri 896 5391 906 5401 se
rect 906 5391 1066 5401
tri 1066 5391 1076 5401 sw
tri 1278 5391 1288 5401 se
rect 1288 5391 1349 5401
rect 145 5321 151 5373
rect 203 5321 220 5373
rect 272 5321 289 5373
rect 341 5321 347 5373
rect 393 5345 445 5351
rect 44 5294 96 5310
rect 44 5236 96 5242
rect 393 5278 445 5293
rect 393 5220 445 5226
rect 394 5218 444 5219
rect 476 5338 528 5369
rect 476 5255 528 5286
rect 476 5197 528 5203
rect 556 5345 1349 5391
rect 1386 5480 1395 5490
rect 1429 5480 1438 5490
rect 1386 5475 1438 5480
rect 1386 5408 1395 5423
rect 1429 5408 1438 5423
rect 394 5181 444 5182
tri 368 5154 393 5179 se
rect 393 5154 445 5180
tri 445 5154 470 5179 sw
tri 531 5154 556 5179 se
rect 556 5154 597 5345
tri 597 5320 622 5345 nw
tri 1364 5320 1386 5342 se
rect 1386 5340 1438 5356
tri 1361 5317 1364 5320 se
rect 1364 5317 1386 5320
rect 749 5311 1217 5317
rect 1269 5311 1287 5317
rect 1339 5311 1386 5317
rect 749 5277 761 5311
rect 795 5277 835 5311
rect 869 5277 909 5311
rect 943 5277 983 5311
rect 1017 5277 1057 5311
rect 1091 5277 1132 5311
rect 1166 5277 1207 5311
rect 1269 5277 1282 5311
rect 1339 5277 1357 5311
rect 1391 5277 1438 5288
rect 749 5265 1217 5277
rect 1269 5265 1287 5277
rect 1339 5265 1438 5277
rect 1640 5335 1701 5377
rect 65 5148 142 5154
rect 117 5108 142 5148
rect 143 5109 144 5153
rect 180 5109 181 5153
rect 182 5148 597 5154
rect 182 5114 229 5148
rect 263 5114 301 5148
rect 335 5114 597 5148
rect 182 5108 597 5114
rect 692 5157 744 5163
rect 65 5027 117 5096
tri 117 5083 142 5108 nw
tri 670 5083 692 5105 se
rect 692 5092 744 5105
tri 667 5080 670 5083 se
rect 670 5080 692 5083
rect 319 5074 692 5080
rect 319 5040 331 5074
rect 365 5040 403 5074
rect 437 5040 692 5074
rect 319 5034 744 5040
tri 117 5005 142 5030 sw
tri 1615 5005 1640 5030 se
rect 1640 5005 1676 5335
tri 1676 5310 1701 5335 nw
rect 117 4975 1676 5005
rect 65 4969 1676 4975
rect -112 4931 99 4937
rect -112 4898 53 4931
rect -112 4846 -106 4898
rect -54 4846 -21 4898
rect 31 4897 53 4898
rect 87 4897 99 4931
rect 31 4859 99 4897
rect 145 4889 151 4941
rect 203 4889 220 4941
rect 272 4889 289 4941
rect 341 4889 347 4941
rect 692 4935 1174 4941
rect 31 4846 53 4859
rect -112 4825 53 4846
rect 87 4825 99 4859
rect -112 4819 99 4825
rect 391 4880 449 4886
rect 744 4883 1174 4935
rect 391 4846 403 4880
rect 437 4846 449 4880
tri 387 4812 391 4816 se
rect 391 4812 449 4846
rect 612 4875 664 4881
tri 449 4812 453 4816 sw
tri 608 4812 612 4816 se
rect 612 4812 664 4823
tri 383 4808 387 4812 se
rect 387 4808 453 4812
tri 366 4791 383 4808 se
rect 383 4791 403 4808
rect -206 4774 403 4791
rect 437 4791 453 4808
tri 453 4791 474 4812 sw
tri 587 4791 608 4812 se
rect 608 4808 664 4812
rect 608 4791 612 4808
rect 437 4774 612 4791
rect -206 4756 612 4774
rect -206 4750 664 4756
rect 692 4825 1174 4883
rect 1482 4825 1488 4941
rect 692 4818 1488 4825
rect 692 4812 1220 4818
rect 692 4808 739 4812
rect 773 4778 822 4812
rect 856 4778 905 4812
rect 939 4778 988 4812
rect 1022 4778 1168 4812
rect 744 4774 1168 4778
rect 744 4772 1119 4774
rect 692 4750 744 4756
tri 744 4750 766 4772 nw
tri 1088 4750 1110 4772 ne
rect 1110 4750 1119 4772
rect -206 4740 -133 4750
tri -133 4740 -123 4750 nw
tri 1110 4747 1113 4750 ne
rect 1113 4740 1119 4750
rect 1153 4760 1168 4774
tri 1220 4793 1245 4818 nw
rect 1153 4747 1220 4760
rect 1153 4740 1168 4747
rect -206 4454 -148 4740
tri -148 4725 -133 4740 nw
rect -206 4420 -194 4454
rect -160 4420 -148 4454
rect -206 4382 -148 4420
rect -206 4348 -194 4382
rect -160 4348 -148 4382
rect -206 4342 -148 4348
tri -120 4713 -111 4722 se
rect -111 4713 145 4722
rect -120 4676 145 4713
rect 157 4676 879 4722
rect 1113 4701 1168 4740
rect -120 4667 -58 4676
tri -58 4667 -49 4676 nw
rect 1113 4667 1119 4701
rect 1153 4695 1168 4701
rect 1153 4682 1220 4695
rect 1153 4667 1168 4682
rect -120 4325 -74 4667
tri -74 4651 -58 4667 nw
rect 319 4642 901 4648
rect 319 4608 331 4642
rect 365 4608 403 4642
rect 437 4608 783 4642
rect 817 4608 855 4642
rect 889 4608 901 4642
rect 319 4602 901 4608
rect 1113 4630 1168 4667
rect 1113 4629 1220 4630
rect 1113 4595 1119 4629
rect 1153 4617 1220 4629
rect 1153 4595 1168 4617
rect 476 4568 528 4574
rect -38 4542 151 4558
rect -38 4490 -34 4542
rect 18 4506 151 4542
rect 203 4506 220 4558
rect 272 4546 289 4558
rect 272 4506 289 4512
rect 341 4506 347 4558
rect 1113 4565 1168 4595
rect 1113 4557 1220 4565
tri 588 4523 611 4546 se
rect 611 4523 674 4546
tri 674 4523 697 4546 sw
rect 1113 4523 1119 4557
rect 1153 4552 1220 4557
rect 1153 4523 1168 4552
rect 393 4516 445 4522
rect 18 4490 24 4506
rect -38 4485 24 4490
tri 24 4485 45 4506 nw
rect -38 4473 20 4485
tri 20 4481 24 4485 nw
rect -38 4421 -34 4473
rect 18 4421 20 4473
rect -38 4420 -26 4421
rect 8 4420 20 4421
rect -38 4404 20 4420
rect -38 4352 -34 4404
rect 18 4352 20 4404
rect -38 4348 -26 4352
rect 8 4348 20 4352
rect -38 4342 20 4348
rect 65 4472 117 4478
rect 476 4509 528 4516
tri 574 4509 588 4523 se
rect 588 4509 697 4523
tri 565 4500 574 4509 se
rect 574 4500 697 4509
tri 697 4500 720 4523 sw
tri 550 4485 565 4500 se
rect 565 4485 609 4500
tri 609 4485 624 4500 nw
tri 658 4485 673 4500 ne
rect 673 4485 720 4500
tri 720 4485 735 4500 sw
tri 529 4464 550 4485 se
rect 550 4464 575 4485
tri 380 4451 393 4464 se
rect 393 4451 445 4464
tri 445 4451 458 4464 sw
tri 516 4451 529 4464 se
rect 529 4451 575 4464
tri 575 4451 609 4485 nw
tri 673 4451 707 4485 ne
rect 707 4451 735 4485
tri 735 4451 769 4485 sw
rect 851 4457 857 4509
rect 909 4457 940 4509
rect 992 4457 1023 4509
rect 1075 4457 1081 4509
rect 1113 4500 1168 4523
rect 1113 4487 1220 4500
rect 1113 4485 1168 4487
rect 1113 4451 1119 4485
rect 1153 4451 1168 4485
tri 368 4439 380 4451 se
rect 380 4449 458 4451
rect 380 4439 393 4449
rect 65 4405 117 4420
rect 314 4427 393 4439
rect 156 4406 286 4412
rect 156 4372 168 4406
rect 202 4372 240 4406
rect 274 4372 286 4406
rect 156 4366 286 4372
rect 314 4393 320 4427
rect 354 4397 393 4427
rect 445 4439 458 4449
tri 458 4439 470 4451 sw
tri 515 4450 516 4451 se
rect 516 4450 574 4451
tri 574 4450 575 4451 nw
tri 707 4450 708 4451 ne
rect 708 4450 769 4451
tri 504 4439 515 4450 se
rect 515 4439 547 4450
rect 445 4423 547 4439
tri 547 4423 574 4450 nw
tri 708 4444 714 4450 ne
rect 714 4444 769 4450
rect 612 4438 664 4444
tri 714 4438 720 4444 ne
rect 720 4443 769 4444
tri 769 4443 777 4451 sw
rect 720 4438 777 4443
rect 445 4397 515 4423
rect 354 4393 515 4397
rect 314 4391 515 4393
tri 515 4391 547 4423 nw
rect 314 4389 383 4391
tri 383 4389 385 4391 nw
rect 314 4379 373 4389
tri 373 4379 383 4389 nw
tri 720 4423 735 4438 ne
rect 735 4429 777 4438
tri 777 4429 791 4443 sw
rect 1113 4435 1168 4451
rect 735 4423 947 4429
tri 735 4389 769 4423 ne
rect 769 4389 803 4423
rect 837 4389 901 4423
rect 935 4389 947 4423
tri 182 4355 193 4366 ne
rect 193 4355 267 4366
tri 267 4355 278 4366 nw
rect 314 4355 360 4379
tri 360 4366 373 4379 nw
rect 612 4374 664 4386
tri 769 4381 777 4389 ne
rect 777 4383 947 4389
rect 1113 4422 1220 4435
rect 1113 4413 1168 4422
rect 65 4347 117 4353
tri 193 4347 201 4355 ne
rect 201 4347 253 4355
tri 201 4346 202 4347 ne
rect 202 4346 253 4347
rect 66 4345 116 4346
tri 202 4345 203 4346 ne
rect 203 4345 253 4346
rect -120 4291 -114 4325
rect -80 4291 -74 4325
rect -120 4253 -74 4291
rect -120 4219 -114 4253
rect -80 4219 -74 4253
rect -120 4207 -74 4219
rect 65 4309 117 4345
tri 203 4341 207 4345 ne
rect 207 4341 253 4345
tri 253 4341 267 4355 nw
rect 66 4308 116 4309
rect 65 4301 117 4307
rect 208 4339 252 4340
rect 207 4303 253 4339
rect 314 4321 320 4355
rect 354 4321 360 4355
rect 314 4309 360 4321
rect 476 4357 528 4363
rect 208 4302 252 4303
tri 117 4286 132 4301 sw
tri 192 4286 207 4301 se
rect 207 4286 253 4301
rect 777 4379 844 4383
tri 844 4379 848 4383 nw
rect 1113 4379 1119 4413
rect 1153 4379 1168 4413
rect 777 4339 823 4379
tri 823 4358 844 4379 nw
rect 1113 4370 1168 4379
rect 778 4337 822 4338
rect 1113 4357 1220 4370
rect 1113 4341 1168 4357
rect 612 4315 664 4322
rect 613 4313 663 4314
rect 117 4276 132 4286
tri 132 4276 142 4286 sw
tri 182 4276 192 4286 se
rect 192 4276 253 4286
rect 117 4249 142 4276
rect 144 4275 180 4276
rect 65 4224 142 4249
rect 143 4225 181 4275
rect 182 4252 253 4276
rect 397 4286 443 4299
rect 476 4298 528 4305
rect 1113 4307 1119 4341
rect 1153 4307 1168 4341
rect 1113 4305 1168 4307
rect 778 4300 822 4301
tri 253 4252 275 4274 sw
tri 375 4252 397 4274 se
rect 397 4252 403 4286
rect 437 4252 443 4286
rect 777 4286 823 4299
rect 613 4276 663 4277
tri 443 4252 466 4275 sw
tri 589 4252 612 4275 se
rect 612 4252 664 4275
tri 664 4252 687 4275 sw
tri 754 4252 777 4275 se
rect 777 4252 783 4286
rect 817 4269 823 4286
rect 1113 4292 1220 4305
tri 823 4269 829 4275 sw
rect 1113 4269 1168 4292
rect 817 4252 829 4269
rect 182 4249 275 4252
tri 275 4249 278 4252 sw
tri 372 4249 375 4252 se
rect 375 4250 466 4252
tri 466 4250 468 4252 sw
tri 587 4250 589 4252 se
rect 589 4250 687 4252
tri 687 4250 689 4252 sw
tri 752 4250 754 4252 se
rect 754 4250 829 4252
tri 829 4250 848 4269 sw
rect 375 4249 871 4250
rect 873 4249 909 4250
rect 144 4224 180 4225
rect 182 4224 871 4249
rect 65 4214 132 4224
tri 132 4214 142 4224 nw
tri 182 4214 192 4224 ne
rect 192 4214 871 4224
tri 117 4199 132 4214 nw
tri 192 4199 207 4214 ne
rect 207 4199 403 4214
tri 372 4180 391 4199 ne
rect 391 4180 403 4199
rect 437 4205 783 4214
rect 437 4180 443 4205
tri 443 4180 468 4205 nw
tri 752 4180 777 4205 ne
rect 777 4180 783 4205
rect 817 4204 871 4214
rect 872 4205 910 4249
rect 911 4244 1077 4250
rect 911 4210 933 4244
rect 967 4210 1031 4244
rect 1065 4210 1077 4244
rect 873 4204 909 4205
rect 911 4204 1077 4210
rect 1113 4235 1119 4269
rect 1153 4240 1168 4269
rect 1153 4235 1220 4240
rect 1113 4227 1220 4235
rect 817 4197 841 4204
tri 841 4197 848 4204 nw
rect 1113 4197 1168 4227
rect 817 4180 823 4197
tri 391 4174 397 4180 ne
rect 397 4168 443 4180
rect 777 4168 823 4180
tri 823 4179 841 4197 nw
tri 117 4163 119 4165 sw
rect 1113 4163 1119 4197
rect 1153 4175 1168 4197
rect 1153 4163 1220 4175
rect 117 4162 119 4163
rect 65 4140 119 4162
tri 119 4140 142 4163 sw
rect 1113 4162 1220 4163
rect 65 4127 142 4140
rect 117 4094 142 4127
rect 143 4095 144 4139
rect 180 4095 181 4139
rect 182 4134 879 4140
rect 182 4100 196 4134
rect 230 4100 294 4134
rect 328 4100 879 4134
rect 182 4094 879 4100
rect 1113 4125 1168 4162
rect 117 4091 139 4094
tri 139 4091 142 4094 nw
tri 372 4091 375 4094 ne
rect 375 4091 465 4094
tri 465 4091 468 4094 nw
tri 587 4091 590 4094 ne
rect 590 4091 686 4094
tri 686 4091 689 4094 nw
tri 752 4091 755 4094 ne
rect 755 4091 845 4094
tri 845 4091 848 4094 nw
rect 1113 4091 1119 4125
rect 1153 4110 1168 4125
rect 1153 4097 1220 4110
rect 1153 4091 1168 4097
rect 65 4069 117 4075
tri 117 4069 139 4091 nw
tri 375 4069 397 4091 ne
rect -354 4006 -308 4018
rect -354 3972 -348 4006
rect -314 3972 -308 4006
rect -354 3864 -308 3972
rect -354 3830 -348 3864
rect -314 3830 -308 3864
rect 16 3887 347 4041
rect 16 3860 151 3887
tri 120 3840 140 3860 ne
rect 140 3840 151 3860
tri 140 3837 143 3840 ne
rect 143 3837 151 3840
tri 143 3835 145 3837 ne
rect 145 3835 151 3837
rect 203 3835 220 3887
rect 272 3835 289 3887
rect 341 3835 347 3887
rect -354 3818 -308 3830
rect 397 3833 443 4091
tri 443 4069 465 4091 nw
tri 590 4069 612 4091 ne
rect 612 4069 664 4091
tri 664 4069 686 4091 nw
tri 755 4069 777 4091 ne
rect 613 4067 663 4068
rect 65 3817 117 3823
rect 65 3752 117 3765
rect 65 3694 117 3700
rect 66 3692 116 3693
rect 397 3799 403 3833
rect 437 3799 443 3833
rect 397 3735 443 3799
rect 397 3701 403 3735
rect 437 3701 443 3735
rect 397 3689 443 3701
rect 476 4052 528 4058
rect 692 4044 744 4050
rect 476 3984 528 4000
rect 476 3926 485 3932
rect 519 3926 528 3932
rect 476 3916 528 3926
rect 476 3848 485 3864
rect 519 3848 528 3864
rect 476 3788 528 3796
rect 476 3781 485 3788
rect 519 3781 528 3788
rect 476 3714 528 3729
rect 613 4030 663 4031
rect 612 4015 664 4029
rect 612 3949 664 3963
rect 612 3884 664 3897
rect 612 3819 664 3832
rect 612 3754 664 3767
rect 612 3694 664 3702
rect 613 3692 663 3693
rect 692 3979 744 3992
rect 692 3922 701 3927
rect 735 3922 744 3927
rect 692 3915 744 3922
rect 692 3851 701 3863
rect 735 3851 744 3863
rect 692 3792 744 3799
rect 692 3787 701 3792
rect 735 3787 744 3792
rect 692 3723 744 3735
rect 777 3833 823 4091
tri 823 4069 845 4091 nw
rect 1113 4053 1168 4091
rect 1113 4019 1119 4053
rect 1153 4045 1168 4053
rect 1153 4032 1220 4045
rect 1153 4019 1168 4032
rect 1113 3981 1168 4019
rect 1113 3947 1119 3981
rect 1153 3980 1168 3981
rect 1153 3967 1220 3980
rect 1153 3947 1168 3967
rect 1113 3915 1168 3947
rect 1113 3909 1220 3915
rect 851 3835 857 3887
rect 909 3835 940 3887
rect 992 3835 1023 3887
rect 1075 3835 1081 3887
rect 1113 3875 1119 3909
rect 1153 3902 1220 3909
rect 1153 3875 1168 3902
rect 1113 3850 1168 3875
rect 1113 3837 1220 3850
rect 777 3799 783 3833
rect 817 3799 823 3833
rect 777 3735 823 3799
rect 777 3701 783 3735
rect 817 3701 823 3735
rect 777 3689 823 3701
rect 1113 3803 1119 3837
rect 1153 3803 1168 3837
rect 1113 3785 1168 3803
rect 1685 3922 1737 3928
rect 1685 3856 1737 3870
rect 1685 3798 1737 3804
rect 1113 3771 1220 3785
rect 1113 3765 1168 3771
rect 1113 3731 1119 3765
rect 1153 3731 1168 3765
rect 1113 3719 1168 3731
rect 1113 3705 1220 3719
rect 1113 3693 1168 3705
rect 692 3665 744 3671
rect 476 3656 528 3662
rect 1113 3659 1119 3693
rect 1153 3659 1168 3693
rect 66 3655 116 3656
rect 65 3628 117 3654
rect 613 3655 663 3656
tri 117 3628 142 3653 sw
tri 587 3628 612 3653 se
rect 612 3628 664 3654
rect 1113 3653 1168 3659
tri 664 3628 689 3653 sw
rect 1113 3639 1220 3653
rect 65 3582 879 3628
rect 1113 3621 1168 3639
rect 1113 3587 1119 3621
rect 1153 3587 1168 3621
rect 1113 3573 1220 3587
rect 1113 3549 1168 3573
rect 65 3472 879 3518
rect 1113 3515 1119 3549
rect 1153 3521 1168 3549
tri 1220 3532 1245 3557 sw
rect 1220 3521 1695 3532
rect 1153 3515 1695 3521
rect 1113 3507 1695 3515
rect 1113 3477 1168 3507
rect 65 3446 117 3472
tri 117 3447 142 3472 nw
tri 372 3447 397 3472 ne
rect 66 3444 116 3445
rect -354 3398 -308 3410
rect -354 3364 -348 3398
rect -314 3364 -308 3398
rect -354 3305 -308 3364
rect -354 3271 -348 3305
rect -314 3271 -308 3305
rect -354 3212 -308 3271
rect -354 3178 -348 3212
rect -314 3178 -308 3212
rect -354 3118 -308 3178
rect -354 3084 -348 3118
rect -314 3084 -308 3118
rect -354 3072 -308 3084
rect 66 3407 116 3408
rect 65 3376 117 3406
rect 65 3302 117 3324
rect 65 3228 117 3250
rect 145 3213 151 3265
rect 203 3213 220 3265
rect 272 3213 289 3265
rect 341 3213 347 3265
rect 65 3155 117 3176
rect 65 3072 117 3103
rect 66 3070 116 3071
rect 397 3211 443 3472
tri 443 3447 468 3472 nw
tri 587 3447 612 3472 ne
rect 612 3446 664 3472
tri 664 3447 689 3472 nw
tri 752 3447 777 3472 ne
rect 613 3444 663 3445
rect 397 3177 403 3211
rect 437 3177 443 3211
rect 397 3113 443 3177
rect 397 3079 403 3113
rect 437 3079 443 3113
rect 397 3067 443 3079
rect 476 3426 528 3432
rect 692 3429 744 3435
rect 476 3359 528 3374
rect 476 3301 485 3307
rect 519 3301 528 3307
rect 476 3292 528 3301
rect 476 3225 485 3240
rect 519 3225 528 3240
rect 476 3165 528 3173
rect 476 3158 485 3165
rect 519 3158 528 3165
rect 476 3092 528 3106
rect 613 3407 663 3408
rect 612 3394 664 3406
rect 612 3328 664 3342
rect 612 3263 664 3276
rect 612 3198 664 3211
rect 612 3133 664 3146
rect 612 3072 664 3081
rect 613 3070 663 3071
rect 692 3363 744 3377
rect 692 3306 701 3311
rect 735 3306 744 3311
rect 692 3297 744 3306
rect 692 3231 701 3245
rect 735 3231 744 3245
rect 692 3173 744 3179
rect 692 3166 701 3173
rect 735 3166 744 3173
rect 692 3101 744 3114
rect 777 3211 823 3472
tri 823 3447 848 3472 nw
rect 1113 3443 1119 3477
rect 1153 3455 1168 3477
rect 1220 3455 1695 3507
rect 1153 3443 1695 3455
rect 1113 3441 1695 3443
rect 1113 3405 1168 3441
rect 1113 3371 1119 3405
rect 1153 3389 1168 3405
rect 1220 3389 1695 3441
rect 1153 3375 1695 3389
rect 1153 3371 1168 3375
rect 1113 3333 1168 3371
rect 1113 3299 1119 3333
rect 1153 3323 1168 3333
rect 1220 3323 1695 3375
rect 1153 3309 1695 3323
rect 1153 3299 1168 3309
rect 851 3213 857 3265
rect 909 3213 940 3265
rect 992 3213 1023 3265
rect 1075 3213 1081 3265
rect 1113 3261 1168 3299
rect 1113 3227 1119 3261
rect 1153 3257 1168 3261
rect 1220 3257 1695 3309
rect 1153 3243 1695 3257
rect 1153 3227 1168 3243
rect 777 3177 783 3211
rect 817 3177 823 3211
rect 777 3113 823 3177
rect 777 3079 783 3113
rect 817 3079 823 3113
rect 777 3067 823 3079
rect 1113 3191 1168 3227
rect 1220 3206 1695 3243
rect 1113 3189 1220 3191
rect 1113 3155 1119 3189
rect 1153 3177 1220 3189
tri 1220 3181 1245 3206 nw
rect 1153 3155 1168 3177
rect 1113 3125 1168 3155
rect 1113 3117 1220 3125
rect 1113 3083 1119 3117
rect 1153 3111 1220 3117
rect 1153 3083 1168 3111
rect 692 3043 744 3049
rect 1113 3059 1168 3083
rect 1113 3045 1220 3059
rect 476 3034 528 3040
rect 66 3033 116 3034
rect 65 3011 117 3032
rect 613 3033 663 3034
tri 117 3011 137 3031 sw
tri 592 3011 612 3031 se
rect 612 3011 664 3032
tri 664 3011 684 3031 sw
rect 1113 3011 1119 3045
rect 1153 3011 1168 3045
rect 65 3006 137 3011
tri 137 3006 142 3011 sw
tri 587 3006 592 3011 se
rect 592 3006 684 3011
tri 684 3006 689 3011 sw
rect 65 3000 1057 3006
rect 65 2966 863 3000
rect 897 2966 937 3000
rect 971 2966 1011 3000
rect 1045 2966 1057 3000
rect 65 2960 1057 2966
rect 1113 2993 1168 3011
rect 1113 2987 1220 2993
tri 1220 2987 1270 3037 sw
rect 1113 2975 1695 2987
rect 1113 2973 1168 2975
rect 1113 2939 1119 2973
rect 1153 2939 1168 2973
rect 1113 2923 1168 2939
rect 1220 2923 1232 2975
rect 1284 2923 1296 2975
rect 1348 2923 1360 2975
rect 1412 2923 1424 2975
rect 1476 2923 1695 2975
rect 1113 2908 1695 2923
rect 1113 2901 1168 2908
rect 65 2890 1057 2896
rect 65 2856 863 2890
rect 897 2856 937 2890
rect 971 2856 1011 2890
rect 1045 2856 1057 2890
rect 65 2850 1057 2856
rect 1113 2867 1119 2901
rect 1153 2867 1168 2901
rect 1113 2856 1168 2867
rect 1220 2856 1232 2908
rect 1284 2856 1296 2908
rect 1348 2856 1360 2908
rect 1412 2856 1424 2908
rect 1476 2856 1695 2908
rect 65 2829 121 2850
tri 121 2829 142 2850 nw
tri 372 2829 393 2850 ne
rect 393 2829 447 2850
tri 447 2829 468 2850 nw
tri 587 2829 608 2850 ne
rect 608 2829 668 2850
tri 668 2829 689 2850 nw
tri 752 2829 773 2850 ne
rect 773 2829 827 2850
tri 827 2829 848 2850 nw
rect 1113 2841 1695 2856
rect 1113 2829 1168 2841
rect -354 2814 -308 2826
rect 65 2824 117 2829
tri 117 2825 121 2829 nw
tri 393 2825 397 2829 ne
rect 66 2822 116 2823
rect -354 2780 -348 2814
rect -314 2780 -308 2814
rect -354 2737 -308 2780
rect -354 2703 -348 2737
rect -314 2703 -308 2737
rect -354 2691 -308 2703
rect 66 2785 116 2786
rect 65 2753 117 2784
rect 65 2682 117 2701
rect 65 2610 117 2630
rect 145 2591 151 2643
rect 203 2591 220 2643
rect 272 2591 289 2643
rect 341 2591 347 2643
rect 65 2538 117 2558
rect 65 2450 117 2486
rect 66 2448 116 2449
rect 397 2589 443 2829
tri 443 2825 447 2829 nw
tri 608 2825 612 2829 ne
rect 612 2823 664 2829
tri 664 2825 668 2829 nw
tri 773 2825 777 2829 ne
rect 613 2821 663 2822
rect 692 2807 744 2813
rect 397 2555 403 2589
rect 437 2555 443 2589
rect 397 2491 443 2555
rect 397 2457 403 2491
rect 437 2457 443 2491
rect 397 2445 443 2457
rect 476 2801 528 2807
rect 476 2734 528 2749
rect 476 2677 485 2682
rect 519 2677 528 2682
rect 476 2668 528 2677
rect 613 2784 663 2785
rect 612 2752 664 2783
rect 612 2685 664 2700
rect 612 2627 664 2633
rect 692 2742 744 2755
rect 692 2685 701 2690
rect 735 2685 744 2690
rect 692 2677 744 2685
rect 476 2602 485 2616
rect 519 2602 528 2616
rect 476 2543 528 2550
rect 476 2536 485 2543
rect 519 2536 528 2543
rect 476 2470 528 2484
rect 476 2412 528 2418
rect 692 2613 701 2625
rect 735 2613 744 2625
rect 692 2555 744 2561
rect 692 2549 701 2555
rect 735 2549 744 2555
rect 692 2485 744 2497
rect 777 2524 823 2829
tri 823 2825 827 2829 nw
rect 1113 2795 1119 2829
rect 1153 2795 1168 2829
rect 1113 2789 1168 2795
rect 1220 2789 1232 2841
rect 1284 2789 1296 2841
rect 1348 2789 1360 2841
rect 1412 2789 1424 2841
rect 1476 2789 1695 2841
rect 1113 2783 1695 2789
rect 863 2749 1695 2755
rect 915 2697 927 2749
rect 979 2697 991 2749
rect 1043 2697 1055 2749
rect 1107 2697 1695 2749
rect 863 2680 1695 2697
rect 915 2628 927 2680
rect 979 2634 991 2680
rect 1043 2634 1055 2680
rect 1043 2628 1048 2634
rect 1107 2628 1695 2680
rect 863 2610 875 2628
rect 909 2610 962 2628
rect 996 2610 1048 2628
rect 1082 2610 1695 2628
rect 915 2558 927 2610
rect 1043 2600 1048 2610
rect 979 2558 991 2600
rect 1043 2558 1055 2600
rect 1107 2558 1695 2610
rect 863 2552 1695 2558
tri 823 2524 848 2549 sw
rect 777 2518 943 2524
rect 777 2488 799 2518
tri 777 2484 781 2488 ne
rect 781 2484 799 2488
rect 833 2484 897 2518
rect 931 2484 943 2518
rect 1113 2518 1695 2524
rect 1113 2512 1168 2518
tri 781 2478 787 2484 ne
rect 787 2478 943 2484
tri 1106 2478 1113 2485 se
rect 1113 2478 1119 2512
rect 1153 2478 1168 2512
tri 1103 2475 1106 2478 se
rect 1106 2475 1168 2478
tri 744 2450 769 2475 sw
tri 1078 2450 1103 2475 se
rect 1103 2466 1168 2475
rect 1220 2466 1232 2518
rect 1284 2466 1296 2518
rect 1348 2466 1360 2518
rect 1412 2466 1424 2518
rect 1476 2466 1695 2518
rect 1103 2450 1695 2466
rect 744 2433 1695 2450
rect 692 2429 1695 2433
rect 692 2424 1168 2429
rect 692 2412 1119 2424
rect 66 2411 116 2412
tri 1053 2411 1054 2412 ne
rect 1054 2411 1119 2412
tri 1054 2410 1055 2411 ne
rect 1055 2410 1119 2411
rect 65 2390 117 2410
tri 1055 2409 1056 2410 ne
rect 1056 2409 1119 2410
tri 117 2390 136 2409 sw
tri 1056 2390 1075 2409 ne
rect 1075 2390 1119 2409
rect 1153 2390 1168 2424
rect 65 2384 136 2390
tri 136 2384 142 2390 sw
tri 1075 2384 1081 2390 ne
rect 1081 2384 1168 2390
rect 65 2368 758 2384
tri 758 2368 774 2384 sw
tri 1081 2368 1097 2384 ne
rect 1097 2377 1168 2384
rect 1220 2377 1232 2429
rect 1284 2377 1296 2429
rect 1348 2377 1360 2429
rect 1412 2377 1424 2429
rect 1476 2377 1695 2429
rect 1097 2368 1695 2377
rect 65 2362 1057 2368
rect 65 2338 863 2362
tri 587 2328 597 2338 ne
rect 597 2328 679 2338
tri 679 2328 689 2338 nw
tri 738 2328 748 2338 ne
rect 748 2328 863 2338
rect 897 2328 937 2362
rect 971 2328 1011 2362
rect 1045 2328 1057 2362
tri 1097 2352 1113 2368 ne
tri 597 2313 612 2328 ne
rect 612 2311 664 2328
tri 664 2313 679 2328 nw
tri 748 2322 754 2328 ne
rect 754 2322 1057 2328
rect 1113 2340 1695 2368
tri 1111 2311 1113 2313 se
rect 1113 2311 1168 2340
tri 1110 2310 1111 2311 se
rect 1111 2310 1168 2311
tri -652 2282 -629 2305 se
rect -629 2298 197 2305
rect -629 2282 145 2298
tri -672 2262 -652 2282 se
rect -652 2262 145 2282
tri -706 2228 -672 2262 se
rect -672 2246 145 2262
rect 476 2304 528 2310
tri 465 2282 476 2293 se
tri 451 2268 465 2282 se
rect 465 2268 476 2282
rect -672 2228 197 2246
tri -797 2137 -706 2228 se
rect -706 2226 197 2228
rect -706 2190 145 2226
rect -706 2137 -341 2190
tri -341 2165 -316 2190 nw
tri 120 2165 145 2190 ne
rect -797 1935 -341 2137
rect 145 2154 197 2174
rect 145 2096 197 2102
rect 225 2262 476 2268
rect 225 2249 237 2262
rect 271 2249 315 2262
rect 225 2197 231 2249
rect 283 2228 315 2249
rect 349 2228 394 2262
rect 428 2228 473 2262
rect 507 2229 528 2252
rect 283 2197 476 2228
rect 225 2185 476 2197
rect 225 2133 231 2185
rect 283 2177 476 2185
rect 283 2154 528 2177
rect 283 2136 476 2154
rect 613 2309 663 2310
tri 1109 2309 1110 2310 se
rect 1110 2309 1168 2310
rect 612 2273 664 2309
tri 1088 2288 1109 2309 se
rect 1109 2288 1168 2309
rect 1220 2288 1232 2340
rect 1284 2288 1296 2340
rect 1348 2288 1360 2340
rect 1412 2288 1424 2340
rect 1476 2288 1695 2340
rect 613 2272 663 2273
rect 612 2265 664 2271
rect 695 2282 1695 2288
rect 695 2248 749 2282
rect 783 2248 832 2282
rect 866 2248 915 2282
rect 949 2248 998 2282
rect 1032 2248 1081 2282
rect 1115 2248 1168 2282
rect 695 2242 1168 2248
tri 1168 2242 1208 2282 nw
rect 612 2208 664 2213
tri 664 2208 689 2233 sw
rect 612 2199 1691 2208
rect 664 2147 1691 2199
rect 612 2141 1691 2147
rect 283 2133 315 2136
rect 225 2102 237 2133
rect 271 2102 315 2133
rect 349 2102 394 2136
rect 428 2102 473 2136
rect 225 2096 528 2102
rect -112 2062 1737 2068
rect -112 2034 1685 2062
tri 1660 2009 1685 2034 ne
rect -196 2000 1648 2006
rect -196 1972 1596 2000
tri 1571 1947 1596 1972 ne
rect -280 1929 1568 1935
rect -354 1895 -308 1907
rect -354 1861 -348 1895
rect -314 1861 -308 1895
rect -354 1819 -308 1861
rect -354 1785 -348 1819
rect -314 1785 -308 1819
rect -228 1901 1516 1929
rect -280 1865 -228 1877
tri -228 1876 -203 1901 nw
tri 1491 1876 1516 1901 ne
rect -280 1807 -228 1813
rect 161 1872 528 1873
rect 161 1867 209 1872
rect 261 1867 289 1872
rect 341 1867 528 1872
rect 161 1833 173 1867
rect 207 1833 209 1867
rect 282 1833 289 1867
rect 357 1833 398 1867
rect 432 1833 473 1867
rect 161 1820 209 1833
rect 261 1820 289 1833
rect 341 1820 476 1833
rect 161 1815 476 1820
rect 161 1808 528 1815
rect -354 1742 -308 1785
rect 161 1795 209 1808
rect 261 1795 289 1808
rect 341 1803 528 1808
rect 341 1795 476 1803
rect 161 1761 173 1795
rect 207 1761 209 1795
rect 282 1761 289 1795
rect 357 1761 398 1795
rect 432 1761 473 1795
rect 692 1858 1488 1864
rect 744 1806 1180 1858
rect 1232 1806 1244 1858
rect 1296 1806 1308 1858
rect 1360 1806 1372 1858
rect 1424 1806 1436 1858
rect 692 1792 1488 1806
rect 1516 1863 1568 1877
rect 1516 1805 1568 1811
rect 1596 1934 1648 1948
rect 1685 1996 1737 2010
rect 1685 1938 1737 1944
rect 744 1774 1180 1792
rect 161 1756 209 1761
rect 261 1756 289 1761
rect 341 1756 476 1761
rect 161 1755 476 1756
tri 466 1745 476 1755 ne
rect 476 1745 528 1751
rect 612 1760 664 1766
rect -354 1708 -348 1742
rect -314 1708 -308 1742
rect 397 1709 443 1721
rect -354 1665 -308 1708
rect -354 1631 -348 1665
rect -314 1631 -308 1665
rect 145 1701 347 1708
rect -354 1619 -308 1631
rect -280 1657 -228 1663
tri -283 1603 -280 1606 se
rect -280 1603 -228 1605
tri -305 1581 -283 1603 se
rect -283 1593 -228 1603
rect -283 1581 -280 1593
rect -323 1541 -280 1581
rect -323 1535 -228 1541
rect 197 1699 347 1701
rect 197 1649 209 1699
rect 145 1647 209 1649
rect 261 1647 289 1699
rect 341 1647 347 1699
rect 145 1635 347 1647
rect 145 1629 209 1635
rect 197 1583 209 1629
rect 261 1583 289 1635
rect 341 1583 347 1635
rect 397 1675 403 1709
rect 437 1702 443 1709
tri 443 1702 450 1709 sw
tri 605 1702 612 1709 se
rect 747 1740 795 1774
rect 829 1740 877 1774
rect 911 1740 959 1774
rect 993 1740 1041 1774
rect 1075 1740 1180 1774
rect 1232 1740 1244 1792
rect 1296 1740 1308 1792
rect 1360 1740 1372 1792
rect 1424 1740 1436 1792
rect 692 1736 1488 1740
rect 692 1734 1171 1736
tri 1130 1709 1155 1734 ne
rect 1155 1728 1171 1734
rect 1205 1734 1488 1736
rect 1205 1728 1220 1734
rect 1155 1709 1168 1728
rect 612 1702 664 1708
tri 664 1702 671 1709 sw
tri 1155 1702 1162 1709 ne
rect 1162 1702 1168 1709
rect 437 1684 450 1702
tri 450 1684 468 1702 sw
tri 587 1684 605 1702 se
rect 605 1696 671 1702
rect 605 1684 612 1696
rect 437 1675 612 1684
rect 397 1644 612 1675
rect 664 1684 671 1696
tri 671 1684 689 1702 sw
tri 1162 1699 1165 1702 ne
rect 664 1678 829 1684
rect 664 1644 711 1678
rect 745 1644 783 1678
rect 817 1644 829 1678
rect 397 1638 829 1644
rect 1165 1676 1168 1702
tri 1220 1699 1255 1734 nw
rect 1165 1659 1220 1676
rect 397 1637 448 1638
rect 397 1603 403 1637
rect 437 1618 448 1637
tri 448 1618 468 1638 nw
tri 862 1618 879 1635 se
rect 437 1603 443 1618
tri 443 1613 448 1618 nw
tri 857 1613 862 1618 se
rect 862 1613 879 1618
tri 854 1610 857 1613 se
rect 857 1610 879 1613
rect 397 1590 443 1603
tri 483 1590 503 1610 se
rect 503 1590 1081 1610
tri 476 1583 483 1590 se
rect 483 1583 1081 1590
rect 197 1577 207 1583
rect 145 1568 207 1577
tri 207 1568 222 1583 nw
tri 461 1568 476 1583 se
rect 476 1582 1081 1583
rect 1165 1607 1168 1659
rect 1165 1590 1220 1607
rect 476 1568 529 1582
tri 529 1568 543 1582 nw
rect 145 1557 197 1568
tri 197 1558 207 1568 nw
tri 451 1558 461 1568 se
rect 461 1558 516 1568
rect -354 1495 -308 1507
rect -354 1461 -348 1495
rect -314 1461 -308 1495
rect -354 1415 -308 1461
rect -354 1381 -348 1415
rect -314 1381 -308 1415
rect -354 1369 -308 1381
tri 448 1555 451 1558 se
rect 451 1555 516 1558
tri 516 1555 529 1568 nw
rect 234 1549 495 1555
rect 234 1515 246 1549
rect 280 1515 318 1549
rect 352 1548 495 1549
rect 352 1515 393 1548
rect 234 1509 393 1515
tri 367 1506 370 1509 ne
rect 370 1506 393 1509
rect 145 1485 197 1505
tri 197 1484 219 1506 sw
tri 370 1484 392 1506 ne
rect 392 1496 393 1506
rect 445 1534 495 1548
tri 495 1534 516 1555 nw
rect 556 1548 608 1554
rect 392 1484 445 1496
tri 445 1484 495 1534 nw
tri 534 1484 556 1506 se
rect 1165 1538 1168 1590
rect 1165 1534 1171 1538
rect 1205 1534 1220 1538
rect 1165 1521 1220 1534
rect 556 1484 608 1496
tri 608 1484 630 1506 sw
rect 197 1481 219 1484
tri 219 1481 222 1484 sw
tri 392 1483 393 1484 ne
rect 393 1481 445 1484
rect 197 1433 214 1481
rect 145 1429 214 1433
rect 266 1429 289 1481
rect 341 1429 347 1481
rect 145 1417 347 1429
rect 393 1423 445 1429
tri 531 1481 534 1484 se
rect 534 1481 556 1484
rect 531 1475 556 1481
rect 608 1481 630 1484
tri 630 1481 633 1484 sw
rect 608 1475 662 1481
rect 531 1441 543 1475
rect 608 1441 615 1475
rect 649 1441 662 1475
rect 1165 1469 1168 1521
rect 1165 1452 1171 1469
rect 1205 1452 1220 1469
rect 531 1432 556 1441
rect 608 1432 662 1441
rect 531 1426 662 1432
rect 692 1424 750 1430
rect 145 1413 214 1417
tri 137 1358 145 1366 se
rect 197 1365 214 1413
rect 266 1365 289 1417
rect 341 1365 347 1417
rect 197 1361 215 1365
rect 145 1358 215 1361
tri 215 1358 222 1365 nw
tri 120 1341 137 1358 se
rect 137 1341 197 1358
rect -797 1335 145 1341
rect -797 1283 -95 1335
rect -43 1283 -31 1335
rect 21 1289 145 1335
tri 197 1340 215 1358 nw
rect 476 1346 482 1398
rect 534 1392 606 1398
rect 534 1358 560 1392
rect 594 1358 606 1392
rect 744 1372 750 1424
rect 851 1395 857 1447
rect 909 1395 940 1447
rect 992 1395 1023 1447
rect 1075 1395 1081 1447
rect 1165 1400 1168 1452
rect 692 1366 750 1372
rect 1165 1383 1171 1400
rect 1205 1383 1220 1400
rect 534 1346 606 1358
rect 21 1283 197 1289
rect 229 1326 450 1332
tri 450 1326 456 1332 sw
tri 628 1326 634 1332 se
rect 634 1326 1083 1332
rect 229 1292 241 1326
rect 275 1292 313 1326
rect 347 1318 456 1326
tri 456 1318 464 1326 sw
tri 620 1318 628 1326 se
rect 628 1318 879 1326
rect 347 1311 879 1318
rect 347 1292 612 1311
rect 229 1286 612 1292
tri 587 1283 590 1286 ne
rect 590 1283 612 1286
rect -797 1269 197 1283
tri 590 1274 599 1283 ne
rect 599 1274 612 1283
rect -797 1266 145 1269
rect -797 1214 -95 1266
rect -43 1214 -31 1266
rect 21 1217 145 1266
tri 197 1249 222 1274 sw
tri 599 1261 612 1274 ne
rect 664 1292 879 1311
rect 913 1292 951 1326
rect 985 1292 1023 1326
rect 1057 1292 1083 1326
rect 664 1286 1083 1292
rect 1165 1331 1168 1383
rect 1165 1317 1220 1331
rect 1165 1314 1171 1317
rect 1205 1314 1220 1317
rect 664 1283 686 1286
tri 686 1283 689 1286 nw
tri 664 1261 686 1283 nw
rect 1165 1262 1168 1314
rect 1596 1333 1648 1882
tri 1648 1333 1673 1358 sw
rect 1596 1287 1695 1333
rect 197 1226 347 1249
rect 197 1217 229 1226
rect 21 1214 157 1217
rect -797 1197 157 1214
rect 191 1197 229 1217
rect 263 1197 301 1226
rect -797 1145 -95 1197
rect -43 1145 -31 1197
rect 21 1145 145 1197
rect 197 1145 210 1197
rect 263 1192 274 1197
rect 335 1192 347 1226
rect 262 1145 274 1192
rect 326 1145 347 1192
rect -797 1139 347 1145
rect 381 1206 387 1258
rect 439 1234 445 1258
rect 612 1246 664 1259
tri 445 1234 453 1242 sw
rect 439 1231 453 1234
tri 453 1231 456 1234 sw
rect 439 1217 456 1231
tri 456 1217 470 1231 sw
rect 439 1211 524 1217
rect 381 1194 405 1206
rect 381 1142 387 1194
rect 439 1177 477 1211
rect 511 1177 524 1211
rect 1165 1246 1220 1262
rect 612 1188 664 1194
rect 851 1188 857 1240
rect 909 1231 940 1240
rect 992 1231 1023 1240
rect 909 1197 939 1231
rect 992 1197 1011 1231
rect 909 1188 940 1197
rect 992 1188 1023 1197
rect 1075 1188 1081 1240
rect 1165 1194 1168 1246
rect 1165 1188 1220 1194
rect 439 1171 524 1177
rect 439 1142 445 1171
tri 445 1146 470 1171 nw
rect 476 1131 528 1137
rect -354 1099 -308 1111
rect -354 1065 -348 1099
rect -314 1065 -308 1099
rect -354 1018 -308 1065
rect -354 984 -348 1018
rect -314 984 -308 1018
rect -354 972 -308 984
rect 4 1098 428 1104
rect 4 1064 169 1098
rect 203 1064 241 1098
rect 275 1064 428 1098
rect 476 1073 528 1079
rect 568 1132 1695 1160
rect 4 1058 428 1064
rect 4 1056 75 1058
tri 75 1056 77 1058 nw
tri 359 1056 361 1058 ne
rect 361 1056 428 1058
tri -21 944 4 969 se
rect 4 944 52 1056
tri 52 1033 75 1056 nw
tri 361 1033 384 1056 ne
rect -33 904 52 944
rect 89 984 145 1030
rect 89 978 136 984
tri 136 978 142 984 nw
rect 89 858 117 978
tri 117 959 136 978 nw
tri 380 959 384 963 se
rect 384 959 428 1056
tri 543 1018 568 1043 se
rect 568 1018 596 1132
tri 596 1107 621 1132 nw
rect 692 1098 744 1104
tri 596 1018 621 1043 sw
rect 692 1040 744 1046
rect 783 1098 1081 1104
rect 783 1064 877 1098
rect 911 1064 949 1098
rect 983 1064 1021 1098
rect 1055 1064 1081 1098
rect 783 1058 1081 1064
rect 1165 1098 1220 1104
rect 527 1012 658 1018
rect 527 978 539 1012
rect 573 978 611 1012
rect 645 978 658 1012
rect 527 972 658 978
tri 359 938 380 959 se
rect 380 938 428 959
tri 428 938 453 963 sw
tri 758 938 783 963 se
rect 783 938 836 1058
tri 836 1033 861 1058 nw
rect 1165 1046 1168 1098
rect 1081 984 1137 1030
tri 1084 980 1088 984 ne
rect 1088 980 1137 984
tri 1088 963 1105 980 ne
rect 1105 963 1137 980
tri 836 938 861 963 sw
tri 1105 959 1109 963 ne
rect 347 892 879 938
tri 117 858 130 871 sw
tri 1102 864 1109 871 se
rect 1109 864 1137 963
rect 476 858 528 864
rect 89 852 130 858
tri 130 852 136 858 sw
rect 89 846 136 852
tri 136 846 142 852 sw
rect 89 800 145 846
rect 89 787 129 800
tri 129 787 142 800 nw
rect 393 793 445 799
rect 89 674 117 787
tri 117 775 129 787 nw
rect 145 705 151 757
rect 203 705 220 757
rect 272 705 289 757
rect 341 705 347 757
rect 393 717 445 741
tri 117 674 130 687 sw
rect 89 662 130 674
tri 130 662 142 674 sw
rect 89 616 145 662
rect 393 641 445 665
rect 89 596 122 616
tri 122 596 142 616 nw
rect 89 499 117 596
tri 117 591 122 596 nw
rect 145 521 151 573
rect 203 521 220 573
rect 272 521 289 573
rect 341 521 347 573
rect 393 564 445 589
rect 393 506 445 512
rect 476 791 528 806
rect 476 738 485 739
rect 519 738 528 739
rect 476 724 528 738
rect 689 858 747 864
tri 1096 858 1102 864 se
rect 1102 858 1137 864
rect 689 806 692 858
rect 744 806 747 858
tri 1084 846 1096 858 se
rect 1096 846 1137 858
rect 689 794 747 806
rect 1081 800 1137 846
rect 689 742 692 794
rect 744 742 747 794
tri 1084 780 1104 800 ne
rect 1104 780 1137 800
tri 1104 775 1109 780 ne
rect 689 736 747 742
rect 476 658 485 672
rect 519 658 528 672
rect 476 657 528 658
rect 476 590 485 605
rect 519 590 528 605
rect 612 702 823 708
rect 851 705 857 757
rect 909 705 940 757
rect 992 705 1023 757
rect 1075 705 1081 757
rect 664 696 823 702
rect 664 662 783 696
rect 817 662 823 696
tri 1090 668 1109 687 se
rect 1109 668 1137 780
tri 1084 662 1090 668 se
rect 1090 662 1137 668
rect 664 656 823 662
rect 612 637 664 650
tri 664 631 689 656 nw
tri 752 631 777 656 ne
rect 612 579 664 585
rect 692 610 744 616
rect 476 533 528 538
rect 476 523 485 533
rect 519 523 528 533
tri 117 499 121 503 sw
rect 89 495 121 499
tri 121 495 125 499 sw
rect 89 488 125 495
tri 125 488 132 495 sw
rect 89 478 132 488
tri 132 478 142 488 sw
rect 89 432 145 478
rect 347 432 403 478
tri 350 420 362 432 ne
rect 362 420 403 432
tri 362 407 375 420 ne
rect -354 384 -308 396
rect -354 350 -348 384
rect -314 350 -308 384
rect -354 244 -308 350
rect -256 332 47 386
rect 48 333 49 385
rect 85 333 86 385
rect 87 384 347 386
rect 87 332 151 384
rect 203 332 220 384
rect 272 332 289 384
rect 341 332 347 384
rect -198 326 31 332
rect -198 292 -172 326
rect -138 292 -100 326
rect -66 292 -28 326
rect 6 316 31 326
tri 31 316 47 332 nw
tri 372 316 375 319 se
rect 375 316 403 420
rect 6 309 24 316
tri 24 309 31 316 nw
tri 365 309 372 316 se
rect 372 309 403 316
rect 6 292 22 309
tri 22 307 24 309 nw
tri 363 307 365 309 se
rect 365 307 403 309
tri 362 306 363 307 se
rect 363 306 403 307
tri 352 296 362 306 se
rect 362 296 403 306
tri 350 294 352 296 se
rect 352 294 403 296
rect -198 286 22 292
rect 347 248 403 294
rect 476 456 528 471
rect 476 389 528 404
rect 476 322 528 337
rect 476 262 485 270
rect 519 262 528 270
rect 476 256 528 262
rect -354 210 -348 244
rect -314 210 -308 244
tri -366 196 -354 208 se
rect -354 196 -308 210
tri -308 196 -296 208 sw
tri 464 196 476 208 se
rect 476 196 528 204
tri -370 192 -366 196 se
rect -366 192 -296 196
tri -296 192 -292 196 sw
tri 460 192 464 196 se
rect 464 192 528 196
tri -379 183 -370 192 se
rect -370 183 -292 192
tri -292 183 -283 192 sw
tri 451 183 460 192 se
rect 460 190 528 192
rect 460 183 476 190
rect -487 172 -106 183
rect -54 172 -21 183
rect 31 172 151 183
rect 203 172 220 183
rect -487 138 -461 172
rect -427 138 -386 172
rect -352 138 -311 172
rect -277 138 -236 172
rect -202 138 -161 172
rect -127 138 -106 172
rect -51 138 -21 172
rect 31 138 67 172
rect 101 138 143 172
rect 203 138 219 172
rect -487 131 -106 138
rect -54 131 -21 138
rect 31 131 151 138
rect 203 131 220 138
rect 272 131 289 183
rect 341 172 476 183
rect 341 138 371 172
rect 405 138 447 172
rect 692 543 744 558
rect 692 476 744 491
rect 692 420 701 424
rect 735 420 744 424
rect 692 409 744 420
rect 692 346 701 357
rect 735 346 744 357
rect 692 342 744 346
rect 777 609 823 656
rect 1081 616 1137 662
rect 777 575 783 609
rect 817 575 823 609
tri 1084 591 1109 616 ne
rect 777 522 823 575
rect 777 488 783 522
rect 817 488 823 522
rect 851 521 857 573
rect 909 521 940 573
rect 992 521 1023 573
rect 1075 521 1081 573
rect 777 436 823 488
tri 1084 478 1109 503 se
rect 1109 478 1137 616
rect 777 402 783 436
rect 817 402 823 436
rect 1081 432 1137 478
tri 1084 407 1109 432 ne
rect 777 350 823 402
rect 777 316 783 350
rect 817 316 823 350
rect 851 337 857 389
rect 909 337 940 389
rect 992 337 1023 389
rect 1075 337 1081 389
rect 777 304 823 316
tri 1099 309 1109 319 se
rect 1109 309 1137 432
tri 1094 304 1099 309 se
rect 1099 304 1137 309
tri 1084 294 1094 304 se
rect 1094 294 1137 304
rect 692 276 701 290
rect 735 276 744 290
rect 1081 248 1137 294
rect 1165 1029 1220 1046
rect 1165 977 1168 1029
rect 1165 960 1220 977
rect 1165 908 1168 960
rect 1165 902 1171 908
rect 1205 902 1220 908
rect 1165 891 1220 902
rect 1165 839 1168 891
rect 1165 824 1171 839
rect 1205 824 1220 839
rect 1165 822 1220 824
rect 1165 770 1168 822
rect 1165 754 1171 770
rect 1205 754 1220 770
rect 1165 702 1168 754
rect 1165 686 1171 702
rect 1205 686 1220 702
rect 1165 634 1168 686
rect 1165 624 1220 634
rect 1165 618 1171 624
rect 1205 618 1220 624
rect 1165 566 1168 618
rect 1165 550 1220 566
rect 1165 498 1168 550
rect 1165 482 1220 498
rect 1165 430 1168 482
rect 1165 414 1220 430
rect 1165 362 1168 414
rect 1165 354 1171 362
rect 1205 354 1220 362
rect 1165 346 1220 354
rect 1165 294 1168 346
rect 1165 278 1171 294
rect 1205 278 1220 294
rect 692 210 744 224
rect 1165 226 1168 278
tri 744 198 769 223 sw
tri 1140 198 1165 223 se
rect 1165 210 1171 226
rect 1205 210 1220 226
rect 1165 198 1168 210
rect 744 192 1168 198
rect 773 158 817 192
rect 851 158 895 192
rect 929 158 973 192
rect 1007 158 1051 192
rect 1085 158 1168 192
rect 692 152 1220 158
rect 341 131 528 138
<< rmetal1 >>
rect 393 5651 445 5652
rect 393 5650 394 5651
rect 444 5650 445 5651
rect 393 5613 394 5614
rect 444 5613 445 5614
rect 393 5612 445 5613
rect 393 5219 445 5220
rect 393 5218 394 5219
rect 444 5218 445 5219
rect 393 5181 394 5182
rect 444 5181 445 5182
rect 393 5180 445 5181
rect 142 5153 144 5154
rect 142 5109 143 5153
rect 142 5108 144 5109
rect 180 5153 182 5154
rect 181 5109 182 5153
rect 180 5108 182 5109
rect 65 4346 117 4347
rect 65 4345 66 4346
rect 116 4345 117 4346
rect 65 4308 66 4309
rect 116 4308 117 4309
rect 65 4307 117 4308
rect 207 4340 253 4341
rect 207 4339 208 4340
rect 252 4339 253 4340
rect 207 4302 208 4303
rect 252 4302 253 4303
rect 207 4301 253 4302
rect 777 4338 823 4339
rect 777 4337 778 4338
rect 822 4337 823 4338
rect 612 4314 664 4315
rect 612 4313 613 4314
rect 663 4313 664 4314
rect 142 4275 144 4276
rect 180 4275 182 4276
rect 142 4225 143 4275
rect 181 4225 182 4275
rect 777 4300 778 4301
rect 822 4300 823 4301
rect 777 4299 823 4300
rect 612 4276 613 4277
rect 663 4276 664 4277
rect 612 4275 664 4276
rect 871 4249 873 4250
rect 909 4249 911 4250
rect 142 4224 144 4225
rect 180 4224 182 4225
rect 871 4205 872 4249
rect 910 4205 911 4249
rect 871 4204 873 4205
rect 909 4204 911 4205
rect 142 4139 144 4140
rect 142 4095 143 4139
rect 142 4094 144 4095
rect 180 4139 182 4140
rect 181 4095 182 4139
rect 180 4094 182 4095
rect 612 4068 664 4069
rect 612 4067 613 4068
rect 663 4067 664 4068
rect 65 3693 117 3694
rect 65 3692 66 3693
rect 116 3692 117 3693
rect 612 4030 613 4031
rect 663 4030 664 4031
rect 612 4029 664 4030
rect 612 3693 664 3694
rect 612 3692 613 3693
rect 663 3692 664 3693
rect 65 3655 66 3656
rect 116 3655 117 3656
rect 65 3654 117 3655
rect 612 3655 613 3656
rect 663 3655 664 3656
rect 612 3654 664 3655
rect 65 3445 117 3446
rect 65 3444 66 3445
rect 116 3444 117 3445
rect 65 3407 66 3408
rect 116 3407 117 3408
rect 65 3406 117 3407
rect 65 3071 117 3072
rect 65 3070 66 3071
rect 116 3070 117 3071
rect 612 3445 664 3446
rect 612 3444 613 3445
rect 663 3444 664 3445
rect 612 3407 613 3408
rect 663 3407 664 3408
rect 612 3406 664 3407
rect 612 3071 664 3072
rect 612 3070 613 3071
rect 663 3070 664 3071
rect 65 3033 66 3034
rect 116 3033 117 3034
rect 65 3032 117 3033
rect 612 3033 613 3034
rect 663 3033 664 3034
rect 612 3032 664 3033
rect 65 2823 117 2824
rect 65 2822 66 2823
rect 116 2822 117 2823
rect 65 2785 66 2786
rect 116 2785 117 2786
rect 65 2784 117 2785
rect 65 2449 117 2450
rect 65 2448 66 2449
rect 116 2448 117 2449
rect 612 2822 664 2823
rect 612 2821 613 2822
rect 663 2821 664 2822
rect 612 2784 613 2785
rect 663 2784 664 2785
rect 612 2783 664 2784
rect 65 2411 66 2412
rect 116 2411 117 2412
rect 65 2410 117 2411
rect 612 2310 664 2311
rect 612 2309 613 2310
rect 663 2309 664 2310
rect 612 2272 613 2273
rect 663 2272 664 2273
rect 612 2271 664 2272
rect 47 385 49 386
rect 47 333 48 385
rect 47 332 49 333
rect 85 385 87 386
rect 86 333 87 385
rect 85 332 87 333
<< via1 >>
rect 1522 8505 1574 8557
rect 1592 8505 1644 8557
rect 1662 8505 1714 8557
rect 1732 8505 1784 8557
rect 1803 8505 1855 8557
rect 1522 8441 1574 8493
rect 1592 8441 1644 8493
rect 1662 8441 1714 8493
rect 1732 8441 1784 8493
rect 1803 8441 1855 8493
rect 1522 8377 1574 8429
rect 1592 8377 1644 8429
rect 1662 8377 1714 8429
rect 1732 8377 1784 8429
rect 1803 8377 1855 8429
rect 350 8205 402 8257
rect 420 8205 472 8257
rect 489 8205 541 8257
rect 553 8077 669 8257
rect 1522 8205 1574 8257
rect 1592 8205 1644 8257
rect 1662 8205 1714 8257
rect 1732 8205 1784 8257
rect 1803 8205 1855 8257
rect 2789 8205 2841 8257
rect 2859 8205 2911 8257
rect 2930 8205 2982 8257
rect 3001 8205 3053 8257
rect 1522 8141 1574 8193
rect 1592 8141 1644 8193
rect 1662 8141 1714 8193
rect 1732 8141 1784 8193
rect 1803 8141 1855 8193
rect 2789 8141 2841 8193
rect 2859 8141 2911 8193
rect 2930 8141 2982 8193
rect 3001 8141 3053 8193
rect 1522 8077 1574 8129
rect 1592 8077 1644 8129
rect 1662 8077 1714 8129
rect 1732 8077 1784 8129
rect 1803 8077 1855 8129
rect 2789 8077 2841 8129
rect 2859 8077 2911 8129
rect 2930 8077 2982 8129
rect 3001 8077 3053 8129
rect 3387 8077 3567 8257
rect 4503 8205 4555 8257
rect 4568 8205 4620 8257
rect 4633 8205 4685 8257
rect 4698 8205 4750 8257
rect 4763 8205 4815 8257
rect 4829 8205 4881 8257
rect 4895 8205 4947 8257
rect 4961 8205 5013 8257
rect 5027 8205 5079 8257
rect 5093 8205 5145 8257
rect 5159 8205 5211 8257
rect 4503 8141 4555 8193
rect 4568 8141 4620 8193
rect 4633 8141 4685 8193
rect 4698 8141 4750 8193
rect 4763 8141 4815 8193
rect 4829 8141 4881 8193
rect 4895 8141 4947 8193
rect 4961 8141 5013 8193
rect 5027 8141 5079 8193
rect 5093 8141 5145 8193
rect 5159 8141 5211 8193
rect 4503 8077 4555 8129
rect 4568 8077 4620 8129
rect 4633 8077 4685 8129
rect 4698 8077 4750 8129
rect 4763 8077 4815 8129
rect 4829 8077 4881 8129
rect 4895 8077 4947 8129
rect 4961 8077 5013 8129
rect 5027 8077 5079 8129
rect 5093 8077 5145 8129
rect 5159 8077 5211 8129
rect 388 7935 440 7987
rect 489 7975 541 7987
rect 489 7941 493 7975
rect 493 7941 527 7975
rect 527 7941 541 7975
rect 489 7935 541 7941
rect 3445 7942 3497 7951
rect 3515 7942 3567 7951
rect 2010 7922 2062 7931
rect 2083 7922 2135 7931
rect 2156 7922 2208 7931
rect 2229 7922 2281 7931
rect 2302 7922 2354 7931
rect 2374 7922 2426 7931
rect 2446 7922 2498 7931
rect 2010 7888 2037 7922
rect 2037 7888 2062 7922
rect 2083 7888 2109 7922
rect 2109 7888 2135 7922
rect 2156 7888 2181 7922
rect 2181 7888 2208 7922
rect 2229 7888 2253 7922
rect 2253 7888 2281 7922
rect 2302 7888 2325 7922
rect 2325 7888 2354 7922
rect 2374 7888 2397 7922
rect 2397 7888 2426 7922
rect 2446 7888 2469 7922
rect 2469 7888 2498 7922
rect 2010 7879 2062 7888
rect 2083 7879 2135 7888
rect 2156 7879 2208 7888
rect 2229 7879 2281 7888
rect 2302 7879 2354 7888
rect 2374 7879 2426 7888
rect 2446 7879 2498 7888
rect 1854 7784 1906 7836
rect 1918 7784 1970 7836
rect 1602 7704 1654 7756
rect 1669 7704 1721 7756
rect 2010 7607 2062 7659
rect 2083 7607 2135 7659
rect 2156 7607 2208 7659
rect 2229 7607 2281 7659
rect 2302 7607 2354 7659
rect 2374 7607 2426 7659
rect 2446 7607 2498 7659
rect 3007 7908 3057 7912
rect 3057 7908 3059 7912
rect 3445 7908 3471 7942
rect 3471 7908 3497 7942
rect 3515 7908 3547 7942
rect 3547 7908 3567 7942
rect 3007 7860 3059 7908
rect 3445 7899 3497 7908
rect 3515 7899 3567 7908
rect 3007 7807 3059 7846
rect 3007 7794 3019 7807
rect 3019 7794 3053 7807
rect 3053 7794 3059 7807
rect 3007 7773 3019 7780
rect 3019 7773 3053 7780
rect 3053 7773 3059 7780
rect 3007 7728 3059 7773
rect 3007 7688 3019 7714
rect 3019 7688 3053 7714
rect 3053 7688 3059 7714
rect 3007 7662 3059 7688
rect 3007 7637 3059 7649
rect 3007 7603 3019 7637
rect 3019 7603 3053 7637
rect 3053 7603 3059 7637
rect 3097 7607 3149 7659
rect 3161 7607 3213 7659
rect 3225 7607 3277 7659
rect 3289 7607 3341 7659
rect 3353 7607 3405 7659
rect 3007 7597 3059 7603
rect 350 7444 402 7496
rect 428 7444 480 7496
rect 507 7484 559 7496
rect 507 7450 527 7484
rect 527 7450 559 7484
rect 507 7444 559 7450
rect 350 7380 402 7432
rect 428 7380 480 7432
rect 507 7412 559 7432
rect 507 7380 527 7412
rect 527 7380 559 7412
rect 1691 7511 1743 7563
rect 1758 7511 1810 7563
rect 1854 7431 1906 7483
rect 1918 7431 1970 7483
rect 2937 7466 2989 7475
rect 2937 7432 2941 7466
rect 2941 7432 2975 7466
rect 2975 7432 2989 7466
rect 2937 7423 2989 7432
rect 3001 7466 3053 7475
rect 3001 7432 3013 7466
rect 3013 7432 3047 7466
rect 3047 7432 3053 7466
rect 3001 7423 3053 7432
rect 612 7306 664 7358
rect 3607 7335 3659 7387
rect 3671 7335 3723 7387
rect 612 7239 664 7291
rect 2010 7255 2062 7307
rect 2083 7255 2135 7307
rect 2156 7255 2208 7307
rect 2229 7255 2281 7307
rect 2302 7255 2354 7307
rect 2374 7255 2426 7307
rect 2446 7255 2498 7307
rect 692 7125 744 7177
rect 2567 7165 2619 7217
rect 2631 7165 2683 7217
rect 692 7058 744 7110
rect 1854 7079 1906 7131
rect 1918 7079 1970 7131
rect 3097 7255 3149 7307
rect 3174 7255 3226 7307
rect 3251 7255 3303 7307
rect 3328 7255 3380 7307
rect 3411 7165 3463 7217
rect 3514 7165 3566 7217
rect 44 6838 96 6876
rect 44 6824 53 6838
rect 53 6824 87 6838
rect 87 6824 96 6838
rect 44 6763 96 6775
rect 44 6729 53 6763
rect 53 6729 87 6763
rect 87 6729 96 6763
rect 44 6723 96 6729
rect 151 6717 203 6769
rect 220 6717 272 6769
rect 289 6717 341 6769
rect 612 6835 664 6887
rect 612 6768 664 6820
rect 1516 6894 1568 6946
rect 1516 6827 1568 6879
rect 44 6607 96 6613
rect -119 6419 -67 6471
rect -119 6355 -67 6407
rect 44 6573 53 6607
rect 53 6573 87 6607
rect 87 6573 96 6607
rect 1854 6727 1906 6779
rect 1918 6727 1970 6779
rect 3163 6826 3215 6878
rect 3233 6826 3285 6878
rect 3303 6826 3355 6878
rect 3373 6826 3425 6878
rect 556 6667 608 6719
rect 556 6600 608 6652
rect 2010 6637 2062 6643
rect 2083 6637 2135 6643
rect 2156 6637 2208 6643
rect 2229 6637 2281 6643
rect 2302 6637 2354 6643
rect 2374 6637 2426 6643
rect 2010 6603 2026 6637
rect 2026 6603 2062 6637
rect 2083 6603 2102 6637
rect 2102 6603 2135 6637
rect 2156 6603 2178 6637
rect 2178 6603 2208 6637
rect 2229 6603 2254 6637
rect 2254 6603 2281 6637
rect 2302 6603 2330 6637
rect 2330 6603 2354 6637
rect 2374 6603 2406 6637
rect 2406 6603 2426 6637
rect 44 6561 96 6573
rect 44 6527 96 6544
rect 44 6493 53 6527
rect 53 6493 87 6527
rect 87 6493 96 6527
rect 44 6492 96 6493
rect 612 6490 664 6542
rect 44 6447 96 6475
rect 44 6423 53 6447
rect 53 6423 87 6447
rect 87 6423 96 6447
rect 44 6368 96 6406
rect 151 6405 203 6457
rect 220 6405 272 6457
rect 289 6405 341 6457
rect 612 6423 664 6475
rect 44 6354 53 6368
rect 53 6354 87 6368
rect 87 6354 96 6368
rect 2010 6591 2062 6603
rect 2083 6591 2135 6603
rect 2156 6591 2208 6603
rect 2229 6591 2281 6603
rect 2302 6591 2354 6603
rect 2374 6591 2426 6603
rect 2446 6637 2498 6643
rect 2446 6603 2448 6637
rect 2448 6603 2482 6637
rect 2482 6603 2498 6637
rect 2446 6591 2498 6603
rect 3163 6637 3215 6643
rect 3233 6637 3285 6643
rect 3303 6637 3355 6643
rect 3373 6637 3425 6643
rect 3163 6603 3182 6637
rect 3182 6603 3215 6637
rect 3233 6603 3255 6637
rect 3255 6603 3285 6637
rect 3303 6603 3328 6637
rect 3328 6603 3355 6637
rect 3373 6603 3401 6637
rect 3401 6603 3425 6637
rect 3163 6591 3215 6603
rect 3233 6591 3285 6603
rect 3303 6591 3355 6603
rect 3373 6591 3425 6603
rect 1691 6511 1743 6563
rect 1758 6511 1810 6563
rect 4439 6511 4491 6563
rect 4503 6511 4555 6563
rect 44 6334 53 6337
rect 53 6334 87 6337
rect 87 6334 96 6337
rect 44 6289 96 6334
rect 44 6285 53 6289
rect 53 6285 87 6289
rect 87 6285 96 6289
rect 44 6255 53 6268
rect 53 6255 87 6268
rect 87 6255 96 6268
rect 44 6216 96 6255
rect 44 6176 53 6200
rect 53 6176 87 6200
rect 87 6176 96 6200
rect 44 6148 96 6176
rect 612 6235 664 6287
rect 476 6164 528 6216
rect 44 6131 96 6132
rect 612 6168 664 6220
rect 44 6097 53 6131
rect 53 6097 87 6131
rect 87 6097 96 6131
rect 44 6080 96 6097
rect 151 6079 203 6131
rect 220 6079 272 6131
rect 289 6079 341 6131
rect 44 6052 96 6064
rect 44 6018 53 6052
rect 53 6018 87 6052
rect 87 6018 96 6052
rect 44 6012 96 6018
rect 1178 6028 1230 6037
rect 1270 6028 1322 6037
rect 1178 5994 1201 6028
rect 1201 5994 1230 6028
rect 1270 5994 1277 6028
rect 1277 5994 1311 6028
rect 1311 5994 1322 6028
rect 1178 5985 1230 5994
rect 1270 5985 1322 5994
rect 1363 5990 1415 6037
rect 1363 5985 1395 5990
rect 1395 5985 1415 5990
rect 44 5900 96 5906
rect 44 5866 53 5900
rect 53 5866 87 5900
rect 87 5866 96 5900
rect 44 5854 96 5866
rect 692 5854 744 5906
rect 857 5873 909 5925
rect 940 5919 992 5925
rect 1023 5919 1075 5925
rect 940 5885 967 5919
rect 967 5885 992 5919
rect 1023 5885 1039 5919
rect 1039 5885 1075 5919
rect 940 5873 992 5885
rect 1023 5873 1075 5885
rect 1386 5910 1438 5944
rect 1386 5892 1395 5910
rect 1395 5892 1429 5910
rect 1429 5892 1438 5910
rect 1386 5876 1395 5877
rect 1395 5876 1429 5877
rect 1429 5876 1438 5877
rect 44 5822 96 5838
rect 44 5788 53 5822
rect 53 5788 87 5822
rect 87 5788 96 5822
rect 476 5826 528 5832
rect 44 5786 96 5788
rect 44 5744 96 5770
rect 151 5753 203 5805
rect 220 5753 272 5805
rect 289 5753 341 5805
rect 476 5792 485 5826
rect 485 5792 519 5826
rect 519 5792 528 5826
rect 44 5718 53 5744
rect 53 5718 87 5744
rect 87 5718 96 5744
rect 44 5667 96 5702
rect 44 5650 53 5667
rect 53 5650 87 5667
rect 87 5650 96 5667
rect 44 5633 53 5634
rect 53 5633 87 5634
rect 87 5633 96 5634
rect 44 5590 96 5633
rect 393 5726 445 5778
rect 393 5659 445 5711
rect 476 5780 528 5792
rect 692 5787 744 5839
rect 1386 5830 1438 5876
rect 1386 5825 1395 5830
rect 1395 5825 1429 5830
rect 1429 5825 1438 5830
rect 1386 5796 1395 5810
rect 1395 5796 1429 5810
rect 1429 5796 1438 5810
rect 476 5749 528 5757
rect 1386 5758 1438 5796
rect 476 5715 485 5749
rect 485 5715 519 5749
rect 519 5715 528 5749
rect 476 5705 528 5715
rect 476 5671 528 5683
rect 476 5637 485 5671
rect 485 5637 519 5671
rect 519 5637 528 5671
rect 476 5631 528 5637
rect 1386 5717 1395 5743
rect 1395 5717 1429 5743
rect 1429 5717 1438 5743
rect 1386 5691 1438 5717
rect 1386 5672 1438 5676
rect 1386 5638 1395 5672
rect 1395 5638 1429 5672
rect 1429 5638 1438 5672
rect 1386 5624 1438 5638
rect 1386 5593 1438 5609
rect 44 5582 53 5590
rect 53 5582 87 5590
rect 87 5582 96 5590
rect 44 5556 53 5566
rect 53 5556 87 5566
rect 87 5556 96 5566
rect 44 5514 96 5556
rect 1386 5559 1395 5593
rect 1395 5559 1429 5593
rect 1429 5559 1438 5593
rect 1386 5557 1438 5559
rect 44 5479 53 5498
rect 53 5479 87 5498
rect 87 5479 96 5498
rect 44 5446 96 5479
rect 44 5402 53 5430
rect 53 5402 87 5430
rect 87 5402 96 5430
rect 44 5378 96 5402
rect 476 5499 528 5505
rect 476 5465 485 5499
rect 485 5465 519 5499
rect 519 5465 528 5499
rect 476 5453 528 5465
rect 476 5414 528 5421
rect 476 5380 485 5414
rect 485 5380 519 5414
rect 519 5380 528 5414
rect 44 5359 96 5362
rect 44 5325 53 5359
rect 53 5325 87 5359
rect 87 5325 96 5359
rect 44 5310 96 5325
rect 151 5321 203 5373
rect 220 5321 272 5373
rect 289 5321 341 5373
rect 476 5369 528 5380
rect 44 5282 96 5294
rect 44 5248 53 5282
rect 53 5248 87 5282
rect 87 5248 96 5282
rect 44 5242 96 5248
rect 393 5293 445 5345
rect 393 5226 445 5278
rect 476 5329 528 5338
rect 476 5295 485 5329
rect 485 5295 519 5329
rect 519 5295 528 5329
rect 476 5286 528 5295
rect 476 5243 528 5255
rect 476 5209 485 5243
rect 485 5209 519 5243
rect 519 5209 528 5243
rect 476 5203 528 5209
rect 1386 5514 1438 5542
rect 1386 5490 1395 5514
rect 1395 5490 1429 5514
rect 1429 5490 1438 5514
rect 1386 5435 1438 5475
rect 1386 5423 1395 5435
rect 1395 5423 1429 5435
rect 1429 5423 1438 5435
rect 1386 5401 1395 5408
rect 1395 5401 1429 5408
rect 1429 5401 1438 5408
rect 1386 5356 1438 5401
rect 1217 5311 1269 5317
rect 1287 5311 1339 5317
rect 1386 5311 1438 5340
rect 1217 5277 1241 5311
rect 1241 5277 1269 5311
rect 1287 5277 1316 5311
rect 1316 5277 1339 5311
rect 1386 5288 1391 5311
rect 1391 5288 1438 5311
rect 1217 5265 1269 5277
rect 1287 5265 1339 5277
rect 65 5096 117 5148
rect 692 5105 744 5157
rect 692 5040 744 5092
rect 65 4975 117 5027
rect -106 4846 -54 4898
rect -21 4846 31 4898
rect 151 4889 203 4941
rect 220 4889 272 4941
rect 289 4889 341 4941
rect 692 4883 744 4935
rect 612 4823 664 4875
rect 612 4756 664 4808
rect 1174 4825 1482 4941
rect 692 4778 739 4808
rect 739 4778 744 4808
rect 692 4756 744 4778
rect 1168 4760 1220 4812
rect 1168 4695 1220 4747
rect 1168 4630 1220 4682
rect 151 4546 203 4558
rect -34 4490 18 4542
rect 151 4512 157 4546
rect 157 4512 191 4546
rect 191 4512 203 4546
rect 151 4506 203 4512
rect 220 4546 272 4558
rect 220 4512 255 4546
rect 255 4512 272 4546
rect 220 4506 272 4512
rect 289 4506 341 4558
rect 476 4557 528 4568
rect 476 4523 485 4557
rect 485 4523 519 4557
rect 519 4523 528 4557
rect 1168 4565 1220 4617
rect -34 4454 18 4473
rect -34 4421 -26 4454
rect -26 4421 8 4454
rect 8 4421 18 4454
rect -34 4382 18 4404
rect -34 4352 -26 4382
rect -26 4352 8 4382
rect 8 4352 18 4382
rect 65 4420 117 4472
rect 393 4464 445 4516
rect 476 4516 528 4523
rect 857 4457 909 4509
rect 940 4457 992 4509
rect 1023 4457 1075 4509
rect 1168 4500 1220 4552
rect 65 4353 117 4405
rect 393 4397 445 4449
rect 612 4386 664 4438
rect 1168 4435 1220 4487
rect 476 4348 528 4357
rect 476 4314 485 4348
rect 485 4314 519 4348
rect 519 4314 528 4348
rect 65 4249 117 4301
rect 476 4305 528 4314
rect 612 4322 664 4374
rect 1168 4370 1220 4422
rect 1168 4305 1220 4357
rect 65 4162 117 4214
rect 1168 4240 1220 4292
rect 1168 4175 1220 4227
rect 65 4075 117 4127
rect 1168 4110 1220 4162
rect 151 3835 203 3887
rect 220 3835 272 3887
rect 289 3835 341 3887
rect 65 3765 117 3817
rect 65 3700 117 3752
rect 476 4046 528 4052
rect 476 4012 485 4046
rect 485 4012 519 4046
rect 519 4012 528 4046
rect 692 4038 744 4044
rect 476 4000 528 4012
rect 476 3960 528 3984
rect 476 3932 485 3960
rect 485 3932 519 3960
rect 519 3932 528 3960
rect 476 3874 528 3916
rect 476 3864 485 3874
rect 485 3864 519 3874
rect 519 3864 528 3874
rect 476 3840 485 3848
rect 485 3840 519 3848
rect 519 3840 528 3848
rect 476 3796 528 3840
rect 476 3754 485 3781
rect 485 3754 519 3781
rect 519 3754 528 3781
rect 476 3729 528 3754
rect 476 3702 528 3714
rect 476 3668 485 3702
rect 485 3668 519 3702
rect 519 3668 528 3702
rect 612 3963 664 4015
rect 612 3897 664 3949
rect 612 3832 664 3884
rect 612 3767 664 3819
rect 612 3702 664 3754
rect 692 4004 701 4038
rect 701 4004 735 4038
rect 735 4004 744 4038
rect 692 3992 744 4004
rect 692 3956 744 3979
rect 692 3927 701 3956
rect 701 3927 735 3956
rect 735 3927 744 3956
rect 692 3874 744 3915
rect 692 3863 701 3874
rect 701 3863 735 3874
rect 735 3863 744 3874
rect 692 3840 701 3851
rect 701 3840 735 3851
rect 735 3840 744 3851
rect 692 3799 744 3840
rect 692 3758 701 3787
rect 701 3758 735 3787
rect 735 3758 744 3787
rect 692 3735 744 3758
rect 692 3711 744 3723
rect 476 3662 528 3668
rect 692 3677 701 3711
rect 701 3677 735 3711
rect 735 3677 744 3711
rect 1168 4045 1220 4097
rect 1168 3980 1220 4032
rect 1168 3915 1220 3967
rect 857 3835 909 3887
rect 940 3835 992 3887
rect 1023 3835 1075 3887
rect 1168 3850 1220 3902
rect 1168 3785 1220 3837
rect 1685 3870 1737 3922
rect 1685 3804 1737 3856
rect 1168 3719 1220 3771
rect 692 3671 744 3677
rect 1168 3653 1220 3705
rect 1168 3587 1220 3639
rect 1168 3521 1220 3573
rect 65 3324 117 3376
rect 65 3250 117 3302
rect 65 3176 117 3228
rect 151 3213 203 3265
rect 220 3213 272 3265
rect 289 3213 341 3265
rect 65 3103 117 3155
rect 476 3420 528 3426
rect 476 3386 485 3420
rect 485 3386 519 3420
rect 519 3386 528 3420
rect 692 3423 744 3429
rect 476 3374 528 3386
rect 476 3335 528 3359
rect 476 3307 485 3335
rect 485 3307 519 3335
rect 519 3307 528 3335
rect 476 3250 528 3292
rect 476 3240 485 3250
rect 485 3240 519 3250
rect 519 3240 528 3250
rect 476 3216 485 3225
rect 485 3216 519 3225
rect 519 3216 528 3225
rect 476 3173 528 3216
rect 476 3131 485 3158
rect 485 3131 519 3158
rect 519 3131 528 3158
rect 476 3106 528 3131
rect 476 3080 528 3092
rect 476 3046 485 3080
rect 485 3046 519 3080
rect 519 3046 528 3080
rect 612 3342 664 3394
rect 612 3276 664 3328
rect 612 3211 664 3263
rect 612 3146 664 3198
rect 612 3081 664 3133
rect 692 3389 701 3423
rect 701 3389 735 3423
rect 735 3389 744 3423
rect 692 3377 744 3389
rect 692 3340 744 3363
rect 692 3311 701 3340
rect 701 3311 735 3340
rect 735 3311 744 3340
rect 692 3257 744 3297
rect 692 3245 701 3257
rect 701 3245 735 3257
rect 735 3245 744 3257
rect 692 3223 701 3231
rect 701 3223 735 3231
rect 735 3223 744 3231
rect 692 3179 744 3223
rect 692 3139 701 3166
rect 701 3139 735 3166
rect 735 3139 744 3166
rect 692 3114 744 3139
rect 692 3089 744 3101
rect 476 3040 528 3046
rect 692 3055 701 3089
rect 701 3055 735 3089
rect 735 3055 744 3089
rect 1168 3455 1220 3507
rect 1168 3389 1220 3441
rect 1168 3323 1220 3375
rect 857 3213 909 3265
rect 940 3213 992 3265
rect 1023 3213 1075 3265
rect 1168 3257 1220 3309
rect 1168 3191 1220 3243
rect 1168 3125 1220 3177
rect 692 3049 744 3055
rect 1168 3059 1220 3111
rect 1168 2993 1220 3045
rect 1168 2923 1220 2975
rect 1232 2923 1284 2975
rect 1296 2923 1348 2975
rect 1360 2923 1412 2975
rect 1424 2923 1476 2975
rect 1168 2856 1220 2908
rect 1232 2856 1284 2908
rect 1296 2856 1348 2908
rect 1360 2856 1412 2908
rect 1424 2856 1476 2908
rect 65 2701 117 2753
rect 65 2630 117 2682
rect 65 2558 117 2610
rect 151 2591 203 2643
rect 220 2591 272 2643
rect 289 2591 341 2643
rect 65 2486 117 2538
rect 476 2795 528 2801
rect 476 2761 485 2795
rect 485 2761 519 2795
rect 519 2761 528 2795
rect 692 2801 744 2807
rect 476 2749 528 2761
rect 476 2711 528 2734
rect 476 2682 485 2711
rect 485 2682 519 2711
rect 519 2682 528 2711
rect 476 2627 528 2668
rect 612 2700 664 2752
rect 612 2633 664 2685
rect 692 2767 701 2801
rect 701 2767 735 2801
rect 735 2767 744 2801
rect 692 2755 744 2767
rect 692 2719 744 2742
rect 692 2690 701 2719
rect 701 2690 735 2719
rect 735 2690 744 2719
rect 692 2637 744 2677
rect 476 2616 485 2627
rect 485 2616 519 2627
rect 519 2616 528 2627
rect 476 2593 485 2602
rect 485 2593 519 2602
rect 519 2593 528 2602
rect 476 2550 528 2593
rect 476 2509 485 2536
rect 485 2509 519 2536
rect 519 2509 528 2536
rect 476 2484 528 2509
rect 476 2458 528 2470
rect 476 2424 485 2458
rect 485 2424 519 2458
rect 519 2424 528 2458
rect 476 2418 528 2424
rect 692 2625 701 2637
rect 701 2625 735 2637
rect 735 2625 744 2637
rect 692 2603 701 2613
rect 701 2603 735 2613
rect 735 2603 744 2613
rect 692 2561 744 2603
rect 692 2521 701 2549
rect 701 2521 735 2549
rect 735 2521 744 2549
rect 692 2497 744 2521
rect 692 2473 744 2485
rect 1168 2789 1220 2841
rect 1232 2789 1284 2841
rect 1296 2789 1348 2841
rect 1360 2789 1412 2841
rect 1424 2789 1476 2841
rect 863 2697 915 2749
rect 927 2697 979 2749
rect 991 2697 1043 2749
rect 1055 2697 1107 2749
rect 863 2634 915 2680
rect 863 2628 875 2634
rect 875 2628 909 2634
rect 909 2628 915 2634
rect 927 2634 979 2680
rect 991 2634 1043 2680
rect 1055 2634 1107 2680
rect 927 2628 962 2634
rect 962 2628 979 2634
rect 991 2628 996 2634
rect 996 2628 1043 2634
rect 1055 2628 1082 2634
rect 1082 2628 1107 2634
rect 863 2600 875 2610
rect 875 2600 909 2610
rect 909 2600 915 2610
rect 863 2558 915 2600
rect 927 2600 962 2610
rect 962 2600 979 2610
rect 991 2600 996 2610
rect 996 2600 1043 2610
rect 1055 2600 1082 2610
rect 1082 2600 1107 2610
rect 927 2558 979 2600
rect 991 2558 1043 2600
rect 1055 2558 1107 2600
rect 692 2439 701 2473
rect 701 2439 735 2473
rect 735 2439 744 2473
rect 1168 2466 1220 2518
rect 1232 2466 1284 2518
rect 1296 2466 1348 2518
rect 1360 2466 1412 2518
rect 1424 2466 1476 2518
rect 692 2433 744 2439
rect 1168 2377 1220 2429
rect 1232 2377 1284 2429
rect 1296 2377 1348 2429
rect 1360 2377 1412 2429
rect 1424 2377 1476 2429
rect 145 2246 197 2298
rect 145 2174 197 2226
rect 145 2102 197 2154
rect 476 2262 528 2304
rect 231 2228 237 2249
rect 237 2228 271 2249
rect 271 2228 283 2249
rect 476 2252 507 2262
rect 507 2252 528 2262
rect 476 2228 507 2229
rect 507 2228 528 2229
rect 231 2197 283 2228
rect 231 2136 283 2185
rect 476 2177 528 2228
rect 476 2136 528 2154
rect 1168 2288 1220 2340
rect 1232 2288 1284 2340
rect 1296 2288 1348 2340
rect 1360 2288 1412 2340
rect 1424 2288 1476 2340
rect 612 2213 664 2265
rect 612 2147 664 2199
rect 231 2133 237 2136
rect 237 2133 271 2136
rect 271 2133 283 2136
rect 476 2102 507 2136
rect 507 2102 528 2136
rect 1685 2010 1737 2062
rect 1596 1948 1648 2000
rect -280 1877 -228 1929
rect 1516 1877 1568 1929
rect -280 1813 -228 1865
rect 209 1867 261 1872
rect 289 1867 341 1872
rect 209 1833 248 1867
rect 248 1833 261 1867
rect 289 1833 323 1867
rect 323 1833 341 1867
rect 476 1833 507 1867
rect 507 1833 528 1867
rect 209 1820 261 1833
rect 289 1820 341 1833
rect 476 1815 528 1833
rect 209 1795 261 1808
rect 289 1795 341 1808
rect 476 1795 528 1803
rect 209 1761 248 1795
rect 248 1761 261 1795
rect 289 1761 323 1795
rect 323 1761 341 1795
rect 476 1761 507 1795
rect 507 1761 528 1795
rect 692 1806 744 1858
rect 1180 1806 1232 1858
rect 1244 1806 1296 1858
rect 1308 1806 1360 1858
rect 1372 1806 1424 1858
rect 1436 1806 1488 1858
rect 1516 1811 1568 1863
rect 1685 1944 1737 1996
rect 1596 1882 1648 1934
rect 692 1774 744 1792
rect 209 1756 261 1761
rect 289 1756 341 1761
rect 476 1751 528 1761
rect -280 1605 -228 1657
rect -280 1541 -228 1593
rect 145 1649 197 1701
rect 209 1647 261 1699
rect 289 1647 341 1699
rect 145 1577 197 1629
rect 209 1583 261 1635
rect 289 1583 341 1635
rect 612 1708 664 1760
rect 692 1740 713 1774
rect 713 1740 744 1774
rect 1180 1740 1232 1792
rect 1244 1740 1296 1792
rect 1308 1740 1360 1792
rect 1372 1740 1424 1792
rect 1436 1740 1488 1792
rect 1168 1702 1171 1728
rect 1171 1702 1205 1728
rect 1205 1702 1220 1728
rect 612 1644 664 1696
rect 1168 1676 1220 1702
rect 1168 1652 1220 1659
rect 1168 1618 1171 1652
rect 1171 1618 1205 1652
rect 1205 1618 1220 1652
rect 1168 1607 1220 1618
rect 145 1505 197 1557
rect 145 1433 197 1485
rect 393 1496 445 1548
rect 556 1496 608 1548
rect 1168 1568 1220 1590
rect 1168 1538 1171 1568
rect 1171 1538 1205 1568
rect 1205 1538 1220 1568
rect 214 1429 266 1481
rect 289 1429 341 1481
rect 393 1429 445 1481
rect 556 1475 608 1484
rect 556 1441 577 1475
rect 577 1441 608 1475
rect 1168 1484 1220 1521
rect 1168 1469 1171 1484
rect 1171 1469 1205 1484
rect 1205 1469 1220 1484
rect 556 1432 608 1441
rect 145 1361 197 1413
rect 214 1365 266 1417
rect 289 1365 341 1417
rect 692 1406 744 1424
rect -95 1283 -43 1335
rect -31 1283 21 1335
rect 145 1289 197 1341
rect 482 1392 534 1398
rect 482 1358 488 1392
rect 488 1358 522 1392
rect 522 1358 534 1392
rect 692 1372 704 1406
rect 704 1372 738 1406
rect 738 1372 744 1406
rect 857 1395 909 1447
rect 940 1395 992 1447
rect 1023 1395 1075 1447
rect 1168 1450 1171 1452
rect 1171 1450 1205 1452
rect 1205 1450 1220 1452
rect 1168 1400 1220 1450
rect 482 1346 534 1358
rect -95 1214 -43 1266
rect -31 1214 21 1266
rect 145 1226 197 1269
rect 612 1259 664 1311
rect 1168 1366 1171 1383
rect 1171 1366 1205 1383
rect 1205 1366 1220 1383
rect 1168 1331 1220 1366
rect 1168 1283 1171 1314
rect 1171 1283 1205 1314
rect 1205 1283 1220 1314
rect 1168 1262 1220 1283
rect 145 1217 157 1226
rect 157 1217 191 1226
rect 191 1217 197 1226
rect -95 1145 -43 1197
rect -31 1145 21 1197
rect 145 1192 157 1197
rect 157 1192 191 1197
rect 191 1192 197 1197
rect 145 1145 197 1192
rect 210 1192 229 1197
rect 229 1192 262 1197
rect 274 1192 301 1197
rect 301 1192 326 1197
rect 210 1145 262 1192
rect 274 1145 326 1192
rect 387 1211 439 1258
rect 387 1206 405 1211
rect 405 1206 439 1211
rect 387 1177 405 1194
rect 405 1177 439 1194
rect 612 1194 664 1246
rect 857 1231 909 1240
rect 940 1231 992 1240
rect 1023 1231 1075 1240
rect 857 1197 867 1231
rect 867 1197 901 1231
rect 901 1197 909 1231
rect 940 1197 973 1231
rect 973 1197 992 1231
rect 1023 1197 1045 1231
rect 1045 1197 1075 1231
rect 857 1188 909 1197
rect 940 1188 992 1197
rect 1023 1188 1075 1197
rect 1168 1234 1220 1246
rect 1168 1200 1171 1234
rect 1171 1200 1205 1234
rect 1205 1200 1220 1234
rect 1168 1194 1220 1200
rect 387 1142 439 1177
rect 476 1123 528 1131
rect 476 1089 485 1123
rect 485 1089 519 1123
rect 519 1089 528 1123
rect 476 1079 528 1089
rect 692 1090 744 1098
rect 692 1056 701 1090
rect 701 1056 735 1090
rect 735 1056 744 1090
rect 692 1046 744 1056
rect 1168 1092 1220 1098
rect 1168 1058 1171 1092
rect 1171 1058 1205 1092
rect 1205 1058 1220 1092
rect 1168 1046 1220 1058
rect 476 852 528 858
rect 476 818 485 852
rect 485 818 519 852
rect 519 818 528 852
rect 476 806 528 818
rect 393 787 445 793
rect 151 705 203 757
rect 220 705 272 757
rect 289 705 341 757
rect 393 753 403 787
rect 403 753 437 787
rect 437 753 445 787
rect 393 741 445 753
rect 393 708 445 717
rect 393 674 403 708
rect 403 674 437 708
rect 437 674 445 708
rect 393 665 445 674
rect 393 630 445 641
rect 393 596 403 630
rect 403 596 437 630
rect 437 596 445 630
rect 393 589 445 596
rect 151 521 203 573
rect 220 521 272 573
rect 289 521 341 573
rect 393 552 445 564
rect 393 518 403 552
rect 403 518 437 552
rect 437 518 445 552
rect 393 512 445 518
rect 476 772 528 791
rect 476 739 485 772
rect 485 739 519 772
rect 519 739 528 772
rect 692 824 701 858
rect 701 824 735 858
rect 735 824 744 858
rect 692 806 744 824
rect 692 786 744 794
rect 692 752 701 786
rect 701 752 735 786
rect 735 752 744 786
rect 692 742 744 752
rect 476 692 528 724
rect 476 672 485 692
rect 485 672 519 692
rect 519 672 528 692
rect 476 612 528 657
rect 476 605 485 612
rect 485 605 519 612
rect 519 605 528 612
rect 476 578 485 590
rect 485 578 519 590
rect 519 578 528 590
rect 857 705 909 757
rect 940 705 992 757
rect 1023 705 1075 757
rect 612 650 664 702
rect 612 585 664 637
rect 692 604 744 610
rect 476 538 528 578
rect 476 499 485 523
rect 485 499 519 523
rect 519 499 528 523
rect 151 332 203 384
rect 220 332 272 384
rect 289 332 341 384
rect 476 471 528 499
rect 476 454 528 456
rect 476 420 485 454
rect 485 420 519 454
rect 519 420 528 454
rect 476 404 528 420
rect 476 375 528 389
rect 476 341 485 375
rect 485 341 519 375
rect 519 341 528 375
rect 476 337 528 341
rect 476 296 528 322
rect 476 270 485 296
rect 485 270 519 296
rect 519 270 528 296
rect 476 204 528 256
rect -106 172 -54 183
rect -21 172 31 183
rect 151 172 203 183
rect 220 172 272 183
rect -106 138 -85 172
rect -85 138 -54 172
rect -21 138 -9 172
rect -9 138 25 172
rect 25 138 31 172
rect 151 138 177 172
rect 177 138 203 172
rect 220 138 253 172
rect 253 138 272 172
rect -106 131 -54 138
rect -21 131 31 138
rect 151 131 203 138
rect 220 131 272 138
rect 289 172 341 183
rect 476 172 528 190
rect 289 138 295 172
rect 295 138 329 172
rect 329 138 341 172
rect 476 138 481 172
rect 481 138 528 172
rect 692 570 701 604
rect 701 570 735 604
rect 735 570 744 604
rect 692 558 744 570
rect 692 529 744 543
rect 692 495 701 529
rect 701 495 735 529
rect 735 495 744 529
rect 692 491 744 495
rect 692 454 744 476
rect 692 424 701 454
rect 701 424 735 454
rect 735 424 744 454
rect 692 380 744 409
rect 692 357 701 380
rect 701 357 735 380
rect 735 357 744 380
rect 692 306 744 342
rect 692 290 701 306
rect 701 290 735 306
rect 735 290 744 306
rect 857 521 909 573
rect 940 521 992 573
rect 1023 521 1075 573
rect 857 337 909 389
rect 940 337 992 389
rect 1023 337 1075 389
rect 692 272 701 276
rect 701 272 735 276
rect 735 272 744 276
rect 692 224 744 272
rect 1168 1014 1220 1029
rect 1168 980 1171 1014
rect 1171 980 1205 1014
rect 1205 980 1220 1014
rect 1168 977 1220 980
rect 1168 936 1220 960
rect 1168 908 1171 936
rect 1171 908 1205 936
rect 1205 908 1220 936
rect 1168 858 1220 891
rect 1168 839 1171 858
rect 1171 839 1205 858
rect 1205 839 1220 858
rect 1168 780 1220 822
rect 1168 770 1171 780
rect 1171 770 1205 780
rect 1205 770 1220 780
rect 1168 746 1171 754
rect 1171 746 1205 754
rect 1205 746 1220 754
rect 1168 702 1220 746
rect 1168 668 1171 686
rect 1171 668 1205 686
rect 1205 668 1220 686
rect 1168 634 1220 668
rect 1168 590 1171 618
rect 1171 590 1205 618
rect 1205 590 1220 618
rect 1168 566 1220 590
rect 1168 546 1220 550
rect 1168 512 1171 546
rect 1171 512 1205 546
rect 1205 512 1220 546
rect 1168 498 1220 512
rect 1168 467 1220 482
rect 1168 433 1171 467
rect 1171 433 1205 467
rect 1205 433 1220 467
rect 1168 430 1220 433
rect 1168 388 1220 414
rect 1168 362 1171 388
rect 1171 362 1205 388
rect 1205 362 1220 388
rect 1168 309 1220 346
rect 1168 294 1171 309
rect 1171 294 1205 309
rect 1205 294 1220 309
rect 1168 275 1171 278
rect 1171 275 1205 278
rect 1205 275 1220 278
rect 1168 230 1220 275
rect 1168 226 1171 230
rect 1171 226 1205 230
rect 1205 226 1220 230
rect 692 192 744 210
rect 1168 196 1171 210
rect 1171 196 1205 210
rect 1205 196 1220 210
rect 692 158 739 192
rect 739 158 744 192
rect 1168 158 1220 196
rect 289 131 341 138
<< metal2 >>
rect 598 8997 918 9328
tri 918 8997 950 9029 sw
rect 598 8895 950 8997
tri 598 8863 630 8895 ne
rect 630 8441 950 8895
tri 950 8441 1002 8493 sw
rect 630 8429 1002 8441
tri 1002 8429 1014 8441 sw
rect 1106 8429 1426 9328
rect 1454 8557 1861 8909
rect 1454 8505 1522 8557
rect 1574 8505 1592 8557
rect 1644 8505 1662 8557
rect 1714 8505 1732 8557
rect 1784 8505 1803 8557
rect 1855 8505 1861 8557
rect 1454 8493 1861 8505
rect 1454 8442 1522 8493
tri 1454 8441 1455 8442 ne
rect 1455 8441 1522 8442
rect 1574 8441 1592 8493
rect 1644 8441 1662 8493
rect 1714 8441 1732 8493
rect 1784 8441 1803 8493
rect 1855 8441 1861 8493
rect 2360 8685 2680 9328
tri 2360 8464 2581 8685 ne
rect 2581 8676 2680 8685
tri 2680 8676 2822 8818 sw
rect 2581 8464 3949 8676
tri 1455 8430 1466 8441 ne
rect 1466 8430 1861 8441
tri 1426 8429 1427 8430 sw
tri 1466 8429 1467 8430 ne
rect 1467 8429 1861 8430
rect 630 8423 1014 8429
tri 1014 8423 1020 8429 sw
rect 1106 8423 1427 8429
rect 630 8377 1020 8423
tri 1020 8377 1066 8423 sw
tri 1106 8377 1152 8423 ne
rect 1152 8408 1427 8423
tri 1427 8408 1448 8429 sw
tri 1467 8408 1488 8429 ne
rect 1488 8408 1522 8429
rect 1152 8377 1448 8408
tri 1448 8377 1479 8408 sw
tri 1488 8380 1516 8408 ne
rect 1516 8377 1522 8408
rect 1574 8377 1592 8429
rect 1644 8377 1662 8429
rect 1714 8377 1732 8429
rect 1784 8377 1803 8429
rect 1855 8377 1861 8429
rect 630 8361 1066 8377
tri 1066 8361 1082 8377 sw
tri 1152 8361 1168 8377 ne
rect 1168 8368 1479 8377
tri 1479 8368 1488 8377 sw
rect 630 8359 1082 8361
tri 630 8257 732 8359 ne
rect 732 8336 1082 8359
tri 1082 8336 1107 8361 sw
rect 732 8257 1107 8336
rect 344 8205 350 8257
rect 402 8205 420 8257
rect 472 8205 489 8257
rect 541 8205 553 8257
rect 344 8077 553 8205
rect 669 8077 675 8257
tri 732 8205 784 8257 ne
rect 784 8205 1107 8257
tri 784 8202 787 8205 ne
rect 344 7987 675 8077
rect 344 7935 388 7987
rect 440 7935 489 7987
rect 541 7935 675 7987
tri 314 7607 344 7637 se
rect 344 7607 675 7935
tri 304 7597 314 7607 se
rect 314 7597 675 7607
tri 270 7563 304 7597 se
rect 304 7563 675 7597
tri 218 7511 270 7563 se
rect 270 7511 675 7563
tri 203 7496 218 7511 se
rect 218 7496 675 7511
tri 174 7467 203 7496 se
rect 203 7467 350 7496
tri 151 7444 174 7467 se
rect 174 7444 350 7467
rect 402 7444 428 7496
rect 480 7444 507 7496
rect 559 7467 675 7496
rect 559 7444 639 7467
tri 139 7432 151 7444 se
rect 151 7432 639 7444
tri 87 7380 139 7432 se
rect 139 7380 350 7432
rect 402 7380 428 7432
rect 480 7380 507 7432
rect 559 7431 639 7432
tri 639 7431 675 7467 nw
rect 559 7423 631 7431
tri 631 7423 639 7431 nw
rect 559 7387 595 7423
tri 595 7387 631 7423 nw
rect 559 7380 584 7387
tri 65 7358 87 7380 se
rect 87 7358 584 7380
tri 584 7376 595 7387 nw
tri 13 7306 65 7358 se
rect 65 7306 584 7358
tri -2 7291 13 7306 se
rect 13 7291 584 7306
tri -29 7264 -2 7291 se
rect -2 7264 584 7291
rect -29 6913 584 7264
rect 612 7358 664 7364
rect 612 7291 664 7306
rect 612 7233 664 7239
tri 612 7217 628 7233 ne
rect 628 7217 664 7233
tri 628 7209 636 7217 ne
rect -29 6894 565 6913
tri 565 6894 584 6913 nw
tri 613 6894 636 6917 se
rect 636 6894 664 7217
rect -29 6887 558 6894
tri 558 6887 565 6894 nw
tri 612 6893 613 6894 se
rect 613 6893 664 6894
rect 612 6887 664 6893
rect -29 6876 528 6887
rect -29 6824 44 6876
rect 96 6875 528 6876
rect 96 6824 347 6875
tri 347 6835 387 6875 nw
tri 428 6835 468 6875 ne
rect 468 6835 528 6875
tri 528 6857 558 6887 nw
tri 468 6827 476 6835 ne
rect -29 6775 347 6824
rect -29 6723 44 6775
rect 96 6769 347 6775
rect 96 6723 151 6769
rect -29 6717 151 6723
rect 203 6717 220 6769
rect 272 6717 289 6769
rect 341 6717 347 6769
rect -29 6613 347 6717
rect -29 6561 44 6613
rect 96 6561 347 6613
rect -29 6544 347 6561
rect -29 6492 44 6544
rect 96 6492 347 6544
rect -119 6471 -67 6477
rect -119 6407 -67 6419
tri -138 5446 -119 5465 se
rect -119 5446 -67 6355
tri -154 5430 -138 5446 se
rect -138 5443 -67 5446
rect -138 5430 -80 5443
tri -80 5430 -67 5443 nw
rect -29 6475 347 6492
rect -29 6423 44 6475
rect 96 6457 347 6475
rect 96 6423 151 6457
rect -29 6406 151 6423
rect -29 6354 44 6406
rect 96 6405 151 6406
rect 203 6405 220 6457
rect 272 6405 289 6457
rect 341 6405 347 6457
rect 96 6354 347 6405
rect -29 6337 347 6354
rect -29 6285 44 6337
rect 96 6285 347 6337
rect -29 6268 347 6285
rect -29 6216 44 6268
rect 96 6216 347 6268
rect -29 6200 347 6216
rect -29 6148 44 6200
rect 96 6148 347 6200
rect -29 6132 347 6148
rect -29 6080 44 6132
rect 96 6131 347 6132
rect 96 6080 151 6131
rect -29 6079 151 6080
rect 203 6079 220 6131
rect 272 6079 289 6131
rect 341 6079 347 6131
rect -29 6064 347 6079
rect -29 6012 44 6064
rect 96 6012 347 6064
rect -29 5906 347 6012
rect -29 5854 44 5906
rect 96 5854 347 5906
rect -29 5838 347 5854
rect -29 5786 44 5838
rect 96 5805 347 5838
rect 96 5786 151 5805
rect -29 5770 151 5786
rect -29 5718 44 5770
rect 96 5753 151 5770
rect 203 5753 220 5805
rect 272 5753 289 5805
rect 341 5753 347 5805
rect 476 6216 528 6835
rect 612 6820 664 6835
rect 612 6762 664 6768
tri 612 6738 636 6762 ne
rect 476 5832 528 6164
rect 96 5718 347 5753
rect -29 5702 347 5718
rect -29 5650 44 5702
rect 96 5650 347 5702
rect -29 5634 347 5650
rect -29 5582 44 5634
rect 96 5582 347 5634
rect -29 5566 347 5582
rect -29 5514 44 5566
rect 96 5514 347 5566
rect -29 5498 347 5514
rect -29 5446 44 5498
rect 96 5446 347 5498
rect -29 5430 347 5446
tri -193 5391 -154 5430 se
rect -154 5391 -119 5430
tri -119 5391 -80 5430 nw
tri -206 5378 -193 5391 se
rect -193 5378 -132 5391
tri -132 5378 -119 5391 nw
rect -29 5378 44 5430
rect 96 5378 347 5430
tri -211 5373 -206 5378 se
rect -206 5373 -137 5378
tri -137 5373 -132 5378 nw
rect -29 5373 347 5378
tri -222 5362 -211 5373 se
rect -211 5362 -148 5373
tri -148 5362 -137 5373 nw
rect -29 5362 151 5373
tri -267 5317 -222 5362 se
rect -222 5317 -193 5362
tri -193 5317 -148 5362 nw
tri -274 5310 -267 5317 se
rect -267 5310 -200 5317
tri -200 5310 -193 5317 nw
tri -35 5310 -29 5316 se
rect -29 5310 44 5362
rect 96 5321 151 5362
rect 203 5321 220 5373
rect 272 5321 289 5373
rect 341 5321 347 5373
rect 96 5310 347 5321
tri -290 5294 -274 5310 se
rect -274 5294 -216 5310
tri -216 5294 -200 5310 nw
tri -51 5294 -35 5310 se
rect -35 5294 347 5310
tri -313 5271 -290 5294 se
rect -290 5271 -261 5294
rect -313 2982 -261 5271
tri -261 5249 -216 5294 nw
tri -96 5249 -51 5294 se
rect -51 5249 44 5294
tri -103 5242 -96 5249 se
rect -96 5242 44 5249
rect 96 5242 347 5294
tri -112 5233 -103 5242 se
rect -103 5233 347 5242
rect -112 5217 347 5233
rect -112 5203 68 5217
tri 68 5203 82 5217 nw
tri 111 5203 125 5217 ne
rect 125 5203 347 5217
rect -112 4898 37 5203
tri 37 5172 68 5203 nw
tri 125 5183 145 5203 ne
rect -112 4846 -106 4898
rect -54 4846 -21 4898
rect 31 4846 37 4898
rect -112 4542 37 4846
rect -112 4490 -34 4542
rect 18 4490 37 4542
rect -112 4473 37 4490
rect -112 4421 -34 4473
rect 18 4421 37 4473
rect -112 4404 37 4421
rect -112 4352 -34 4404
rect 18 4352 37 4404
rect -280 1929 -228 1935
rect -280 1865 -228 1877
rect -280 1657 -228 1813
rect -280 1593 -228 1605
rect -280 1535 -228 1541
rect -112 1335 37 4352
rect 65 5148 117 5154
rect 65 5027 117 5096
rect 65 4472 117 4975
rect 65 4405 117 4420
rect 65 4347 117 4353
rect 145 4941 347 5203
rect 145 4889 151 4941
rect 203 4889 220 4941
rect 272 4889 289 4941
rect 341 4889 347 4941
rect 145 4558 347 4889
rect 145 4506 151 4558
rect 203 4506 220 4558
rect 272 4506 289 4558
rect 341 4506 347 4558
rect 65 4301 117 4307
rect 65 4214 117 4249
rect 65 4127 117 4162
rect 65 3817 117 4075
rect 65 3752 117 3765
rect 65 3376 117 3700
rect 65 3302 117 3324
rect 65 3228 117 3250
rect 65 3155 117 3176
rect 65 2753 117 3103
rect 65 2682 117 2701
rect 65 2610 117 2630
rect 65 2538 117 2558
rect 65 2456 117 2486
rect 145 3887 347 4506
rect 393 5778 445 5784
rect 393 5711 445 5726
rect 393 5345 445 5659
rect 393 5278 445 5293
rect 393 4516 445 5226
rect 393 4449 445 4464
rect 393 4391 445 4397
rect 476 5757 528 5780
rect 476 5683 528 5705
rect 476 5505 528 5631
rect 476 5421 528 5453
rect 476 5338 528 5369
rect 476 5255 528 5286
rect 476 4568 528 5203
rect 145 3835 151 3887
rect 203 3835 220 3887
rect 272 3835 289 3887
rect 341 3835 347 3887
rect 145 3265 347 3835
rect 145 3213 151 3265
rect 203 3213 220 3265
rect 272 3213 289 3265
rect 341 3213 347 3265
rect 145 2643 347 3213
rect 145 2591 151 2643
rect 203 2591 220 2643
rect 272 2591 289 2643
rect 341 2591 347 2643
rect -112 1283 -95 1335
rect -43 1283 -31 1335
rect 21 1283 37 1335
rect -112 1266 37 1283
rect -112 1214 -95 1266
rect -43 1214 -31 1266
rect 21 1214 37 1266
rect -112 1197 37 1214
rect -112 1145 -95 1197
rect -43 1145 -31 1197
rect 21 1145 37 1197
rect -112 183 37 1145
rect -112 131 -106 183
rect -54 131 -21 183
rect 31 131 37 183
rect -112 112 37 131
rect 145 2298 347 2591
rect 197 2249 347 2298
rect 197 2246 231 2249
rect 145 2226 231 2246
rect 197 2197 231 2226
rect 283 2197 347 2249
rect 197 2185 347 2197
rect 197 2174 231 2185
rect 145 2154 231 2174
rect 197 2133 231 2154
rect 283 2133 347 2185
rect 197 2102 347 2133
rect 145 1872 347 2102
rect 145 1820 209 1872
rect 261 1820 289 1872
rect 341 1820 347 1872
rect 145 1808 347 1820
rect 145 1756 209 1808
rect 261 1756 289 1808
rect 341 1756 347 1808
rect 145 1701 347 1756
rect 197 1699 347 1701
rect 197 1649 209 1699
rect 145 1647 209 1649
rect 261 1647 289 1699
rect 341 1647 347 1699
rect 145 1635 347 1647
rect 145 1629 209 1635
rect 197 1583 209 1629
rect 261 1583 289 1635
rect 341 1583 347 1635
rect 197 1577 347 1583
rect 145 1557 347 1577
rect 197 1505 347 1557
rect 476 4357 528 4516
rect 476 4052 528 4305
rect 476 3984 528 4000
rect 476 3916 528 3932
rect 476 3848 528 3864
rect 476 3781 528 3796
rect 476 3714 528 3729
rect 476 3426 528 3662
rect 476 3359 528 3374
rect 476 3292 528 3307
rect 476 3225 528 3240
rect 476 3158 528 3173
rect 476 3092 528 3106
rect 476 2801 528 3040
rect 476 2734 528 2749
rect 476 2668 528 2682
rect 476 2602 528 2616
rect 476 2536 528 2550
rect 476 2470 528 2484
rect 476 2304 528 2418
rect 476 2229 528 2252
rect 476 2154 528 2177
rect 476 1867 528 2102
rect 476 1803 528 1815
rect 145 1485 347 1505
rect 197 1481 347 1485
rect 197 1433 214 1481
rect 145 1429 214 1433
rect 266 1429 289 1481
rect 341 1429 347 1481
rect 145 1417 347 1429
rect 145 1413 214 1417
rect 197 1365 214 1413
rect 266 1365 289 1417
rect 341 1365 347 1417
rect 197 1361 347 1365
rect 145 1341 347 1361
rect 197 1289 347 1341
rect 145 1269 347 1289
rect 197 1217 347 1269
rect 145 1197 347 1217
rect 197 1145 210 1197
rect 262 1145 274 1197
rect 326 1145 347 1197
rect 145 757 347 1145
rect 145 705 151 757
rect 203 705 220 757
rect 272 705 289 757
rect 341 705 347 757
rect 145 573 347 705
rect 145 521 151 573
rect 203 521 220 573
rect 272 521 289 573
rect 341 521 347 573
rect 145 384 347 521
rect 381 1548 445 1554
rect 381 1496 393 1548
rect 381 1481 445 1496
rect 381 1429 393 1481
rect 381 1258 445 1429
rect 381 1206 387 1258
rect 439 1206 445 1258
rect 381 1194 445 1206
rect 381 1142 387 1194
rect 439 1142 445 1194
rect 381 793 445 1142
rect 381 741 393 793
rect 381 717 445 741
rect 381 665 393 717
rect 381 641 445 665
rect 381 589 393 641
rect 381 564 445 589
rect 381 512 393 564
rect 381 506 445 512
rect 476 1398 528 1751
rect 556 6719 608 6725
rect 556 6652 608 6667
rect 556 6594 608 6600
rect 556 6591 600 6594
tri 600 6591 603 6594 nw
rect 556 1554 584 6591
tri 584 6575 600 6591 nw
tri 627 6563 636 6572 se
rect 636 6563 664 6762
tri 612 6548 627 6563 se
rect 627 6548 664 6563
rect 612 6542 664 6548
rect 612 6475 664 6490
rect 612 6417 664 6423
tri 612 6393 636 6417 ne
tri 612 6293 636 6317 se
rect 636 6293 664 6417
rect 612 6287 664 6293
rect 612 6220 664 6235
rect 612 6162 664 6168
tri 612 6138 636 6162 ne
tri 614 4883 636 4905 se
rect 636 4883 664 6162
rect 692 7177 744 7183
rect 692 7110 744 7125
rect 692 5906 744 7058
rect 787 6712 1107 8205
tri 787 6689 810 6712 ne
rect 692 5839 744 5854
rect 692 5157 744 5787
rect 810 5925 1107 6712
rect 810 5873 857 5925
rect 909 5873 940 5925
rect 992 5873 1023 5925
rect 1075 5873 1107 5925
rect 692 5092 744 5105
rect 692 5034 744 5040
tri 787 5650 810 5673 se
rect 810 5650 1107 5873
tri 612 4881 614 4883 se
rect 614 4881 664 4883
rect 612 4875 664 4881
rect 612 4808 664 4823
rect 612 4750 664 4756
rect 692 4935 744 4941
rect 692 4808 744 4883
rect 612 4438 664 4444
rect 612 4374 664 4386
rect 612 4015 664 4322
rect 612 3949 664 3963
rect 612 3884 664 3897
rect 612 3819 664 3832
rect 612 3754 664 3767
rect 612 3394 664 3702
rect 612 3328 664 3342
rect 612 3263 664 3276
rect 612 3198 664 3211
rect 612 3133 664 3146
rect 612 2752 664 3081
rect 612 2685 664 2700
rect 612 2265 664 2633
rect 612 2199 664 2213
rect 612 1760 664 2147
rect 612 1696 664 1708
rect 612 1638 664 1644
rect 692 4044 744 4756
rect 692 3979 744 3992
rect 692 3915 744 3927
rect 692 3851 744 3863
rect 692 3787 744 3799
rect 692 3723 744 3735
rect 692 3429 744 3671
rect 692 3363 744 3377
rect 692 3297 744 3311
rect 692 3231 744 3245
rect 692 3166 744 3179
rect 692 3101 744 3114
rect 692 2807 744 3049
rect 692 2742 744 2755
rect 692 2677 744 2690
rect 692 2613 744 2625
rect 692 2549 744 2561
rect 692 2485 744 2497
rect 692 1858 744 2433
rect 692 1792 744 1806
tri 584 1554 608 1578 sw
rect 556 1548 608 1554
rect 556 1484 608 1496
rect 556 1426 608 1432
rect 692 1424 744 1740
tri 528 1398 540 1410 sw
rect 476 1346 482 1398
rect 534 1346 540 1398
rect 476 1131 528 1346
tri 528 1334 540 1346 nw
rect 476 858 528 1079
rect 476 791 528 806
rect 476 724 528 739
rect 476 657 528 672
rect 476 590 528 605
rect 612 1311 664 1317
rect 612 1246 664 1259
rect 612 702 664 1194
rect 612 637 664 650
rect 612 579 664 585
rect 692 1098 744 1372
rect 692 858 744 1046
rect 692 794 744 806
rect 692 610 744 742
rect 476 523 528 538
rect 145 332 151 384
rect 203 332 220 384
rect 272 332 289 384
rect 341 332 347 384
rect 145 183 347 332
rect 145 131 151 183
rect 203 131 220 183
rect 272 131 289 183
rect 341 131 347 183
rect 145 112 347 131
rect 476 456 528 471
rect 476 389 528 404
rect 476 322 528 337
rect 476 256 528 270
rect 476 190 528 204
rect 476 112 528 138
rect 692 543 744 558
rect 692 476 744 491
rect 692 409 744 424
rect 692 342 744 357
rect 692 276 744 290
rect 692 210 744 224
rect 692 112 744 158
rect 787 4509 1107 5650
rect 787 4457 857 4509
rect 909 4457 940 4509
rect 992 4457 1023 4509
rect 1075 4457 1107 4509
rect 787 3887 1107 4457
rect 787 3835 857 3887
rect 909 3835 940 3887
rect 992 3835 1023 3887
rect 1075 3835 1107 3887
rect 787 3265 1107 3835
rect 787 3213 857 3265
rect 909 3213 940 3265
rect 992 3213 1023 3265
rect 1075 3213 1107 3265
rect 787 2749 1107 3213
rect 787 2697 863 2749
rect 915 2697 927 2749
rect 979 2697 991 2749
rect 1043 2697 1055 2749
rect 787 2680 1107 2697
rect 787 2628 863 2680
rect 915 2628 927 2680
rect 979 2628 991 2680
rect 1043 2628 1055 2680
rect 787 2610 1107 2628
rect 787 2558 863 2610
rect 915 2558 927 2610
rect 979 2558 991 2610
rect 1043 2558 1055 2610
rect 787 1447 1107 2558
rect 787 1395 857 1447
rect 909 1395 940 1447
rect 992 1395 1023 1447
rect 1075 1395 1107 1447
rect 787 1240 1107 1395
rect 787 1188 857 1240
rect 909 1188 940 1240
rect 992 1188 1023 1240
rect 1075 1188 1107 1240
rect 787 757 1107 1188
rect 787 705 857 757
rect 909 705 940 757
rect 992 705 1023 757
rect 1075 705 1107 757
rect 787 573 1107 705
rect 787 521 857 573
rect 909 521 940 573
rect 992 521 1023 573
rect 1075 521 1107 573
rect 787 389 1107 521
rect 787 337 857 389
rect 909 337 940 389
rect 992 337 1023 389
rect 1075 337 1107 389
rect 787 112 1107 337
rect 1168 6713 1488 8368
rect 1516 8257 1861 8377
rect 1516 8205 1522 8257
rect 1574 8205 1592 8257
rect 1644 8205 1662 8257
rect 1714 8205 1732 8257
rect 1784 8205 1803 8257
rect 1855 8205 1861 8257
rect 1516 8193 1861 8205
rect 1516 8141 1522 8193
rect 1574 8141 1592 8193
rect 1644 8141 1662 8193
rect 1714 8141 1732 8193
rect 1784 8141 1803 8193
rect 1855 8141 1861 8193
rect 1516 8129 1861 8141
rect 1516 8077 1522 8129
rect 1574 8077 1592 8129
rect 1644 8077 1662 8129
rect 1714 8077 1732 8129
rect 1784 8077 1803 8129
rect 1855 8077 1861 8129
rect 2004 7931 2504 8464
tri 2581 8365 2680 8464 ne
rect 2680 8365 3949 8464
tri 2680 8356 2689 8365 ne
rect 2689 8356 3949 8365
tri 3816 8257 3915 8356 ne
rect 3915 8257 3949 8356
tri 3949 8257 4368 8676 sw
rect 4369 8385 5217 9328
tri 4369 8257 4497 8385 ne
rect 4497 8257 5217 8385
rect 2004 7879 2010 7931
rect 2062 7879 2083 7931
rect 2135 7879 2156 7931
rect 2208 7879 2229 7931
rect 2281 7879 2302 7931
rect 2354 7879 2374 7931
rect 2426 7879 2446 7931
rect 2498 7879 2504 7931
rect 1848 7784 1854 7836
rect 1906 7784 1918 7836
rect 1970 7784 1976 7836
rect 1596 7704 1602 7756
rect 1654 7704 1669 7756
rect 1721 7704 1727 7756
rect 1168 6037 1452 6713
tri 1452 6677 1488 6713 nw
rect 1516 6946 1568 6952
rect 1516 6879 1568 6894
rect 1168 5985 1178 6037
rect 1230 5985 1270 6037
rect 1322 5985 1363 6037
rect 1415 5985 1452 6037
rect 1168 5944 1452 5985
rect 1168 5892 1386 5944
rect 1438 5892 1452 5944
rect 1168 5877 1452 5892
rect 1168 5825 1386 5877
rect 1438 5825 1452 5877
rect 1168 5810 1452 5825
rect 1168 5758 1386 5810
rect 1438 5758 1452 5810
rect 1168 5743 1452 5758
rect 1168 5691 1386 5743
rect 1438 5691 1452 5743
rect 1168 5676 1452 5691
rect 1168 5624 1386 5676
rect 1438 5635 1452 5676
tri 1452 5635 1488 5671 sw
rect 1438 5624 1488 5635
rect 1168 5609 1488 5624
rect 1168 5557 1386 5609
rect 1438 5557 1488 5609
rect 1168 5542 1488 5557
rect 1168 5490 1386 5542
rect 1438 5490 1488 5542
rect 1168 5475 1488 5490
rect 1168 5423 1386 5475
rect 1438 5423 1488 5475
rect 1168 5408 1488 5423
rect 1168 5356 1386 5408
rect 1438 5356 1488 5408
rect 1168 5340 1488 5356
rect 1168 5317 1386 5340
rect 1168 5265 1217 5317
rect 1269 5265 1287 5317
rect 1339 5288 1386 5317
rect 1438 5288 1488 5340
rect 1339 5265 1488 5288
rect 1168 4941 1488 5265
rect 1168 4825 1174 4941
rect 1482 4825 1488 4941
rect 1168 4812 1488 4825
rect 1220 4760 1488 4812
rect 1168 4747 1488 4760
rect 1220 4695 1488 4747
rect 1168 4682 1488 4695
rect 1220 4630 1488 4682
rect 1168 4617 1488 4630
rect 1220 4565 1488 4617
rect 1168 4552 1488 4565
rect 1220 4500 1488 4552
rect 1168 4487 1488 4500
rect 1220 4435 1488 4487
rect 1168 4422 1488 4435
rect 1220 4370 1488 4422
rect 1168 4357 1488 4370
rect 1220 4305 1488 4357
rect 1168 4292 1488 4305
rect 1220 4240 1488 4292
rect 1168 4227 1488 4240
rect 1220 4175 1488 4227
rect 1168 4162 1488 4175
rect 1220 4110 1488 4162
rect 1168 4097 1488 4110
rect 1220 4045 1488 4097
rect 1168 4032 1488 4045
rect 1220 3980 1488 4032
rect 1168 3967 1488 3980
rect 1220 3915 1488 3967
rect 1168 3902 1488 3915
rect 1220 3850 1488 3902
rect 1168 3837 1488 3850
rect 1220 3785 1488 3837
rect 1168 3771 1488 3785
rect 1220 3719 1488 3771
rect 1168 3705 1488 3719
rect 1220 3653 1488 3705
rect 1168 3639 1488 3653
rect 1220 3587 1488 3639
rect 1168 3573 1488 3587
rect 1220 3521 1488 3573
rect 1168 3507 1488 3521
rect 1220 3455 1488 3507
rect 1168 3441 1488 3455
rect 1220 3389 1488 3441
rect 1168 3375 1488 3389
rect 1220 3323 1488 3375
rect 1168 3309 1488 3323
rect 1220 3257 1488 3309
rect 1168 3243 1488 3257
rect 1220 3191 1488 3243
rect 1168 3177 1488 3191
rect 1220 3125 1488 3177
rect 1168 3111 1488 3125
rect 1220 3059 1488 3111
rect 1168 3045 1488 3059
rect 1220 2993 1488 3045
rect 1168 2975 1488 2993
rect 1220 2923 1232 2975
rect 1284 2923 1296 2975
rect 1348 2923 1360 2975
rect 1412 2923 1424 2975
rect 1476 2923 1488 2975
rect 1168 2908 1488 2923
rect 1220 2856 1232 2908
rect 1284 2856 1296 2908
rect 1348 2856 1360 2908
rect 1412 2856 1424 2908
rect 1476 2856 1488 2908
rect 1168 2841 1488 2856
rect 1220 2789 1232 2841
rect 1284 2789 1296 2841
rect 1348 2789 1360 2841
rect 1412 2789 1424 2841
rect 1476 2789 1488 2841
rect 1168 2518 1488 2789
rect 1220 2466 1232 2518
rect 1284 2466 1296 2518
rect 1348 2466 1360 2518
rect 1412 2466 1424 2518
rect 1476 2466 1488 2518
rect 1168 2429 1488 2466
rect 1220 2377 1232 2429
rect 1284 2377 1296 2429
rect 1348 2377 1360 2429
rect 1412 2377 1424 2429
rect 1476 2377 1488 2429
rect 1168 2340 1488 2377
rect 1220 2288 1232 2340
rect 1284 2288 1296 2340
rect 1348 2288 1360 2340
rect 1412 2288 1424 2340
rect 1476 2288 1488 2340
rect 1168 1858 1488 2288
rect 1168 1806 1180 1858
rect 1232 1806 1244 1858
rect 1296 1806 1308 1858
rect 1360 1806 1372 1858
rect 1424 1806 1436 1858
rect 1168 1792 1488 1806
rect 1516 1929 1568 6827
rect 1516 1863 1568 1877
rect 1596 2000 1648 7704
tri 1648 7679 1673 7704 nw
rect 1596 1934 1648 1948
rect 1685 7511 1691 7563
rect 1743 7511 1758 7563
rect 1810 7511 1816 7563
rect 1685 6563 1737 7511
tri 1737 7486 1762 7511 nw
rect 1848 7483 1976 7784
rect 1848 7431 1854 7483
rect 1906 7431 1918 7483
rect 1970 7431 1976 7483
rect 1848 7131 1976 7431
rect 1848 7079 1854 7131
rect 1906 7079 1918 7131
rect 1970 7079 1976 7131
rect 1848 6779 1976 7079
rect 1848 6727 1854 6779
rect 1906 6727 1918 6779
rect 1970 6727 1976 6779
rect 2004 7659 2504 7879
rect 2004 7607 2010 7659
rect 2062 7607 2083 7659
rect 2135 7607 2156 7659
rect 2208 7607 2229 7659
rect 2281 7607 2302 7659
rect 2354 7607 2374 7659
rect 2426 7607 2446 7659
rect 2498 7607 2504 7659
rect 2004 7307 2504 7607
rect 2004 7255 2010 7307
rect 2062 7255 2083 7307
rect 2135 7255 2156 7307
rect 2208 7255 2229 7307
rect 2281 7255 2302 7307
rect 2354 7255 2374 7307
rect 2426 7255 2446 7307
rect 2498 7255 2504 7307
rect 2783 8205 2789 8257
rect 2841 8205 2859 8257
rect 2911 8205 2930 8257
rect 2982 8205 3001 8257
rect 3053 8205 3059 8257
rect 2783 8193 3059 8205
rect 2783 8141 2789 8193
rect 2841 8141 2859 8193
rect 2911 8141 2930 8193
rect 2982 8141 3001 8193
rect 3053 8141 3059 8193
rect 2783 8129 3059 8141
rect 2783 8077 2789 8129
rect 2841 8077 2859 8129
rect 2911 8077 2930 8129
rect 2982 8077 3001 8129
rect 3053 8077 3059 8129
rect 2783 7912 3059 8077
rect 3381 8077 3387 8257
rect 3567 8077 3573 8257
tri 3915 8223 3949 8257 ne
rect 3949 8239 4368 8257
tri 4368 8239 4386 8257 sw
rect 3949 8223 4386 8239
tri 3949 8205 3967 8223 ne
rect 3967 8205 4386 8223
tri 3967 8193 3979 8205 ne
rect 3979 8193 4386 8205
tri 3979 8186 3986 8193 ne
tri 3381 8019 3439 8077 ne
rect 2783 7860 3007 7912
rect 2783 7846 3059 7860
rect 2783 7794 3007 7846
rect 2783 7780 3059 7794
rect 2783 7728 3007 7780
rect 2783 7714 3059 7728
rect 2783 7662 3007 7714
rect 2783 7649 3059 7662
rect 3439 7951 3573 8077
rect 3439 7899 3445 7951
rect 3497 7899 3515 7951
rect 3567 7899 3573 7951
rect 2783 7597 3007 7649
rect 2783 7475 3059 7597
rect 2783 7423 2937 7475
rect 2989 7423 3001 7475
rect 3053 7423 3059 7475
rect 2783 7415 3051 7423
tri 3051 7415 3059 7423 nw
rect 3091 7607 3097 7659
rect 3149 7607 3161 7659
rect 3213 7607 3225 7659
rect 3277 7607 3289 7659
rect 3341 7607 3353 7659
rect 3405 7607 3411 7659
rect 2783 7387 3023 7415
tri 3023 7387 3051 7415 nw
tri 3063 7387 3091 7415 se
rect 3091 7387 3411 7607
rect 2783 7375 3011 7387
tri 3011 7375 3023 7387 nw
tri 3051 7375 3063 7387 se
rect 3063 7375 3411 7387
rect 2783 7335 2971 7375
tri 2971 7335 3011 7375 nw
tri 3011 7335 3051 7375 se
rect 3051 7335 3411 7375
rect 2783 7307 2943 7335
tri 2943 7307 2971 7335 nw
tri 2983 7307 3011 7335 se
rect 3011 7307 3411 7335
rect 2783 7295 2931 7307
tri 2931 7295 2943 7307 nw
tri 2971 7295 2983 7307 se
rect 2983 7295 3097 7307
rect 2004 6643 2504 7255
tri 2613 7255 2651 7293 sw
rect 2783 7291 2927 7295
tri 2927 7291 2931 7295 nw
tri 2967 7291 2971 7295 se
rect 2971 7291 3097 7295
rect 2783 7255 2891 7291
tri 2891 7255 2927 7291 nw
tri 2931 7255 2967 7291 se
rect 2967 7255 3097 7291
rect 3149 7255 3174 7307
rect 3226 7255 3251 7307
rect 3303 7255 3328 7307
rect 3380 7280 3411 7307
rect 3380 7255 3386 7280
tri 3386 7255 3411 7280 nw
rect 2613 7217 2651 7255
tri 2651 7217 2689 7255 sw
rect 2783 7251 2887 7255
tri 2887 7251 2891 7255 nw
tri 2927 7251 2931 7255 se
rect 2931 7251 3354 7255
tri 2781 7217 2783 7219 se
rect 2783 7217 2853 7251
tri 2853 7217 2887 7251 nw
tri 2893 7217 2927 7251 se
rect 2927 7223 3354 7251
tri 3354 7223 3386 7255 nw
tri 3411 7223 3439 7251 se
rect 3439 7223 3573 7899
rect 3986 7704 4386 8193
rect 4497 8205 4503 8257
rect 4555 8205 4568 8257
rect 4620 8205 4633 8257
rect 4685 8205 4698 8257
rect 4750 8205 4763 8257
rect 4815 8205 4829 8257
rect 4881 8205 4895 8257
rect 4947 8205 4961 8257
rect 5013 8205 5027 8257
rect 5079 8205 5093 8257
rect 5145 8205 5159 8257
rect 5211 8205 5217 8257
rect 4497 8193 5217 8205
rect 4497 8141 4503 8193
rect 4555 8141 4568 8193
rect 4620 8141 4633 8193
rect 4685 8141 4698 8193
rect 4750 8141 4763 8193
rect 4815 8141 4829 8193
rect 4881 8141 4895 8193
rect 4947 8141 4961 8193
rect 5013 8141 5027 8193
rect 5079 8141 5093 8193
rect 5145 8141 5159 8193
rect 5211 8141 5217 8193
rect 4497 8129 5217 8141
rect 4497 8077 4503 8129
rect 4555 8077 4568 8129
rect 4620 8077 4633 8129
rect 4685 8077 4698 8129
rect 4750 8077 4763 8129
rect 4815 8077 4829 8129
rect 4881 8077 4895 8129
rect 4947 8077 4961 8129
rect 5013 8077 5027 8129
rect 5079 8077 5093 8129
rect 5145 8077 5159 8129
rect 5211 8077 5217 8129
rect 3601 7335 3607 7387
rect 3659 7335 3671 7387
rect 3723 7335 3729 7387
tri 3601 7307 3629 7335 ne
rect 2927 7217 3348 7223
tri 3348 7217 3354 7223 nw
tri 3405 7217 3411 7223 se
rect 3411 7217 3573 7223
rect 2004 6591 2010 6643
rect 2062 6591 2083 6643
rect 2135 6591 2156 6643
rect 2208 6591 2229 6643
rect 2281 6591 2302 6643
rect 2354 6591 2374 6643
rect 2426 6591 2446 6643
rect 2498 6591 2504 6643
tri 1737 6563 1762 6588 sw
rect 1685 6511 1691 6563
rect 1743 6511 1758 6563
rect 1810 6511 1816 6563
rect 1685 3922 1737 6511
tri 1737 6486 1762 6511 nw
rect 2004 6503 2504 6591
rect 2561 7165 2567 7217
rect 2619 7165 2631 7217
rect 2683 7165 2689 7217
tri 2729 7165 2781 7217 se
rect 2781 7211 2847 7217
tri 2847 7211 2853 7217 nw
tri 2887 7211 2893 7217 se
rect 2893 7211 3296 7217
rect 2781 7171 2807 7211
tri 2807 7171 2847 7211 nw
tri 2847 7171 2887 7211 se
rect 2887 7171 3296 7211
rect 2781 7165 2801 7171
tri 2801 7165 2807 7171 nw
tri 2841 7165 2847 7171 se
rect 2847 7165 3296 7171
tri 3296 7165 3348 7217 nw
tri 3353 7165 3405 7217 se
rect 3405 7165 3411 7217
rect 3463 7165 3514 7217
rect 3566 7165 3573 7217
rect 2561 7147 2671 7165
tri 2671 7147 2689 7165 nw
tri 2711 7147 2729 7165 se
rect 2729 7147 2783 7165
tri 2783 7147 2801 7165 nw
tri 2823 7147 2841 7165 se
rect 2841 7160 3291 7165
tri 3291 7160 3296 7165 nw
tri 3348 7160 3353 7165 se
rect 3353 7160 3573 7165
rect 2841 7147 3240 7160
rect 2561 7117 2641 7147
tri 2641 7117 2671 7147 nw
tri 2681 7117 2711 7147 se
rect 2711 7117 2713 7147
rect 2561 6503 2613 7117
tri 2613 7089 2641 7117 nw
tri 2653 7089 2681 7117 se
rect 2681 7089 2713 7117
tri 2641 7077 2653 7089 se
rect 2653 7077 2713 7089
tri 2713 7077 2783 7147 nw
tri 2807 7131 2823 7147 se
rect 2823 7131 3240 7147
rect 2807 7109 3240 7131
tri 3240 7109 3291 7160 nw
tri 3297 7109 3348 7160 se
rect 3348 7109 3573 7160
rect 2641 6503 2693 7077
tri 2693 7057 2713 7077 nw
rect 2807 7052 3183 7109
tri 3183 7052 3240 7109 nw
tri 3240 7052 3297 7109 se
rect 3297 7058 3573 7109
rect 3297 7052 3481 7058
rect 2807 6503 3126 7052
tri 3126 6995 3183 7052 nw
tri 3183 6995 3240 7052 se
rect 3240 6995 3481 7052
tri 3154 6966 3183 6995 se
rect 3183 6966 3481 6995
tri 3481 6966 3573 7058 nw
rect 3154 6878 3431 6966
tri 3431 6916 3481 6966 nw
rect 3154 6826 3163 6878
rect 3215 6826 3233 6878
rect 3285 6826 3303 6878
rect 3355 6826 3373 6878
rect 3425 6826 3431 6878
rect 3154 6643 3431 6826
rect 3154 6591 3163 6643
rect 3215 6591 3233 6643
rect 3285 6591 3303 6643
rect 3355 6591 3373 6643
rect 3425 6591 3431 6643
rect 3154 6503 3206 6591
tri 3206 6566 3231 6591 nw
rect 3629 6503 3681 7335
tri 3681 7287 3729 7335 nw
rect 4497 6867 5217 8077
tri 4497 6563 4801 6867 ne
rect 4801 6563 5217 6867
rect 4433 6511 4439 6563
rect 4491 6511 4503 6563
rect 4555 6511 4561 6563
tri 4801 6511 4853 6563 ne
rect 4853 6511 5217 6563
rect 4433 6486 4485 6511
tri 4485 6486 4510 6511 nw
tri 4853 6503 4861 6511 ne
rect 4861 6503 5217 6511
rect 1685 3856 1737 3870
rect 1685 2062 1737 3804
rect 1685 1996 1737 2010
rect 1685 1938 1737 1944
rect 1596 1876 1648 1882
rect 1516 1805 1568 1811
rect 1168 1740 1180 1792
rect 1232 1740 1244 1792
rect 1296 1740 1308 1792
rect 1360 1740 1372 1792
rect 1424 1740 1436 1792
rect 1168 1728 1488 1740
rect 1220 1676 1488 1728
rect 1168 1659 1488 1676
rect 1220 1607 1488 1659
rect 1168 1590 1488 1607
rect 1220 1538 1488 1590
rect 1168 1521 1488 1538
rect 1220 1469 1488 1521
rect 1168 1452 1488 1469
rect 1220 1400 1488 1452
rect 1168 1383 1488 1400
rect 1220 1331 1488 1383
rect 1168 1314 1488 1331
rect 1220 1262 1488 1314
rect 1168 1246 1488 1262
rect 1220 1194 1488 1246
rect 1168 1098 1488 1194
rect 1220 1046 1488 1098
rect 1168 1029 1488 1046
rect 1220 977 1488 1029
rect 1168 960 1488 977
rect 1220 908 1488 960
rect 1168 891 1488 908
rect 1220 839 1488 891
rect 1168 822 1488 839
rect 1220 770 1488 822
rect 1168 754 1488 770
rect 1220 702 1488 754
rect 1168 686 1488 702
rect 1220 634 1488 686
rect 1168 618 1488 634
rect 1220 566 1488 618
rect 1168 550 1488 566
rect 1220 498 1488 550
rect 1168 482 1488 498
rect 1220 430 1488 482
rect 1168 414 1488 430
rect 1220 362 1488 414
rect 1168 346 1488 362
rect 1220 294 1488 346
rect 1168 278 1488 294
rect 1220 226 1488 278
rect 1168 210 1488 226
rect 1220 158 1488 210
rect 1168 112 1488 158
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_0
timestamp 1704896540
transform 0 1 -12 1 0 4340
box 0 0 1 1
use DFL1_CDNS_5246887918578  DFL1_CDNS_5246887918578_1
timestamp 1704896540
transform 0 -1 -182 1 0 4340
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_0
timestamp 1704896540
transform 1 0 701 0 -1 858
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_1
timestamp 1704896540
transform 1 0 403 0 -1 4880
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_2
timestamp 1704896540
transform 1 0 -26 0 1 4348
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_3
timestamp 1704896540
transform 1 0 -194 0 1 4348
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1704896540
transform 0 1 403 -1 0 6281
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1704896540
transform 0 1 403 -1 0 6713
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1704896540
transform -1 0 1243 0 1 5546
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1704896540
transform -1 0 1039 0 1 5885
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_4
timestamp 1704896540
transform -1 0 1039 0 1 5435
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_5
timestamp 1704896540
transform -1 0 1243 0 1 5885
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_6
timestamp 1704896540
transform -1 0 594 0 1 1358
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_7
timestamp 1704896540
transform 0 1 1309 1 0 5403
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_8
timestamp 1704896540
transform 1 0 331 0 -1 4642
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_9
timestamp 1704896540
transform 1 0 783 0 -1 4642
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_10
timestamp 1704896540
transform 1 0 331 0 -1 5074
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_11
timestamp 1704896540
transform 1 0 854 0 -1 5580
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_12
timestamp 1704896540
transform 1 0 309 0 1 6011
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_13
timestamp 1704896540
transform 1 0 229 0 1 5114
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1704896540
transform 1 0 -172 0 1 292
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_0
timestamp 1704896540
transform -1 0 738 0 -1 1406
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_1
timestamp 1704896540
transform 0 -1 735 1 0 1056
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_2
timestamp 1704896540
transform 0 -1 519 1 0 1089
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_3
timestamp 1704896540
transform 0 -1 519 1 0 4314
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_4
timestamp 1704896540
transform 0 -1 519 1 0 4523
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_5
timestamp 1704896540
transform 0 -1 519 1 0 6121
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1704896540
transform 0 -1 744 -1 0 864
box 0 0 1 1
use M1M2_CDNS_52468879185200  M1M2_CDNS_52468879185200_0
timestamp 1704896540
transform 1 0 547 0 1 8077
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_0
timestamp 1704896540
transform 1 0 381 0 -1 1258
box 0 0 1 1
use M1M2_CDNS_52468879185970  M1M2_CDNS_52468879185970_0
timestamp 1704896540
transform -1 0 540 0 -1 1398
box 0 0 1 1
use M1M2_CDNS_52468879185970  M1M2_CDNS_52468879185970_1
timestamp 1704896540
transform 0 -1 744 1 0 1040
box 0 0 1 1
use M1M2_CDNS_52468879185970  M1M2_CDNS_52468879185970_2
timestamp 1704896540
transform 0 -1 744 1 0 1366
box 0 0 1 1
use M1M2_CDNS_52468879185970  M1M2_CDNS_52468879185970_3
timestamp 1704896540
transform 0 -1 528 1 0 1073
box 0 0 1 1
use nfet_CDNS_524688791851356  nfet_CDNS_524688791851356_0
timestamp 1704896540
transform 0 1 161 -1 0 3833
box -79 -26 279 226
use nfet_CDNS_524688791851356  nfet_CDNS_524688791851356_1
timestamp 1704896540
transform 0 1 161 -1 0 3211
box -79 -26 279 226
use nfet_CDNS_524688791851356  nfet_CDNS_524688791851356_2
timestamp 1704896540
transform 0 1 161 -1 0 2589
box -79 -26 279 226
use nfet_CDNS_524688791851356  nfet_CDNS_524688791851356_3
timestamp 1704896540
transform 0 1 161 1 0 3267
box -79 -26 279 226
use nfet_CDNS_524688791851356  nfet_CDNS_524688791851356_4
timestamp 1704896540
transform 0 1 161 1 0 2645
box -79 -26 279 226
use nfet_CDNS_524688791851357  nfet_CDNS_524688791851357_0
timestamp 1704896540
transform 0 1 161 -1 0 6715
box -79 -26 335 226
use nfet_CDNS_524688791851358  nfet_CDNS_524688791851358_0
timestamp 1704896540
transform 0 1 161 -1 0 795
box -79 -26 575 226
use nfet_CDNS_524688791851359  nfet_CDNS_524688791851359_0
timestamp 1704896540
transform 0 1 161 -1 0 5751
box -79 -26 455 226
use nfet_CDNS_524688791851360  nfet_CDNS_524688791851360_0
timestamp 1704896540
transform 0 1 3183 -1 0 7781
box -79 -26 727 626
use nfet_CDNS_524688791851361  nfet_CDNS_524688791851361_0
timestamp 1704896540
transform 0 1 3183 -1 0 7077
box -79 -26 375 626
use nfet_CDNS_524688791851362  nfet_CDNS_524688791851362_0
timestamp 1704896540
transform 0 1 161 -1 0 6077
box -79 -26 239 226
use nfet_CDNS_524688791851362  nfet_CDNS_524688791851362_1
timestamp 1704896540
transform 0 1 161 1 0 6133
box -79 -26 239 226
use nfet_CDNS_524688791851363  nfet_CDNS_524688791851363_0
timestamp 1704896540
transform 0 1 161 1 0 851
box -79 -26 299 226
use nfet_CDNS_524688791851364  nfet_CDNS_524688791851364_0
timestamp 1704896540
transform 0 1 161 -1 0 4455
box -79 -26 279 226
use nfet_CDNS_524688791851365  nfet_CDNS_524688791851365_0
timestamp 1704896540
transform 0 1 161 -1 0 4887
box -79 -26 455 226
use nfet_CDNS_524688791851366  nfet_CDNS_524688791851366_0
timestamp 1704896540
transform 0 1 161 1 0 3889
box -79 -26 279 226
use nfet_CDNS_524688791851367  nfet_CDNS_524688791851367_0
timestamp 1704896540
transform 0 -1 46 -1 0 4337
box -79 -26 4079 110
use nfet_CDNS_524688791851368  nfet_CDNS_524688791851368_0
timestamp 1704896540
transform 0 1 161 -1 0 5319
box -79 -26 455 226
use nfet_CDNS_524688791851369  nfet_CDNS_524688791851369_0
timestamp 1704896540
transform 0 1 161 1 0 1237
box -79 -26 129 226
use nfet_CDNS_524688791851370  nfet_CDNS_524688791851370_0
timestamp 1704896540
transform 0 1 -240 -1 0 4337
box -79 -26 4079 110
use nfet_CDNS_524688791851371  nfet_CDNS_524688791851371_0
timestamp 1704896540
transform 0 1 161 1 0 1453
box -79 -26 129 226
use nfet_CDNS_524688791851372  nfet_CDNS_524688791851372_0
timestamp 1704896540
transform 0 1 161 -1 0 1609
box -79 -26 129 226
use pfet_CDNS_524688791851373  pfet_CDNS_524688791851373_0
timestamp 1704896540
transform 0 -1 1065 -1 0 3833
box -119 -66 319 266
use pfet_CDNS_524688791851373  pfet_CDNS_524688791851373_1
timestamp 1704896540
transform 0 -1 1065 1 0 3889
box -119 -66 319 266
use pfet_CDNS_524688791851373  pfet_CDNS_524688791851373_2
timestamp 1704896540
transform 0 -1 1065 1 0 3267
box -119 -66 319 266
use pfet_CDNS_524688791851374  pfet_CDNS_524688791851374_0
timestamp 1704896540
transform 0 1 835 -1 0 6831
box -119 -66 279 266
use pfet_CDNS_524688791851374  pfet_CDNS_524688791851374_1
timestamp 1704896540
transform 0 1 835 1 0 6887
box -119 -66 279 266
use pfet_CDNS_524688791851374  pfet_CDNS_524688791851374_2
timestamp 1704896540
transform 0 -1 1065 1 0 4511
box -119 -66 279 266
use pfet_CDNS_524688791851375  pfet_CDNS_524688791851375_0
timestamp 1704896540
transform 0 1 835 1 0 7213
box -119 -66 375 366
use pfet_CDNS_524688791851376  pfet_CDNS_524688791851376_0
timestamp 1704896540
transform 0 -1 1065 1 0 299
box -89 -36 585 236
use pfet_CDNS_524688791851379  pfet_CDNS_524688791851379_0
timestamp 1704896540
transform 0 -1 1065 1 0 1449
box -89 -36 139 236
use pfet_CDNS_524688791851380  pfet_CDNS_524688791851380_0
timestamp 1704896540
transform 0 -1 1065 -1 0 1605
box -89 -36 139 236
use pfet_CDNS_524688791851381  pfet_CDNS_524688791851381_0
timestamp 1704896540
transform 0 1 1373 1 0 7133
box -119 -66 767 666
use pfet_CDNS_524688791851381  pfet_CDNS_524688791851381_1
timestamp 1704896540
transform 0 1 2103 1 0 7133
box -119 -66 767 666
use pfet_CDNS_524688791851382  pfet_CDNS_524688791851382_0
timestamp 1704896540
transform 0 1 1373 1 0 6781
box -119 -66 415 666
use pfet_CDNS_524688791851382  pfet_CDNS_524688791851382_1
timestamp 1704896540
transform 0 1 2103 1 0 6781
box -119 -66 415 666
use pfet_CDNS_524688791851383  pfet_CDNS_524688791851383_0
timestamp 1704896540
transform 0 1 835 1 0 7525
box -119 -66 375 366
use pfet_CDNS_524688791851384  pfet_CDNS_524688791851384_0
timestamp 1704896540
transform 0 -1 1065 1 0 851
box -89 -36 309 236
use pfet_CDNS_524688791851385  pfet_CDNS_524688791851385_0
timestamp 1704896540
transform 0 -1 1065 -1 0 4455
box -119 -66 319 266
use pfet_CDNS_524688791851385  pfet_CDNS_524688791851385_1
timestamp 1704896540
transform 0 -1 1065 -1 0 3211
box -119 -66 319 266
use pfet_CDNS_524688791851386  pfet_CDNS_524688791851386_0
timestamp 1704896540
transform 0 1 1129 -1 0 5871
box -89 -36 489 146
use pfet_CDNS_524688791851386  pfet_CDNS_524688791851386_1
timestamp 1704896540
transform 0 1 925 -1 0 5871
box -89 -36 489 146
use pfet_CDNS_524688791851388  pfet_CDNS_524688791851388_0
timestamp 1704896540
transform 0 -1 1065 -1 0 1393
box -89 -36 245 236
use pfet_CDNS_524688791851389  pfet_CDNS_524688791851389_0
timestamp 1704896540
transform 0 -1 1065 -1 0 2589
box -119 -66 319 266
use pfet_CDNS_524688791851389  pfet_CDNS_524688791851389_1
timestamp 1704896540
transform 0 -1 1065 1 0 2645
box -119 -66 319 266
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_0
timestamp 1704896540
transform 0 1 699 -1 0 1501
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185315  sky130_fd_io__tk_em1o_CDNS_52468879185315_0
timestamp 1704896540
transform 0 -1 664 -1 0 2875
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185315  sky130_fd_io__tk_em1o_CDNS_52468879185315_1
timestamp 1704896540
transform 0 -1 117 -1 0 2876
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185315  sky130_fd_io__tk_em1o_CDNS_52468879185315_2
timestamp 1704896540
transform 0 1 393 -1 0 5272
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185315  sky130_fd_io__tk_em1o_CDNS_52468879185315_3
timestamp 1704896540
transform 0 1 612 -1 0 4121
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185315  sky130_fd_io__tk_em1o_CDNS_52468879185315_4
timestamp 1704896540
transform 0 1 612 -1 0 3498
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185315  sky130_fd_io__tk_em1o_CDNS_52468879185315_5
timestamp 1704896540
transform 0 1 65 -1 0 3498
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185315  sky130_fd_io__tk_em1o_CDNS_52468879185315_6
timestamp 1704896540
transform 0 1 612 1 0 3602
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185315  sky130_fd_io__tk_em1o_CDNS_52468879185315_7
timestamp 1704896540
transform 0 1 65 1 0 2358
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185315  sky130_fd_io__tk_em1o_CDNS_52468879185315_8
timestamp 1704896540
transform 0 -1 664 1 0 4223
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185315  sky130_fd_io__tk_em1o_CDNS_52468879185315_9
timestamp 1704896540
transform 0 -1 664 1 0 2980
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185315  sky130_fd_io__tk_em1o_CDNS_52468879185315_10
timestamp 1704896540
transform 0 -1 117 1 0 3602
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185315  sky130_fd_io__tk_em1o_CDNS_52468879185315_11
timestamp 1704896540
transform 0 -1 117 1 0 2980
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185340  sky130_fd_io__tk_em1o_CDNS_52468879185340_0
timestamp 1704896540
transform -1 0 234 0 1 4094
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185340  sky130_fd_io__tk_em1o_CDNS_52468879185340_1
timestamp 1704896540
transform 0 -1 823 1 0 4247
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185340  sky130_fd_io__tk_em1o_CDNS_52468879185340_2
timestamp 1704896540
transform 1 0 90 0 1 5108
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_524688791851353  sky130_fd_io__tk_em1o_CDNS_524688791851353_0
timestamp 1704896540
transform 1 0 -5 0 -1 386
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185314  sky130_fd_io__tk_em1s_CDNS_52468879185314_0
timestamp 1704896540
transform 0 1 65 -1 0 4399
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185314  sky130_fd_io__tk_em1s_CDNS_52468879185314_1
timestamp 1704896540
transform 0 1 393 -1 0 5704
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185314  sky130_fd_io__tk_em1s_CDNS_52468879185314_2
timestamp 1704896540
transform -1 0 234 0 1 4224
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185341  sky130_fd_io__tk_em1s_CDNS_52468879185341_0
timestamp 1704896540
transform -1 0 963 0 1 4204
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_524688791851354  sky130_fd_io__tk_em1s_CDNS_524688791851354_0
timestamp 1704896540
transform 0 1 612 -1 0 2363
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_524688791851355  sky130_fd_io__tk_em1s_CDNS_524688791851355_0
timestamp 1704896540
transform 0 -1 253 -1 0 4393
box 0 0 1 1
<< labels >>
flabel comment s 109 5963 109 5963 0 FreeSans 200 0 0 0 sio_diff_hyst_en_h
flabel comment s 1469 6470 1469 6470 0 FreeSans 200 0 0 0 m1_float
flabel comment s 950 2112 950 2112 0 FreeSans 200 0 0 0 vpwr_ka
flabel comment s 940 6243 940 6243 0 FreeSans 200 0 0 0 vpwr_ka
flabel comment s 940 7967 940 7967 0 FreeSans 200 0 0 0 vpwr_ka
flabel comment s 1343 1478 1343 1478 0 FreeSans 200 0 0 0 vpb_ka
flabel comment s 1388 4384 1388 4384 0 FreeSans 200 0 0 0 vpb_ka
flabel comment s 1310 7954 1310 7954 0 FreeSans 200 0 0 0 vpb_ka
flabel comment s 1310 6229 1310 6229 0 FreeSans 200 0 0 0 vpb_ka
flabel comment s -200 1925 -200 1925 0 FreeSans 200 0 0 0 out_h_n
flabel comment s 1146 1925 1146 1925 0 FreeSans 200 0 0 0 out_h_n
flabel comment s 1548 2419 1548 2419 0 FreeSans 200 270 0 0 out_h_n
flabel comment s 1551 4385 1551 4385 0 FreeSans 200 270 0 0 out_h_n
flabel comment s 1550 6161 1550 6161 0 FreeSans 200 270 0 0 out_h_n
flabel comment s 1629 6166 1629 6166 0 FreeSans 200 270 0 0 ie_diff_sel_h_n
flabel comment s 1629 4385 1629 4385 0 FreeSans 200 270 0 0 ie_diff_sel_h_n
flabel comment s 1631 2409 1631 2409 0 FreeSans 200 270 0 0 ie_diff_sel_h_n
flabel comment s 1153 1986 1153 1986 0 FreeSans 200 180 0 0 ie_diff_sel_h_n
flabel comment s 1143 2045 1143 2045 0 FreeSans 200 180 0 0 ie_diff_sel_h
flabel comment s 1718 2421 1718 2421 0 FreeSans 200 90 0 0 ie_diff_sel_h
flabel comment s 1710 4394 1710 4394 0 FreeSans 200 90 0 0 ie_diff_sel_h
flabel comment s 1712 6172 1712 6172 0 FreeSans 200 90 0 0 ie_diff_sel_h
flabel comment s -753 4186 -753 4186 0 FreeSans 200 0 0 0 vgnd
flabel comment s -751 1238 -751 1238 0 FreeSans 200 0 0 0 vgnd
flabel comment s -733 2002 -733 2002 0 FreeSans 200 0 0 0 vgnd
flabel comment s 719 6348 719 6348 0 FreeSans 400 270 0 0 m1_int<4>
flabel comment s 254 6312 254 6312 0 FreeSans 400 180 0 0 int<4>
flabel comment s 402 5058 402 5058 0 FreeSans 400 0 0 0 int<5>
flabel comment s 278 5583 278 5583 0 FreeSans 400 0 0 0 int<9>
flabel comment s 419 4401 419 4401 0 FreeSans 400 180 0 0 int<8>
flabel comment s 837 4401 837 4401 0 FreeSans 400 180 0 0 int<8>
flabel comment s 906 2267 906 2267 0 FreeSans 400 0 0 0 lv_net
flabel comment s 741 6348 741 6348 0 FreeSans 400 270 0 0 m2_int<5>
flabel comment s 229 5877 229 5877 0 FreeSans 400 180 0 0 int<5>
flabel comment s 713 2733 713 2733 0 FreeSans 400 90 0 0 lv_net
flabel comment s 713 3328 713 3328 0 FreeSans 400 90 0 0 lv_net
flabel comment s 716 3888 716 3888 0 FreeSans 400 90 0 0 lv_net
flabel comment s 709 4352 709 4352 0 FreeSans 400 90 0 0 lv_net
flabel comment s 936 4786 936 4786 0 FreeSans 400 180 0 0 lv_net
flabel comment s -144 4829 -144 4829 0 FreeSans 400 180 0 0 int<1>
flabel comment s -52 4680 -52 4680 0 FreeSans 400 180 0 0 int<3>
flabel comment s 1132 6985 1132 6985 0 FreeSans 400 270 0 0 int<4>
flabel comment s 923 7053 923 7053 0 FreeSans 400 180 0 0 int<5>
flabel comment s 923 6614 923 6614 0 FreeSans 400 180 0 0 int<4>
flabel comment s 1131 6767 1131 6767 0 FreeSans 400 270 0 0 int<1>
flabel comment s 642 5354 642 5354 0 FreeSans 400 90 0 0 int<1>
flabel comment s 579 5399 579 5399 0 FreeSans 400 270 0 0 ie_diff_sel_n
flabel comment s 650 1938 650 1938 0 FreeSans 400 270 0 0 ie_diff_dly_n
flabel comment s 888 6855 888 6855 0 FreeSans 400 180 0 0 vcc_io
flabel comment s 613 4228 613 4228 0 FreeSans 400 0 0 0 invout<1>
flabel comment s 592 4122 592 4122 0 FreeSans 400 0 0 0 invout<2>
flabel comment s 594 3610 594 3610 0 FreeSans 400 0 0 0 invout<3>
flabel comment s 562 3499 562 3499 0 FreeSans 400 0 0 0 invout<4>
flabel comment s 562 2985 562 2985 0 FreeSans 400 0 0 0 invout<5>
flabel comment s 562 2879 562 2879 0 FreeSans 400 0 0 0 invout<6>
flabel comment s 602 2364 602 2364 0 FreeSans 400 0 0 0 invout<7>
flabel comment s 579 1981 579 1981 0 FreeSans 400 270 0 0 ie_diff_sel_n
flabel comment s 292 6569 292 6569 0 FreeSans 400 180 0 0 int<1>
flabel comment s 784 4586 784 4586 0 FreeSans 400 90 0 0 int<1>
flabel comment s 447 4765 447 4765 0 FreeSans 400 90 0 0 int<1>
flabel comment s 447 5996 447 5996 0 FreeSans 400 90 0 0 int<4>
flabel comment s 447 6215 447 6215 0 FreeSans 400 90 0 0 int<1>
flabel comment s 3772 6474 3772 6474 0 FreeSans 200 0 0 0 sio_diff_hyst_en_h
flabel comment s 1545 6096 1545 6096 0 FreeSans 200 0 0 0 sio_diff_hyst_en_h
flabel comment s 736 5712 736 5712 0 FreeSans 400 270 0 0 int<5>
flabel comment s 975 7325 975 7325 0 FreeSans 400 180 0 0 int<1>
flabel comment s 270 5109 270 5109 0 FreeSans 400 0 0 0 int<6>
flabel comment s 447 5573 447 5573 0 FreeSans 400 270 0 0 int<4>
flabel comment s 445 5148 445 5148 0 FreeSans 400 270 0 0 int<5>
flabel comment s 3095 7384 3095 7384 0 FreeSans 400 270 0 0 ie_diff_sel_h
flabel comment s 2061 7536 2061 7536 0 FreeSans 400 90 0 0 ie_diff_sel_h_n
flabel comment s 2059 6948 2059 6948 0 FreeSans 400 90 0 0 out_hv
flabel comment s 790 973 790 973 0 FreeSans 400 90 0 0 out_lv
flabel comment s 233 2596 233 2596 0 FreeSans 400 180 0 0 vgnd
flabel comment s 233 3841 233 3841 0 FreeSans 400 180 0 0 vgnd
flabel comment s 256 4515 256 4515 0 FreeSans 400 180 0 0 vgnd
flabel comment s 1123 4476 1123 4476 0 FreeSans 400 180 0 0 vpwr
flabel comment s 1123 3851 1123 3851 0 FreeSans 400 180 0 0 vpwr
flabel comment s 233 3217 233 3217 0 FreeSans 400 180 0 0 vgnd
flabel comment s 105 4907 105 4907 0 FreeSans 400 180 0 0 vgnd
flabel comment s 2960 6935 2960 6935 0 FreeSans 400 0 0 0 out_h_n
flabel comment s 177 6663 177 6663 0 FreeSans 200 0 0 0 ie_diff_sel_n
flabel comment s 874 5420 874 5420 0 FreeSans 400 0 0 0 int<6>
flabel comment s 218 5343 218 5343 0 FreeSans 400 180 0 0 vgnd
flabel comment s 593 1647 593 1647 0 FreeSans 400 180 0 0 ie_diff_dly_n
flabel comment s 586 1439 586 1439 0 FreeSans 400 180 0 0 ie_diff_sel_n
flabel comment s 342 1321 342 1321 0 FreeSans 400 0 0 0 int<11>
flabel comment s 804 550 804 550 0 FreeSans 400 90 0 0 int<11>
flabel comment s 431 550 431 550 0 FreeSans 400 90 0 0 int<10>
flabel comment s 436 973 436 973 0 FreeSans 400 90 0 0 out_lv
flabel comment s 319 1542 319 1542 0 FreeSans 400 0 0 0 int<10>
flabel comment s 259 1204 259 1204 0 FreeSans 400 180 0 0 vgnd
flabel comment s 100 1626 100 1626 0 FreeSans 400 180 0 0 vgnd
flabel comment s 246 1401 246 1401 0 FreeSans 400 180 0 0 vgnd
flabel comment s 1002 1528 1002 1528 0 FreeSans 400 0 0 0 int1_nor
flabel comment s 986 1321 986 1321 0 FreeSans 400 0 0 0 int<11>
flabel comment s 1108 1191 1108 1191 0 FreeSans 400 180 0 0 vpwr
flabel comment s 1108 1406 1108 1406 0 FreeSans 400 180 0 0 vpwr
flabel comment s 993 1624 993 1624 0 FreeSans 400 180 0 0 int<10>
flabel comment s 933 716 933 716 0 FreeSans 400 180 0 0 vpwr
flabel comment s 116 484 116 484 0 FreeSans 400 270 0 0 en_lv_inv_n1
flabel comment s 1132 712 1132 712 0 FreeSans 400 270 0 0 en_lv_inv_n0
flabel comment s 1286 5674 1286 5674 0 FreeSans 400 270 0 0 int<6>
flabel comment s 913 5658 913 5658 0 FreeSans 400 270 0 0 int<9>
flabel comment s 1194 5419 1194 5419 0 FreeSans 400 0 0 0 int<9>
flabel comment s 218 5770 218 5770 0 FreeSans 400 180 0 0 vgnd
flabel comment s 933 539 933 539 0 FreeSans 400 180 0 0 vpwr
flabel comment s 933 347 933 347 0 FreeSans 400 180 0 0 vpwr
flabel comment s 438 6683 438 6683 0 FreeSans 400 270 0 0 ie_diff_sel_n
flabel comment s -113 3426 -113 3426 0 FreeSans 400 90 0 0 int<3>
flabel comment s 1123 3217 1123 3217 0 FreeSans 400 180 0 0 vpwr
flabel comment s 1123 2596 1123 2596 0 FreeSans 400 180 0 0 vpwr
flabel comment s -196 4398 -196 4398 0 FreeSans 400 0 0 0 int<1>
flabel comment s 3332 7618 3332 7618 0 FreeSans 400 180 0 0 vgnd
flabel comment s 1793 7281 1793 7281 0 FreeSans 400 180 0 0 vcc_io
flabel comment s 1793 7613 1793 7613 0 FreeSans 400 180 0 0 vcc_io
flabel comment s 3332 7267 3332 7267 0 FreeSans 400 180 0 0 vgnd
flabel comment s 984 7643 984 7643 0 FreeSans 400 180 0 0 vcc_io
flabel comment s 956 7805 956 7805 0 FreeSans 400 180 0 0 int<0>
flabel comment s 937 7493 937 7493 0 FreeSans 400 180 0 0 int<0>
flabel comment s 942 7173 942 7173 0 FreeSans 400 180 0 0 int<0>
flabel comment s 22 4446 22 4446 0 FreeSans 400 0 0 0 vgnd
flabel metal1 s -311 1535 -273 1581 7 FreeSans 400 0 0 0 out_h_n
port 8 nsew
flabel metal1 s -196 1972 -153 2006 3 FreeSans 400 0 0 0 ie_diff_sel_h_n
port 2 nsew
flabel metal1 s 1665 2141 1691 2208 7 FreeSans 400 0 0 0 ie_diff_dly_n
port 3 nsew
flabel metal1 s 1676 5335 1695 5377 7 FreeSans 400 0 0 0 ie_diff_n
port 4 nsew
flabel metal1 s 1649 2783 1695 2987 3 FreeSans 400 180 0 0 vpb_ka
port 5 nsew
flabel metal1 s 1649 3206 1695 3532 3 FreeSans 400 180 0 0 vpb_ka
port 5 nsew
flabel metal1 s -33 904 4 944 7 FreeSans 400 0 0 0 out_n
port 7 nsew
flabel metal1 s -112 2034 -69 2068 3 FreeSans 400 0 0 0 ie_diff_sel_h
port 6 nsew
flabel metal1 s 1665 1132 1695 1160 7 FreeSans 400 0 0 0 out_lv
port 9 nsew
flabel metal1 s 1685 3798 1737 3832 3 FreeSans 400 270 0 0 ie_diff_sel_h
port 6 nsew
flabel metal1 s 1685 2034 1737 2068 3 FreeSans 400 270 0 0 ie_diff_sel_h
port 6 nsew
flabel metal1 s 1652 1287 1695 1333 7 FreeSans 400 0 0 0 ie_diff_sel_h_n
port 2 nsew
flabel metal2 s 2641 6503 2693 6539 0 FreeSans 400 0 0 0 vgnd
port 10 nsew
flabel metal2 s 3154 6503 3206 6539 0 FreeSans 400 0 0 0 vgnd
port 10 nsew
flabel metal2 s 476 112 528 158 0 FreeSans 400 0 0 0 vgnd
port 10 nsew
flabel metal2 s 1106 8863 1426 8909 0 FreeSans 400 0 0 0 vpb_ka
port 5 nsew
flabel metal2 s 630 8863 950 8909 0 FreeSans 400 0 0 0 vpwr_ka
port 11 nsew
flabel metal2 s 145 112 347 158 0 FreeSans 400 0 0 0 vgnd
port 10 nsew
flabel metal2 s 2004 6503 2504 6539 0 FreeSans 400 0 0 0 vcc_io
port 12 nsew
flabel metal2 s 2807 6503 3126 6539 0 FreeSans 400 0 0 0 vgnd
port 10 nsew
flabel metal2 s 692 112 744 158 0 FreeSans 400 90 0 0 vpb_ka
port 5 nsew
flabel metal2 s 2561 6503 2613 6539 0 FreeSans 400 90 0 0 out_hv
port 13 nsew
flabel metal2 s 3629 6503 3681 6539 0 FreeSans 400 0 0 0 pcasc
port 14 nsew
<< properties >>
string GDS_END 86199234
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86002098
string path 5.075 45.350 8.675 45.350 
<< end >>
