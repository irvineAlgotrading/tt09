magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< dnwell >>
tri -700 6714 -614 6800 se
rect -614 6714 764 6800
tri 764 6714 850 6800 sw
rect -700 -714 850 6714
tri -700 -800 -614 -714 ne
rect -614 -800 764 -714
tri 764 -800 850 -714 nw
<< nwell >>
rect -10 0 160 6000
<< pwell >>
rect -1166 7074 1316 7208
rect -1166 6026 -1032 7074
rect 1182 6026 1316 7074
rect -1166 -26 -574 6026
rect 724 -26 1316 6026
rect -1166 -1074 -1032 -26
rect 1182 -1074 1316 -26
rect -1166 -1208 1316 -1074
<< mvnmos >>
rect -900 0 -730 6000
rect 880 0 1050 6000
<< mvnnmos >>
rect -730 0 -600 6000
rect 750 0 880 6000
<< mvndiff >>
rect -958 5975 -900 6000
rect -958 5941 -946 5975
rect -912 5941 -900 5975
rect -958 5907 -900 5941
rect -958 5873 -946 5907
rect -912 5873 -900 5907
rect -958 5839 -900 5873
rect -958 5805 -946 5839
rect -912 5805 -900 5839
rect -958 5771 -900 5805
rect -958 5737 -946 5771
rect -912 5737 -900 5771
rect -958 5703 -900 5737
rect -958 5669 -946 5703
rect -912 5669 -900 5703
rect -958 5635 -900 5669
rect -958 5601 -946 5635
rect -912 5601 -900 5635
rect -958 5567 -900 5601
rect -958 5533 -946 5567
rect -912 5533 -900 5567
rect -958 5499 -900 5533
rect -958 5465 -946 5499
rect -912 5465 -900 5499
rect -958 5431 -900 5465
rect -958 5397 -946 5431
rect -912 5397 -900 5431
rect -958 5363 -900 5397
rect -958 5329 -946 5363
rect -912 5329 -900 5363
rect -958 5295 -900 5329
rect -958 5261 -946 5295
rect -912 5261 -900 5295
rect -958 5227 -900 5261
rect -958 5193 -946 5227
rect -912 5193 -900 5227
rect -958 5159 -900 5193
rect -958 5125 -946 5159
rect -912 5125 -900 5159
rect -958 5091 -900 5125
rect -958 5057 -946 5091
rect -912 5057 -900 5091
rect -958 5023 -900 5057
rect -958 4989 -946 5023
rect -912 4989 -900 5023
rect -958 4955 -900 4989
rect -958 4921 -946 4955
rect -912 4921 -900 4955
rect -958 4887 -900 4921
rect -958 4853 -946 4887
rect -912 4853 -900 4887
rect -958 4819 -900 4853
rect -958 4785 -946 4819
rect -912 4785 -900 4819
rect -958 4751 -900 4785
rect -958 4717 -946 4751
rect -912 4717 -900 4751
rect -958 4683 -900 4717
rect -958 4649 -946 4683
rect -912 4649 -900 4683
rect -958 4615 -900 4649
rect -958 4581 -946 4615
rect -912 4581 -900 4615
rect -958 4547 -900 4581
rect -958 4513 -946 4547
rect -912 4513 -900 4547
rect -958 4479 -900 4513
rect -958 4445 -946 4479
rect -912 4445 -900 4479
rect -958 4411 -900 4445
rect -958 4377 -946 4411
rect -912 4377 -900 4411
rect -958 4343 -900 4377
rect -958 4309 -946 4343
rect -912 4309 -900 4343
rect -958 4275 -900 4309
rect -958 4241 -946 4275
rect -912 4241 -900 4275
rect -958 4207 -900 4241
rect -958 4173 -946 4207
rect -912 4173 -900 4207
rect -958 4139 -900 4173
rect -958 4105 -946 4139
rect -912 4105 -900 4139
rect -958 4071 -900 4105
rect -958 4037 -946 4071
rect -912 4037 -900 4071
rect -958 4003 -900 4037
rect -958 3969 -946 4003
rect -912 3969 -900 4003
rect -958 3935 -900 3969
rect -958 3901 -946 3935
rect -912 3901 -900 3935
rect -958 3867 -900 3901
rect -958 3833 -946 3867
rect -912 3833 -900 3867
rect -958 3799 -900 3833
rect -958 3765 -946 3799
rect -912 3765 -900 3799
rect -958 3731 -900 3765
rect -958 3697 -946 3731
rect -912 3697 -900 3731
rect -958 3663 -900 3697
rect -958 3629 -946 3663
rect -912 3629 -900 3663
rect -958 3595 -900 3629
rect -958 3561 -946 3595
rect -912 3561 -900 3595
rect -958 3527 -900 3561
rect -958 3493 -946 3527
rect -912 3493 -900 3527
rect -958 3459 -900 3493
rect -958 3425 -946 3459
rect -912 3425 -900 3459
rect -958 3391 -900 3425
rect -958 3357 -946 3391
rect -912 3357 -900 3391
rect -958 3323 -900 3357
rect -958 3289 -946 3323
rect -912 3289 -900 3323
rect -958 3255 -900 3289
rect -958 3221 -946 3255
rect -912 3221 -900 3255
rect -958 3187 -900 3221
rect -958 3153 -946 3187
rect -912 3153 -900 3187
rect -958 3119 -900 3153
rect -958 3085 -946 3119
rect -912 3085 -900 3119
rect -958 3051 -900 3085
rect -958 3017 -946 3051
rect -912 3017 -900 3051
rect -958 2983 -900 3017
rect -958 2949 -946 2983
rect -912 2949 -900 2983
rect -958 2915 -900 2949
rect -958 2881 -946 2915
rect -912 2881 -900 2915
rect -958 2847 -900 2881
rect -958 2813 -946 2847
rect -912 2813 -900 2847
rect -958 2779 -900 2813
rect -958 2745 -946 2779
rect -912 2745 -900 2779
rect -958 2711 -900 2745
rect -958 2677 -946 2711
rect -912 2677 -900 2711
rect -958 2643 -900 2677
rect -958 2609 -946 2643
rect -912 2609 -900 2643
rect -958 2575 -900 2609
rect -958 2541 -946 2575
rect -912 2541 -900 2575
rect -958 2507 -900 2541
rect -958 2473 -946 2507
rect -912 2473 -900 2507
rect -958 2439 -900 2473
rect -958 2405 -946 2439
rect -912 2405 -900 2439
rect -958 2371 -900 2405
rect -958 2337 -946 2371
rect -912 2337 -900 2371
rect -958 2303 -900 2337
rect -958 2269 -946 2303
rect -912 2269 -900 2303
rect -958 2235 -900 2269
rect -958 2201 -946 2235
rect -912 2201 -900 2235
rect -958 2167 -900 2201
rect -958 2133 -946 2167
rect -912 2133 -900 2167
rect -958 2099 -900 2133
rect -958 2065 -946 2099
rect -912 2065 -900 2099
rect -958 2031 -900 2065
rect -958 1997 -946 2031
rect -912 1997 -900 2031
rect -958 1963 -900 1997
rect -958 1929 -946 1963
rect -912 1929 -900 1963
rect -958 1895 -900 1929
rect -958 1861 -946 1895
rect -912 1861 -900 1895
rect -958 1827 -900 1861
rect -958 1793 -946 1827
rect -912 1793 -900 1827
rect -958 1759 -900 1793
rect -958 1725 -946 1759
rect -912 1725 -900 1759
rect -958 1691 -900 1725
rect -958 1657 -946 1691
rect -912 1657 -900 1691
rect -958 1623 -900 1657
rect -958 1589 -946 1623
rect -912 1589 -900 1623
rect -958 1555 -900 1589
rect -958 1521 -946 1555
rect -912 1521 -900 1555
rect -958 1487 -900 1521
rect -958 1453 -946 1487
rect -912 1453 -900 1487
rect -958 1419 -900 1453
rect -958 1385 -946 1419
rect -912 1385 -900 1419
rect -958 1351 -900 1385
rect -958 1317 -946 1351
rect -912 1317 -900 1351
rect -958 1283 -900 1317
rect -958 1249 -946 1283
rect -912 1249 -900 1283
rect -958 1215 -900 1249
rect -958 1181 -946 1215
rect -912 1181 -900 1215
rect -958 1147 -900 1181
rect -958 1113 -946 1147
rect -912 1113 -900 1147
rect -958 1079 -900 1113
rect -958 1045 -946 1079
rect -912 1045 -900 1079
rect -958 1011 -900 1045
rect -958 977 -946 1011
rect -912 977 -900 1011
rect -958 943 -900 977
rect -958 909 -946 943
rect -912 909 -900 943
rect -958 875 -900 909
rect -958 841 -946 875
rect -912 841 -900 875
rect -958 807 -900 841
rect -958 773 -946 807
rect -912 773 -900 807
rect -958 739 -900 773
rect -958 705 -946 739
rect -912 705 -900 739
rect -958 671 -900 705
rect -958 637 -946 671
rect -912 637 -900 671
rect -958 603 -900 637
rect -958 569 -946 603
rect -912 569 -900 603
rect -958 535 -900 569
rect -958 501 -946 535
rect -912 501 -900 535
rect -958 467 -900 501
rect -958 433 -946 467
rect -912 433 -900 467
rect -958 399 -900 433
rect -958 365 -946 399
rect -912 365 -900 399
rect -958 331 -900 365
rect -958 297 -946 331
rect -912 297 -900 331
rect -958 263 -900 297
rect -958 229 -946 263
rect -912 229 -900 263
rect -958 195 -900 229
rect -958 161 -946 195
rect -912 161 -900 195
rect -958 127 -900 161
rect -958 93 -946 127
rect -912 93 -900 127
rect -958 59 -900 93
rect -958 25 -946 59
rect -912 25 -900 59
rect -958 0 -900 25
rect 1050 5975 1108 6000
rect 1050 5941 1062 5975
rect 1096 5941 1108 5975
rect 1050 5907 1108 5941
rect 1050 5873 1062 5907
rect 1096 5873 1108 5907
rect 1050 5839 1108 5873
rect 1050 5805 1062 5839
rect 1096 5805 1108 5839
rect 1050 5771 1108 5805
rect 1050 5737 1062 5771
rect 1096 5737 1108 5771
rect 1050 5703 1108 5737
rect 1050 5669 1062 5703
rect 1096 5669 1108 5703
rect 1050 5635 1108 5669
rect 1050 5601 1062 5635
rect 1096 5601 1108 5635
rect 1050 5567 1108 5601
rect 1050 5533 1062 5567
rect 1096 5533 1108 5567
rect 1050 5499 1108 5533
rect 1050 5465 1062 5499
rect 1096 5465 1108 5499
rect 1050 5431 1108 5465
rect 1050 5397 1062 5431
rect 1096 5397 1108 5431
rect 1050 5363 1108 5397
rect 1050 5329 1062 5363
rect 1096 5329 1108 5363
rect 1050 5295 1108 5329
rect 1050 5261 1062 5295
rect 1096 5261 1108 5295
rect 1050 5227 1108 5261
rect 1050 5193 1062 5227
rect 1096 5193 1108 5227
rect 1050 5159 1108 5193
rect 1050 5125 1062 5159
rect 1096 5125 1108 5159
rect 1050 5091 1108 5125
rect 1050 5057 1062 5091
rect 1096 5057 1108 5091
rect 1050 5023 1108 5057
rect 1050 4989 1062 5023
rect 1096 4989 1108 5023
rect 1050 4955 1108 4989
rect 1050 4921 1062 4955
rect 1096 4921 1108 4955
rect 1050 4887 1108 4921
rect 1050 4853 1062 4887
rect 1096 4853 1108 4887
rect 1050 4819 1108 4853
rect 1050 4785 1062 4819
rect 1096 4785 1108 4819
rect 1050 4751 1108 4785
rect 1050 4717 1062 4751
rect 1096 4717 1108 4751
rect 1050 4683 1108 4717
rect 1050 4649 1062 4683
rect 1096 4649 1108 4683
rect 1050 4615 1108 4649
rect 1050 4581 1062 4615
rect 1096 4581 1108 4615
rect 1050 4547 1108 4581
rect 1050 4513 1062 4547
rect 1096 4513 1108 4547
rect 1050 4479 1108 4513
rect 1050 4445 1062 4479
rect 1096 4445 1108 4479
rect 1050 4411 1108 4445
rect 1050 4377 1062 4411
rect 1096 4377 1108 4411
rect 1050 4343 1108 4377
rect 1050 4309 1062 4343
rect 1096 4309 1108 4343
rect 1050 4275 1108 4309
rect 1050 4241 1062 4275
rect 1096 4241 1108 4275
rect 1050 4207 1108 4241
rect 1050 4173 1062 4207
rect 1096 4173 1108 4207
rect 1050 4139 1108 4173
rect 1050 4105 1062 4139
rect 1096 4105 1108 4139
rect 1050 4071 1108 4105
rect 1050 4037 1062 4071
rect 1096 4037 1108 4071
rect 1050 4003 1108 4037
rect 1050 3969 1062 4003
rect 1096 3969 1108 4003
rect 1050 3935 1108 3969
rect 1050 3901 1062 3935
rect 1096 3901 1108 3935
rect 1050 3867 1108 3901
rect 1050 3833 1062 3867
rect 1096 3833 1108 3867
rect 1050 3799 1108 3833
rect 1050 3765 1062 3799
rect 1096 3765 1108 3799
rect 1050 3731 1108 3765
rect 1050 3697 1062 3731
rect 1096 3697 1108 3731
rect 1050 3663 1108 3697
rect 1050 3629 1062 3663
rect 1096 3629 1108 3663
rect 1050 3595 1108 3629
rect 1050 3561 1062 3595
rect 1096 3561 1108 3595
rect 1050 3527 1108 3561
rect 1050 3493 1062 3527
rect 1096 3493 1108 3527
rect 1050 3459 1108 3493
rect 1050 3425 1062 3459
rect 1096 3425 1108 3459
rect 1050 3391 1108 3425
rect 1050 3357 1062 3391
rect 1096 3357 1108 3391
rect 1050 3323 1108 3357
rect 1050 3289 1062 3323
rect 1096 3289 1108 3323
rect 1050 3255 1108 3289
rect 1050 3221 1062 3255
rect 1096 3221 1108 3255
rect 1050 3187 1108 3221
rect 1050 3153 1062 3187
rect 1096 3153 1108 3187
rect 1050 3119 1108 3153
rect 1050 3085 1062 3119
rect 1096 3085 1108 3119
rect 1050 3051 1108 3085
rect 1050 3017 1062 3051
rect 1096 3017 1108 3051
rect 1050 2983 1108 3017
rect 1050 2949 1062 2983
rect 1096 2949 1108 2983
rect 1050 2915 1108 2949
rect 1050 2881 1062 2915
rect 1096 2881 1108 2915
rect 1050 2847 1108 2881
rect 1050 2813 1062 2847
rect 1096 2813 1108 2847
rect 1050 2779 1108 2813
rect 1050 2745 1062 2779
rect 1096 2745 1108 2779
rect 1050 2711 1108 2745
rect 1050 2677 1062 2711
rect 1096 2677 1108 2711
rect 1050 2643 1108 2677
rect 1050 2609 1062 2643
rect 1096 2609 1108 2643
rect 1050 2575 1108 2609
rect 1050 2541 1062 2575
rect 1096 2541 1108 2575
rect 1050 2507 1108 2541
rect 1050 2473 1062 2507
rect 1096 2473 1108 2507
rect 1050 2439 1108 2473
rect 1050 2405 1062 2439
rect 1096 2405 1108 2439
rect 1050 2371 1108 2405
rect 1050 2337 1062 2371
rect 1096 2337 1108 2371
rect 1050 2303 1108 2337
rect 1050 2269 1062 2303
rect 1096 2269 1108 2303
rect 1050 2235 1108 2269
rect 1050 2201 1062 2235
rect 1096 2201 1108 2235
rect 1050 2167 1108 2201
rect 1050 2133 1062 2167
rect 1096 2133 1108 2167
rect 1050 2099 1108 2133
rect 1050 2065 1062 2099
rect 1096 2065 1108 2099
rect 1050 2031 1108 2065
rect 1050 1997 1062 2031
rect 1096 1997 1108 2031
rect 1050 1963 1108 1997
rect 1050 1929 1062 1963
rect 1096 1929 1108 1963
rect 1050 1895 1108 1929
rect 1050 1861 1062 1895
rect 1096 1861 1108 1895
rect 1050 1827 1108 1861
rect 1050 1793 1062 1827
rect 1096 1793 1108 1827
rect 1050 1759 1108 1793
rect 1050 1725 1062 1759
rect 1096 1725 1108 1759
rect 1050 1691 1108 1725
rect 1050 1657 1062 1691
rect 1096 1657 1108 1691
rect 1050 1623 1108 1657
rect 1050 1589 1062 1623
rect 1096 1589 1108 1623
rect 1050 1555 1108 1589
rect 1050 1521 1062 1555
rect 1096 1521 1108 1555
rect 1050 1487 1108 1521
rect 1050 1453 1062 1487
rect 1096 1453 1108 1487
rect 1050 1419 1108 1453
rect 1050 1385 1062 1419
rect 1096 1385 1108 1419
rect 1050 1351 1108 1385
rect 1050 1317 1062 1351
rect 1096 1317 1108 1351
rect 1050 1283 1108 1317
rect 1050 1249 1062 1283
rect 1096 1249 1108 1283
rect 1050 1215 1108 1249
rect 1050 1181 1062 1215
rect 1096 1181 1108 1215
rect 1050 1147 1108 1181
rect 1050 1113 1062 1147
rect 1096 1113 1108 1147
rect 1050 1079 1108 1113
rect 1050 1045 1062 1079
rect 1096 1045 1108 1079
rect 1050 1011 1108 1045
rect 1050 977 1062 1011
rect 1096 977 1108 1011
rect 1050 943 1108 977
rect 1050 909 1062 943
rect 1096 909 1108 943
rect 1050 875 1108 909
rect 1050 841 1062 875
rect 1096 841 1108 875
rect 1050 807 1108 841
rect 1050 773 1062 807
rect 1096 773 1108 807
rect 1050 739 1108 773
rect 1050 705 1062 739
rect 1096 705 1108 739
rect 1050 671 1108 705
rect 1050 637 1062 671
rect 1096 637 1108 671
rect 1050 603 1108 637
rect 1050 569 1062 603
rect 1096 569 1108 603
rect 1050 535 1108 569
rect 1050 501 1062 535
rect 1096 501 1108 535
rect 1050 467 1108 501
rect 1050 433 1062 467
rect 1096 433 1108 467
rect 1050 399 1108 433
rect 1050 365 1062 399
rect 1096 365 1108 399
rect 1050 331 1108 365
rect 1050 297 1062 331
rect 1096 297 1108 331
rect 1050 263 1108 297
rect 1050 229 1062 263
rect 1096 229 1108 263
rect 1050 195 1108 229
rect 1050 161 1062 195
rect 1096 161 1108 195
rect 1050 127 1108 161
rect 1050 93 1062 127
rect 1096 93 1108 127
rect 1050 59 1108 93
rect 1050 25 1062 59
rect 1096 25 1108 59
rect 1050 0 1108 25
<< mvndiffc >>
rect -946 5941 -912 5975
rect -946 5873 -912 5907
rect -946 5805 -912 5839
rect -946 5737 -912 5771
rect -946 5669 -912 5703
rect -946 5601 -912 5635
rect -946 5533 -912 5567
rect -946 5465 -912 5499
rect -946 5397 -912 5431
rect -946 5329 -912 5363
rect -946 5261 -912 5295
rect -946 5193 -912 5227
rect -946 5125 -912 5159
rect -946 5057 -912 5091
rect -946 4989 -912 5023
rect -946 4921 -912 4955
rect -946 4853 -912 4887
rect -946 4785 -912 4819
rect -946 4717 -912 4751
rect -946 4649 -912 4683
rect -946 4581 -912 4615
rect -946 4513 -912 4547
rect -946 4445 -912 4479
rect -946 4377 -912 4411
rect -946 4309 -912 4343
rect -946 4241 -912 4275
rect -946 4173 -912 4207
rect -946 4105 -912 4139
rect -946 4037 -912 4071
rect -946 3969 -912 4003
rect -946 3901 -912 3935
rect -946 3833 -912 3867
rect -946 3765 -912 3799
rect -946 3697 -912 3731
rect -946 3629 -912 3663
rect -946 3561 -912 3595
rect -946 3493 -912 3527
rect -946 3425 -912 3459
rect -946 3357 -912 3391
rect -946 3289 -912 3323
rect -946 3221 -912 3255
rect -946 3153 -912 3187
rect -946 3085 -912 3119
rect -946 3017 -912 3051
rect -946 2949 -912 2983
rect -946 2881 -912 2915
rect -946 2813 -912 2847
rect -946 2745 -912 2779
rect -946 2677 -912 2711
rect -946 2609 -912 2643
rect -946 2541 -912 2575
rect -946 2473 -912 2507
rect -946 2405 -912 2439
rect -946 2337 -912 2371
rect -946 2269 -912 2303
rect -946 2201 -912 2235
rect -946 2133 -912 2167
rect -946 2065 -912 2099
rect -946 1997 -912 2031
rect -946 1929 -912 1963
rect -946 1861 -912 1895
rect -946 1793 -912 1827
rect -946 1725 -912 1759
rect -946 1657 -912 1691
rect -946 1589 -912 1623
rect -946 1521 -912 1555
rect -946 1453 -912 1487
rect -946 1385 -912 1419
rect -946 1317 -912 1351
rect -946 1249 -912 1283
rect -946 1181 -912 1215
rect -946 1113 -912 1147
rect -946 1045 -912 1079
rect -946 977 -912 1011
rect -946 909 -912 943
rect -946 841 -912 875
rect -946 773 -912 807
rect -946 705 -912 739
rect -946 637 -912 671
rect -946 569 -912 603
rect -946 501 -912 535
rect -946 433 -912 467
rect -946 365 -912 399
rect -946 297 -912 331
rect -946 229 -912 263
rect -946 161 -912 195
rect -946 93 -912 127
rect -946 25 -912 59
rect 1062 5941 1096 5975
rect 1062 5873 1096 5907
rect 1062 5805 1096 5839
rect 1062 5737 1096 5771
rect 1062 5669 1096 5703
rect 1062 5601 1096 5635
rect 1062 5533 1096 5567
rect 1062 5465 1096 5499
rect 1062 5397 1096 5431
rect 1062 5329 1096 5363
rect 1062 5261 1096 5295
rect 1062 5193 1096 5227
rect 1062 5125 1096 5159
rect 1062 5057 1096 5091
rect 1062 4989 1096 5023
rect 1062 4921 1096 4955
rect 1062 4853 1096 4887
rect 1062 4785 1096 4819
rect 1062 4717 1096 4751
rect 1062 4649 1096 4683
rect 1062 4581 1096 4615
rect 1062 4513 1096 4547
rect 1062 4445 1096 4479
rect 1062 4377 1096 4411
rect 1062 4309 1096 4343
rect 1062 4241 1096 4275
rect 1062 4173 1096 4207
rect 1062 4105 1096 4139
rect 1062 4037 1096 4071
rect 1062 3969 1096 4003
rect 1062 3901 1096 3935
rect 1062 3833 1096 3867
rect 1062 3765 1096 3799
rect 1062 3697 1096 3731
rect 1062 3629 1096 3663
rect 1062 3561 1096 3595
rect 1062 3493 1096 3527
rect 1062 3425 1096 3459
rect 1062 3357 1096 3391
rect 1062 3289 1096 3323
rect 1062 3221 1096 3255
rect 1062 3153 1096 3187
rect 1062 3085 1096 3119
rect 1062 3017 1096 3051
rect 1062 2949 1096 2983
rect 1062 2881 1096 2915
rect 1062 2813 1096 2847
rect 1062 2745 1096 2779
rect 1062 2677 1096 2711
rect 1062 2609 1096 2643
rect 1062 2541 1096 2575
rect 1062 2473 1096 2507
rect 1062 2405 1096 2439
rect 1062 2337 1096 2371
rect 1062 2269 1096 2303
rect 1062 2201 1096 2235
rect 1062 2133 1096 2167
rect 1062 2065 1096 2099
rect 1062 1997 1096 2031
rect 1062 1929 1096 1963
rect 1062 1861 1096 1895
rect 1062 1793 1096 1827
rect 1062 1725 1096 1759
rect 1062 1657 1096 1691
rect 1062 1589 1096 1623
rect 1062 1521 1096 1555
rect 1062 1453 1096 1487
rect 1062 1385 1096 1419
rect 1062 1317 1096 1351
rect 1062 1249 1096 1283
rect 1062 1181 1096 1215
rect 1062 1113 1096 1147
rect 1062 1045 1096 1079
rect 1062 977 1096 1011
rect 1062 909 1096 943
rect 1062 841 1096 875
rect 1062 773 1096 807
rect 1062 705 1096 739
rect 1062 637 1096 671
rect 1062 569 1096 603
rect 1062 501 1096 535
rect 1062 433 1096 467
rect 1062 365 1096 399
rect 1062 297 1096 331
rect 1062 229 1096 263
rect 1062 161 1096 195
rect 1062 93 1096 127
rect 1062 25 1096 59
<< mvpsubdiff >>
rect -1140 7158 1290 7182
rect -1140 7124 -866 7158
rect -832 7124 -798 7158
rect -764 7124 -730 7158
rect -696 7124 -662 7158
rect -628 7124 -594 7158
rect -560 7124 -526 7158
rect -492 7124 -458 7158
rect -424 7124 -390 7158
rect -356 7124 -322 7158
rect -288 7124 -254 7158
rect -220 7124 -186 7158
rect -152 7124 -118 7158
rect -84 7124 -50 7158
rect -16 7124 18 7158
rect 52 7124 86 7158
rect 120 7124 154 7158
rect 188 7124 222 7158
rect 256 7124 290 7158
rect 324 7124 358 7158
rect 392 7124 426 7158
rect 460 7124 494 7158
rect 528 7124 562 7158
rect 596 7124 630 7158
rect 664 7124 698 7158
rect 732 7124 766 7158
rect 800 7124 834 7158
rect 868 7124 902 7158
rect 936 7124 970 7158
rect 1004 7124 1290 7158
rect -1140 7100 1290 7124
rect -1140 7029 -1058 7100
rect -1140 6995 -1116 7029
rect -1082 6995 -1058 7029
rect 1208 7029 1290 7100
rect -1140 6961 -1058 6995
rect -1140 6927 -1116 6961
rect -1082 6927 -1058 6961
rect -1140 6893 -1058 6927
rect -1140 6859 -1116 6893
rect -1082 6859 -1058 6893
rect -1140 6825 -1058 6859
rect -1140 6791 -1116 6825
rect -1082 6791 -1058 6825
rect -1140 6757 -1058 6791
rect -1140 6723 -1116 6757
rect -1082 6723 -1058 6757
rect -1140 6689 -1058 6723
rect -1140 6655 -1116 6689
rect -1082 6655 -1058 6689
rect -1140 6621 -1058 6655
rect -1140 6587 -1116 6621
rect -1082 6587 -1058 6621
rect -1140 6553 -1058 6587
rect -1140 6519 -1116 6553
rect -1082 6519 -1058 6553
rect -1140 6485 -1058 6519
rect -1140 6451 -1116 6485
rect -1082 6451 -1058 6485
rect -1140 6417 -1058 6451
rect -1140 6383 -1116 6417
rect -1082 6383 -1058 6417
rect -1140 6349 -1058 6383
rect -1140 6315 -1116 6349
rect -1082 6315 -1058 6349
rect -1140 6281 -1058 6315
rect -1140 6247 -1116 6281
rect -1082 6247 -1058 6281
rect -1140 6213 -1058 6247
rect -1140 6179 -1116 6213
rect -1082 6179 -1058 6213
rect -1140 6145 -1058 6179
rect -1140 6111 -1116 6145
rect -1082 6111 -1058 6145
rect -1140 6077 -1058 6111
rect -1140 6043 -1116 6077
rect -1082 6043 -1058 6077
rect -1140 6009 -1058 6043
rect -1140 5975 -1116 6009
rect -1082 5975 -1058 6009
rect 1208 6995 1232 7029
rect 1266 6995 1290 7029
rect 1208 6961 1290 6995
rect 1208 6927 1232 6961
rect 1266 6927 1290 6961
rect 1208 6893 1290 6927
rect 1208 6859 1232 6893
rect 1266 6859 1290 6893
rect 1208 6825 1290 6859
rect 1208 6791 1232 6825
rect 1266 6791 1290 6825
rect 1208 6757 1290 6791
rect 1208 6723 1232 6757
rect 1266 6723 1290 6757
rect 1208 6689 1290 6723
rect 1208 6655 1232 6689
rect 1266 6655 1290 6689
rect 1208 6621 1290 6655
rect 1208 6587 1232 6621
rect 1266 6587 1290 6621
rect 1208 6553 1290 6587
rect 1208 6519 1232 6553
rect 1266 6519 1290 6553
rect 1208 6485 1290 6519
rect 1208 6451 1232 6485
rect 1266 6451 1290 6485
rect 1208 6417 1290 6451
rect 1208 6383 1232 6417
rect 1266 6383 1290 6417
rect 1208 6349 1290 6383
rect 1208 6315 1232 6349
rect 1266 6315 1290 6349
rect 1208 6281 1290 6315
rect 1208 6247 1232 6281
rect 1266 6247 1290 6281
rect 1208 6213 1290 6247
rect 1208 6179 1232 6213
rect 1266 6179 1290 6213
rect 1208 6145 1290 6179
rect 1208 6111 1232 6145
rect 1266 6111 1290 6145
rect 1208 6077 1290 6111
rect 1208 6043 1232 6077
rect 1266 6043 1290 6077
rect 1208 6009 1290 6043
rect -1140 5941 -1058 5975
rect -1140 5907 -1116 5941
rect -1082 5907 -1058 5941
rect -1140 5873 -1058 5907
rect -1140 5839 -1116 5873
rect -1082 5839 -1058 5873
rect -1140 5805 -1058 5839
rect -1140 5771 -1116 5805
rect -1082 5771 -1058 5805
rect -1140 5737 -1058 5771
rect -1140 5703 -1116 5737
rect -1082 5703 -1058 5737
rect -1140 5669 -1058 5703
rect -1140 5635 -1116 5669
rect -1082 5635 -1058 5669
rect -1140 5601 -1058 5635
rect -1140 5567 -1116 5601
rect -1082 5567 -1058 5601
rect -1140 5533 -1058 5567
rect -1140 5499 -1116 5533
rect -1082 5499 -1058 5533
rect -1140 5465 -1058 5499
rect -1140 5431 -1116 5465
rect -1082 5431 -1058 5465
rect -1140 5397 -1058 5431
rect -1140 5363 -1116 5397
rect -1082 5363 -1058 5397
rect -1140 5329 -1058 5363
rect -1140 5295 -1116 5329
rect -1082 5295 -1058 5329
rect -1140 5261 -1058 5295
rect -1140 5227 -1116 5261
rect -1082 5227 -1058 5261
rect -1140 5193 -1058 5227
rect -1140 5159 -1116 5193
rect -1082 5159 -1058 5193
rect -1140 5125 -1058 5159
rect -1140 5091 -1116 5125
rect -1082 5091 -1058 5125
rect -1140 5057 -1058 5091
rect -1140 5023 -1116 5057
rect -1082 5023 -1058 5057
rect -1140 4989 -1058 5023
rect -1140 4955 -1116 4989
rect -1082 4955 -1058 4989
rect -1140 4921 -1058 4955
rect -1140 4887 -1116 4921
rect -1082 4887 -1058 4921
rect -1140 4853 -1058 4887
rect -1140 4819 -1116 4853
rect -1082 4819 -1058 4853
rect -1140 4785 -1058 4819
rect -1140 4751 -1116 4785
rect -1082 4751 -1058 4785
rect -1140 4717 -1058 4751
rect -1140 4683 -1116 4717
rect -1082 4683 -1058 4717
rect -1140 4649 -1058 4683
rect -1140 4615 -1116 4649
rect -1082 4615 -1058 4649
rect -1140 4581 -1058 4615
rect -1140 4547 -1116 4581
rect -1082 4547 -1058 4581
rect -1140 4513 -1058 4547
rect -1140 4479 -1116 4513
rect -1082 4479 -1058 4513
rect -1140 4445 -1058 4479
rect -1140 4411 -1116 4445
rect -1082 4411 -1058 4445
rect -1140 4377 -1058 4411
rect -1140 4343 -1116 4377
rect -1082 4343 -1058 4377
rect -1140 4309 -1058 4343
rect -1140 4275 -1116 4309
rect -1082 4275 -1058 4309
rect -1140 4241 -1058 4275
rect -1140 4207 -1116 4241
rect -1082 4207 -1058 4241
rect -1140 4173 -1058 4207
rect -1140 4139 -1116 4173
rect -1082 4139 -1058 4173
rect -1140 4105 -1058 4139
rect -1140 4071 -1116 4105
rect -1082 4071 -1058 4105
rect -1140 4037 -1058 4071
rect -1140 4003 -1116 4037
rect -1082 4003 -1058 4037
rect -1140 3969 -1058 4003
rect -1140 3935 -1116 3969
rect -1082 3935 -1058 3969
rect -1140 3901 -1058 3935
rect -1140 3867 -1116 3901
rect -1082 3867 -1058 3901
rect -1140 3833 -1058 3867
rect -1140 3799 -1116 3833
rect -1082 3799 -1058 3833
rect -1140 3765 -1058 3799
rect -1140 3731 -1116 3765
rect -1082 3731 -1058 3765
rect -1140 3697 -1058 3731
rect -1140 3663 -1116 3697
rect -1082 3663 -1058 3697
rect -1140 3629 -1058 3663
rect -1140 3595 -1116 3629
rect -1082 3595 -1058 3629
rect -1140 3561 -1058 3595
rect -1140 3527 -1116 3561
rect -1082 3527 -1058 3561
rect -1140 3493 -1058 3527
rect -1140 3459 -1116 3493
rect -1082 3459 -1058 3493
rect -1140 3425 -1058 3459
rect -1140 3391 -1116 3425
rect -1082 3391 -1058 3425
rect -1140 3357 -1058 3391
rect -1140 3323 -1116 3357
rect -1082 3323 -1058 3357
rect -1140 3289 -1058 3323
rect -1140 3255 -1116 3289
rect -1082 3255 -1058 3289
rect -1140 3221 -1058 3255
rect -1140 3187 -1116 3221
rect -1082 3187 -1058 3221
rect -1140 3153 -1058 3187
rect -1140 3119 -1116 3153
rect -1082 3119 -1058 3153
rect -1140 3085 -1058 3119
rect -1140 3051 -1116 3085
rect -1082 3051 -1058 3085
rect -1140 3017 -1058 3051
rect -1140 2983 -1116 3017
rect -1082 2983 -1058 3017
rect -1140 2949 -1058 2983
rect -1140 2915 -1116 2949
rect -1082 2915 -1058 2949
rect -1140 2881 -1058 2915
rect -1140 2847 -1116 2881
rect -1082 2847 -1058 2881
rect -1140 2813 -1058 2847
rect -1140 2779 -1116 2813
rect -1082 2779 -1058 2813
rect -1140 2745 -1058 2779
rect -1140 2711 -1116 2745
rect -1082 2711 -1058 2745
rect -1140 2677 -1058 2711
rect -1140 2643 -1116 2677
rect -1082 2643 -1058 2677
rect -1140 2609 -1058 2643
rect -1140 2575 -1116 2609
rect -1082 2575 -1058 2609
rect -1140 2541 -1058 2575
rect -1140 2507 -1116 2541
rect -1082 2507 -1058 2541
rect -1140 2473 -1058 2507
rect -1140 2439 -1116 2473
rect -1082 2439 -1058 2473
rect -1140 2405 -1058 2439
rect -1140 2371 -1116 2405
rect -1082 2371 -1058 2405
rect -1140 2337 -1058 2371
rect -1140 2303 -1116 2337
rect -1082 2303 -1058 2337
rect -1140 2269 -1058 2303
rect -1140 2235 -1116 2269
rect -1082 2235 -1058 2269
rect -1140 2201 -1058 2235
rect -1140 2167 -1116 2201
rect -1082 2167 -1058 2201
rect -1140 2133 -1058 2167
rect -1140 2099 -1116 2133
rect -1082 2099 -1058 2133
rect -1140 2065 -1058 2099
rect -1140 2031 -1116 2065
rect -1082 2031 -1058 2065
rect -1140 1997 -1058 2031
rect -1140 1963 -1116 1997
rect -1082 1963 -1058 1997
rect -1140 1929 -1058 1963
rect -1140 1895 -1116 1929
rect -1082 1895 -1058 1929
rect -1140 1861 -1058 1895
rect -1140 1827 -1116 1861
rect -1082 1827 -1058 1861
rect -1140 1793 -1058 1827
rect -1140 1759 -1116 1793
rect -1082 1759 -1058 1793
rect -1140 1725 -1058 1759
rect -1140 1691 -1116 1725
rect -1082 1691 -1058 1725
rect -1140 1657 -1058 1691
rect -1140 1623 -1116 1657
rect -1082 1623 -1058 1657
rect -1140 1589 -1058 1623
rect -1140 1555 -1116 1589
rect -1082 1555 -1058 1589
rect -1140 1521 -1058 1555
rect -1140 1487 -1116 1521
rect -1082 1487 -1058 1521
rect -1140 1453 -1058 1487
rect -1140 1419 -1116 1453
rect -1082 1419 -1058 1453
rect -1140 1385 -1058 1419
rect -1140 1351 -1116 1385
rect -1082 1351 -1058 1385
rect -1140 1317 -1058 1351
rect -1140 1283 -1116 1317
rect -1082 1283 -1058 1317
rect -1140 1249 -1058 1283
rect -1140 1215 -1116 1249
rect -1082 1215 -1058 1249
rect -1140 1181 -1058 1215
rect -1140 1147 -1116 1181
rect -1082 1147 -1058 1181
rect -1140 1113 -1058 1147
rect -1140 1079 -1116 1113
rect -1082 1079 -1058 1113
rect -1140 1045 -1058 1079
rect -1140 1011 -1116 1045
rect -1082 1011 -1058 1045
rect -1140 977 -1058 1011
rect -1140 943 -1116 977
rect -1082 943 -1058 977
rect -1140 909 -1058 943
rect -1140 875 -1116 909
rect -1082 875 -1058 909
rect -1140 841 -1058 875
rect -1140 807 -1116 841
rect -1082 807 -1058 841
rect -1140 773 -1058 807
rect -1140 739 -1116 773
rect -1082 739 -1058 773
rect -1140 705 -1058 739
rect -1140 671 -1116 705
rect -1082 671 -1058 705
rect -1140 637 -1058 671
rect -1140 603 -1116 637
rect -1082 603 -1058 637
rect -1140 569 -1058 603
rect -1140 535 -1116 569
rect -1082 535 -1058 569
rect -1140 501 -1058 535
rect -1140 467 -1116 501
rect -1082 467 -1058 501
rect -1140 433 -1058 467
rect -1140 399 -1116 433
rect -1082 399 -1058 433
rect -1140 365 -1058 399
rect -1140 331 -1116 365
rect -1082 331 -1058 365
rect -1140 297 -1058 331
rect -1140 263 -1116 297
rect -1082 263 -1058 297
rect -1140 229 -1058 263
rect -1140 195 -1116 229
rect -1082 195 -1058 229
rect -1140 161 -1058 195
rect -1140 127 -1116 161
rect -1082 127 -1058 161
rect -1140 93 -1058 127
rect -1140 59 -1116 93
rect -1082 59 -1058 93
rect -1140 25 -1058 59
rect -1140 -9 -1116 25
rect -1082 -9 -1058 25
rect 1208 5975 1232 6009
rect 1266 5975 1290 6009
rect 1208 5941 1290 5975
rect 1208 5907 1232 5941
rect 1266 5907 1290 5941
rect 1208 5873 1290 5907
rect 1208 5839 1232 5873
rect 1266 5839 1290 5873
rect 1208 5805 1290 5839
rect 1208 5771 1232 5805
rect 1266 5771 1290 5805
rect 1208 5737 1290 5771
rect 1208 5703 1232 5737
rect 1266 5703 1290 5737
rect 1208 5669 1290 5703
rect 1208 5635 1232 5669
rect 1266 5635 1290 5669
rect 1208 5601 1290 5635
rect 1208 5567 1232 5601
rect 1266 5567 1290 5601
rect 1208 5533 1290 5567
rect 1208 5499 1232 5533
rect 1266 5499 1290 5533
rect 1208 5465 1290 5499
rect 1208 5431 1232 5465
rect 1266 5431 1290 5465
rect 1208 5397 1290 5431
rect 1208 5363 1232 5397
rect 1266 5363 1290 5397
rect 1208 5329 1290 5363
rect 1208 5295 1232 5329
rect 1266 5295 1290 5329
rect 1208 5261 1290 5295
rect 1208 5227 1232 5261
rect 1266 5227 1290 5261
rect 1208 5193 1290 5227
rect 1208 5159 1232 5193
rect 1266 5159 1290 5193
rect 1208 5125 1290 5159
rect 1208 5091 1232 5125
rect 1266 5091 1290 5125
rect 1208 5057 1290 5091
rect 1208 5023 1232 5057
rect 1266 5023 1290 5057
rect 1208 4989 1290 5023
rect 1208 4955 1232 4989
rect 1266 4955 1290 4989
rect 1208 4921 1290 4955
rect 1208 4887 1232 4921
rect 1266 4887 1290 4921
rect 1208 4853 1290 4887
rect 1208 4819 1232 4853
rect 1266 4819 1290 4853
rect 1208 4785 1290 4819
rect 1208 4751 1232 4785
rect 1266 4751 1290 4785
rect 1208 4717 1290 4751
rect 1208 4683 1232 4717
rect 1266 4683 1290 4717
rect 1208 4649 1290 4683
rect 1208 4615 1232 4649
rect 1266 4615 1290 4649
rect 1208 4581 1290 4615
rect 1208 4547 1232 4581
rect 1266 4547 1290 4581
rect 1208 4513 1290 4547
rect 1208 4479 1232 4513
rect 1266 4479 1290 4513
rect 1208 4445 1290 4479
rect 1208 4411 1232 4445
rect 1266 4411 1290 4445
rect 1208 4377 1290 4411
rect 1208 4343 1232 4377
rect 1266 4343 1290 4377
rect 1208 4309 1290 4343
rect 1208 4275 1232 4309
rect 1266 4275 1290 4309
rect 1208 4241 1290 4275
rect 1208 4207 1232 4241
rect 1266 4207 1290 4241
rect 1208 4173 1290 4207
rect 1208 4139 1232 4173
rect 1266 4139 1290 4173
rect 1208 4105 1290 4139
rect 1208 4071 1232 4105
rect 1266 4071 1290 4105
rect 1208 4037 1290 4071
rect 1208 4003 1232 4037
rect 1266 4003 1290 4037
rect 1208 3969 1290 4003
rect 1208 3935 1232 3969
rect 1266 3935 1290 3969
rect 1208 3901 1290 3935
rect 1208 3867 1232 3901
rect 1266 3867 1290 3901
rect 1208 3833 1290 3867
rect 1208 3799 1232 3833
rect 1266 3799 1290 3833
rect 1208 3765 1290 3799
rect 1208 3731 1232 3765
rect 1266 3731 1290 3765
rect 1208 3697 1290 3731
rect 1208 3663 1232 3697
rect 1266 3663 1290 3697
rect 1208 3629 1290 3663
rect 1208 3595 1232 3629
rect 1266 3595 1290 3629
rect 1208 3561 1290 3595
rect 1208 3527 1232 3561
rect 1266 3527 1290 3561
rect 1208 3493 1290 3527
rect 1208 3459 1232 3493
rect 1266 3459 1290 3493
rect 1208 3425 1290 3459
rect 1208 3391 1232 3425
rect 1266 3391 1290 3425
rect 1208 3357 1290 3391
rect 1208 3323 1232 3357
rect 1266 3323 1290 3357
rect 1208 3289 1290 3323
rect 1208 3255 1232 3289
rect 1266 3255 1290 3289
rect 1208 3221 1290 3255
rect 1208 3187 1232 3221
rect 1266 3187 1290 3221
rect 1208 3153 1290 3187
rect 1208 3119 1232 3153
rect 1266 3119 1290 3153
rect 1208 3085 1290 3119
rect 1208 3051 1232 3085
rect 1266 3051 1290 3085
rect 1208 3017 1290 3051
rect 1208 2983 1232 3017
rect 1266 2983 1290 3017
rect 1208 2949 1290 2983
rect 1208 2915 1232 2949
rect 1266 2915 1290 2949
rect 1208 2881 1290 2915
rect 1208 2847 1232 2881
rect 1266 2847 1290 2881
rect 1208 2813 1290 2847
rect 1208 2779 1232 2813
rect 1266 2779 1290 2813
rect 1208 2745 1290 2779
rect 1208 2711 1232 2745
rect 1266 2711 1290 2745
rect 1208 2677 1290 2711
rect 1208 2643 1232 2677
rect 1266 2643 1290 2677
rect 1208 2609 1290 2643
rect 1208 2575 1232 2609
rect 1266 2575 1290 2609
rect 1208 2541 1290 2575
rect 1208 2507 1232 2541
rect 1266 2507 1290 2541
rect 1208 2473 1290 2507
rect 1208 2439 1232 2473
rect 1266 2439 1290 2473
rect 1208 2405 1290 2439
rect 1208 2371 1232 2405
rect 1266 2371 1290 2405
rect 1208 2337 1290 2371
rect 1208 2303 1232 2337
rect 1266 2303 1290 2337
rect 1208 2269 1290 2303
rect 1208 2235 1232 2269
rect 1266 2235 1290 2269
rect 1208 2201 1290 2235
rect 1208 2167 1232 2201
rect 1266 2167 1290 2201
rect 1208 2133 1290 2167
rect 1208 2099 1232 2133
rect 1266 2099 1290 2133
rect 1208 2065 1290 2099
rect 1208 2031 1232 2065
rect 1266 2031 1290 2065
rect 1208 1997 1290 2031
rect 1208 1963 1232 1997
rect 1266 1963 1290 1997
rect 1208 1929 1290 1963
rect 1208 1895 1232 1929
rect 1266 1895 1290 1929
rect 1208 1861 1290 1895
rect 1208 1827 1232 1861
rect 1266 1827 1290 1861
rect 1208 1793 1290 1827
rect 1208 1759 1232 1793
rect 1266 1759 1290 1793
rect 1208 1725 1290 1759
rect 1208 1691 1232 1725
rect 1266 1691 1290 1725
rect 1208 1657 1290 1691
rect 1208 1623 1232 1657
rect 1266 1623 1290 1657
rect 1208 1589 1290 1623
rect 1208 1555 1232 1589
rect 1266 1555 1290 1589
rect 1208 1521 1290 1555
rect 1208 1487 1232 1521
rect 1266 1487 1290 1521
rect 1208 1453 1290 1487
rect 1208 1419 1232 1453
rect 1266 1419 1290 1453
rect 1208 1385 1290 1419
rect 1208 1351 1232 1385
rect 1266 1351 1290 1385
rect 1208 1317 1290 1351
rect 1208 1283 1232 1317
rect 1266 1283 1290 1317
rect 1208 1249 1290 1283
rect 1208 1215 1232 1249
rect 1266 1215 1290 1249
rect 1208 1181 1290 1215
rect 1208 1147 1232 1181
rect 1266 1147 1290 1181
rect 1208 1113 1290 1147
rect 1208 1079 1232 1113
rect 1266 1079 1290 1113
rect 1208 1045 1290 1079
rect 1208 1011 1232 1045
rect 1266 1011 1290 1045
rect 1208 977 1290 1011
rect 1208 943 1232 977
rect 1266 943 1290 977
rect 1208 909 1290 943
rect 1208 875 1232 909
rect 1266 875 1290 909
rect 1208 841 1290 875
rect 1208 807 1232 841
rect 1266 807 1290 841
rect 1208 773 1290 807
rect 1208 739 1232 773
rect 1266 739 1290 773
rect 1208 705 1290 739
rect 1208 671 1232 705
rect 1266 671 1290 705
rect 1208 637 1290 671
rect 1208 603 1232 637
rect 1266 603 1290 637
rect 1208 569 1290 603
rect 1208 535 1232 569
rect 1266 535 1290 569
rect 1208 501 1290 535
rect 1208 467 1232 501
rect 1266 467 1290 501
rect 1208 433 1290 467
rect 1208 399 1232 433
rect 1266 399 1290 433
rect 1208 365 1290 399
rect 1208 331 1232 365
rect 1266 331 1290 365
rect 1208 297 1290 331
rect 1208 263 1232 297
rect 1266 263 1290 297
rect 1208 229 1290 263
rect 1208 195 1232 229
rect 1266 195 1290 229
rect 1208 161 1290 195
rect 1208 127 1232 161
rect 1266 127 1290 161
rect 1208 93 1290 127
rect 1208 59 1232 93
rect 1266 59 1290 93
rect 1208 25 1290 59
rect -1140 -43 -1058 -9
rect -1140 -77 -1116 -43
rect -1082 -77 -1058 -43
rect -1140 -111 -1058 -77
rect -1140 -145 -1116 -111
rect -1082 -145 -1058 -111
rect -1140 -179 -1058 -145
rect -1140 -213 -1116 -179
rect -1082 -213 -1058 -179
rect -1140 -247 -1058 -213
rect -1140 -281 -1116 -247
rect -1082 -281 -1058 -247
rect -1140 -315 -1058 -281
rect -1140 -349 -1116 -315
rect -1082 -349 -1058 -315
rect -1140 -383 -1058 -349
rect -1140 -417 -1116 -383
rect -1082 -417 -1058 -383
rect -1140 -451 -1058 -417
rect -1140 -485 -1116 -451
rect -1082 -485 -1058 -451
rect -1140 -519 -1058 -485
rect -1140 -553 -1116 -519
rect -1082 -553 -1058 -519
rect -1140 -587 -1058 -553
rect -1140 -621 -1116 -587
rect -1082 -621 -1058 -587
rect -1140 -655 -1058 -621
rect -1140 -689 -1116 -655
rect -1082 -689 -1058 -655
rect -1140 -723 -1058 -689
rect -1140 -757 -1116 -723
rect -1082 -757 -1058 -723
rect -1140 -791 -1058 -757
rect -1140 -825 -1116 -791
rect -1082 -825 -1058 -791
rect -1140 -859 -1058 -825
rect -1140 -893 -1116 -859
rect -1082 -893 -1058 -859
rect -1140 -927 -1058 -893
rect -1140 -961 -1116 -927
rect -1082 -961 -1058 -927
rect -1140 -995 -1058 -961
rect -1140 -1029 -1116 -995
rect -1082 -1029 -1058 -995
rect 1208 -9 1232 25
rect 1266 -9 1290 25
rect 1208 -43 1290 -9
rect 1208 -77 1232 -43
rect 1266 -77 1290 -43
rect 1208 -111 1290 -77
rect 1208 -145 1232 -111
rect 1266 -145 1290 -111
rect 1208 -179 1290 -145
rect 1208 -213 1232 -179
rect 1266 -213 1290 -179
rect 1208 -247 1290 -213
rect 1208 -281 1232 -247
rect 1266 -281 1290 -247
rect 1208 -315 1290 -281
rect 1208 -349 1232 -315
rect 1266 -349 1290 -315
rect 1208 -383 1290 -349
rect 1208 -417 1232 -383
rect 1266 -417 1290 -383
rect 1208 -451 1290 -417
rect 1208 -485 1232 -451
rect 1266 -485 1290 -451
rect 1208 -519 1290 -485
rect 1208 -553 1232 -519
rect 1266 -553 1290 -519
rect 1208 -587 1290 -553
rect 1208 -621 1232 -587
rect 1266 -621 1290 -587
rect 1208 -655 1290 -621
rect 1208 -689 1232 -655
rect 1266 -689 1290 -655
rect 1208 -723 1290 -689
rect 1208 -757 1232 -723
rect 1266 -757 1290 -723
rect 1208 -791 1290 -757
rect 1208 -825 1232 -791
rect 1266 -825 1290 -791
rect 1208 -859 1290 -825
rect 1208 -893 1232 -859
rect 1266 -893 1290 -859
rect 1208 -927 1290 -893
rect 1208 -961 1232 -927
rect 1266 -961 1290 -927
rect 1208 -995 1290 -961
rect -1140 -1100 -1058 -1029
rect 1208 -1029 1232 -995
rect 1266 -1029 1290 -995
rect 1208 -1100 1290 -1029
rect -1140 -1124 1290 -1100
rect -1140 -1158 -866 -1124
rect -832 -1158 -798 -1124
rect -764 -1158 -730 -1124
rect -696 -1158 -662 -1124
rect -628 -1158 -594 -1124
rect -560 -1158 -526 -1124
rect -492 -1158 -458 -1124
rect -424 -1158 -390 -1124
rect -356 -1158 -322 -1124
rect -288 -1158 -254 -1124
rect -220 -1158 -186 -1124
rect -152 -1158 -118 -1124
rect -84 -1158 -50 -1124
rect -16 -1158 18 -1124
rect 52 -1158 86 -1124
rect 120 -1158 154 -1124
rect 188 -1158 222 -1124
rect 256 -1158 290 -1124
rect 324 -1158 358 -1124
rect 392 -1158 426 -1124
rect 460 -1158 494 -1124
rect 528 -1158 562 -1124
rect 596 -1158 630 -1124
rect 664 -1158 698 -1124
rect 732 -1158 766 -1124
rect 800 -1158 834 -1124
rect 868 -1158 902 -1124
rect 936 -1158 970 -1124
rect 1004 -1158 1290 -1124
rect -1140 -1182 1290 -1158
<< mvnsubdiff >>
tri 0 5970 30 6000 se
rect 30 5970 120 6000
tri 120 5970 150 6000 sw
rect 0 5941 150 5970
rect 0 59 24 5941
rect 126 59 150 5941
rect 0 30 150 59
tri 0 0 30 30 ne
rect 30 0 120 30
tri 120 0 150 30 nw
<< mvpsubdiffcont >>
rect -866 7124 -832 7158
rect -798 7124 -764 7158
rect -730 7124 -696 7158
rect -662 7124 -628 7158
rect -594 7124 -560 7158
rect -526 7124 -492 7158
rect -458 7124 -424 7158
rect -390 7124 -356 7158
rect -322 7124 -288 7158
rect -254 7124 -220 7158
rect -186 7124 -152 7158
rect -118 7124 -84 7158
rect -50 7124 -16 7158
rect 18 7124 52 7158
rect 86 7124 120 7158
rect 154 7124 188 7158
rect 222 7124 256 7158
rect 290 7124 324 7158
rect 358 7124 392 7158
rect 426 7124 460 7158
rect 494 7124 528 7158
rect 562 7124 596 7158
rect 630 7124 664 7158
rect 698 7124 732 7158
rect 766 7124 800 7158
rect 834 7124 868 7158
rect 902 7124 936 7158
rect 970 7124 1004 7158
rect -1116 6995 -1082 7029
rect -1116 6927 -1082 6961
rect -1116 6859 -1082 6893
rect -1116 6791 -1082 6825
rect -1116 6723 -1082 6757
rect -1116 6655 -1082 6689
rect -1116 6587 -1082 6621
rect -1116 6519 -1082 6553
rect -1116 6451 -1082 6485
rect -1116 6383 -1082 6417
rect -1116 6315 -1082 6349
rect -1116 6247 -1082 6281
rect -1116 6179 -1082 6213
rect -1116 6111 -1082 6145
rect -1116 6043 -1082 6077
rect -1116 5975 -1082 6009
rect 1232 6995 1266 7029
rect 1232 6927 1266 6961
rect 1232 6859 1266 6893
rect 1232 6791 1266 6825
rect 1232 6723 1266 6757
rect 1232 6655 1266 6689
rect 1232 6587 1266 6621
rect 1232 6519 1266 6553
rect 1232 6451 1266 6485
rect 1232 6383 1266 6417
rect 1232 6315 1266 6349
rect 1232 6247 1266 6281
rect 1232 6179 1266 6213
rect 1232 6111 1266 6145
rect 1232 6043 1266 6077
rect -1116 5907 -1082 5941
rect -1116 5839 -1082 5873
rect -1116 5771 -1082 5805
rect -1116 5703 -1082 5737
rect -1116 5635 -1082 5669
rect -1116 5567 -1082 5601
rect -1116 5499 -1082 5533
rect -1116 5431 -1082 5465
rect -1116 5363 -1082 5397
rect -1116 5295 -1082 5329
rect -1116 5227 -1082 5261
rect -1116 5159 -1082 5193
rect -1116 5091 -1082 5125
rect -1116 5023 -1082 5057
rect -1116 4955 -1082 4989
rect -1116 4887 -1082 4921
rect -1116 4819 -1082 4853
rect -1116 4751 -1082 4785
rect -1116 4683 -1082 4717
rect -1116 4615 -1082 4649
rect -1116 4547 -1082 4581
rect -1116 4479 -1082 4513
rect -1116 4411 -1082 4445
rect -1116 4343 -1082 4377
rect -1116 4275 -1082 4309
rect -1116 4207 -1082 4241
rect -1116 4139 -1082 4173
rect -1116 4071 -1082 4105
rect -1116 4003 -1082 4037
rect -1116 3935 -1082 3969
rect -1116 3867 -1082 3901
rect -1116 3799 -1082 3833
rect -1116 3731 -1082 3765
rect -1116 3663 -1082 3697
rect -1116 3595 -1082 3629
rect -1116 3527 -1082 3561
rect -1116 3459 -1082 3493
rect -1116 3391 -1082 3425
rect -1116 3323 -1082 3357
rect -1116 3255 -1082 3289
rect -1116 3187 -1082 3221
rect -1116 3119 -1082 3153
rect -1116 3051 -1082 3085
rect -1116 2983 -1082 3017
rect -1116 2915 -1082 2949
rect -1116 2847 -1082 2881
rect -1116 2779 -1082 2813
rect -1116 2711 -1082 2745
rect -1116 2643 -1082 2677
rect -1116 2575 -1082 2609
rect -1116 2507 -1082 2541
rect -1116 2439 -1082 2473
rect -1116 2371 -1082 2405
rect -1116 2303 -1082 2337
rect -1116 2235 -1082 2269
rect -1116 2167 -1082 2201
rect -1116 2099 -1082 2133
rect -1116 2031 -1082 2065
rect -1116 1963 -1082 1997
rect -1116 1895 -1082 1929
rect -1116 1827 -1082 1861
rect -1116 1759 -1082 1793
rect -1116 1691 -1082 1725
rect -1116 1623 -1082 1657
rect -1116 1555 -1082 1589
rect -1116 1487 -1082 1521
rect -1116 1419 -1082 1453
rect -1116 1351 -1082 1385
rect -1116 1283 -1082 1317
rect -1116 1215 -1082 1249
rect -1116 1147 -1082 1181
rect -1116 1079 -1082 1113
rect -1116 1011 -1082 1045
rect -1116 943 -1082 977
rect -1116 875 -1082 909
rect -1116 807 -1082 841
rect -1116 739 -1082 773
rect -1116 671 -1082 705
rect -1116 603 -1082 637
rect -1116 535 -1082 569
rect -1116 467 -1082 501
rect -1116 399 -1082 433
rect -1116 331 -1082 365
rect -1116 263 -1082 297
rect -1116 195 -1082 229
rect -1116 127 -1082 161
rect -1116 59 -1082 93
rect -1116 -9 -1082 25
rect 1232 5975 1266 6009
rect 1232 5907 1266 5941
rect 1232 5839 1266 5873
rect 1232 5771 1266 5805
rect 1232 5703 1266 5737
rect 1232 5635 1266 5669
rect 1232 5567 1266 5601
rect 1232 5499 1266 5533
rect 1232 5431 1266 5465
rect 1232 5363 1266 5397
rect 1232 5295 1266 5329
rect 1232 5227 1266 5261
rect 1232 5159 1266 5193
rect 1232 5091 1266 5125
rect 1232 5023 1266 5057
rect 1232 4955 1266 4989
rect 1232 4887 1266 4921
rect 1232 4819 1266 4853
rect 1232 4751 1266 4785
rect 1232 4683 1266 4717
rect 1232 4615 1266 4649
rect 1232 4547 1266 4581
rect 1232 4479 1266 4513
rect 1232 4411 1266 4445
rect 1232 4343 1266 4377
rect 1232 4275 1266 4309
rect 1232 4207 1266 4241
rect 1232 4139 1266 4173
rect 1232 4071 1266 4105
rect 1232 4003 1266 4037
rect 1232 3935 1266 3969
rect 1232 3867 1266 3901
rect 1232 3799 1266 3833
rect 1232 3731 1266 3765
rect 1232 3663 1266 3697
rect 1232 3595 1266 3629
rect 1232 3527 1266 3561
rect 1232 3459 1266 3493
rect 1232 3391 1266 3425
rect 1232 3323 1266 3357
rect 1232 3255 1266 3289
rect 1232 3187 1266 3221
rect 1232 3119 1266 3153
rect 1232 3051 1266 3085
rect 1232 2983 1266 3017
rect 1232 2915 1266 2949
rect 1232 2847 1266 2881
rect 1232 2779 1266 2813
rect 1232 2711 1266 2745
rect 1232 2643 1266 2677
rect 1232 2575 1266 2609
rect 1232 2507 1266 2541
rect 1232 2439 1266 2473
rect 1232 2371 1266 2405
rect 1232 2303 1266 2337
rect 1232 2235 1266 2269
rect 1232 2167 1266 2201
rect 1232 2099 1266 2133
rect 1232 2031 1266 2065
rect 1232 1963 1266 1997
rect 1232 1895 1266 1929
rect 1232 1827 1266 1861
rect 1232 1759 1266 1793
rect 1232 1691 1266 1725
rect 1232 1623 1266 1657
rect 1232 1555 1266 1589
rect 1232 1487 1266 1521
rect 1232 1419 1266 1453
rect 1232 1351 1266 1385
rect 1232 1283 1266 1317
rect 1232 1215 1266 1249
rect 1232 1147 1266 1181
rect 1232 1079 1266 1113
rect 1232 1011 1266 1045
rect 1232 943 1266 977
rect 1232 875 1266 909
rect 1232 807 1266 841
rect 1232 739 1266 773
rect 1232 671 1266 705
rect 1232 603 1266 637
rect 1232 535 1266 569
rect 1232 467 1266 501
rect 1232 399 1266 433
rect 1232 331 1266 365
rect 1232 263 1266 297
rect 1232 195 1266 229
rect 1232 127 1266 161
rect 1232 59 1266 93
rect -1116 -77 -1082 -43
rect -1116 -145 -1082 -111
rect -1116 -213 -1082 -179
rect -1116 -281 -1082 -247
rect -1116 -349 -1082 -315
rect -1116 -417 -1082 -383
rect -1116 -485 -1082 -451
rect -1116 -553 -1082 -519
rect -1116 -621 -1082 -587
rect -1116 -689 -1082 -655
rect -1116 -757 -1082 -723
rect -1116 -825 -1082 -791
rect -1116 -893 -1082 -859
rect -1116 -961 -1082 -927
rect -1116 -1029 -1082 -995
rect 1232 -9 1266 25
rect 1232 -77 1266 -43
rect 1232 -145 1266 -111
rect 1232 -213 1266 -179
rect 1232 -281 1266 -247
rect 1232 -349 1266 -315
rect 1232 -417 1266 -383
rect 1232 -485 1266 -451
rect 1232 -553 1266 -519
rect 1232 -621 1266 -587
rect 1232 -689 1266 -655
rect 1232 -757 1266 -723
rect 1232 -825 1266 -791
rect 1232 -893 1266 -859
rect 1232 -961 1266 -927
rect 1232 -1029 1266 -995
rect -866 -1158 -832 -1124
rect -798 -1158 -764 -1124
rect -730 -1158 -696 -1124
rect -662 -1158 -628 -1124
rect -594 -1158 -560 -1124
rect -526 -1158 -492 -1124
rect -458 -1158 -424 -1124
rect -390 -1158 -356 -1124
rect -322 -1158 -288 -1124
rect -254 -1158 -220 -1124
rect -186 -1158 -152 -1124
rect -118 -1158 -84 -1124
rect -50 -1158 -16 -1124
rect 18 -1158 52 -1124
rect 86 -1158 120 -1124
rect 154 -1158 188 -1124
rect 222 -1158 256 -1124
rect 290 -1158 324 -1124
rect 358 -1158 392 -1124
rect 426 -1158 460 -1124
rect 494 -1158 528 -1124
rect 562 -1158 596 -1124
rect 630 -1158 664 -1124
rect 698 -1158 732 -1124
rect 766 -1158 800 -1124
rect 834 -1158 868 -1124
rect 902 -1158 936 -1124
rect 970 -1158 1004 -1124
<< mvnsubdiffcont >>
rect 24 59 126 5941
<< poly >>
rect -900 6400 1050 7000
rect -900 6000 -300 6400
rect 450 6000 1050 6400
rect -600 0 -300 6000
rect 450 0 750 6000
rect -900 -400 -300 0
rect 450 -400 1050 0
rect -900 -659 1050 -400
rect -900 -693 -280 -659
rect -246 -693 -206 -659
rect -172 -693 -132 -659
rect -98 -693 -58 -659
rect -24 -693 16 -659
rect 50 -693 90 -659
rect 124 -693 164 -659
rect 198 -693 238 -659
rect 272 -693 312 -659
rect 346 -693 386 -659
rect 420 -693 1050 -659
rect -900 -733 1050 -693
rect -900 -767 -280 -733
rect -246 -767 -206 -733
rect -172 -767 -132 -733
rect -98 -767 -58 -733
rect -24 -767 16 -733
rect 50 -767 90 -733
rect 124 -767 164 -733
rect 198 -767 238 -733
rect 272 -767 312 -733
rect 346 -767 386 -733
rect 420 -767 1050 -733
rect -900 -807 1050 -767
rect -900 -841 -280 -807
rect -246 -841 -206 -807
rect -172 -841 -132 -807
rect -98 -841 -58 -807
rect -24 -841 16 -807
rect 50 -841 90 -807
rect 124 -841 164 -807
rect 198 -841 238 -807
rect 272 -841 312 -807
rect 346 -841 386 -807
rect 420 -841 1050 -807
rect -900 -1000 1050 -841
<< polycont >>
rect -280 -693 -246 -659
rect -206 -693 -172 -659
rect -132 -693 -98 -659
rect -58 -693 -24 -659
rect 16 -693 50 -659
rect 90 -693 124 -659
rect 164 -693 198 -659
rect 238 -693 272 -659
rect 312 -693 346 -659
rect 386 -693 420 -659
rect -280 -767 -246 -733
rect -206 -767 -172 -733
rect -132 -767 -98 -733
rect -58 -767 -24 -733
rect 16 -767 50 -733
rect 90 -767 124 -733
rect 164 -767 198 -733
rect 238 -767 272 -733
rect 312 -767 346 -733
rect 386 -767 420 -733
rect -280 -841 -246 -807
rect -206 -841 -172 -807
rect -132 -841 -98 -807
rect -58 -841 -24 -807
rect 16 -841 50 -807
rect 90 -841 124 -807
rect 164 -841 198 -807
rect 238 -841 272 -807
rect 312 -841 346 -807
rect 386 -841 420 -807
<< locali >>
rect -1140 7158 1290 7182
rect -1140 7124 -986 7158
rect -952 7124 -914 7158
rect -880 7124 -866 7158
rect -808 7124 -798 7158
rect -736 7124 -730 7158
rect -664 7124 -662 7158
rect -628 7124 -626 7158
rect -560 7124 -554 7158
rect -492 7124 -482 7158
rect -424 7124 -410 7158
rect -356 7124 -338 7158
rect -288 7124 -266 7158
rect -220 7124 -194 7158
rect -152 7124 -122 7158
rect -84 7124 -50 7158
rect -16 7124 18 7158
rect 56 7124 86 7158
rect 128 7124 154 7158
rect 200 7124 222 7158
rect 272 7124 290 7158
rect 344 7124 358 7158
rect 416 7124 426 7158
rect 488 7124 494 7158
rect 560 7124 562 7158
rect 596 7124 598 7158
rect 664 7124 670 7158
rect 732 7124 742 7158
rect 800 7124 814 7158
rect 868 7124 886 7158
rect 936 7124 958 7158
rect 1004 7124 1030 7158
rect 1064 7124 1102 7158
rect 1136 7124 1290 7158
rect -1140 7100 1290 7124
rect -1140 7085 -1058 7100
rect -1140 7051 -1116 7085
rect -1082 7051 -1058 7085
rect -1140 7029 -1058 7051
rect -1140 6979 -1116 7029
rect -1082 6979 -1058 7029
rect -1140 6961 -1058 6979
rect -1140 6907 -1116 6961
rect -1082 6907 -1058 6961
rect -1140 6893 -1058 6907
rect -1140 6835 -1116 6893
rect -1082 6835 -1058 6893
rect -1140 6825 -1058 6835
rect -1140 6763 -1116 6825
rect -1082 6763 -1058 6825
rect -1140 6757 -1058 6763
rect -1140 6691 -1116 6757
rect -1082 6691 -1058 6757
rect -1140 6689 -1058 6691
rect -1140 6655 -1116 6689
rect -1082 6655 -1058 6689
rect -1140 6653 -1058 6655
rect -1140 6587 -1116 6653
rect -1082 6587 -1058 6653
rect -1140 6581 -1058 6587
rect -1140 6519 -1116 6581
rect -1082 6519 -1058 6581
rect -1140 6509 -1058 6519
rect -1140 6451 -1116 6509
rect -1082 6451 -1058 6509
rect -1140 6437 -1058 6451
rect -1140 6383 -1116 6437
rect -1082 6383 -1058 6437
rect -1140 6365 -1058 6383
rect -1140 6315 -1116 6365
rect -1082 6315 -1058 6365
rect -1140 6293 -1058 6315
rect -1140 6247 -1116 6293
rect -1082 6247 -1058 6293
rect -1140 6221 -1058 6247
rect -1140 6179 -1116 6221
rect -1082 6179 -1058 6221
rect -1140 6149 -1058 6179
rect -1140 6111 -1116 6149
rect -1082 6111 -1058 6149
rect -1140 6077 -1058 6111
rect -1140 6043 -1116 6077
rect -1082 6043 -1058 6077
rect -1140 6009 -1058 6043
rect -1140 5971 -1116 6009
rect -1082 5971 -1058 6009
rect 1208 7085 1290 7100
rect 1208 7051 1232 7085
rect 1266 7051 1290 7085
rect 1208 7029 1290 7051
rect 1208 6979 1232 7029
rect 1266 6979 1290 7029
rect 1208 6961 1290 6979
rect 1208 6907 1232 6961
rect 1266 6907 1290 6961
rect 1208 6893 1290 6907
rect 1208 6835 1232 6893
rect 1266 6835 1290 6893
rect 1208 6825 1290 6835
rect 1208 6763 1232 6825
rect 1266 6763 1290 6825
rect 1208 6757 1290 6763
rect 1208 6691 1232 6757
rect 1266 6691 1290 6757
rect 1208 6689 1290 6691
rect 1208 6655 1232 6689
rect 1266 6655 1290 6689
rect 1208 6653 1290 6655
rect 1208 6587 1232 6653
rect 1266 6587 1290 6653
rect 1208 6581 1290 6587
rect 1208 6519 1232 6581
rect 1266 6519 1290 6581
rect 1208 6509 1290 6519
rect 1208 6451 1232 6509
rect 1266 6451 1290 6509
rect 1208 6437 1290 6451
rect 1208 6383 1232 6437
rect 1266 6383 1290 6437
rect 1208 6365 1290 6383
rect 1208 6315 1232 6365
rect 1266 6315 1290 6365
rect 1208 6293 1290 6315
rect 1208 6247 1232 6293
rect 1266 6247 1290 6293
rect 1208 6221 1290 6247
rect 1208 6179 1232 6221
rect 1266 6179 1290 6221
rect 1208 6149 1290 6179
rect 1208 6111 1232 6149
rect 1266 6111 1290 6149
rect 1208 6077 1290 6111
rect 1208 6043 1232 6077
rect 1266 6043 1290 6077
rect 1208 6009 1290 6043
rect -1140 5941 -1058 5971
rect -1140 5899 -1116 5941
rect -1082 5899 -1058 5941
rect -1140 5873 -1058 5899
rect -1140 5827 -1116 5873
rect -1082 5827 -1058 5873
rect -1140 5805 -1058 5827
rect -1140 5755 -1116 5805
rect -1082 5755 -1058 5805
rect -1140 5737 -1058 5755
rect -1140 5683 -1116 5737
rect -1082 5683 -1058 5737
rect -1140 5669 -1058 5683
rect -1140 5611 -1116 5669
rect -1082 5611 -1058 5669
rect -1140 5601 -1058 5611
rect -1140 5539 -1116 5601
rect -1082 5539 -1058 5601
rect -1140 5533 -1058 5539
rect -1140 5467 -1116 5533
rect -1082 5467 -1058 5533
rect -1140 5465 -1058 5467
rect -1140 5431 -1116 5465
rect -1082 5431 -1058 5465
rect -1140 5429 -1058 5431
rect -1140 5363 -1116 5429
rect -1082 5363 -1058 5429
rect -1140 5357 -1058 5363
rect -1140 5295 -1116 5357
rect -1082 5295 -1058 5357
rect -1140 5285 -1058 5295
rect -1140 5227 -1116 5285
rect -1082 5227 -1058 5285
rect -1140 5213 -1058 5227
rect -1140 5159 -1116 5213
rect -1082 5159 -1058 5213
rect -1140 5141 -1058 5159
rect -1140 5091 -1116 5141
rect -1082 5091 -1058 5141
rect -1140 5069 -1058 5091
rect -1140 5023 -1116 5069
rect -1082 5023 -1058 5069
rect -1140 4997 -1058 5023
rect -1140 4955 -1116 4997
rect -1082 4955 -1058 4997
rect -1140 4925 -1058 4955
rect -1140 4887 -1116 4925
rect -1082 4887 -1058 4925
rect -1140 4853 -1058 4887
rect -1140 4819 -1116 4853
rect -1082 4819 -1058 4853
rect -1140 4785 -1058 4819
rect -1140 4747 -1116 4785
rect -1082 4747 -1058 4785
rect -1140 4717 -1058 4747
rect -1140 4675 -1116 4717
rect -1082 4675 -1058 4717
rect -1140 4649 -1058 4675
rect -1140 4603 -1116 4649
rect -1082 4603 -1058 4649
rect -1140 4581 -1058 4603
rect -1140 4531 -1116 4581
rect -1082 4531 -1058 4581
rect -1140 4513 -1058 4531
rect -1140 4459 -1116 4513
rect -1082 4459 -1058 4513
rect -1140 4445 -1058 4459
rect -1140 4387 -1116 4445
rect -1082 4387 -1058 4445
rect -1140 4377 -1058 4387
rect -1140 4315 -1116 4377
rect -1082 4315 -1058 4377
rect -1140 4309 -1058 4315
rect -1140 4243 -1116 4309
rect -1082 4243 -1058 4309
rect -1140 4241 -1058 4243
rect -1140 4207 -1116 4241
rect -1082 4207 -1058 4241
rect -1140 4205 -1058 4207
rect -1140 4139 -1116 4205
rect -1082 4139 -1058 4205
rect -1140 4133 -1058 4139
rect -1140 4071 -1116 4133
rect -1082 4071 -1058 4133
rect -1140 4061 -1058 4071
rect -1140 4003 -1116 4061
rect -1082 4003 -1058 4061
rect -1140 3989 -1058 4003
rect -1140 3935 -1116 3989
rect -1082 3935 -1058 3989
rect -1140 3917 -1058 3935
rect -1140 3867 -1116 3917
rect -1082 3867 -1058 3917
rect -1140 3845 -1058 3867
rect -1140 3799 -1116 3845
rect -1082 3799 -1058 3845
rect -1140 3773 -1058 3799
rect -1140 3731 -1116 3773
rect -1082 3731 -1058 3773
rect -1140 3701 -1058 3731
rect -1140 3663 -1116 3701
rect -1082 3663 -1058 3701
rect -1140 3629 -1058 3663
rect -1140 3595 -1116 3629
rect -1082 3595 -1058 3629
rect -1140 3561 -1058 3595
rect -1140 3523 -1116 3561
rect -1082 3523 -1058 3561
rect -1140 3493 -1058 3523
rect -1140 3451 -1116 3493
rect -1082 3451 -1058 3493
rect -1140 3425 -1058 3451
rect -1140 3379 -1116 3425
rect -1082 3379 -1058 3425
rect -1140 3357 -1058 3379
rect -1140 3307 -1116 3357
rect -1082 3307 -1058 3357
rect -1140 3289 -1058 3307
rect -1140 3235 -1116 3289
rect -1082 3235 -1058 3289
rect -1140 3221 -1058 3235
rect -1140 3163 -1116 3221
rect -1082 3163 -1058 3221
rect -1140 3153 -1058 3163
rect -1140 3091 -1116 3153
rect -1082 3091 -1058 3153
rect -1140 3085 -1058 3091
rect -1140 3019 -1116 3085
rect -1082 3019 -1058 3085
rect -1140 3017 -1058 3019
rect -1140 2983 -1116 3017
rect -1082 2983 -1058 3017
rect -1140 2981 -1058 2983
rect -1140 2915 -1116 2981
rect -1082 2915 -1058 2981
rect -1140 2909 -1058 2915
rect -1140 2847 -1116 2909
rect -1082 2847 -1058 2909
rect -1140 2837 -1058 2847
rect -1140 2779 -1116 2837
rect -1082 2779 -1058 2837
rect -1140 2765 -1058 2779
rect -1140 2711 -1116 2765
rect -1082 2711 -1058 2765
rect -1140 2693 -1058 2711
rect -1140 2643 -1116 2693
rect -1082 2643 -1058 2693
rect -1140 2621 -1058 2643
rect -1140 2575 -1116 2621
rect -1082 2575 -1058 2621
rect -1140 2549 -1058 2575
rect -1140 2507 -1116 2549
rect -1082 2507 -1058 2549
rect -1140 2477 -1058 2507
rect -1140 2439 -1116 2477
rect -1082 2439 -1058 2477
rect -1140 2405 -1058 2439
rect -1140 2371 -1116 2405
rect -1082 2371 -1058 2405
rect -1140 2337 -1058 2371
rect -1140 2299 -1116 2337
rect -1082 2299 -1058 2337
rect -1140 2269 -1058 2299
rect -1140 2227 -1116 2269
rect -1082 2227 -1058 2269
rect -1140 2201 -1058 2227
rect -1140 2155 -1116 2201
rect -1082 2155 -1058 2201
rect -1140 2133 -1058 2155
rect -1140 2083 -1116 2133
rect -1082 2083 -1058 2133
rect -1140 2065 -1058 2083
rect -1140 2011 -1116 2065
rect -1082 2011 -1058 2065
rect -1140 1997 -1058 2011
rect -1140 1939 -1116 1997
rect -1082 1939 -1058 1997
rect -1140 1929 -1058 1939
rect -1140 1867 -1116 1929
rect -1082 1867 -1058 1929
rect -1140 1861 -1058 1867
rect -1140 1795 -1116 1861
rect -1082 1795 -1058 1861
rect -1140 1793 -1058 1795
rect -1140 1759 -1116 1793
rect -1082 1759 -1058 1793
rect -1140 1757 -1058 1759
rect -1140 1691 -1116 1757
rect -1082 1691 -1058 1757
rect -1140 1685 -1058 1691
rect -1140 1623 -1116 1685
rect -1082 1623 -1058 1685
rect -1140 1613 -1058 1623
rect -1140 1555 -1116 1613
rect -1082 1555 -1058 1613
rect -1140 1541 -1058 1555
rect -1140 1487 -1116 1541
rect -1082 1487 -1058 1541
rect -1140 1469 -1058 1487
rect -1140 1419 -1116 1469
rect -1082 1419 -1058 1469
rect -1140 1397 -1058 1419
rect -1140 1351 -1116 1397
rect -1082 1351 -1058 1397
rect -1140 1325 -1058 1351
rect -1140 1283 -1116 1325
rect -1082 1283 -1058 1325
rect -1140 1253 -1058 1283
rect -1140 1215 -1116 1253
rect -1082 1215 -1058 1253
rect -1140 1181 -1058 1215
rect -1140 1147 -1116 1181
rect -1082 1147 -1058 1181
rect -1140 1113 -1058 1147
rect -1140 1075 -1116 1113
rect -1082 1075 -1058 1113
rect -1140 1045 -1058 1075
rect -1140 1003 -1116 1045
rect -1082 1003 -1058 1045
rect -1140 977 -1058 1003
rect -1140 931 -1116 977
rect -1082 931 -1058 977
rect -1140 909 -1058 931
rect -1140 859 -1116 909
rect -1082 859 -1058 909
rect -1140 841 -1058 859
rect -1140 787 -1116 841
rect -1082 787 -1058 841
rect -1140 773 -1058 787
rect -1140 715 -1116 773
rect -1082 715 -1058 773
rect -1140 705 -1058 715
rect -1140 643 -1116 705
rect -1082 643 -1058 705
rect -1140 637 -1058 643
rect -1140 571 -1116 637
rect -1082 571 -1058 637
rect -1140 569 -1058 571
rect -1140 535 -1116 569
rect -1082 535 -1058 569
rect -1140 533 -1058 535
rect -1140 467 -1116 533
rect -1082 467 -1058 533
rect -1140 461 -1058 467
rect -1140 399 -1116 461
rect -1082 399 -1058 461
rect -1140 389 -1058 399
rect -1140 331 -1116 389
rect -1082 331 -1058 389
rect -1140 317 -1058 331
rect -1140 263 -1116 317
rect -1082 263 -1058 317
rect -1140 245 -1058 263
rect -1140 195 -1116 245
rect -1082 195 -1058 245
rect -1140 173 -1058 195
rect -1140 127 -1116 173
rect -1082 127 -1058 173
rect -1140 101 -1058 127
rect -1140 59 -1116 101
rect -1082 59 -1058 101
rect -1140 29 -1058 59
rect -1140 -9 -1116 29
rect -1082 -9 -1058 29
rect -962 5975 -896 5991
rect -962 5935 -946 5975
rect -912 5935 -896 5975
rect 1046 5975 1112 5991
rect -962 5907 -896 5935
rect -962 5863 -946 5907
rect -912 5863 -896 5907
rect -962 5839 -896 5863
rect -962 5791 -946 5839
rect -912 5791 -896 5839
rect -962 5771 -896 5791
rect -962 5719 -946 5771
rect -912 5719 -896 5771
rect -962 5703 -896 5719
rect -962 5647 -946 5703
rect -912 5647 -896 5703
rect -962 5635 -896 5647
rect -962 5575 -946 5635
rect -912 5575 -896 5635
rect -962 5567 -896 5575
rect -962 5503 -946 5567
rect -912 5503 -896 5567
rect -962 5499 -896 5503
rect -962 5397 -946 5499
rect -912 5397 -896 5499
rect -962 5393 -896 5397
rect -962 5329 -946 5393
rect -912 5329 -896 5393
rect -962 5321 -896 5329
rect -962 5261 -946 5321
rect -912 5261 -896 5321
rect -962 5249 -896 5261
rect -962 5193 -946 5249
rect -912 5193 -896 5249
rect -962 5177 -896 5193
rect -962 5125 -946 5177
rect -912 5125 -896 5177
rect -962 5105 -896 5125
rect -962 5057 -946 5105
rect -912 5057 -896 5105
rect -962 5033 -896 5057
rect -962 4989 -946 5033
rect -912 4989 -896 5033
rect -962 4961 -896 4989
rect -962 4921 -946 4961
rect -912 4921 -896 4961
rect -962 4889 -896 4921
rect -962 4853 -946 4889
rect -912 4853 -896 4889
rect -962 4819 -896 4853
rect -962 4783 -946 4819
rect -912 4783 -896 4819
rect -962 4751 -896 4783
rect -962 4711 -946 4751
rect -912 4711 -896 4751
rect -962 4683 -896 4711
rect -962 4639 -946 4683
rect -912 4639 -896 4683
rect -962 4615 -896 4639
rect -962 4567 -946 4615
rect -912 4567 -896 4615
rect -962 4547 -896 4567
rect -962 4495 -946 4547
rect -912 4495 -896 4547
rect -962 4479 -896 4495
rect -962 4423 -946 4479
rect -912 4423 -896 4479
rect -962 4411 -896 4423
rect -962 4351 -946 4411
rect -912 4351 -896 4411
rect -962 4343 -896 4351
rect -962 4279 -946 4343
rect -912 4279 -896 4343
rect -962 4275 -896 4279
rect -962 4173 -946 4275
rect -912 4173 -896 4275
rect -962 4169 -896 4173
rect -962 4105 -946 4169
rect -912 4105 -896 4169
rect -962 4097 -896 4105
rect -962 4037 -946 4097
rect -912 4037 -896 4097
rect -962 4025 -896 4037
rect -962 3969 -946 4025
rect -912 3969 -896 4025
rect -962 3953 -896 3969
rect -962 3901 -946 3953
rect -912 3901 -896 3953
rect -962 3881 -896 3901
rect -962 3833 -946 3881
rect -912 3833 -896 3881
rect -962 3809 -896 3833
rect -962 3765 -946 3809
rect -912 3765 -896 3809
rect -962 3737 -896 3765
rect -962 3697 -946 3737
rect -912 3697 -896 3737
rect -962 3665 -896 3697
rect -962 3629 -946 3665
rect -912 3629 -896 3665
rect -962 3595 -896 3629
rect -962 3559 -946 3595
rect -912 3559 -896 3595
rect -962 3527 -896 3559
rect -962 3487 -946 3527
rect -912 3487 -896 3527
rect -962 3459 -896 3487
rect -962 3415 -946 3459
rect -912 3415 -896 3459
rect -962 3391 -896 3415
rect -962 3343 -946 3391
rect -912 3343 -896 3391
rect -962 3323 -896 3343
rect -962 3271 -946 3323
rect -912 3271 -896 3323
rect -962 3255 -896 3271
rect -962 3199 -946 3255
rect -912 3199 -896 3255
rect -962 3187 -896 3199
rect -962 3127 -946 3187
rect -912 3127 -896 3187
rect -962 3119 -896 3127
rect -962 3055 -946 3119
rect -912 3055 -896 3119
rect -962 3051 -896 3055
rect -962 2949 -946 3051
rect -912 2949 -896 3051
rect -962 2945 -896 2949
rect -962 2881 -946 2945
rect -912 2881 -896 2945
rect -962 2873 -896 2881
rect -962 2813 -946 2873
rect -912 2813 -896 2873
rect -962 2801 -896 2813
rect -962 2745 -946 2801
rect -912 2745 -896 2801
rect -962 2729 -896 2745
rect -962 2677 -946 2729
rect -912 2677 -896 2729
rect -962 2657 -896 2677
rect -962 2609 -946 2657
rect -912 2609 -896 2657
rect -962 2585 -896 2609
rect -962 2541 -946 2585
rect -912 2541 -896 2585
rect -962 2513 -896 2541
rect -962 2473 -946 2513
rect -912 2473 -896 2513
rect -962 2441 -896 2473
rect -962 2405 -946 2441
rect -912 2405 -896 2441
rect -962 2371 -896 2405
rect -962 2335 -946 2371
rect -912 2335 -896 2371
rect -962 2303 -896 2335
rect -962 2263 -946 2303
rect -912 2263 -896 2303
rect -962 2235 -896 2263
rect -962 2191 -946 2235
rect -912 2191 -896 2235
rect -962 2167 -896 2191
rect -962 2119 -946 2167
rect -912 2119 -896 2167
rect -962 2099 -896 2119
rect -962 2047 -946 2099
rect -912 2047 -896 2099
rect -962 2031 -896 2047
rect -962 1975 -946 2031
rect -912 1975 -896 2031
rect -962 1963 -896 1975
rect -962 1903 -946 1963
rect -912 1903 -896 1963
rect -962 1895 -896 1903
rect -962 1831 -946 1895
rect -912 1831 -896 1895
rect -962 1827 -896 1831
rect -962 1725 -946 1827
rect -912 1725 -896 1827
rect -962 1721 -896 1725
rect -962 1657 -946 1721
rect -912 1657 -896 1721
rect -962 1649 -896 1657
rect -962 1589 -946 1649
rect -912 1589 -896 1649
rect -962 1577 -896 1589
rect -962 1521 -946 1577
rect -912 1521 -896 1577
rect -962 1505 -896 1521
rect -962 1453 -946 1505
rect -912 1453 -896 1505
rect -962 1433 -896 1453
rect -962 1385 -946 1433
rect -912 1385 -896 1433
rect -962 1361 -896 1385
rect -962 1317 -946 1361
rect -912 1317 -896 1361
rect -962 1289 -896 1317
rect -962 1249 -946 1289
rect -912 1249 -896 1289
rect -962 1217 -896 1249
rect -962 1181 -946 1217
rect -912 1181 -896 1217
rect -962 1147 -896 1181
rect -962 1111 -946 1147
rect -912 1111 -896 1147
rect -962 1079 -896 1111
rect -962 1039 -946 1079
rect -912 1039 -896 1079
rect -962 1011 -896 1039
rect -962 967 -946 1011
rect -912 967 -896 1011
rect -962 943 -896 967
rect -962 895 -946 943
rect -912 895 -896 943
rect -962 875 -896 895
rect -962 823 -946 875
rect -912 823 -896 875
rect -962 807 -896 823
rect -962 751 -946 807
rect -912 751 -896 807
rect -962 739 -896 751
rect -962 679 -946 739
rect -912 679 -896 739
rect -962 671 -896 679
rect -962 607 -946 671
rect -912 607 -896 671
rect -962 603 -896 607
rect -962 501 -946 603
rect -912 501 -896 603
rect -962 497 -896 501
rect -962 433 -946 497
rect -912 433 -896 497
rect -962 425 -896 433
rect -962 365 -946 425
rect -912 365 -896 425
rect -962 353 -896 365
rect -962 297 -946 353
rect -912 297 -896 353
rect -962 281 -896 297
rect -962 229 -946 281
rect -912 229 -896 281
rect -962 209 -896 229
rect -962 161 -946 209
rect -912 161 -896 209
rect -962 137 -896 161
rect -962 93 -946 137
rect -912 93 -896 137
rect -962 65 -896 93
rect -962 25 -946 65
rect -912 25 -896 65
rect 8 5941 142 5957
rect 8 5933 24 5941
rect 126 5933 142 5941
rect 8 67 22 5933
rect 128 67 142 5933
rect 8 59 24 67
rect 126 59 142 67
rect 8 43 142 59
rect 1046 5935 1062 5975
rect 1096 5935 1112 5975
rect 1046 5907 1112 5935
rect 1046 5863 1062 5907
rect 1096 5863 1112 5907
rect 1046 5839 1112 5863
rect 1046 5791 1062 5839
rect 1096 5791 1112 5839
rect 1046 5771 1112 5791
rect 1046 5719 1062 5771
rect 1096 5719 1112 5771
rect 1046 5703 1112 5719
rect 1046 5647 1062 5703
rect 1096 5647 1112 5703
rect 1046 5635 1112 5647
rect 1046 5575 1062 5635
rect 1096 5575 1112 5635
rect 1046 5567 1112 5575
rect 1046 5503 1062 5567
rect 1096 5503 1112 5567
rect 1046 5499 1112 5503
rect 1046 5397 1062 5499
rect 1096 5397 1112 5499
rect 1046 5393 1112 5397
rect 1046 5329 1062 5393
rect 1096 5329 1112 5393
rect 1046 5321 1112 5329
rect 1046 5261 1062 5321
rect 1096 5261 1112 5321
rect 1046 5249 1112 5261
rect 1046 5193 1062 5249
rect 1096 5193 1112 5249
rect 1046 5177 1112 5193
rect 1046 5125 1062 5177
rect 1096 5125 1112 5177
rect 1046 5105 1112 5125
rect 1046 5057 1062 5105
rect 1096 5057 1112 5105
rect 1046 5033 1112 5057
rect 1046 4989 1062 5033
rect 1096 4989 1112 5033
rect 1046 4961 1112 4989
rect 1046 4921 1062 4961
rect 1096 4921 1112 4961
rect 1046 4889 1112 4921
rect 1046 4853 1062 4889
rect 1096 4853 1112 4889
rect 1046 4819 1112 4853
rect 1046 4783 1062 4819
rect 1096 4783 1112 4819
rect 1046 4751 1112 4783
rect 1046 4711 1062 4751
rect 1096 4711 1112 4751
rect 1046 4683 1112 4711
rect 1046 4639 1062 4683
rect 1096 4639 1112 4683
rect 1046 4615 1112 4639
rect 1046 4567 1062 4615
rect 1096 4567 1112 4615
rect 1046 4547 1112 4567
rect 1046 4495 1062 4547
rect 1096 4495 1112 4547
rect 1046 4479 1112 4495
rect 1046 4423 1062 4479
rect 1096 4423 1112 4479
rect 1046 4411 1112 4423
rect 1046 4351 1062 4411
rect 1096 4351 1112 4411
rect 1046 4343 1112 4351
rect 1046 4279 1062 4343
rect 1096 4279 1112 4343
rect 1046 4275 1112 4279
rect 1046 4173 1062 4275
rect 1096 4173 1112 4275
rect 1046 4169 1112 4173
rect 1046 4105 1062 4169
rect 1096 4105 1112 4169
rect 1046 4097 1112 4105
rect 1046 4037 1062 4097
rect 1096 4037 1112 4097
rect 1046 4025 1112 4037
rect 1046 3969 1062 4025
rect 1096 3969 1112 4025
rect 1046 3953 1112 3969
rect 1046 3901 1062 3953
rect 1096 3901 1112 3953
rect 1046 3881 1112 3901
rect 1046 3833 1062 3881
rect 1096 3833 1112 3881
rect 1046 3809 1112 3833
rect 1046 3765 1062 3809
rect 1096 3765 1112 3809
rect 1046 3737 1112 3765
rect 1046 3697 1062 3737
rect 1096 3697 1112 3737
rect 1046 3665 1112 3697
rect 1046 3629 1062 3665
rect 1096 3629 1112 3665
rect 1046 3595 1112 3629
rect 1046 3559 1062 3595
rect 1096 3559 1112 3595
rect 1046 3527 1112 3559
rect 1046 3487 1062 3527
rect 1096 3487 1112 3527
rect 1046 3459 1112 3487
rect 1046 3415 1062 3459
rect 1096 3415 1112 3459
rect 1046 3391 1112 3415
rect 1046 3343 1062 3391
rect 1096 3343 1112 3391
rect 1046 3323 1112 3343
rect 1046 3271 1062 3323
rect 1096 3271 1112 3323
rect 1046 3255 1112 3271
rect 1046 3199 1062 3255
rect 1096 3199 1112 3255
rect 1046 3187 1112 3199
rect 1046 3127 1062 3187
rect 1096 3127 1112 3187
rect 1046 3119 1112 3127
rect 1046 3055 1062 3119
rect 1096 3055 1112 3119
rect 1046 3051 1112 3055
rect 1046 2949 1062 3051
rect 1096 2949 1112 3051
rect 1046 2945 1112 2949
rect 1046 2881 1062 2945
rect 1096 2881 1112 2945
rect 1046 2873 1112 2881
rect 1046 2813 1062 2873
rect 1096 2813 1112 2873
rect 1046 2801 1112 2813
rect 1046 2745 1062 2801
rect 1096 2745 1112 2801
rect 1046 2729 1112 2745
rect 1046 2677 1062 2729
rect 1096 2677 1112 2729
rect 1046 2657 1112 2677
rect 1046 2609 1062 2657
rect 1096 2609 1112 2657
rect 1046 2585 1112 2609
rect 1046 2541 1062 2585
rect 1096 2541 1112 2585
rect 1046 2513 1112 2541
rect 1046 2473 1062 2513
rect 1096 2473 1112 2513
rect 1046 2441 1112 2473
rect 1046 2405 1062 2441
rect 1096 2405 1112 2441
rect 1046 2371 1112 2405
rect 1046 2335 1062 2371
rect 1096 2335 1112 2371
rect 1046 2303 1112 2335
rect 1046 2263 1062 2303
rect 1096 2263 1112 2303
rect 1046 2235 1112 2263
rect 1046 2191 1062 2235
rect 1096 2191 1112 2235
rect 1046 2167 1112 2191
rect 1046 2119 1062 2167
rect 1096 2119 1112 2167
rect 1046 2099 1112 2119
rect 1046 2047 1062 2099
rect 1096 2047 1112 2099
rect 1046 2031 1112 2047
rect 1046 1975 1062 2031
rect 1096 1975 1112 2031
rect 1046 1963 1112 1975
rect 1046 1903 1062 1963
rect 1096 1903 1112 1963
rect 1046 1895 1112 1903
rect 1046 1831 1062 1895
rect 1096 1831 1112 1895
rect 1046 1827 1112 1831
rect 1046 1725 1062 1827
rect 1096 1725 1112 1827
rect 1046 1721 1112 1725
rect 1046 1657 1062 1721
rect 1096 1657 1112 1721
rect 1046 1649 1112 1657
rect 1046 1589 1062 1649
rect 1096 1589 1112 1649
rect 1046 1577 1112 1589
rect 1046 1521 1062 1577
rect 1096 1521 1112 1577
rect 1046 1505 1112 1521
rect 1046 1453 1062 1505
rect 1096 1453 1112 1505
rect 1046 1433 1112 1453
rect 1046 1385 1062 1433
rect 1096 1385 1112 1433
rect 1046 1361 1112 1385
rect 1046 1317 1062 1361
rect 1096 1317 1112 1361
rect 1046 1289 1112 1317
rect 1046 1249 1062 1289
rect 1096 1249 1112 1289
rect 1046 1217 1112 1249
rect 1046 1181 1062 1217
rect 1096 1181 1112 1217
rect 1046 1147 1112 1181
rect 1046 1111 1062 1147
rect 1096 1111 1112 1147
rect 1046 1079 1112 1111
rect 1046 1039 1062 1079
rect 1096 1039 1112 1079
rect 1046 1011 1112 1039
rect 1046 967 1062 1011
rect 1096 967 1112 1011
rect 1046 943 1112 967
rect 1046 895 1062 943
rect 1096 895 1112 943
rect 1046 875 1112 895
rect 1046 823 1062 875
rect 1096 823 1112 875
rect 1046 807 1112 823
rect 1046 751 1062 807
rect 1096 751 1112 807
rect 1046 739 1112 751
rect 1046 679 1062 739
rect 1096 679 1112 739
rect 1046 671 1112 679
rect 1046 607 1062 671
rect 1096 607 1112 671
rect 1046 603 1112 607
rect 1046 501 1062 603
rect 1096 501 1112 603
rect 1046 497 1112 501
rect 1046 433 1062 497
rect 1096 433 1112 497
rect 1046 425 1112 433
rect 1046 365 1062 425
rect 1096 365 1112 425
rect 1046 353 1112 365
rect 1046 297 1062 353
rect 1096 297 1112 353
rect 1046 281 1112 297
rect 1046 229 1062 281
rect 1096 229 1112 281
rect 1046 209 1112 229
rect 1046 161 1062 209
rect 1096 161 1112 209
rect 1046 137 1112 161
rect 1046 93 1062 137
rect 1096 93 1112 137
rect 1046 65 1112 93
rect -962 9 -896 25
rect 1046 25 1062 65
rect 1096 25 1112 65
rect 1046 9 1112 25
rect 1208 5971 1232 6009
rect 1266 5971 1290 6009
rect 1208 5941 1290 5971
rect 1208 5899 1232 5941
rect 1266 5899 1290 5941
rect 1208 5873 1290 5899
rect 1208 5827 1232 5873
rect 1266 5827 1290 5873
rect 1208 5805 1290 5827
rect 1208 5755 1232 5805
rect 1266 5755 1290 5805
rect 1208 5737 1290 5755
rect 1208 5683 1232 5737
rect 1266 5683 1290 5737
rect 1208 5669 1290 5683
rect 1208 5611 1232 5669
rect 1266 5611 1290 5669
rect 1208 5601 1290 5611
rect 1208 5539 1232 5601
rect 1266 5539 1290 5601
rect 1208 5533 1290 5539
rect 1208 5467 1232 5533
rect 1266 5467 1290 5533
rect 1208 5465 1290 5467
rect 1208 5431 1232 5465
rect 1266 5431 1290 5465
rect 1208 5429 1290 5431
rect 1208 5363 1232 5429
rect 1266 5363 1290 5429
rect 1208 5357 1290 5363
rect 1208 5295 1232 5357
rect 1266 5295 1290 5357
rect 1208 5285 1290 5295
rect 1208 5227 1232 5285
rect 1266 5227 1290 5285
rect 1208 5213 1290 5227
rect 1208 5159 1232 5213
rect 1266 5159 1290 5213
rect 1208 5141 1290 5159
rect 1208 5091 1232 5141
rect 1266 5091 1290 5141
rect 1208 5069 1290 5091
rect 1208 5023 1232 5069
rect 1266 5023 1290 5069
rect 1208 4997 1290 5023
rect 1208 4955 1232 4997
rect 1266 4955 1290 4997
rect 1208 4925 1290 4955
rect 1208 4887 1232 4925
rect 1266 4887 1290 4925
rect 1208 4853 1290 4887
rect 1208 4819 1232 4853
rect 1266 4819 1290 4853
rect 1208 4785 1290 4819
rect 1208 4747 1232 4785
rect 1266 4747 1290 4785
rect 1208 4717 1290 4747
rect 1208 4675 1232 4717
rect 1266 4675 1290 4717
rect 1208 4649 1290 4675
rect 1208 4603 1232 4649
rect 1266 4603 1290 4649
rect 1208 4581 1290 4603
rect 1208 4531 1232 4581
rect 1266 4531 1290 4581
rect 1208 4513 1290 4531
rect 1208 4459 1232 4513
rect 1266 4459 1290 4513
rect 1208 4445 1290 4459
rect 1208 4387 1232 4445
rect 1266 4387 1290 4445
rect 1208 4377 1290 4387
rect 1208 4315 1232 4377
rect 1266 4315 1290 4377
rect 1208 4309 1290 4315
rect 1208 4243 1232 4309
rect 1266 4243 1290 4309
rect 1208 4241 1290 4243
rect 1208 4207 1232 4241
rect 1266 4207 1290 4241
rect 1208 4205 1290 4207
rect 1208 4139 1232 4205
rect 1266 4139 1290 4205
rect 1208 4133 1290 4139
rect 1208 4071 1232 4133
rect 1266 4071 1290 4133
rect 1208 4061 1290 4071
rect 1208 4003 1232 4061
rect 1266 4003 1290 4061
rect 1208 3989 1290 4003
rect 1208 3935 1232 3989
rect 1266 3935 1290 3989
rect 1208 3917 1290 3935
rect 1208 3867 1232 3917
rect 1266 3867 1290 3917
rect 1208 3845 1290 3867
rect 1208 3799 1232 3845
rect 1266 3799 1290 3845
rect 1208 3773 1290 3799
rect 1208 3731 1232 3773
rect 1266 3731 1290 3773
rect 1208 3701 1290 3731
rect 1208 3663 1232 3701
rect 1266 3663 1290 3701
rect 1208 3629 1290 3663
rect 1208 3595 1232 3629
rect 1266 3595 1290 3629
rect 1208 3561 1290 3595
rect 1208 3523 1232 3561
rect 1266 3523 1290 3561
rect 1208 3493 1290 3523
rect 1208 3451 1232 3493
rect 1266 3451 1290 3493
rect 1208 3425 1290 3451
rect 1208 3379 1232 3425
rect 1266 3379 1290 3425
rect 1208 3357 1290 3379
rect 1208 3307 1232 3357
rect 1266 3307 1290 3357
rect 1208 3289 1290 3307
rect 1208 3235 1232 3289
rect 1266 3235 1290 3289
rect 1208 3221 1290 3235
rect 1208 3163 1232 3221
rect 1266 3163 1290 3221
rect 1208 3153 1290 3163
rect 1208 3091 1232 3153
rect 1266 3091 1290 3153
rect 1208 3085 1290 3091
rect 1208 3019 1232 3085
rect 1266 3019 1290 3085
rect 1208 3017 1290 3019
rect 1208 2983 1232 3017
rect 1266 2983 1290 3017
rect 1208 2981 1290 2983
rect 1208 2915 1232 2981
rect 1266 2915 1290 2981
rect 1208 2909 1290 2915
rect 1208 2847 1232 2909
rect 1266 2847 1290 2909
rect 1208 2837 1290 2847
rect 1208 2779 1232 2837
rect 1266 2779 1290 2837
rect 1208 2765 1290 2779
rect 1208 2711 1232 2765
rect 1266 2711 1290 2765
rect 1208 2693 1290 2711
rect 1208 2643 1232 2693
rect 1266 2643 1290 2693
rect 1208 2621 1290 2643
rect 1208 2575 1232 2621
rect 1266 2575 1290 2621
rect 1208 2549 1290 2575
rect 1208 2507 1232 2549
rect 1266 2507 1290 2549
rect 1208 2477 1290 2507
rect 1208 2439 1232 2477
rect 1266 2439 1290 2477
rect 1208 2405 1290 2439
rect 1208 2371 1232 2405
rect 1266 2371 1290 2405
rect 1208 2337 1290 2371
rect 1208 2299 1232 2337
rect 1266 2299 1290 2337
rect 1208 2269 1290 2299
rect 1208 2227 1232 2269
rect 1266 2227 1290 2269
rect 1208 2201 1290 2227
rect 1208 2155 1232 2201
rect 1266 2155 1290 2201
rect 1208 2133 1290 2155
rect 1208 2083 1232 2133
rect 1266 2083 1290 2133
rect 1208 2065 1290 2083
rect 1208 2011 1232 2065
rect 1266 2011 1290 2065
rect 1208 1997 1290 2011
rect 1208 1939 1232 1997
rect 1266 1939 1290 1997
rect 1208 1929 1290 1939
rect 1208 1867 1232 1929
rect 1266 1867 1290 1929
rect 1208 1861 1290 1867
rect 1208 1795 1232 1861
rect 1266 1795 1290 1861
rect 1208 1793 1290 1795
rect 1208 1759 1232 1793
rect 1266 1759 1290 1793
rect 1208 1757 1290 1759
rect 1208 1691 1232 1757
rect 1266 1691 1290 1757
rect 1208 1685 1290 1691
rect 1208 1623 1232 1685
rect 1266 1623 1290 1685
rect 1208 1613 1290 1623
rect 1208 1555 1232 1613
rect 1266 1555 1290 1613
rect 1208 1541 1290 1555
rect 1208 1487 1232 1541
rect 1266 1487 1290 1541
rect 1208 1469 1290 1487
rect 1208 1419 1232 1469
rect 1266 1419 1290 1469
rect 1208 1397 1290 1419
rect 1208 1351 1232 1397
rect 1266 1351 1290 1397
rect 1208 1325 1290 1351
rect 1208 1283 1232 1325
rect 1266 1283 1290 1325
rect 1208 1253 1290 1283
rect 1208 1215 1232 1253
rect 1266 1215 1290 1253
rect 1208 1181 1290 1215
rect 1208 1147 1232 1181
rect 1266 1147 1290 1181
rect 1208 1113 1290 1147
rect 1208 1075 1232 1113
rect 1266 1075 1290 1113
rect 1208 1045 1290 1075
rect 1208 1003 1232 1045
rect 1266 1003 1290 1045
rect 1208 977 1290 1003
rect 1208 931 1232 977
rect 1266 931 1290 977
rect 1208 909 1290 931
rect 1208 859 1232 909
rect 1266 859 1290 909
rect 1208 841 1290 859
rect 1208 787 1232 841
rect 1266 787 1290 841
rect 1208 773 1290 787
rect 1208 715 1232 773
rect 1266 715 1290 773
rect 1208 705 1290 715
rect 1208 643 1232 705
rect 1266 643 1290 705
rect 1208 637 1290 643
rect 1208 571 1232 637
rect 1266 571 1290 637
rect 1208 569 1290 571
rect 1208 535 1232 569
rect 1266 535 1290 569
rect 1208 533 1290 535
rect 1208 467 1232 533
rect 1266 467 1290 533
rect 1208 461 1290 467
rect 1208 399 1232 461
rect 1266 399 1290 461
rect 1208 389 1290 399
rect 1208 331 1232 389
rect 1266 331 1290 389
rect 1208 317 1290 331
rect 1208 263 1232 317
rect 1266 263 1290 317
rect 1208 245 1290 263
rect 1208 195 1232 245
rect 1266 195 1290 245
rect 1208 173 1290 195
rect 1208 127 1232 173
rect 1266 127 1290 173
rect 1208 101 1290 127
rect 1208 59 1232 101
rect 1266 59 1290 101
rect 1208 29 1290 59
rect -1140 -43 -1058 -9
rect -1140 -77 -1116 -43
rect -1082 -77 -1058 -43
rect -1140 -111 -1058 -77
rect -1140 -149 -1116 -111
rect -1082 -149 -1058 -111
rect -1140 -179 -1058 -149
rect -1140 -221 -1116 -179
rect -1082 -221 -1058 -179
rect -1140 -247 -1058 -221
rect -1140 -293 -1116 -247
rect -1082 -293 -1058 -247
rect -1140 -315 -1058 -293
rect -1140 -365 -1116 -315
rect -1082 -365 -1058 -315
rect -1140 -383 -1058 -365
rect -1140 -437 -1116 -383
rect -1082 -437 -1058 -383
rect -1140 -451 -1058 -437
rect -1140 -509 -1116 -451
rect -1082 -509 -1058 -451
rect -1140 -519 -1058 -509
rect -1140 -581 -1116 -519
rect -1082 -581 -1058 -519
rect -1140 -587 -1058 -581
rect -1140 -653 -1116 -587
rect -1082 -653 -1058 -587
rect 1208 -9 1232 29
rect 1266 -9 1290 29
rect 1208 -43 1290 -9
rect 1208 -77 1232 -43
rect 1266 -77 1290 -43
rect 1208 -111 1290 -77
rect 1208 -149 1232 -111
rect 1266 -149 1290 -111
rect 1208 -179 1290 -149
rect 1208 -221 1232 -179
rect 1266 -221 1290 -179
rect 1208 -247 1290 -221
rect 1208 -293 1232 -247
rect 1266 -293 1290 -247
rect 1208 -315 1290 -293
rect 1208 -365 1232 -315
rect 1266 -365 1290 -315
rect 1208 -383 1290 -365
rect 1208 -437 1232 -383
rect 1266 -437 1290 -383
rect 1208 -451 1290 -437
rect 1208 -509 1232 -451
rect 1266 -509 1290 -451
rect 1208 -519 1290 -509
rect 1208 -581 1232 -519
rect 1266 -581 1290 -519
rect 1208 -587 1290 -581
rect -1140 -655 -1058 -653
rect -1140 -689 -1116 -655
rect -1082 -689 -1058 -655
rect -1140 -691 -1058 -689
rect -1140 -757 -1116 -691
rect -1082 -757 -1058 -691
rect -1140 -763 -1058 -757
rect -1140 -825 -1116 -763
rect -1082 -825 -1058 -763
rect -1140 -835 -1058 -825
rect -1140 -893 -1116 -835
rect -1082 -893 -1058 -835
rect -296 -659 460 -643
rect -296 -693 -280 -659
rect -246 -693 -206 -659
rect -172 -693 -132 -659
rect -98 -693 -58 -659
rect -24 -693 16 -659
rect 50 -693 90 -659
rect 124 -693 164 -659
rect 198 -693 238 -659
rect 272 -693 312 -659
rect 346 -693 386 -659
rect 420 -693 460 -659
rect -296 -733 460 -693
rect -296 -767 -280 -733
rect -246 -767 -206 -733
rect -172 -767 -132 -733
rect -98 -767 -58 -733
rect -24 -767 16 -733
rect 50 -767 90 -733
rect 124 -767 164 -733
rect 198 -767 238 -733
rect 272 -767 312 -733
rect 346 -767 386 -733
rect 420 -767 460 -733
rect -296 -807 460 -767
rect -296 -841 -280 -807
rect -246 -841 -206 -807
rect -172 -841 -132 -807
rect -98 -841 -58 -807
rect -24 -841 16 -807
rect 50 -841 90 -807
rect 124 -841 164 -807
rect 198 -841 238 -807
rect 272 -841 312 -807
rect 346 -841 386 -807
rect 420 -841 460 -807
rect -296 -857 460 -841
rect 1208 -653 1232 -587
rect 1266 -653 1290 -587
rect 1208 -655 1290 -653
rect 1208 -689 1232 -655
rect 1266 -689 1290 -655
rect 1208 -691 1290 -689
rect 1208 -757 1232 -691
rect 1266 -757 1290 -691
rect 1208 -763 1290 -757
rect 1208 -825 1232 -763
rect 1266 -825 1290 -763
rect 1208 -835 1290 -825
rect -1140 -907 -1058 -893
rect -1140 -961 -1116 -907
rect -1082 -961 -1058 -907
rect -1140 -979 -1058 -961
rect -1140 -1029 -1116 -979
rect -1082 -1029 -1058 -979
rect -1140 -1051 -1058 -1029
rect -1140 -1085 -1116 -1051
rect -1082 -1085 -1058 -1051
rect -1140 -1100 -1058 -1085
rect 1208 -893 1232 -835
rect 1266 -893 1290 -835
rect 1208 -907 1290 -893
rect 1208 -961 1232 -907
rect 1266 -961 1290 -907
rect 1208 -979 1290 -961
rect 1208 -1029 1232 -979
rect 1266 -1029 1290 -979
rect 1208 -1051 1290 -1029
rect 1208 -1085 1232 -1051
rect 1266 -1085 1290 -1051
rect 1208 -1100 1290 -1085
rect -1140 -1124 1290 -1100
rect -1140 -1158 -986 -1124
rect -952 -1158 -914 -1124
rect -880 -1158 -866 -1124
rect -808 -1158 -798 -1124
rect -736 -1158 -730 -1124
rect -664 -1158 -662 -1124
rect -628 -1158 -626 -1124
rect -560 -1158 -554 -1124
rect -492 -1158 -482 -1124
rect -424 -1158 -410 -1124
rect -356 -1158 -338 -1124
rect -288 -1158 -266 -1124
rect -220 -1158 -194 -1124
rect -152 -1158 -122 -1124
rect -84 -1158 -50 -1124
rect -16 -1158 18 -1124
rect 56 -1158 86 -1124
rect 128 -1158 154 -1124
rect 200 -1158 222 -1124
rect 272 -1158 290 -1124
rect 344 -1158 358 -1124
rect 416 -1158 426 -1124
rect 488 -1158 494 -1124
rect 560 -1158 562 -1124
rect 596 -1158 598 -1124
rect 664 -1158 670 -1124
rect 732 -1158 742 -1124
rect 800 -1158 814 -1124
rect 868 -1158 886 -1124
rect 936 -1158 958 -1124
rect 1004 -1158 1030 -1124
rect 1064 -1158 1102 -1124
rect 1136 -1158 1290 -1124
rect -1140 -1182 1290 -1158
<< viali >>
rect -986 7124 -952 7158
rect -914 7124 -880 7158
rect -842 7124 -832 7158
rect -832 7124 -808 7158
rect -770 7124 -764 7158
rect -764 7124 -736 7158
rect -698 7124 -696 7158
rect -696 7124 -664 7158
rect -626 7124 -594 7158
rect -594 7124 -592 7158
rect -554 7124 -526 7158
rect -526 7124 -520 7158
rect -482 7124 -458 7158
rect -458 7124 -448 7158
rect -410 7124 -390 7158
rect -390 7124 -376 7158
rect -338 7124 -322 7158
rect -322 7124 -304 7158
rect -266 7124 -254 7158
rect -254 7124 -232 7158
rect -194 7124 -186 7158
rect -186 7124 -160 7158
rect -122 7124 -118 7158
rect -118 7124 -88 7158
rect -50 7124 -16 7158
rect 22 7124 52 7158
rect 52 7124 56 7158
rect 94 7124 120 7158
rect 120 7124 128 7158
rect 166 7124 188 7158
rect 188 7124 200 7158
rect 238 7124 256 7158
rect 256 7124 272 7158
rect 310 7124 324 7158
rect 324 7124 344 7158
rect 382 7124 392 7158
rect 392 7124 416 7158
rect 454 7124 460 7158
rect 460 7124 488 7158
rect 526 7124 528 7158
rect 528 7124 560 7158
rect 598 7124 630 7158
rect 630 7124 632 7158
rect 670 7124 698 7158
rect 698 7124 704 7158
rect 742 7124 766 7158
rect 766 7124 776 7158
rect 814 7124 834 7158
rect 834 7124 848 7158
rect 886 7124 902 7158
rect 902 7124 920 7158
rect 958 7124 970 7158
rect 970 7124 992 7158
rect 1030 7124 1064 7158
rect 1102 7124 1136 7158
rect -1116 7051 -1082 7085
rect -1116 6995 -1082 7013
rect -1116 6979 -1082 6995
rect -1116 6927 -1082 6941
rect -1116 6907 -1082 6927
rect -1116 6859 -1082 6869
rect -1116 6835 -1082 6859
rect -1116 6791 -1082 6797
rect -1116 6763 -1082 6791
rect -1116 6723 -1082 6725
rect -1116 6691 -1082 6723
rect -1116 6621 -1082 6653
rect -1116 6619 -1082 6621
rect -1116 6553 -1082 6581
rect -1116 6547 -1082 6553
rect -1116 6485 -1082 6509
rect -1116 6475 -1082 6485
rect -1116 6417 -1082 6437
rect -1116 6403 -1082 6417
rect -1116 6349 -1082 6365
rect -1116 6331 -1082 6349
rect -1116 6281 -1082 6293
rect -1116 6259 -1082 6281
rect -1116 6213 -1082 6221
rect -1116 6187 -1082 6213
rect -1116 6145 -1082 6149
rect -1116 6115 -1082 6145
rect -1116 6043 -1082 6077
rect -1116 5975 -1082 6005
rect -1116 5971 -1082 5975
rect 1232 7051 1266 7085
rect 1232 6995 1266 7013
rect 1232 6979 1266 6995
rect 1232 6927 1266 6941
rect 1232 6907 1266 6927
rect 1232 6859 1266 6869
rect 1232 6835 1266 6859
rect 1232 6791 1266 6797
rect 1232 6763 1266 6791
rect 1232 6723 1266 6725
rect 1232 6691 1266 6723
rect 1232 6621 1266 6653
rect 1232 6619 1266 6621
rect 1232 6553 1266 6581
rect 1232 6547 1266 6553
rect 1232 6485 1266 6509
rect 1232 6475 1266 6485
rect 1232 6417 1266 6437
rect 1232 6403 1266 6417
rect 1232 6349 1266 6365
rect 1232 6331 1266 6349
rect 1232 6281 1266 6293
rect 1232 6259 1266 6281
rect 1232 6213 1266 6221
rect 1232 6187 1266 6213
rect 1232 6145 1266 6149
rect 1232 6115 1266 6145
rect 1232 6043 1266 6077
rect -1116 5907 -1082 5933
rect -1116 5899 -1082 5907
rect -1116 5839 -1082 5861
rect -1116 5827 -1082 5839
rect -1116 5771 -1082 5789
rect -1116 5755 -1082 5771
rect -1116 5703 -1082 5717
rect -1116 5683 -1082 5703
rect -1116 5635 -1082 5645
rect -1116 5611 -1082 5635
rect -1116 5567 -1082 5573
rect -1116 5539 -1082 5567
rect -1116 5499 -1082 5501
rect -1116 5467 -1082 5499
rect -1116 5397 -1082 5429
rect -1116 5395 -1082 5397
rect -1116 5329 -1082 5357
rect -1116 5323 -1082 5329
rect -1116 5261 -1082 5285
rect -1116 5251 -1082 5261
rect -1116 5193 -1082 5213
rect -1116 5179 -1082 5193
rect -1116 5125 -1082 5141
rect -1116 5107 -1082 5125
rect -1116 5057 -1082 5069
rect -1116 5035 -1082 5057
rect -1116 4989 -1082 4997
rect -1116 4963 -1082 4989
rect -1116 4921 -1082 4925
rect -1116 4891 -1082 4921
rect -1116 4819 -1082 4853
rect -1116 4751 -1082 4781
rect -1116 4747 -1082 4751
rect -1116 4683 -1082 4709
rect -1116 4675 -1082 4683
rect -1116 4615 -1082 4637
rect -1116 4603 -1082 4615
rect -1116 4547 -1082 4565
rect -1116 4531 -1082 4547
rect -1116 4479 -1082 4493
rect -1116 4459 -1082 4479
rect -1116 4411 -1082 4421
rect -1116 4387 -1082 4411
rect -1116 4343 -1082 4349
rect -1116 4315 -1082 4343
rect -1116 4275 -1082 4277
rect -1116 4243 -1082 4275
rect -1116 4173 -1082 4205
rect -1116 4171 -1082 4173
rect -1116 4105 -1082 4133
rect -1116 4099 -1082 4105
rect -1116 4037 -1082 4061
rect -1116 4027 -1082 4037
rect -1116 3969 -1082 3989
rect -1116 3955 -1082 3969
rect -1116 3901 -1082 3917
rect -1116 3883 -1082 3901
rect -1116 3833 -1082 3845
rect -1116 3811 -1082 3833
rect -1116 3765 -1082 3773
rect -1116 3739 -1082 3765
rect -1116 3697 -1082 3701
rect -1116 3667 -1082 3697
rect -1116 3595 -1082 3629
rect -1116 3527 -1082 3557
rect -1116 3523 -1082 3527
rect -1116 3459 -1082 3485
rect -1116 3451 -1082 3459
rect -1116 3391 -1082 3413
rect -1116 3379 -1082 3391
rect -1116 3323 -1082 3341
rect -1116 3307 -1082 3323
rect -1116 3255 -1082 3269
rect -1116 3235 -1082 3255
rect -1116 3187 -1082 3197
rect -1116 3163 -1082 3187
rect -1116 3119 -1082 3125
rect -1116 3091 -1082 3119
rect -1116 3051 -1082 3053
rect -1116 3019 -1082 3051
rect -1116 2949 -1082 2981
rect -1116 2947 -1082 2949
rect -1116 2881 -1082 2909
rect -1116 2875 -1082 2881
rect -1116 2813 -1082 2837
rect -1116 2803 -1082 2813
rect -1116 2745 -1082 2765
rect -1116 2731 -1082 2745
rect -1116 2677 -1082 2693
rect -1116 2659 -1082 2677
rect -1116 2609 -1082 2621
rect -1116 2587 -1082 2609
rect -1116 2541 -1082 2549
rect -1116 2515 -1082 2541
rect -1116 2473 -1082 2477
rect -1116 2443 -1082 2473
rect -1116 2371 -1082 2405
rect -1116 2303 -1082 2333
rect -1116 2299 -1082 2303
rect -1116 2235 -1082 2261
rect -1116 2227 -1082 2235
rect -1116 2167 -1082 2189
rect -1116 2155 -1082 2167
rect -1116 2099 -1082 2117
rect -1116 2083 -1082 2099
rect -1116 2031 -1082 2045
rect -1116 2011 -1082 2031
rect -1116 1963 -1082 1973
rect -1116 1939 -1082 1963
rect -1116 1895 -1082 1901
rect -1116 1867 -1082 1895
rect -1116 1827 -1082 1829
rect -1116 1795 -1082 1827
rect -1116 1725 -1082 1757
rect -1116 1723 -1082 1725
rect -1116 1657 -1082 1685
rect -1116 1651 -1082 1657
rect -1116 1589 -1082 1613
rect -1116 1579 -1082 1589
rect -1116 1521 -1082 1541
rect -1116 1507 -1082 1521
rect -1116 1453 -1082 1469
rect -1116 1435 -1082 1453
rect -1116 1385 -1082 1397
rect -1116 1363 -1082 1385
rect -1116 1317 -1082 1325
rect -1116 1291 -1082 1317
rect -1116 1249 -1082 1253
rect -1116 1219 -1082 1249
rect -1116 1147 -1082 1181
rect -1116 1079 -1082 1109
rect -1116 1075 -1082 1079
rect -1116 1011 -1082 1037
rect -1116 1003 -1082 1011
rect -1116 943 -1082 965
rect -1116 931 -1082 943
rect -1116 875 -1082 893
rect -1116 859 -1082 875
rect -1116 807 -1082 821
rect -1116 787 -1082 807
rect -1116 739 -1082 749
rect -1116 715 -1082 739
rect -1116 671 -1082 677
rect -1116 643 -1082 671
rect -1116 603 -1082 605
rect -1116 571 -1082 603
rect -1116 501 -1082 533
rect -1116 499 -1082 501
rect -1116 433 -1082 461
rect -1116 427 -1082 433
rect -1116 365 -1082 389
rect -1116 355 -1082 365
rect -1116 297 -1082 317
rect -1116 283 -1082 297
rect -1116 229 -1082 245
rect -1116 211 -1082 229
rect -1116 161 -1082 173
rect -1116 139 -1082 161
rect -1116 93 -1082 101
rect -1116 67 -1082 93
rect -1116 25 -1082 29
rect -1116 -5 -1082 25
rect -946 5941 -912 5969
rect -946 5935 -912 5941
rect -946 5873 -912 5897
rect -946 5863 -912 5873
rect -946 5805 -912 5825
rect -946 5791 -912 5805
rect -946 5737 -912 5753
rect -946 5719 -912 5737
rect -946 5669 -912 5681
rect -946 5647 -912 5669
rect -946 5601 -912 5609
rect -946 5575 -912 5601
rect -946 5533 -912 5537
rect -946 5503 -912 5533
rect -946 5431 -912 5465
rect -946 5363 -912 5393
rect -946 5359 -912 5363
rect -946 5295 -912 5321
rect -946 5287 -912 5295
rect -946 5227 -912 5249
rect -946 5215 -912 5227
rect -946 5159 -912 5177
rect -946 5143 -912 5159
rect -946 5091 -912 5105
rect -946 5071 -912 5091
rect -946 5023 -912 5033
rect -946 4999 -912 5023
rect -946 4955 -912 4961
rect -946 4927 -912 4955
rect -946 4887 -912 4889
rect -946 4855 -912 4887
rect -946 4785 -912 4817
rect -946 4783 -912 4785
rect -946 4717 -912 4745
rect -946 4711 -912 4717
rect -946 4649 -912 4673
rect -946 4639 -912 4649
rect -946 4581 -912 4601
rect -946 4567 -912 4581
rect -946 4513 -912 4529
rect -946 4495 -912 4513
rect -946 4445 -912 4457
rect -946 4423 -912 4445
rect -946 4377 -912 4385
rect -946 4351 -912 4377
rect -946 4309 -912 4313
rect -946 4279 -912 4309
rect -946 4207 -912 4241
rect -946 4139 -912 4169
rect -946 4135 -912 4139
rect -946 4071 -912 4097
rect -946 4063 -912 4071
rect -946 4003 -912 4025
rect -946 3991 -912 4003
rect -946 3935 -912 3953
rect -946 3919 -912 3935
rect -946 3867 -912 3881
rect -946 3847 -912 3867
rect -946 3799 -912 3809
rect -946 3775 -912 3799
rect -946 3731 -912 3737
rect -946 3703 -912 3731
rect -946 3663 -912 3665
rect -946 3631 -912 3663
rect -946 3561 -912 3593
rect -946 3559 -912 3561
rect -946 3493 -912 3521
rect -946 3487 -912 3493
rect -946 3425 -912 3449
rect -946 3415 -912 3425
rect -946 3357 -912 3377
rect -946 3343 -912 3357
rect -946 3289 -912 3305
rect -946 3271 -912 3289
rect -946 3221 -912 3233
rect -946 3199 -912 3221
rect -946 3153 -912 3161
rect -946 3127 -912 3153
rect -946 3085 -912 3089
rect -946 3055 -912 3085
rect -946 2983 -912 3017
rect -946 2915 -912 2945
rect -946 2911 -912 2915
rect -946 2847 -912 2873
rect -946 2839 -912 2847
rect -946 2779 -912 2801
rect -946 2767 -912 2779
rect -946 2711 -912 2729
rect -946 2695 -912 2711
rect -946 2643 -912 2657
rect -946 2623 -912 2643
rect -946 2575 -912 2585
rect -946 2551 -912 2575
rect -946 2507 -912 2513
rect -946 2479 -912 2507
rect -946 2439 -912 2441
rect -946 2407 -912 2439
rect -946 2337 -912 2369
rect -946 2335 -912 2337
rect -946 2269 -912 2297
rect -946 2263 -912 2269
rect -946 2201 -912 2225
rect -946 2191 -912 2201
rect -946 2133 -912 2153
rect -946 2119 -912 2133
rect -946 2065 -912 2081
rect -946 2047 -912 2065
rect -946 1997 -912 2009
rect -946 1975 -912 1997
rect -946 1929 -912 1937
rect -946 1903 -912 1929
rect -946 1861 -912 1865
rect -946 1831 -912 1861
rect -946 1759 -912 1793
rect -946 1691 -912 1721
rect -946 1687 -912 1691
rect -946 1623 -912 1649
rect -946 1615 -912 1623
rect -946 1555 -912 1577
rect -946 1543 -912 1555
rect -946 1487 -912 1505
rect -946 1471 -912 1487
rect -946 1419 -912 1433
rect -946 1399 -912 1419
rect -946 1351 -912 1361
rect -946 1327 -912 1351
rect -946 1283 -912 1289
rect -946 1255 -912 1283
rect -946 1215 -912 1217
rect -946 1183 -912 1215
rect -946 1113 -912 1145
rect -946 1111 -912 1113
rect -946 1045 -912 1073
rect -946 1039 -912 1045
rect -946 977 -912 1001
rect -946 967 -912 977
rect -946 909 -912 929
rect -946 895 -912 909
rect -946 841 -912 857
rect -946 823 -912 841
rect -946 773 -912 785
rect -946 751 -912 773
rect -946 705 -912 713
rect -946 679 -912 705
rect -946 637 -912 641
rect -946 607 -912 637
rect -946 535 -912 569
rect -946 467 -912 497
rect -946 463 -912 467
rect -946 399 -912 425
rect -946 391 -912 399
rect -946 331 -912 353
rect -946 319 -912 331
rect -946 263 -912 281
rect -946 247 -912 263
rect -946 195 -912 209
rect -946 175 -912 195
rect -946 127 -912 137
rect -946 103 -912 127
rect -946 59 -912 65
rect -946 31 -912 59
rect 22 67 24 5933
rect 24 67 126 5933
rect 126 67 128 5933
rect 1062 5941 1096 5969
rect 1062 5935 1096 5941
rect 1062 5873 1096 5897
rect 1062 5863 1096 5873
rect 1062 5805 1096 5825
rect 1062 5791 1096 5805
rect 1062 5737 1096 5753
rect 1062 5719 1096 5737
rect 1062 5669 1096 5681
rect 1062 5647 1096 5669
rect 1062 5601 1096 5609
rect 1062 5575 1096 5601
rect 1062 5533 1096 5537
rect 1062 5503 1096 5533
rect 1062 5431 1096 5465
rect 1062 5363 1096 5393
rect 1062 5359 1096 5363
rect 1062 5295 1096 5321
rect 1062 5287 1096 5295
rect 1062 5227 1096 5249
rect 1062 5215 1096 5227
rect 1062 5159 1096 5177
rect 1062 5143 1096 5159
rect 1062 5091 1096 5105
rect 1062 5071 1096 5091
rect 1062 5023 1096 5033
rect 1062 4999 1096 5023
rect 1062 4955 1096 4961
rect 1062 4927 1096 4955
rect 1062 4887 1096 4889
rect 1062 4855 1096 4887
rect 1062 4785 1096 4817
rect 1062 4783 1096 4785
rect 1062 4717 1096 4745
rect 1062 4711 1096 4717
rect 1062 4649 1096 4673
rect 1062 4639 1096 4649
rect 1062 4581 1096 4601
rect 1062 4567 1096 4581
rect 1062 4513 1096 4529
rect 1062 4495 1096 4513
rect 1062 4445 1096 4457
rect 1062 4423 1096 4445
rect 1062 4377 1096 4385
rect 1062 4351 1096 4377
rect 1062 4309 1096 4313
rect 1062 4279 1096 4309
rect 1062 4207 1096 4241
rect 1062 4139 1096 4169
rect 1062 4135 1096 4139
rect 1062 4071 1096 4097
rect 1062 4063 1096 4071
rect 1062 4003 1096 4025
rect 1062 3991 1096 4003
rect 1062 3935 1096 3953
rect 1062 3919 1096 3935
rect 1062 3867 1096 3881
rect 1062 3847 1096 3867
rect 1062 3799 1096 3809
rect 1062 3775 1096 3799
rect 1062 3731 1096 3737
rect 1062 3703 1096 3731
rect 1062 3663 1096 3665
rect 1062 3631 1096 3663
rect 1062 3561 1096 3593
rect 1062 3559 1096 3561
rect 1062 3493 1096 3521
rect 1062 3487 1096 3493
rect 1062 3425 1096 3449
rect 1062 3415 1096 3425
rect 1062 3357 1096 3377
rect 1062 3343 1096 3357
rect 1062 3289 1096 3305
rect 1062 3271 1096 3289
rect 1062 3221 1096 3233
rect 1062 3199 1096 3221
rect 1062 3153 1096 3161
rect 1062 3127 1096 3153
rect 1062 3085 1096 3089
rect 1062 3055 1096 3085
rect 1062 2983 1096 3017
rect 1062 2915 1096 2945
rect 1062 2911 1096 2915
rect 1062 2847 1096 2873
rect 1062 2839 1096 2847
rect 1062 2779 1096 2801
rect 1062 2767 1096 2779
rect 1062 2711 1096 2729
rect 1062 2695 1096 2711
rect 1062 2643 1096 2657
rect 1062 2623 1096 2643
rect 1062 2575 1096 2585
rect 1062 2551 1096 2575
rect 1062 2507 1096 2513
rect 1062 2479 1096 2507
rect 1062 2439 1096 2441
rect 1062 2407 1096 2439
rect 1062 2337 1096 2369
rect 1062 2335 1096 2337
rect 1062 2269 1096 2297
rect 1062 2263 1096 2269
rect 1062 2201 1096 2225
rect 1062 2191 1096 2201
rect 1062 2133 1096 2153
rect 1062 2119 1096 2133
rect 1062 2065 1096 2081
rect 1062 2047 1096 2065
rect 1062 1997 1096 2009
rect 1062 1975 1096 1997
rect 1062 1929 1096 1937
rect 1062 1903 1096 1929
rect 1062 1861 1096 1865
rect 1062 1831 1096 1861
rect 1062 1759 1096 1793
rect 1062 1691 1096 1721
rect 1062 1687 1096 1691
rect 1062 1623 1096 1649
rect 1062 1615 1096 1623
rect 1062 1555 1096 1577
rect 1062 1543 1096 1555
rect 1062 1487 1096 1505
rect 1062 1471 1096 1487
rect 1062 1419 1096 1433
rect 1062 1399 1096 1419
rect 1062 1351 1096 1361
rect 1062 1327 1096 1351
rect 1062 1283 1096 1289
rect 1062 1255 1096 1283
rect 1062 1215 1096 1217
rect 1062 1183 1096 1215
rect 1062 1113 1096 1145
rect 1062 1111 1096 1113
rect 1062 1045 1096 1073
rect 1062 1039 1096 1045
rect 1062 977 1096 1001
rect 1062 967 1096 977
rect 1062 909 1096 929
rect 1062 895 1096 909
rect 1062 841 1096 857
rect 1062 823 1096 841
rect 1062 773 1096 785
rect 1062 751 1096 773
rect 1062 705 1096 713
rect 1062 679 1096 705
rect 1062 637 1096 641
rect 1062 607 1096 637
rect 1062 535 1096 569
rect 1062 467 1096 497
rect 1062 463 1096 467
rect 1062 399 1096 425
rect 1062 391 1096 399
rect 1062 331 1096 353
rect 1062 319 1096 331
rect 1062 263 1096 281
rect 1062 247 1096 263
rect 1062 195 1096 209
rect 1062 175 1096 195
rect 1062 127 1096 137
rect 1062 103 1096 127
rect 1062 59 1096 65
rect 1062 31 1096 59
rect 1232 5975 1266 6005
rect 1232 5971 1266 5975
rect 1232 5907 1266 5933
rect 1232 5899 1266 5907
rect 1232 5839 1266 5861
rect 1232 5827 1266 5839
rect 1232 5771 1266 5789
rect 1232 5755 1266 5771
rect 1232 5703 1266 5717
rect 1232 5683 1266 5703
rect 1232 5635 1266 5645
rect 1232 5611 1266 5635
rect 1232 5567 1266 5573
rect 1232 5539 1266 5567
rect 1232 5499 1266 5501
rect 1232 5467 1266 5499
rect 1232 5397 1266 5429
rect 1232 5395 1266 5397
rect 1232 5329 1266 5357
rect 1232 5323 1266 5329
rect 1232 5261 1266 5285
rect 1232 5251 1266 5261
rect 1232 5193 1266 5213
rect 1232 5179 1266 5193
rect 1232 5125 1266 5141
rect 1232 5107 1266 5125
rect 1232 5057 1266 5069
rect 1232 5035 1266 5057
rect 1232 4989 1266 4997
rect 1232 4963 1266 4989
rect 1232 4921 1266 4925
rect 1232 4891 1266 4921
rect 1232 4819 1266 4853
rect 1232 4751 1266 4781
rect 1232 4747 1266 4751
rect 1232 4683 1266 4709
rect 1232 4675 1266 4683
rect 1232 4615 1266 4637
rect 1232 4603 1266 4615
rect 1232 4547 1266 4565
rect 1232 4531 1266 4547
rect 1232 4479 1266 4493
rect 1232 4459 1266 4479
rect 1232 4411 1266 4421
rect 1232 4387 1266 4411
rect 1232 4343 1266 4349
rect 1232 4315 1266 4343
rect 1232 4275 1266 4277
rect 1232 4243 1266 4275
rect 1232 4173 1266 4205
rect 1232 4171 1266 4173
rect 1232 4105 1266 4133
rect 1232 4099 1266 4105
rect 1232 4037 1266 4061
rect 1232 4027 1266 4037
rect 1232 3969 1266 3989
rect 1232 3955 1266 3969
rect 1232 3901 1266 3917
rect 1232 3883 1266 3901
rect 1232 3833 1266 3845
rect 1232 3811 1266 3833
rect 1232 3765 1266 3773
rect 1232 3739 1266 3765
rect 1232 3697 1266 3701
rect 1232 3667 1266 3697
rect 1232 3595 1266 3629
rect 1232 3527 1266 3557
rect 1232 3523 1266 3527
rect 1232 3459 1266 3485
rect 1232 3451 1266 3459
rect 1232 3391 1266 3413
rect 1232 3379 1266 3391
rect 1232 3323 1266 3341
rect 1232 3307 1266 3323
rect 1232 3255 1266 3269
rect 1232 3235 1266 3255
rect 1232 3187 1266 3197
rect 1232 3163 1266 3187
rect 1232 3119 1266 3125
rect 1232 3091 1266 3119
rect 1232 3051 1266 3053
rect 1232 3019 1266 3051
rect 1232 2949 1266 2981
rect 1232 2947 1266 2949
rect 1232 2881 1266 2909
rect 1232 2875 1266 2881
rect 1232 2813 1266 2837
rect 1232 2803 1266 2813
rect 1232 2745 1266 2765
rect 1232 2731 1266 2745
rect 1232 2677 1266 2693
rect 1232 2659 1266 2677
rect 1232 2609 1266 2621
rect 1232 2587 1266 2609
rect 1232 2541 1266 2549
rect 1232 2515 1266 2541
rect 1232 2473 1266 2477
rect 1232 2443 1266 2473
rect 1232 2371 1266 2405
rect 1232 2303 1266 2333
rect 1232 2299 1266 2303
rect 1232 2235 1266 2261
rect 1232 2227 1266 2235
rect 1232 2167 1266 2189
rect 1232 2155 1266 2167
rect 1232 2099 1266 2117
rect 1232 2083 1266 2099
rect 1232 2031 1266 2045
rect 1232 2011 1266 2031
rect 1232 1963 1266 1973
rect 1232 1939 1266 1963
rect 1232 1895 1266 1901
rect 1232 1867 1266 1895
rect 1232 1827 1266 1829
rect 1232 1795 1266 1827
rect 1232 1725 1266 1757
rect 1232 1723 1266 1725
rect 1232 1657 1266 1685
rect 1232 1651 1266 1657
rect 1232 1589 1266 1613
rect 1232 1579 1266 1589
rect 1232 1521 1266 1541
rect 1232 1507 1266 1521
rect 1232 1453 1266 1469
rect 1232 1435 1266 1453
rect 1232 1385 1266 1397
rect 1232 1363 1266 1385
rect 1232 1317 1266 1325
rect 1232 1291 1266 1317
rect 1232 1249 1266 1253
rect 1232 1219 1266 1249
rect 1232 1147 1266 1181
rect 1232 1079 1266 1109
rect 1232 1075 1266 1079
rect 1232 1011 1266 1037
rect 1232 1003 1266 1011
rect 1232 943 1266 965
rect 1232 931 1266 943
rect 1232 875 1266 893
rect 1232 859 1266 875
rect 1232 807 1266 821
rect 1232 787 1266 807
rect 1232 739 1266 749
rect 1232 715 1266 739
rect 1232 671 1266 677
rect 1232 643 1266 671
rect 1232 603 1266 605
rect 1232 571 1266 603
rect 1232 501 1266 533
rect 1232 499 1266 501
rect 1232 433 1266 461
rect 1232 427 1266 433
rect 1232 365 1266 389
rect 1232 355 1266 365
rect 1232 297 1266 317
rect 1232 283 1266 297
rect 1232 229 1266 245
rect 1232 211 1266 229
rect 1232 161 1266 173
rect 1232 139 1266 161
rect 1232 93 1266 101
rect 1232 67 1266 93
rect -1116 -77 -1082 -43
rect -1116 -145 -1082 -115
rect -1116 -149 -1082 -145
rect -1116 -213 -1082 -187
rect -1116 -221 -1082 -213
rect -1116 -281 -1082 -259
rect -1116 -293 -1082 -281
rect -1116 -349 -1082 -331
rect -1116 -365 -1082 -349
rect -1116 -417 -1082 -403
rect -1116 -437 -1082 -417
rect -1116 -485 -1082 -475
rect -1116 -509 -1082 -485
rect -1116 -553 -1082 -547
rect -1116 -581 -1082 -553
rect -1116 -621 -1082 -619
rect -1116 -653 -1082 -621
rect 1232 25 1266 29
rect 1232 -5 1266 25
rect 1232 -77 1266 -43
rect 1232 -145 1266 -115
rect 1232 -149 1266 -145
rect 1232 -213 1266 -187
rect 1232 -221 1266 -213
rect 1232 -281 1266 -259
rect 1232 -293 1266 -281
rect 1232 -349 1266 -331
rect 1232 -365 1266 -349
rect 1232 -417 1266 -403
rect 1232 -437 1266 -417
rect 1232 -485 1266 -475
rect 1232 -509 1266 -485
rect 1232 -553 1266 -547
rect 1232 -581 1266 -553
rect -1116 -723 -1082 -691
rect -1116 -725 -1082 -723
rect -1116 -791 -1082 -763
rect -1116 -797 -1082 -791
rect -1116 -859 -1082 -835
rect -1116 -869 -1082 -859
rect -280 -693 -246 -659
rect -206 -693 -172 -659
rect -132 -693 -98 -659
rect -58 -693 -24 -659
rect 16 -693 50 -659
rect 90 -693 124 -659
rect 164 -693 198 -659
rect 238 -693 272 -659
rect 312 -693 346 -659
rect 386 -693 420 -659
rect -280 -767 -246 -733
rect -206 -767 -172 -733
rect -132 -767 -98 -733
rect -58 -767 -24 -733
rect 16 -767 50 -733
rect 90 -767 124 -733
rect 164 -767 198 -733
rect 238 -767 272 -733
rect 312 -767 346 -733
rect 386 -767 420 -733
rect -280 -841 -246 -807
rect -206 -841 -172 -807
rect -132 -841 -98 -807
rect -58 -841 -24 -807
rect 16 -841 50 -807
rect 90 -841 124 -807
rect 164 -841 198 -807
rect 238 -841 272 -807
rect 312 -841 346 -807
rect 386 -841 420 -807
rect 1232 -621 1266 -619
rect 1232 -653 1266 -621
rect 1232 -723 1266 -691
rect 1232 -725 1266 -723
rect 1232 -791 1266 -763
rect 1232 -797 1266 -791
rect -1116 -927 -1082 -907
rect -1116 -941 -1082 -927
rect -1116 -995 -1082 -979
rect -1116 -1013 -1082 -995
rect -1116 -1085 -1082 -1051
rect 1232 -859 1266 -835
rect 1232 -869 1266 -859
rect 1232 -927 1266 -907
rect 1232 -941 1266 -927
rect 1232 -995 1266 -979
rect 1232 -1013 1266 -995
rect 1232 -1085 1266 -1051
rect -986 -1158 -952 -1124
rect -914 -1158 -880 -1124
rect -842 -1158 -832 -1124
rect -832 -1158 -808 -1124
rect -770 -1158 -764 -1124
rect -764 -1158 -736 -1124
rect -698 -1158 -696 -1124
rect -696 -1158 -664 -1124
rect -626 -1158 -594 -1124
rect -594 -1158 -592 -1124
rect -554 -1158 -526 -1124
rect -526 -1158 -520 -1124
rect -482 -1158 -458 -1124
rect -458 -1158 -448 -1124
rect -410 -1158 -390 -1124
rect -390 -1158 -376 -1124
rect -338 -1158 -322 -1124
rect -322 -1158 -304 -1124
rect -266 -1158 -254 -1124
rect -254 -1158 -232 -1124
rect -194 -1158 -186 -1124
rect -186 -1158 -160 -1124
rect -122 -1158 -118 -1124
rect -118 -1158 -88 -1124
rect -50 -1158 -16 -1124
rect 22 -1158 52 -1124
rect 52 -1158 56 -1124
rect 94 -1158 120 -1124
rect 120 -1158 128 -1124
rect 166 -1158 188 -1124
rect 188 -1158 200 -1124
rect 238 -1158 256 -1124
rect 256 -1158 272 -1124
rect 310 -1158 324 -1124
rect 324 -1158 344 -1124
rect 382 -1158 392 -1124
rect 392 -1158 416 -1124
rect 454 -1158 460 -1124
rect 460 -1158 488 -1124
rect 526 -1158 528 -1124
rect 528 -1158 560 -1124
rect 598 -1158 630 -1124
rect 630 -1158 632 -1124
rect 670 -1158 698 -1124
rect 698 -1158 704 -1124
rect 742 -1158 766 -1124
rect 766 -1158 776 -1124
rect 814 -1158 834 -1124
rect 834 -1158 848 -1124
rect 886 -1158 902 -1124
rect 902 -1158 920 -1124
rect 958 -1158 970 -1124
rect 970 -1158 992 -1124
rect 1030 -1158 1064 -1124
rect 1102 -1158 1136 -1124
<< metal1 >>
rect -1140 7158 1290 7182
rect -1140 7124 -986 7158
rect -952 7124 -914 7158
rect -880 7124 -842 7158
rect -808 7124 -770 7158
rect -736 7124 -698 7158
rect -664 7124 -626 7158
rect -592 7124 -554 7158
rect -520 7124 -482 7158
rect -448 7124 -410 7158
rect -376 7124 -338 7158
rect -304 7124 -266 7158
rect -232 7124 -194 7158
rect -160 7124 -122 7158
rect -88 7124 -50 7158
rect -16 7124 22 7158
rect 56 7124 94 7158
rect 128 7124 166 7158
rect 200 7124 238 7158
rect 272 7124 310 7158
rect 344 7124 382 7158
rect 416 7124 454 7158
rect 488 7124 526 7158
rect 560 7124 598 7158
rect 632 7124 670 7158
rect 704 7124 742 7158
rect 776 7124 814 7158
rect 848 7124 886 7158
rect 920 7124 958 7158
rect 992 7124 1030 7158
rect 1064 7124 1102 7158
rect 1136 7124 1290 7158
rect -1140 7100 1290 7124
rect -1140 7085 -1058 7100
rect -1140 7051 -1116 7085
rect -1082 7051 -1058 7085
rect -1140 7013 -1058 7051
rect -1140 6979 -1116 7013
rect -1082 6979 -1058 7013
rect -1140 6941 -1058 6979
rect -1140 6907 -1116 6941
rect -1082 6907 -1058 6941
rect -1140 6869 -1058 6907
rect -1140 6835 -1116 6869
rect -1082 6835 -1058 6869
rect -1140 6797 -1058 6835
rect -1140 6763 -1116 6797
rect -1082 6763 -1058 6797
rect -1140 6725 -1058 6763
rect -1140 6691 -1116 6725
rect -1082 6691 -1058 6725
rect -1140 6653 -1058 6691
rect -1140 6619 -1116 6653
rect -1082 6619 -1058 6653
rect -1140 6581 -1058 6619
rect -1140 6547 -1116 6581
rect -1082 6547 -1058 6581
rect -1140 6509 -1058 6547
rect -1140 6475 -1116 6509
rect -1082 6475 -1058 6509
rect -1140 6437 -1058 6475
rect -1140 6403 -1116 6437
rect -1082 6403 -1058 6437
rect -1140 6365 -1058 6403
rect -1140 6331 -1116 6365
rect -1082 6331 -1058 6365
rect -1140 6293 -1058 6331
rect -1140 6259 -1116 6293
rect -1082 6259 -1058 6293
rect -1140 6221 -1058 6259
rect -1140 6187 -1116 6221
rect -1082 6187 -1058 6221
rect -1140 6149 -1058 6187
rect -1140 6115 -1116 6149
rect -1082 6115 -1058 6149
rect -1140 6077 -1058 6115
rect -1140 6043 -1116 6077
rect -1082 6043 -1058 6077
rect -1140 6005 -1058 6043
rect -1140 5971 -1116 6005
rect -1082 5971 -1058 6005
rect 1208 7085 1290 7100
rect 1208 7051 1232 7085
rect 1266 7051 1290 7085
rect 1208 7013 1290 7051
rect 1208 6979 1232 7013
rect 1266 6979 1290 7013
rect 1208 6941 1290 6979
rect 1208 6907 1232 6941
rect 1266 6907 1290 6941
rect 1208 6869 1290 6907
rect 1208 6835 1232 6869
rect 1266 6835 1290 6869
rect 1208 6797 1290 6835
rect 1208 6763 1232 6797
rect 1266 6763 1290 6797
rect 1208 6725 1290 6763
rect 1208 6691 1232 6725
rect 1266 6691 1290 6725
rect 1208 6653 1290 6691
rect 1208 6619 1232 6653
rect 1266 6619 1290 6653
rect 1208 6581 1290 6619
rect 1208 6547 1232 6581
rect 1266 6547 1290 6581
rect 1208 6509 1290 6547
rect 1208 6475 1232 6509
rect 1266 6475 1290 6509
rect 1208 6437 1290 6475
rect 1208 6403 1232 6437
rect 1266 6403 1290 6437
rect 1208 6365 1290 6403
rect 1208 6331 1232 6365
rect 1266 6331 1290 6365
rect 1208 6293 1290 6331
rect 1208 6259 1232 6293
rect 1266 6259 1290 6293
rect 1208 6221 1290 6259
rect 1208 6187 1232 6221
rect 1266 6187 1290 6221
rect 1208 6149 1290 6187
rect 1208 6115 1232 6149
rect 1266 6115 1290 6149
rect 1208 6077 1290 6115
rect 1208 6043 1232 6077
rect 1266 6043 1290 6077
rect 1208 6005 1290 6043
rect -1140 5933 -1058 5971
rect -1140 5899 -1116 5933
rect -1082 5899 -1058 5933
rect -1140 5861 -1058 5899
rect -1140 5827 -1116 5861
rect -1082 5827 -1058 5861
rect -1140 5789 -1058 5827
rect -1140 5755 -1116 5789
rect -1082 5755 -1058 5789
rect -1140 5717 -1058 5755
rect -1140 5683 -1116 5717
rect -1082 5683 -1058 5717
rect -1140 5645 -1058 5683
rect -1140 5611 -1116 5645
rect -1082 5611 -1058 5645
rect -1140 5573 -1058 5611
rect -1140 5539 -1116 5573
rect -1082 5539 -1058 5573
rect -1140 5501 -1058 5539
rect -1140 5467 -1116 5501
rect -1082 5467 -1058 5501
rect -1140 5429 -1058 5467
rect -1140 5395 -1116 5429
rect -1082 5395 -1058 5429
rect -1140 5357 -1058 5395
rect -1140 5323 -1116 5357
rect -1082 5323 -1058 5357
rect -1140 5285 -1058 5323
rect -1140 5251 -1116 5285
rect -1082 5251 -1058 5285
rect -1140 5213 -1058 5251
rect -1140 5179 -1116 5213
rect -1082 5179 -1058 5213
rect -1140 5141 -1058 5179
rect -1140 5107 -1116 5141
rect -1082 5107 -1058 5141
rect -1140 5069 -1058 5107
rect -1140 5035 -1116 5069
rect -1082 5035 -1058 5069
rect -1140 4997 -1058 5035
rect -1140 4963 -1116 4997
rect -1082 4963 -1058 4997
rect -1140 4925 -1058 4963
rect -1140 4891 -1116 4925
rect -1082 4891 -1058 4925
rect -1140 4853 -1058 4891
rect -1140 4819 -1116 4853
rect -1082 4819 -1058 4853
rect -1140 4781 -1058 4819
rect -1140 4747 -1116 4781
rect -1082 4747 -1058 4781
rect -1140 4709 -1058 4747
rect -1140 4675 -1116 4709
rect -1082 4675 -1058 4709
rect -1140 4637 -1058 4675
rect -1140 4603 -1116 4637
rect -1082 4603 -1058 4637
rect -1140 4565 -1058 4603
rect -1140 4531 -1116 4565
rect -1082 4531 -1058 4565
rect -1140 4493 -1058 4531
rect -1140 4459 -1116 4493
rect -1082 4459 -1058 4493
rect -1140 4421 -1058 4459
rect -1140 4387 -1116 4421
rect -1082 4387 -1058 4421
rect -1140 4349 -1058 4387
rect -1140 4315 -1116 4349
rect -1082 4315 -1058 4349
rect -1140 4277 -1058 4315
rect -1140 4243 -1116 4277
rect -1082 4243 -1058 4277
rect -1140 4205 -1058 4243
rect -1140 4171 -1116 4205
rect -1082 4171 -1058 4205
rect -1140 4133 -1058 4171
rect -1140 4099 -1116 4133
rect -1082 4099 -1058 4133
rect -1140 4061 -1058 4099
rect -1140 4027 -1116 4061
rect -1082 4027 -1058 4061
rect -1140 3989 -1058 4027
rect -1140 3955 -1116 3989
rect -1082 3955 -1058 3989
rect -1140 3917 -1058 3955
rect -1140 3883 -1116 3917
rect -1082 3883 -1058 3917
rect -1140 3845 -1058 3883
rect -1140 3811 -1116 3845
rect -1082 3811 -1058 3845
rect -1140 3773 -1058 3811
rect -1140 3739 -1116 3773
rect -1082 3739 -1058 3773
rect -1140 3701 -1058 3739
rect -1140 3667 -1116 3701
rect -1082 3667 -1058 3701
rect -1140 3629 -1058 3667
rect -1140 3595 -1116 3629
rect -1082 3595 -1058 3629
rect -1140 3557 -1058 3595
rect -1140 3523 -1116 3557
rect -1082 3523 -1058 3557
rect -1140 3485 -1058 3523
rect -1140 3451 -1116 3485
rect -1082 3451 -1058 3485
rect -1140 3413 -1058 3451
rect -1140 3379 -1116 3413
rect -1082 3379 -1058 3413
rect -1140 3341 -1058 3379
rect -1140 3307 -1116 3341
rect -1082 3307 -1058 3341
rect -1140 3269 -1058 3307
rect -1140 3235 -1116 3269
rect -1082 3235 -1058 3269
rect -1140 3197 -1058 3235
rect -1140 3163 -1116 3197
rect -1082 3163 -1058 3197
rect -1140 3125 -1058 3163
rect -1140 3091 -1116 3125
rect -1082 3091 -1058 3125
rect -1140 3053 -1058 3091
rect -1140 3019 -1116 3053
rect -1082 3019 -1058 3053
rect -1140 2981 -1058 3019
rect -1140 2947 -1116 2981
rect -1082 2947 -1058 2981
rect -1140 2909 -1058 2947
rect -1140 2875 -1116 2909
rect -1082 2875 -1058 2909
rect -1140 2837 -1058 2875
rect -1140 2803 -1116 2837
rect -1082 2803 -1058 2837
rect -1140 2765 -1058 2803
rect -1140 2731 -1116 2765
rect -1082 2731 -1058 2765
rect -1140 2693 -1058 2731
rect -1140 2659 -1116 2693
rect -1082 2659 -1058 2693
rect -1140 2621 -1058 2659
rect -1140 2587 -1116 2621
rect -1082 2587 -1058 2621
rect -1140 2549 -1058 2587
rect -1140 2515 -1116 2549
rect -1082 2515 -1058 2549
rect -1140 2477 -1058 2515
rect -1140 2443 -1116 2477
rect -1082 2443 -1058 2477
rect -1140 2405 -1058 2443
rect -1140 2371 -1116 2405
rect -1082 2371 -1058 2405
rect -1140 2333 -1058 2371
rect -1140 2299 -1116 2333
rect -1082 2299 -1058 2333
rect -1140 2261 -1058 2299
rect -1140 2227 -1116 2261
rect -1082 2227 -1058 2261
rect -1140 2189 -1058 2227
rect -1140 2155 -1116 2189
rect -1082 2155 -1058 2189
rect -1140 2117 -1058 2155
rect -1140 2083 -1116 2117
rect -1082 2083 -1058 2117
rect -1140 2045 -1058 2083
rect -1140 2011 -1116 2045
rect -1082 2011 -1058 2045
rect -1140 1973 -1058 2011
rect -1140 1939 -1116 1973
rect -1082 1939 -1058 1973
rect -1140 1901 -1058 1939
rect -1140 1867 -1116 1901
rect -1082 1867 -1058 1901
rect -1140 1829 -1058 1867
rect -1140 1795 -1116 1829
rect -1082 1795 -1058 1829
rect -1140 1757 -1058 1795
rect -1140 1723 -1116 1757
rect -1082 1723 -1058 1757
rect -1140 1685 -1058 1723
rect -1140 1651 -1116 1685
rect -1082 1651 -1058 1685
rect -1140 1613 -1058 1651
rect -1140 1579 -1116 1613
rect -1082 1579 -1058 1613
rect -1140 1541 -1058 1579
rect -1140 1507 -1116 1541
rect -1082 1507 -1058 1541
rect -1140 1469 -1058 1507
rect -1140 1435 -1116 1469
rect -1082 1435 -1058 1469
rect -1140 1397 -1058 1435
rect -1140 1363 -1116 1397
rect -1082 1363 -1058 1397
rect -1140 1325 -1058 1363
rect -1140 1291 -1116 1325
rect -1082 1291 -1058 1325
rect -1140 1253 -1058 1291
rect -1140 1219 -1116 1253
rect -1082 1219 -1058 1253
rect -1140 1181 -1058 1219
rect -1140 1147 -1116 1181
rect -1082 1147 -1058 1181
rect -1140 1109 -1058 1147
rect -1140 1075 -1116 1109
rect -1082 1075 -1058 1109
rect -1140 1037 -1058 1075
rect -1140 1003 -1116 1037
rect -1082 1003 -1058 1037
rect -1140 965 -1058 1003
rect -1140 931 -1116 965
rect -1082 931 -1058 965
rect -1140 893 -1058 931
rect -1140 859 -1116 893
rect -1082 859 -1058 893
rect -1140 821 -1058 859
rect -1140 787 -1116 821
rect -1082 787 -1058 821
rect -1140 749 -1058 787
rect -1140 715 -1116 749
rect -1082 715 -1058 749
rect -1140 677 -1058 715
rect -1140 643 -1116 677
rect -1082 643 -1058 677
rect -1140 605 -1058 643
rect -1140 571 -1116 605
rect -1082 571 -1058 605
rect -1140 533 -1058 571
rect -1140 499 -1116 533
rect -1082 499 -1058 533
rect -1140 461 -1058 499
rect -1140 427 -1116 461
rect -1082 427 -1058 461
rect -1140 389 -1058 427
rect -1140 355 -1116 389
rect -1082 355 -1058 389
rect -1140 317 -1058 355
rect -1140 283 -1116 317
rect -1082 283 -1058 317
rect -1140 245 -1058 283
rect -1140 211 -1116 245
rect -1082 211 -1058 245
rect -1140 173 -1058 211
rect -1140 139 -1116 173
rect -1082 139 -1058 173
rect -1140 101 -1058 139
rect -1140 67 -1116 101
rect -1082 67 -1058 101
rect -1140 29 -1058 67
rect -1140 -5 -1116 29
rect -1082 -5 -1058 29
rect -958 5969 -900 5981
rect -958 5935 -946 5969
rect -912 5935 -900 5969
rect 1050 5969 1108 5981
rect -958 5897 -900 5935
rect -958 5863 -946 5897
rect -912 5863 -900 5897
rect -958 5825 -900 5863
rect -958 5791 -946 5825
rect -912 5791 -900 5825
rect -958 5753 -900 5791
rect -958 5719 -946 5753
rect -912 5719 -900 5753
rect -958 5681 -900 5719
rect -958 5647 -946 5681
rect -912 5647 -900 5681
rect -958 5609 -900 5647
rect -958 5575 -946 5609
rect -912 5575 -900 5609
rect -958 5537 -900 5575
rect -958 5503 -946 5537
rect -912 5503 -900 5537
rect -958 5465 -900 5503
rect -958 5431 -946 5465
rect -912 5431 -900 5465
rect -958 5393 -900 5431
rect -958 5359 -946 5393
rect -912 5359 -900 5393
rect -958 5321 -900 5359
rect -958 5287 -946 5321
rect -912 5287 -900 5321
rect -958 5249 -900 5287
rect -958 5215 -946 5249
rect -912 5215 -900 5249
rect -958 5177 -900 5215
rect -958 5143 -946 5177
rect -912 5143 -900 5177
rect -958 5105 -900 5143
rect -958 5071 -946 5105
rect -912 5071 -900 5105
rect -958 5033 -900 5071
rect -958 4999 -946 5033
rect -912 4999 -900 5033
rect -958 4961 -900 4999
rect -958 4927 -946 4961
rect -912 4927 -900 4961
rect -958 4889 -900 4927
rect -958 4855 -946 4889
rect -912 4855 -900 4889
rect -958 4817 -900 4855
rect -958 4783 -946 4817
rect -912 4783 -900 4817
rect -958 4745 -900 4783
rect -958 4711 -946 4745
rect -912 4711 -900 4745
rect -958 4673 -900 4711
rect -958 4639 -946 4673
rect -912 4639 -900 4673
rect -958 4601 -900 4639
rect -958 4567 -946 4601
rect -912 4567 -900 4601
rect -958 4529 -900 4567
rect -958 4495 -946 4529
rect -912 4495 -900 4529
rect -958 4457 -900 4495
rect -958 4423 -946 4457
rect -912 4423 -900 4457
rect -958 4385 -900 4423
rect -958 4351 -946 4385
rect -912 4351 -900 4385
rect -958 4313 -900 4351
rect -958 4279 -946 4313
rect -912 4279 -900 4313
rect -958 4241 -900 4279
rect -958 4207 -946 4241
rect -912 4207 -900 4241
rect -958 4169 -900 4207
rect -958 4135 -946 4169
rect -912 4135 -900 4169
rect -958 4097 -900 4135
rect -958 4063 -946 4097
rect -912 4063 -900 4097
rect -958 4025 -900 4063
rect -958 3991 -946 4025
rect -912 3991 -900 4025
rect -958 3953 -900 3991
rect -958 3919 -946 3953
rect -912 3919 -900 3953
rect -958 3881 -900 3919
rect -958 3847 -946 3881
rect -912 3847 -900 3881
rect -958 3809 -900 3847
rect -958 3775 -946 3809
rect -912 3775 -900 3809
rect -958 3737 -900 3775
rect -958 3703 -946 3737
rect -912 3703 -900 3737
rect -958 3665 -900 3703
rect -958 3631 -946 3665
rect -912 3631 -900 3665
rect -958 3593 -900 3631
rect -958 3559 -946 3593
rect -912 3559 -900 3593
rect -958 3521 -900 3559
rect -958 3487 -946 3521
rect -912 3487 -900 3521
rect -958 3449 -900 3487
rect -958 3415 -946 3449
rect -912 3415 -900 3449
rect -958 3377 -900 3415
rect -958 3343 -946 3377
rect -912 3343 -900 3377
rect -958 3305 -900 3343
rect -958 3271 -946 3305
rect -912 3271 -900 3305
rect -958 3233 -900 3271
rect -958 3199 -946 3233
rect -912 3199 -900 3233
rect -958 3161 -900 3199
rect -958 3127 -946 3161
rect -912 3127 -900 3161
rect -958 3089 -900 3127
rect -958 3055 -946 3089
rect -912 3055 -900 3089
rect -958 3017 -900 3055
rect -958 2983 -946 3017
rect -912 2983 -900 3017
rect -958 2945 -900 2983
rect -958 2911 -946 2945
rect -912 2911 -900 2945
rect -958 2873 -900 2911
rect -958 2839 -946 2873
rect -912 2839 -900 2873
rect -958 2801 -900 2839
rect -958 2767 -946 2801
rect -912 2767 -900 2801
rect -958 2729 -900 2767
rect -958 2695 -946 2729
rect -912 2695 -900 2729
rect -958 2657 -900 2695
rect -958 2623 -946 2657
rect -912 2623 -900 2657
rect -958 2585 -900 2623
rect -958 2551 -946 2585
rect -912 2551 -900 2585
rect -958 2513 -900 2551
rect -958 2479 -946 2513
rect -912 2479 -900 2513
rect -958 2441 -900 2479
rect -958 2407 -946 2441
rect -912 2407 -900 2441
rect -958 2369 -900 2407
rect -958 2335 -946 2369
rect -912 2335 -900 2369
rect -958 2297 -900 2335
rect -958 2263 -946 2297
rect -912 2263 -900 2297
rect -958 2225 -900 2263
rect -958 2191 -946 2225
rect -912 2191 -900 2225
rect -958 2153 -900 2191
rect -958 2119 -946 2153
rect -912 2119 -900 2153
rect -958 2081 -900 2119
rect -958 2047 -946 2081
rect -912 2047 -900 2081
rect -958 2009 -900 2047
rect -958 1975 -946 2009
rect -912 1975 -900 2009
rect -958 1937 -900 1975
rect -958 1903 -946 1937
rect -912 1903 -900 1937
rect -958 1865 -900 1903
rect -958 1831 -946 1865
rect -912 1831 -900 1865
rect -958 1793 -900 1831
rect -958 1759 -946 1793
rect -912 1759 -900 1793
rect -958 1721 -900 1759
rect -958 1687 -946 1721
rect -912 1687 -900 1721
rect -958 1649 -900 1687
rect -958 1615 -946 1649
rect -912 1615 -900 1649
rect -958 1577 -900 1615
rect -958 1543 -946 1577
rect -912 1543 -900 1577
rect -958 1505 -900 1543
rect -958 1471 -946 1505
rect -912 1471 -900 1505
rect -958 1433 -900 1471
rect -958 1399 -946 1433
rect -912 1399 -900 1433
rect -958 1361 -900 1399
rect -958 1327 -946 1361
rect -912 1327 -900 1361
rect -958 1289 -900 1327
rect -958 1255 -946 1289
rect -912 1255 -900 1289
rect -958 1217 -900 1255
rect -958 1183 -946 1217
rect -912 1183 -900 1217
rect -958 1145 -900 1183
rect -958 1111 -946 1145
rect -912 1111 -900 1145
rect -958 1073 -900 1111
rect -958 1039 -946 1073
rect -912 1039 -900 1073
rect -958 1001 -900 1039
rect -958 967 -946 1001
rect -912 967 -900 1001
rect -958 929 -900 967
rect -958 895 -946 929
rect -912 895 -900 929
rect -958 857 -900 895
rect -958 823 -946 857
rect -912 823 -900 857
rect -958 785 -900 823
rect -958 751 -946 785
rect -912 751 -900 785
rect -958 713 -900 751
rect -958 679 -946 713
rect -912 679 -900 713
rect -958 641 -900 679
rect -958 607 -946 641
rect -912 607 -900 641
rect -958 569 -900 607
rect -958 535 -946 569
rect -912 535 -900 569
rect -958 497 -900 535
rect -958 463 -946 497
rect -912 463 -900 497
rect -958 425 -900 463
rect -958 391 -946 425
rect -912 391 -900 425
rect -958 353 -900 391
rect -958 319 -946 353
rect -912 319 -900 353
rect -958 281 -900 319
rect -958 247 -946 281
rect -912 247 -900 281
rect -958 209 -900 247
rect -958 175 -946 209
rect -912 175 -900 209
rect -958 137 -900 175
rect -958 103 -946 137
rect -912 103 -900 137
rect -958 65 -900 103
rect -958 31 -946 65
rect -912 31 -900 65
rect 10 5939 140 5945
rect 10 63 17 5939
rect 133 63 140 5939
rect 10 55 140 63
rect 1050 5935 1062 5969
rect 1096 5935 1108 5969
rect 1050 5897 1108 5935
rect 1050 5863 1062 5897
rect 1096 5863 1108 5897
rect 1050 5825 1108 5863
rect 1050 5791 1062 5825
rect 1096 5791 1108 5825
rect 1050 5753 1108 5791
rect 1050 5719 1062 5753
rect 1096 5719 1108 5753
rect 1050 5681 1108 5719
rect 1050 5647 1062 5681
rect 1096 5647 1108 5681
rect 1050 5609 1108 5647
rect 1050 5575 1062 5609
rect 1096 5575 1108 5609
rect 1050 5537 1108 5575
rect 1050 5503 1062 5537
rect 1096 5503 1108 5537
rect 1050 5465 1108 5503
rect 1050 5431 1062 5465
rect 1096 5431 1108 5465
rect 1050 5393 1108 5431
rect 1050 5359 1062 5393
rect 1096 5359 1108 5393
rect 1050 5321 1108 5359
rect 1050 5287 1062 5321
rect 1096 5287 1108 5321
rect 1050 5249 1108 5287
rect 1050 5215 1062 5249
rect 1096 5215 1108 5249
rect 1050 5177 1108 5215
rect 1050 5143 1062 5177
rect 1096 5143 1108 5177
rect 1050 5105 1108 5143
rect 1050 5071 1062 5105
rect 1096 5071 1108 5105
rect 1050 5033 1108 5071
rect 1050 4999 1062 5033
rect 1096 4999 1108 5033
rect 1050 4961 1108 4999
rect 1050 4927 1062 4961
rect 1096 4927 1108 4961
rect 1050 4889 1108 4927
rect 1050 4855 1062 4889
rect 1096 4855 1108 4889
rect 1050 4817 1108 4855
rect 1050 4783 1062 4817
rect 1096 4783 1108 4817
rect 1050 4745 1108 4783
rect 1050 4711 1062 4745
rect 1096 4711 1108 4745
rect 1050 4673 1108 4711
rect 1050 4639 1062 4673
rect 1096 4639 1108 4673
rect 1050 4601 1108 4639
rect 1050 4567 1062 4601
rect 1096 4567 1108 4601
rect 1050 4529 1108 4567
rect 1050 4495 1062 4529
rect 1096 4495 1108 4529
rect 1050 4457 1108 4495
rect 1050 4423 1062 4457
rect 1096 4423 1108 4457
rect 1050 4385 1108 4423
rect 1050 4351 1062 4385
rect 1096 4351 1108 4385
rect 1050 4313 1108 4351
rect 1050 4279 1062 4313
rect 1096 4279 1108 4313
rect 1050 4241 1108 4279
rect 1050 4207 1062 4241
rect 1096 4207 1108 4241
rect 1050 4169 1108 4207
rect 1050 4135 1062 4169
rect 1096 4135 1108 4169
rect 1050 4097 1108 4135
rect 1050 4063 1062 4097
rect 1096 4063 1108 4097
rect 1050 4025 1108 4063
rect 1050 3991 1062 4025
rect 1096 3991 1108 4025
rect 1050 3953 1108 3991
rect 1050 3919 1062 3953
rect 1096 3919 1108 3953
rect 1050 3881 1108 3919
rect 1050 3847 1062 3881
rect 1096 3847 1108 3881
rect 1050 3809 1108 3847
rect 1050 3775 1062 3809
rect 1096 3775 1108 3809
rect 1050 3737 1108 3775
rect 1050 3703 1062 3737
rect 1096 3703 1108 3737
rect 1050 3665 1108 3703
rect 1050 3631 1062 3665
rect 1096 3631 1108 3665
rect 1050 3593 1108 3631
rect 1050 3559 1062 3593
rect 1096 3559 1108 3593
rect 1050 3521 1108 3559
rect 1050 3487 1062 3521
rect 1096 3487 1108 3521
rect 1050 3449 1108 3487
rect 1050 3415 1062 3449
rect 1096 3415 1108 3449
rect 1050 3377 1108 3415
rect 1050 3343 1062 3377
rect 1096 3343 1108 3377
rect 1050 3305 1108 3343
rect 1050 3271 1062 3305
rect 1096 3271 1108 3305
rect 1050 3233 1108 3271
rect 1050 3199 1062 3233
rect 1096 3199 1108 3233
rect 1050 3161 1108 3199
rect 1050 3127 1062 3161
rect 1096 3127 1108 3161
rect 1050 3089 1108 3127
rect 1050 3055 1062 3089
rect 1096 3055 1108 3089
rect 1050 3017 1108 3055
rect 1050 2983 1062 3017
rect 1096 2983 1108 3017
rect 1050 2945 1108 2983
rect 1050 2911 1062 2945
rect 1096 2911 1108 2945
rect 1050 2873 1108 2911
rect 1050 2839 1062 2873
rect 1096 2839 1108 2873
rect 1050 2801 1108 2839
rect 1050 2767 1062 2801
rect 1096 2767 1108 2801
rect 1050 2729 1108 2767
rect 1050 2695 1062 2729
rect 1096 2695 1108 2729
rect 1050 2657 1108 2695
rect 1050 2623 1062 2657
rect 1096 2623 1108 2657
rect 1050 2585 1108 2623
rect 1050 2551 1062 2585
rect 1096 2551 1108 2585
rect 1050 2513 1108 2551
rect 1050 2479 1062 2513
rect 1096 2479 1108 2513
rect 1050 2441 1108 2479
rect 1050 2407 1062 2441
rect 1096 2407 1108 2441
rect 1050 2369 1108 2407
rect 1050 2335 1062 2369
rect 1096 2335 1108 2369
rect 1050 2297 1108 2335
rect 1050 2263 1062 2297
rect 1096 2263 1108 2297
rect 1050 2225 1108 2263
rect 1050 2191 1062 2225
rect 1096 2191 1108 2225
rect 1050 2153 1108 2191
rect 1050 2119 1062 2153
rect 1096 2119 1108 2153
rect 1050 2081 1108 2119
rect 1050 2047 1062 2081
rect 1096 2047 1108 2081
rect 1050 2009 1108 2047
rect 1050 1975 1062 2009
rect 1096 1975 1108 2009
rect 1050 1937 1108 1975
rect 1050 1903 1062 1937
rect 1096 1903 1108 1937
rect 1050 1865 1108 1903
rect 1050 1831 1062 1865
rect 1096 1831 1108 1865
rect 1050 1793 1108 1831
rect 1050 1759 1062 1793
rect 1096 1759 1108 1793
rect 1050 1721 1108 1759
rect 1050 1687 1062 1721
rect 1096 1687 1108 1721
rect 1050 1649 1108 1687
rect 1050 1615 1062 1649
rect 1096 1615 1108 1649
rect 1050 1577 1108 1615
rect 1050 1543 1062 1577
rect 1096 1543 1108 1577
rect 1050 1505 1108 1543
rect 1050 1471 1062 1505
rect 1096 1471 1108 1505
rect 1050 1433 1108 1471
rect 1050 1399 1062 1433
rect 1096 1399 1108 1433
rect 1050 1361 1108 1399
rect 1050 1327 1062 1361
rect 1096 1327 1108 1361
rect 1050 1289 1108 1327
rect 1050 1255 1062 1289
rect 1096 1255 1108 1289
rect 1050 1217 1108 1255
rect 1050 1183 1062 1217
rect 1096 1183 1108 1217
rect 1050 1145 1108 1183
rect 1050 1111 1062 1145
rect 1096 1111 1108 1145
rect 1050 1073 1108 1111
rect 1050 1039 1062 1073
rect 1096 1039 1108 1073
rect 1050 1001 1108 1039
rect 1050 967 1062 1001
rect 1096 967 1108 1001
rect 1050 929 1108 967
rect 1050 895 1062 929
rect 1096 895 1108 929
rect 1050 857 1108 895
rect 1050 823 1062 857
rect 1096 823 1108 857
rect 1050 785 1108 823
rect 1050 751 1062 785
rect 1096 751 1108 785
rect 1050 713 1108 751
rect 1050 679 1062 713
rect 1096 679 1108 713
rect 1050 641 1108 679
rect 1050 607 1062 641
rect 1096 607 1108 641
rect 1050 569 1108 607
rect 1050 535 1062 569
rect 1096 535 1108 569
rect 1050 497 1108 535
rect 1050 463 1062 497
rect 1096 463 1108 497
rect 1050 425 1108 463
rect 1050 391 1062 425
rect 1096 391 1108 425
rect 1050 353 1108 391
rect 1050 319 1062 353
rect 1096 319 1108 353
rect 1050 281 1108 319
rect 1050 247 1062 281
rect 1096 247 1108 281
rect 1050 209 1108 247
rect 1050 175 1062 209
rect 1096 175 1108 209
rect 1050 137 1108 175
rect 1050 103 1062 137
rect 1096 103 1108 137
rect 1050 65 1108 103
rect -958 19 -900 31
rect 1050 31 1062 65
rect 1096 31 1108 65
rect 1050 19 1108 31
rect 1208 5971 1232 6005
rect 1266 5971 1290 6005
rect 1208 5933 1290 5971
rect 1208 5899 1232 5933
rect 1266 5899 1290 5933
rect 1208 5861 1290 5899
rect 1208 5827 1232 5861
rect 1266 5827 1290 5861
rect 1208 5789 1290 5827
rect 1208 5755 1232 5789
rect 1266 5755 1290 5789
rect 1208 5717 1290 5755
rect 1208 5683 1232 5717
rect 1266 5683 1290 5717
rect 1208 5645 1290 5683
rect 1208 5611 1232 5645
rect 1266 5611 1290 5645
rect 1208 5573 1290 5611
rect 1208 5539 1232 5573
rect 1266 5539 1290 5573
rect 1208 5501 1290 5539
rect 1208 5467 1232 5501
rect 1266 5467 1290 5501
rect 1208 5429 1290 5467
rect 1208 5395 1232 5429
rect 1266 5395 1290 5429
rect 1208 5357 1290 5395
rect 1208 5323 1232 5357
rect 1266 5323 1290 5357
rect 1208 5285 1290 5323
rect 1208 5251 1232 5285
rect 1266 5251 1290 5285
rect 1208 5213 1290 5251
rect 1208 5179 1232 5213
rect 1266 5179 1290 5213
rect 1208 5141 1290 5179
rect 1208 5107 1232 5141
rect 1266 5107 1290 5141
rect 1208 5069 1290 5107
rect 1208 5035 1232 5069
rect 1266 5035 1290 5069
rect 1208 4997 1290 5035
rect 1208 4963 1232 4997
rect 1266 4963 1290 4997
rect 1208 4925 1290 4963
rect 1208 4891 1232 4925
rect 1266 4891 1290 4925
rect 1208 4853 1290 4891
rect 1208 4819 1232 4853
rect 1266 4819 1290 4853
rect 1208 4781 1290 4819
rect 1208 4747 1232 4781
rect 1266 4747 1290 4781
rect 1208 4709 1290 4747
rect 1208 4675 1232 4709
rect 1266 4675 1290 4709
rect 1208 4637 1290 4675
rect 1208 4603 1232 4637
rect 1266 4603 1290 4637
rect 1208 4565 1290 4603
rect 1208 4531 1232 4565
rect 1266 4531 1290 4565
rect 1208 4493 1290 4531
rect 1208 4459 1232 4493
rect 1266 4459 1290 4493
rect 1208 4421 1290 4459
rect 1208 4387 1232 4421
rect 1266 4387 1290 4421
rect 1208 4349 1290 4387
rect 1208 4315 1232 4349
rect 1266 4315 1290 4349
rect 1208 4277 1290 4315
rect 1208 4243 1232 4277
rect 1266 4243 1290 4277
rect 1208 4205 1290 4243
rect 1208 4171 1232 4205
rect 1266 4171 1290 4205
rect 1208 4133 1290 4171
rect 1208 4099 1232 4133
rect 1266 4099 1290 4133
rect 1208 4061 1290 4099
rect 1208 4027 1232 4061
rect 1266 4027 1290 4061
rect 1208 3989 1290 4027
rect 1208 3955 1232 3989
rect 1266 3955 1290 3989
rect 1208 3917 1290 3955
rect 1208 3883 1232 3917
rect 1266 3883 1290 3917
rect 1208 3845 1290 3883
rect 1208 3811 1232 3845
rect 1266 3811 1290 3845
rect 1208 3773 1290 3811
rect 1208 3739 1232 3773
rect 1266 3739 1290 3773
rect 1208 3701 1290 3739
rect 1208 3667 1232 3701
rect 1266 3667 1290 3701
rect 1208 3629 1290 3667
rect 1208 3595 1232 3629
rect 1266 3595 1290 3629
rect 1208 3557 1290 3595
rect 1208 3523 1232 3557
rect 1266 3523 1290 3557
rect 1208 3485 1290 3523
rect 1208 3451 1232 3485
rect 1266 3451 1290 3485
rect 1208 3413 1290 3451
rect 1208 3379 1232 3413
rect 1266 3379 1290 3413
rect 1208 3341 1290 3379
rect 1208 3307 1232 3341
rect 1266 3307 1290 3341
rect 1208 3269 1290 3307
rect 1208 3235 1232 3269
rect 1266 3235 1290 3269
rect 1208 3197 1290 3235
rect 1208 3163 1232 3197
rect 1266 3163 1290 3197
rect 1208 3125 1290 3163
rect 1208 3091 1232 3125
rect 1266 3091 1290 3125
rect 1208 3053 1290 3091
rect 1208 3019 1232 3053
rect 1266 3019 1290 3053
rect 1208 2981 1290 3019
rect 1208 2947 1232 2981
rect 1266 2947 1290 2981
rect 1208 2909 1290 2947
rect 1208 2875 1232 2909
rect 1266 2875 1290 2909
rect 1208 2837 1290 2875
rect 1208 2803 1232 2837
rect 1266 2803 1290 2837
rect 1208 2765 1290 2803
rect 1208 2731 1232 2765
rect 1266 2731 1290 2765
rect 1208 2693 1290 2731
rect 1208 2659 1232 2693
rect 1266 2659 1290 2693
rect 1208 2621 1290 2659
rect 1208 2587 1232 2621
rect 1266 2587 1290 2621
rect 1208 2549 1290 2587
rect 1208 2515 1232 2549
rect 1266 2515 1290 2549
rect 1208 2477 1290 2515
rect 1208 2443 1232 2477
rect 1266 2443 1290 2477
rect 1208 2405 1290 2443
rect 1208 2371 1232 2405
rect 1266 2371 1290 2405
rect 1208 2333 1290 2371
rect 1208 2299 1232 2333
rect 1266 2299 1290 2333
rect 1208 2261 1290 2299
rect 1208 2227 1232 2261
rect 1266 2227 1290 2261
rect 1208 2189 1290 2227
rect 1208 2155 1232 2189
rect 1266 2155 1290 2189
rect 1208 2117 1290 2155
rect 1208 2083 1232 2117
rect 1266 2083 1290 2117
rect 1208 2045 1290 2083
rect 1208 2011 1232 2045
rect 1266 2011 1290 2045
rect 1208 1973 1290 2011
rect 1208 1939 1232 1973
rect 1266 1939 1290 1973
rect 1208 1901 1290 1939
rect 1208 1867 1232 1901
rect 1266 1867 1290 1901
rect 1208 1829 1290 1867
rect 1208 1795 1232 1829
rect 1266 1795 1290 1829
rect 1208 1757 1290 1795
rect 1208 1723 1232 1757
rect 1266 1723 1290 1757
rect 1208 1685 1290 1723
rect 1208 1651 1232 1685
rect 1266 1651 1290 1685
rect 1208 1613 1290 1651
rect 1208 1579 1232 1613
rect 1266 1579 1290 1613
rect 1208 1541 1290 1579
rect 1208 1507 1232 1541
rect 1266 1507 1290 1541
rect 1208 1469 1290 1507
rect 1208 1435 1232 1469
rect 1266 1435 1290 1469
rect 1208 1397 1290 1435
rect 1208 1363 1232 1397
rect 1266 1363 1290 1397
rect 1208 1325 1290 1363
rect 1208 1291 1232 1325
rect 1266 1291 1290 1325
rect 1208 1253 1290 1291
rect 1208 1219 1232 1253
rect 1266 1219 1290 1253
rect 1208 1181 1290 1219
rect 1208 1147 1232 1181
rect 1266 1147 1290 1181
rect 1208 1109 1290 1147
rect 1208 1075 1232 1109
rect 1266 1075 1290 1109
rect 1208 1037 1290 1075
rect 1208 1003 1232 1037
rect 1266 1003 1290 1037
rect 1208 965 1290 1003
rect 1208 931 1232 965
rect 1266 931 1290 965
rect 1208 893 1290 931
rect 1208 859 1232 893
rect 1266 859 1290 893
rect 1208 821 1290 859
rect 1208 787 1232 821
rect 1266 787 1290 821
rect 1208 749 1290 787
rect 1208 715 1232 749
rect 1266 715 1290 749
rect 1208 677 1290 715
rect 1208 643 1232 677
rect 1266 643 1290 677
rect 1208 605 1290 643
rect 1208 571 1232 605
rect 1266 571 1290 605
rect 1208 533 1290 571
rect 1208 499 1232 533
rect 1266 499 1290 533
rect 1208 461 1290 499
rect 1208 427 1232 461
rect 1266 427 1290 461
rect 1208 389 1290 427
rect 1208 355 1232 389
rect 1266 355 1290 389
rect 1208 317 1290 355
rect 1208 283 1232 317
rect 1266 283 1290 317
rect 1208 245 1290 283
rect 1208 211 1232 245
rect 1266 211 1290 245
rect 1208 173 1290 211
rect 1208 139 1232 173
rect 1266 139 1290 173
rect 1208 101 1290 139
rect 1208 67 1232 101
rect 1266 67 1290 101
rect 1208 29 1290 67
rect -1140 -43 -1058 -5
rect -1140 -77 -1116 -43
rect -1082 -77 -1058 -43
rect -1140 -115 -1058 -77
rect -1140 -149 -1116 -115
rect -1082 -149 -1058 -115
rect -1140 -187 -1058 -149
rect -1140 -221 -1116 -187
rect -1082 -221 -1058 -187
rect -1140 -259 -1058 -221
rect -1140 -293 -1116 -259
rect -1082 -293 -1058 -259
rect -1140 -331 -1058 -293
rect -1140 -365 -1116 -331
rect -1082 -365 -1058 -331
rect -1140 -403 -1058 -365
rect -1140 -437 -1116 -403
rect -1082 -437 -1058 -403
rect -1140 -475 -1058 -437
rect -1140 -509 -1116 -475
rect -1082 -509 -1058 -475
rect -1140 -547 -1058 -509
rect -1140 -581 -1116 -547
rect -1082 -581 -1058 -547
rect -1140 -619 -1058 -581
rect -1140 -653 -1116 -619
rect -1082 -653 -1058 -619
rect 1208 -5 1232 29
rect 1266 -5 1290 29
rect 1208 -43 1290 -5
rect 1208 -77 1232 -43
rect 1266 -77 1290 -43
rect 1208 -115 1290 -77
rect 1208 -149 1232 -115
rect 1266 -149 1290 -115
rect 1208 -187 1290 -149
rect 1208 -221 1232 -187
rect 1266 -221 1290 -187
rect 1208 -259 1290 -221
rect 1208 -293 1232 -259
rect 1266 -293 1290 -259
rect 1208 -331 1290 -293
rect 1208 -365 1232 -331
rect 1266 -365 1290 -331
rect 1208 -403 1290 -365
rect 1208 -437 1232 -403
rect 1266 -437 1290 -403
rect 1208 -475 1290 -437
rect 1208 -509 1232 -475
rect 1266 -509 1290 -475
rect 1208 -547 1290 -509
rect 1208 -581 1232 -547
rect 1266 -581 1290 -547
rect 1208 -619 1290 -581
rect -1140 -691 -1058 -653
rect -1140 -725 -1116 -691
rect -1082 -725 -1058 -691
rect -1140 -763 -1058 -725
rect -1140 -797 -1116 -763
rect -1082 -797 -1058 -763
rect -1140 -835 -1058 -797
rect -1140 -869 -1116 -835
rect -1082 -869 -1058 -835
rect -296 -650 460 -643
rect -296 -702 -289 -650
rect -237 -702 -215 -650
rect -163 -702 -141 -650
rect -89 -702 -67 -650
rect -15 -702 7 -650
rect 59 -702 81 -650
rect 133 -702 155 -650
rect 207 -702 229 -650
rect 281 -702 303 -650
rect 355 -702 377 -650
rect 429 -702 460 -650
rect -296 -724 460 -702
rect -296 -776 -289 -724
rect -237 -776 -215 -724
rect -163 -776 -141 -724
rect -89 -776 -67 -724
rect -15 -776 7 -724
rect 59 -776 81 -724
rect 133 -776 155 -724
rect 207 -776 229 -724
rect 281 -776 303 -724
rect 355 -776 377 -724
rect 429 -776 460 -724
rect -296 -798 460 -776
rect -296 -850 -289 -798
rect -237 -850 -215 -798
rect -163 -850 -141 -798
rect -89 -850 -67 -798
rect -15 -850 7 -798
rect 59 -850 81 -798
rect 133 -850 155 -798
rect 207 -850 229 -798
rect 281 -850 303 -798
rect 355 -850 377 -798
rect 429 -850 460 -798
rect -296 -857 460 -850
rect 1208 -653 1232 -619
rect 1266 -653 1290 -619
rect 1208 -691 1290 -653
rect 1208 -725 1232 -691
rect 1266 -725 1290 -691
rect 1208 -763 1290 -725
rect 1208 -797 1232 -763
rect 1266 -797 1290 -763
rect 1208 -835 1290 -797
rect -1140 -907 -1058 -869
rect -1140 -941 -1116 -907
rect -1082 -941 -1058 -907
rect -1140 -979 -1058 -941
rect -1140 -1013 -1116 -979
rect -1082 -1013 -1058 -979
rect -1140 -1051 -1058 -1013
rect -1140 -1085 -1116 -1051
rect -1082 -1085 -1058 -1051
rect -1140 -1100 -1058 -1085
rect 1208 -869 1232 -835
rect 1266 -869 1290 -835
rect 1208 -907 1290 -869
rect 1208 -941 1232 -907
rect 1266 -941 1290 -907
rect 1208 -979 1290 -941
rect 1208 -1013 1232 -979
rect 1266 -1013 1290 -979
rect 1208 -1051 1290 -1013
rect 1208 -1085 1232 -1051
rect 1266 -1085 1290 -1051
rect 1208 -1100 1290 -1085
rect -1140 -1124 1290 -1100
rect -1140 -1158 -986 -1124
rect -952 -1158 -914 -1124
rect -880 -1158 -842 -1124
rect -808 -1158 -770 -1124
rect -736 -1158 -698 -1124
rect -664 -1158 -626 -1124
rect -592 -1158 -554 -1124
rect -520 -1158 -482 -1124
rect -448 -1158 -410 -1124
rect -376 -1158 -338 -1124
rect -304 -1158 -266 -1124
rect -232 -1158 -194 -1124
rect -160 -1158 -122 -1124
rect -88 -1158 -50 -1124
rect -16 -1158 22 -1124
rect 56 -1158 94 -1124
rect 128 -1158 166 -1124
rect 200 -1158 238 -1124
rect 272 -1158 310 -1124
rect 344 -1158 382 -1124
rect 416 -1158 454 -1124
rect 488 -1158 526 -1124
rect 560 -1158 598 -1124
rect 632 -1158 670 -1124
rect 704 -1158 742 -1124
rect 776 -1158 814 -1124
rect 848 -1158 886 -1124
rect 920 -1158 958 -1124
rect 992 -1158 1030 -1124
rect 1064 -1158 1102 -1124
rect 1136 -1158 1290 -1124
rect -1140 -1182 1290 -1158
<< via1 >>
rect 17 5933 133 5939
rect 17 67 22 5933
rect 22 67 128 5933
rect 128 67 133 5933
rect 17 63 133 67
rect -289 -659 -237 -650
rect -289 -693 -280 -659
rect -280 -693 -246 -659
rect -246 -693 -237 -659
rect -289 -702 -237 -693
rect -215 -659 -163 -650
rect -215 -693 -206 -659
rect -206 -693 -172 -659
rect -172 -693 -163 -659
rect -215 -702 -163 -693
rect -141 -659 -89 -650
rect -141 -693 -132 -659
rect -132 -693 -98 -659
rect -98 -693 -89 -659
rect -141 -702 -89 -693
rect -67 -659 -15 -650
rect -67 -693 -58 -659
rect -58 -693 -24 -659
rect -24 -693 -15 -659
rect -67 -702 -15 -693
rect 7 -659 59 -650
rect 7 -693 16 -659
rect 16 -693 50 -659
rect 50 -693 59 -659
rect 7 -702 59 -693
rect 81 -659 133 -650
rect 81 -693 90 -659
rect 90 -693 124 -659
rect 124 -693 133 -659
rect 81 -702 133 -693
rect 155 -659 207 -650
rect 155 -693 164 -659
rect 164 -693 198 -659
rect 198 -693 207 -659
rect 155 -702 207 -693
rect 229 -659 281 -650
rect 229 -693 238 -659
rect 238 -693 272 -659
rect 272 -693 281 -659
rect 229 -702 281 -693
rect 303 -659 355 -650
rect 303 -693 312 -659
rect 312 -693 346 -659
rect 346 -693 355 -659
rect 303 -702 355 -693
rect 377 -659 429 -650
rect 377 -693 386 -659
rect 386 -693 420 -659
rect 420 -693 429 -659
rect 377 -702 429 -693
rect -289 -733 -237 -724
rect -289 -767 -280 -733
rect -280 -767 -246 -733
rect -246 -767 -237 -733
rect -289 -776 -237 -767
rect -215 -733 -163 -724
rect -215 -767 -206 -733
rect -206 -767 -172 -733
rect -172 -767 -163 -733
rect -215 -776 -163 -767
rect -141 -733 -89 -724
rect -141 -767 -132 -733
rect -132 -767 -98 -733
rect -98 -767 -89 -733
rect -141 -776 -89 -767
rect -67 -733 -15 -724
rect -67 -767 -58 -733
rect -58 -767 -24 -733
rect -24 -767 -15 -733
rect -67 -776 -15 -767
rect 7 -733 59 -724
rect 7 -767 16 -733
rect 16 -767 50 -733
rect 50 -767 59 -733
rect 7 -776 59 -767
rect 81 -733 133 -724
rect 81 -767 90 -733
rect 90 -767 124 -733
rect 124 -767 133 -733
rect 81 -776 133 -767
rect 155 -733 207 -724
rect 155 -767 164 -733
rect 164 -767 198 -733
rect 198 -767 207 -733
rect 155 -776 207 -767
rect 229 -733 281 -724
rect 229 -767 238 -733
rect 238 -767 272 -733
rect 272 -767 281 -733
rect 229 -776 281 -767
rect 303 -733 355 -724
rect 303 -767 312 -733
rect 312 -767 346 -733
rect 346 -767 355 -733
rect 303 -776 355 -767
rect 377 -733 429 -724
rect 377 -767 386 -733
rect 386 -767 420 -733
rect 420 -767 429 -733
rect 377 -776 429 -767
rect -289 -807 -237 -798
rect -289 -841 -280 -807
rect -280 -841 -246 -807
rect -246 -841 -237 -807
rect -289 -850 -237 -841
rect -215 -807 -163 -798
rect -215 -841 -206 -807
rect -206 -841 -172 -807
rect -172 -841 -163 -807
rect -215 -850 -163 -841
rect -141 -807 -89 -798
rect -141 -841 -132 -807
rect -132 -841 -98 -807
rect -98 -841 -89 -807
rect -141 -850 -89 -841
rect -67 -807 -15 -798
rect -67 -841 -58 -807
rect -58 -841 -24 -807
rect -24 -841 -15 -807
rect -67 -850 -15 -841
rect 7 -807 59 -798
rect 7 -841 16 -807
rect 16 -841 50 -807
rect 50 -841 59 -807
rect 7 -850 59 -841
rect 81 -807 133 -798
rect 81 -841 90 -807
rect 90 -841 124 -807
rect 124 -841 133 -807
rect 81 -850 133 -841
rect 155 -807 207 -798
rect 155 -841 164 -807
rect 164 -841 198 -807
rect 198 -841 207 -807
rect 155 -850 207 -841
rect 229 -807 281 -798
rect 229 -841 238 -807
rect 238 -841 272 -807
rect 272 -841 281 -807
rect 229 -850 281 -841
rect 303 -807 355 -798
rect 303 -841 312 -807
rect 312 -841 346 -807
rect 346 -841 355 -807
rect 303 -850 355 -841
rect 377 -807 429 -798
rect 377 -841 386 -807
rect 386 -841 420 -807
rect 420 -841 429 -807
rect 377 -850 429 -841
<< metal2 >>
rect 11 5939 139 5945
rect 11 63 17 5939
rect 133 63 139 5939
rect 11 57 139 63
rect -296 -650 460 -643
rect -296 -702 -289 -650
rect -237 -702 -215 -650
rect -163 -702 -141 -650
rect -89 -702 -67 -650
rect -15 -702 7 -650
rect 59 -702 81 -650
rect 133 -702 155 -650
rect 207 -702 229 -650
rect 281 -702 303 -650
rect 355 -702 377 -650
rect 429 -702 460 -650
rect -296 -724 460 -702
rect -296 -776 -289 -724
rect -237 -776 -215 -724
rect -163 -776 -141 -724
rect -89 -776 -67 -724
rect -15 -776 7 -724
rect 59 -776 81 -724
rect 133 -776 155 -724
rect 207 -776 229 -724
rect 281 -776 303 -724
rect 355 -776 377 -724
rect 429 -776 460 -724
rect -296 -798 460 -776
rect -296 -850 -289 -798
rect -237 -850 -215 -798
rect -163 -850 -141 -798
rect -89 -850 -67 -798
rect -15 -850 7 -798
rect 59 -850 81 -798
rect 133 -850 155 -798
rect 207 -850 229 -798
rect 281 -850 303 -798
rect 355 -850 377 -798
rect 429 -850 460 -798
rect -296 -857 460 -850
<< labels >>
flabel comment s 1085 159 1085 159 0 FreeSans 1600 0 0 0 S
flabel comment s -925 159 -925 159 0 FreeSans 1600 0 0 0 S
flabel comment s 67 159 67 159 0 FreeSans 1600 0 0 0 D
<< properties >>
string GDS_END 7253944
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 7133936
<< end >>
