magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -83 -161 1111 619
<< pwell >>
rect -147 1208 1123 1332
rect -147 788 -59 1208
rect 1035 788 1123 1208
<< pdiff >>
rect 61 373 73 441
rect 579 373 591 441
rect 61 361 111 373
rect 61 327 69 361
rect 103 327 111 361
rect 61 315 111 327
rect 541 361 591 373
rect 541 327 549 361
rect 583 327 591 361
rect 541 315 591 327
rect 61 97 111 109
rect 61 63 69 97
rect 103 63 111 97
rect 61 51 111 63
rect 541 97 591 109
rect 541 63 549 97
rect 583 63 591 97
rect 541 51 591 63
rect 61 -17 73 51
rect 579 -17 591 51
<< pdiffc >>
rect 69 327 103 361
rect 549 327 583 361
rect 69 63 103 97
rect 549 63 583 97
<< psubdiff >>
rect -121 1269 1097 1306
rect -121 1235 -87 1269
rect -53 1235 -19 1269
rect 15 1235 49 1269
rect 83 1235 117 1269
rect 151 1235 185 1269
rect 219 1235 253 1269
rect 287 1235 321 1269
rect 355 1235 389 1269
rect 423 1235 457 1269
rect 491 1235 525 1269
rect 559 1235 593 1269
rect 627 1235 661 1269
rect 695 1235 729 1269
rect 763 1235 797 1269
rect 831 1235 865 1269
rect 899 1235 933 1269
rect 967 1236 1097 1269
rect 967 1235 1062 1236
rect -121 1234 1062 1235
rect -121 1154 -85 1234
rect 1061 1202 1062 1234
rect 1096 1202 1097 1236
rect 1061 1168 1097 1202
rect -121 1120 -120 1154
rect -86 1120 -85 1154
rect -121 1086 -85 1120
rect -121 1052 -120 1086
rect -86 1052 -85 1086
rect -121 1018 -85 1052
rect -121 984 -120 1018
rect -86 984 -85 1018
rect -121 950 -85 984
rect -121 916 -120 950
rect -86 916 -85 950
rect -121 882 -85 916
rect 1061 1134 1062 1168
rect 1096 1134 1097 1168
rect 1061 1100 1097 1134
rect 1061 1066 1062 1100
rect 1096 1066 1097 1100
rect 1061 1032 1097 1066
rect 1061 998 1062 1032
rect 1096 998 1097 1032
rect 1061 964 1097 998
rect 1061 930 1062 964
rect 1096 930 1097 964
rect -121 848 -120 882
rect -86 848 -85 882
rect -121 814 -85 848
rect 1061 896 1097 930
rect 1061 862 1062 896
rect 1096 862 1097 896
rect 1061 814 1097 862
<< nsubdiff >>
rect -47 559 -13 583
rect -47 487 -13 525
rect -47 415 -13 453
rect 665 559 699 583
rect 665 487 699 525
rect -47 343 -13 381
rect 665 415 699 453
rect 665 343 699 381
rect -47 271 -13 309
rect -47 199 -13 237
rect 665 271 699 309
rect 665 199 699 237
rect -47 127 -13 165
rect 665 127 699 165
rect -47 55 -13 93
rect -47 -17 -13 21
rect 665 55 699 93
rect 665 -17 699 21
rect -47 -91 -13 -51
rect 665 -91 699 -51
rect 1041 559 1075 583
rect 1041 487 1075 525
rect 1041 415 1075 453
rect 1041 343 1075 381
rect 1041 271 1075 309
rect 1041 199 1075 237
rect 1041 127 1075 165
rect 1041 55 1075 93
rect 1041 -17 1075 21
rect 1041 -91 1075 -51
rect -47 -125 -23 -91
rect 11 -125 46 -91
rect 80 -125 115 -91
rect 149 -125 184 -91
rect 218 -125 253 -91
rect 287 -125 322 -91
rect 356 -125 391 -91
rect 425 -125 460 -91
rect 494 -125 529 -91
rect 563 -125 598 -91
rect 632 -125 667 -91
rect 701 -125 737 -91
rect 771 -125 807 -91
rect 841 -125 877 -91
rect 911 -125 947 -91
rect 981 -125 1017 -91
rect 1051 -125 1075 -91
<< psubdiffcont >>
rect -87 1235 -53 1269
rect -19 1235 15 1269
rect 49 1235 83 1269
rect 117 1235 151 1269
rect 185 1235 219 1269
rect 253 1235 287 1269
rect 321 1235 355 1269
rect 389 1235 423 1269
rect 457 1235 491 1269
rect 525 1235 559 1269
rect 593 1235 627 1269
rect 661 1235 695 1269
rect 729 1235 763 1269
rect 797 1235 831 1269
rect 865 1235 899 1269
rect 933 1235 967 1269
rect 1062 1202 1096 1236
rect -120 1120 -86 1154
rect -120 1052 -86 1086
rect -120 984 -86 1018
rect -120 916 -86 950
rect 1062 1134 1096 1168
rect 1062 1066 1096 1100
rect 1062 998 1096 1032
rect 1062 930 1096 964
rect -120 848 -86 882
rect 1062 862 1096 896
<< nsubdiffcont >>
rect -47 525 -13 559
rect -47 453 -13 487
rect 665 525 699 559
rect 665 453 699 487
rect -47 381 -13 415
rect -47 309 -13 343
rect 665 381 699 415
rect 665 309 699 343
rect -47 237 -13 271
rect 665 237 699 271
rect -47 165 -13 199
rect -47 93 -13 127
rect 665 165 699 199
rect -47 21 -13 55
rect 665 93 699 127
rect 665 21 699 55
rect -47 -51 -13 -17
rect 665 -51 699 -17
rect 1041 525 1075 559
rect 1041 453 1075 487
rect 1041 381 1075 415
rect 1041 309 1075 343
rect 1041 237 1075 271
rect 1041 165 1075 199
rect 1041 93 1075 127
rect 1041 21 1075 55
rect 1041 -51 1075 -17
rect -23 -125 11 -91
rect 46 -125 80 -91
rect 115 -125 149 -91
rect 184 -125 218 -91
rect 253 -125 287 -91
rect 322 -125 356 -91
rect 391 -125 425 -91
rect 460 -125 494 -91
rect 529 -125 563 -91
rect 598 -125 632 -91
rect 667 -125 701 -91
rect 737 -125 771 -91
rect 807 -125 841 -91
rect 877 -125 911 -91
rect 947 -125 981 -91
rect 1017 -125 1051 -91
<< poly >>
rect 806 1161 842 1167
rect 898 1161 934 1167
rect 42 868 142 909
rect 198 868 298 909
rect 42 802 298 868
rect 354 868 454 909
rect 510 868 610 909
rect 806 868 934 909
rect 354 802 610 868
rect 685 852 934 868
rect 685 818 701 852
rect 735 818 769 852
rect 803 818 934 852
rect 685 802 934 818
rect 42 784 142 802
rect 42 750 69 784
rect 103 750 142 784
rect 42 716 142 750
rect 42 682 69 716
rect 103 682 142 716
rect 42 666 142 682
rect 510 784 610 802
rect 510 750 549 784
rect 583 750 610 784
rect 510 716 610 750
rect 510 682 549 716
rect 583 682 610 716
rect 510 666 610 682
rect 806 609 934 802
rect 126 283 526 305
rect 126 249 169 283
rect 203 249 237 283
rect 271 249 305 283
rect 339 249 526 283
rect 126 233 526 249
rect 126 175 526 191
rect 126 141 313 175
rect 347 141 381 175
rect 415 141 449 175
rect 483 141 526 175
rect 126 119 526 141
<< polycont >>
rect 701 818 735 852
rect 769 818 803 852
rect 69 750 103 784
rect 69 682 103 716
rect 549 750 583 784
rect 549 682 583 716
rect 169 249 203 283
rect 237 249 271 283
rect 305 249 339 283
rect 313 141 347 175
rect 381 141 415 175
rect 449 141 483 175
<< locali >>
rect -121 1269 1097 1270
rect -121 1235 -87 1269
rect -53 1235 -19 1269
rect 15 1235 49 1269
rect 83 1235 117 1269
rect 151 1235 185 1269
rect 219 1235 253 1269
rect 287 1235 321 1269
rect 355 1235 389 1269
rect 423 1235 457 1269
rect 491 1235 525 1269
rect 559 1235 593 1269
rect 627 1235 661 1269
rect 695 1235 729 1269
rect 763 1235 797 1269
rect 831 1235 865 1269
rect 899 1235 933 1269
rect 967 1236 1097 1269
rect 967 1235 1062 1236
rect -121 1234 1062 1235
rect -121 1187 -85 1234
rect -121 1120 -120 1187
rect -86 1120 -85 1187
rect 1061 1202 1062 1234
rect 1096 1202 1097 1236
rect 1061 1187 1097 1202
rect -121 1086 -85 1120
rect -121 1052 -120 1086
rect -86 1052 -85 1086
rect -121 1018 -85 1052
rect -121 984 -120 1018
rect -86 984 -85 1018
rect -121 950 -85 984
rect -121 916 -120 950
rect -86 916 -85 950
rect -3 1029 31 1067
rect -3 957 31 995
rect -121 882 -85 916
rect -121 877 -120 882
rect -86 877 -85 882
rect -86 848 -49 877
rect -87 843 -49 848
rect -121 814 -85 843
rect 53 750 69 784
rect 103 750 119 784
rect 53 716 119 750
rect 53 682 69 716
rect 103 682 119 716
rect -47 559 -13 583
rect -47 487 -13 525
rect -47 415 -13 453
rect -47 351 -13 381
rect -47 279 -13 309
rect -47 207 -13 237
rect 51 361 115 461
rect 51 317 69 361
rect 103 317 115 361
rect 51 279 115 317
rect 51 245 69 279
rect 103 245 115 279
rect 51 207 115 245
rect 51 173 69 207
rect 103 173 115 207
rect 51 167 115 173
rect 153 283 263 1139
rect 309 1029 343 1067
rect 309 957 343 995
rect 389 852 499 1139
rect 1061 1134 1062 1187
rect 1096 1134 1097 1187
rect 621 1029 655 1067
rect 621 957 655 995
rect 761 1029 795 1067
rect 761 957 795 995
rect 945 1029 979 1067
rect 945 957 979 995
rect 389 818 701 852
rect 735 818 769 852
rect 803 818 819 852
rect 389 445 499 818
rect 533 750 549 784
rect 583 750 599 784
rect 533 716 599 750
rect 533 682 549 716
rect 583 682 599 716
rect 665 559 699 583
rect 665 487 699 525
rect 853 521 887 937
rect 1061 1100 1097 1134
rect 1061 1066 1062 1100
rect 1096 1066 1097 1100
rect 1061 1032 1097 1066
rect 1061 998 1062 1032
rect 1096 998 1097 1032
rect 1061 964 1097 998
rect 1061 930 1062 964
rect 1096 930 1097 964
rect 1061 896 1097 930
rect 1061 877 1062 896
rect 1024 843 1062 877
rect 1096 843 1097 896
rect 1061 814 1097 843
rect 1041 559 1075 583
rect 389 361 583 445
rect 389 327 549 361
rect 389 311 583 327
rect 665 415 699 453
rect 665 351 699 381
rect 1041 487 1075 525
rect 1041 415 1075 453
rect 1041 351 1075 381
rect 153 249 169 283
rect 203 249 237 283
rect 271 249 305 283
rect 339 249 355 283
rect -47 135 -13 165
rect 153 113 263 249
rect 389 175 499 311
rect 665 279 699 309
rect 297 141 313 175
rect 347 141 381 175
rect 415 141 449 175
rect 483 141 499 175
rect 537 251 599 257
rect 537 217 549 251
rect 583 217 599 251
rect 537 179 599 217
rect 537 145 549 179
rect 583 145 599 179
rect -47 63 -13 93
rect -47 -9 -13 21
rect 69 97 263 113
rect 103 63 263 97
rect 69 -21 263 63
rect 537 107 599 145
rect 537 63 549 107
rect 583 63 599 107
rect 537 -21 599 63
rect 665 207 699 237
rect 665 135 699 165
rect 761 279 795 317
rect 761 207 795 245
rect 761 135 795 173
rect 945 279 979 317
rect 945 207 979 245
rect 945 135 979 173
rect 1041 279 1075 309
rect 1041 207 1075 237
rect 1041 135 1075 165
rect 665 63 699 93
rect 665 -9 699 21
rect -47 -91 -13 -51
rect 665 -91 699 -51
rect 1041 63 1075 93
rect 1041 -9 1075 21
rect 1041 -91 1075 -51
rect -47 -125 -23 -91
rect 11 -125 46 -91
rect 80 -125 115 -91
rect 149 -125 184 -91
rect 218 -125 253 -91
rect 287 -125 322 -91
rect 356 -125 391 -91
rect 425 -125 460 -91
rect 494 -125 529 -91
rect 563 -125 598 -91
rect 632 -125 667 -91
rect 701 -125 737 -91
rect 771 -125 807 -91
rect 841 -125 877 -91
rect 911 -125 947 -91
rect 981 -125 1017 -91
rect 1051 -125 1075 -91
<< viali >>
rect -120 1154 -86 1187
rect -120 1153 -86 1154
rect -3 1067 31 1101
rect -3 995 31 1029
rect -3 923 31 957
rect -121 848 -120 877
rect -120 848 -87 877
rect -121 843 -87 848
rect -49 843 -15 877
rect -47 343 -13 351
rect -47 317 -13 343
rect -47 271 -13 279
rect -47 245 -13 271
rect -47 199 -13 207
rect -47 173 -13 199
rect 69 327 103 351
rect 69 317 103 327
rect 69 245 103 279
rect 69 173 103 207
rect 309 1067 343 1101
rect 309 995 343 1029
rect 309 923 343 957
rect 1062 1168 1096 1187
rect 1062 1153 1096 1168
rect 621 1067 655 1101
rect 621 995 655 1029
rect 621 923 655 957
rect 761 1067 795 1101
rect 761 995 795 1029
rect 761 923 795 957
rect 945 1067 979 1101
rect 945 995 979 1029
rect 945 923 979 957
rect 990 843 1024 877
rect 1062 862 1096 877
rect 1062 843 1096 862
rect 665 343 699 351
rect 665 317 699 343
rect -47 127 -13 135
rect -47 101 -13 127
rect 665 271 699 279
rect 549 217 583 251
rect 549 145 583 179
rect -47 55 -13 63
rect -47 29 -13 55
rect -47 -17 -13 -9
rect -47 -43 -13 -17
rect 549 97 583 107
rect 549 73 583 97
rect 665 245 699 271
rect 665 199 699 207
rect 665 173 699 199
rect 665 127 699 135
rect 665 101 699 127
rect 761 317 795 351
rect 761 245 795 279
rect 761 173 795 207
rect 761 101 795 135
rect 945 317 979 351
rect 945 245 979 279
rect 945 173 979 207
rect 945 101 979 135
rect 1041 343 1075 351
rect 1041 317 1075 343
rect 1041 271 1075 279
rect 1041 245 1075 271
rect 1041 199 1075 207
rect 1041 173 1075 199
rect 1041 127 1075 135
rect 1041 101 1075 127
rect 665 55 699 63
rect 665 29 699 55
rect 665 -17 699 -9
rect 665 -43 699 -17
rect 1041 55 1075 63
rect 1041 29 1075 55
rect 1041 -17 1075 -9
rect 1041 -43 1075 -17
<< metal1 >>
rect -132 1187 1108 1193
rect -132 1153 -120 1187
rect -86 1153 1062 1187
rect 1096 1153 1108 1187
rect -132 1141 1108 1153
rect -133 1101 1111 1113
rect -133 1067 -3 1101
rect 31 1067 309 1101
rect 343 1067 621 1101
rect 655 1067 761 1101
rect 795 1067 945 1101
rect 979 1067 1111 1101
rect -133 1029 1111 1067
rect -133 995 -3 1029
rect 31 995 309 1029
rect 343 995 621 1029
rect 655 995 761 1029
rect 795 995 945 1029
rect 979 995 1111 1029
rect -133 957 1111 995
rect -133 923 -3 957
rect 31 923 309 957
rect 343 923 621 957
rect 655 923 761 957
rect 795 923 945 957
rect 979 923 1111 957
rect -133 911 1111 923
rect -133 877 1111 883
rect -133 843 -121 877
rect -87 843 -49 877
rect -15 843 990 877
rect 1024 843 1062 877
rect 1096 843 1111 877
rect -133 837 1111 843
rect -83 385 1101 587
rect -83 351 1112 357
rect -83 317 -47 351
rect -13 317 69 351
rect 103 317 665 351
rect 699 317 761 351
rect 795 317 945 351
rect 979 317 1041 351
rect 1075 317 1112 351
rect -83 279 1112 317
rect -83 245 -47 279
rect -13 245 69 279
rect 103 251 665 279
rect 103 245 549 251
rect -83 217 549 245
rect 583 245 665 251
rect 699 245 761 279
rect 795 245 945 279
rect 979 245 1041 279
rect 1075 245 1112 279
rect 583 217 1112 245
rect -83 207 1112 217
rect -83 173 -47 207
rect -13 173 69 207
rect 103 179 665 207
rect 103 173 549 179
rect -83 145 549 173
rect 583 173 665 179
rect 699 173 761 207
rect 795 173 945 207
rect 979 173 1041 207
rect 1075 173 1112 207
rect 583 145 1112 173
rect -83 135 1112 145
rect -83 101 -47 135
rect -13 107 665 135
rect -13 101 549 107
rect -83 73 549 101
rect 583 101 665 107
rect 699 101 761 135
rect 795 101 945 135
rect 979 101 1041 135
rect 1075 101 1112 135
rect 583 73 1112 101
rect -83 67 1112 73
tri -84 63 -80 67 ne
rect -80 63 20 67
tri 20 63 24 67 nw
tri 628 63 632 67 ne
rect 632 63 732 67
tri 732 63 736 67 nw
tri 1004 63 1008 67 ne
rect 1008 63 1087 67
tri -80 42 -59 63 ne
rect -59 29 -47 63
rect -13 29 -1 63
tri -1 42 20 63 nw
tri 632 42 653 63 ne
rect -59 -9 -1 29
rect -59 -43 -47 -9
rect -13 -43 -1 -9
rect -59 -137 -1 -43
rect 653 29 665 63
rect 699 29 711 63
tri 711 42 732 63 nw
tri 1008 42 1029 63 ne
rect 653 -9 711 29
rect 653 -43 665 -9
rect 699 -43 711 -9
tri -1 -79 24 -54 sw
tri 629 -79 653 -55 se
rect 653 -79 711 -43
rect 1029 29 1041 63
rect 1075 29 1087 63
tri 1087 42 1112 67 nw
rect 1029 -9 1087 29
rect 1029 -43 1041 -9
rect 1075 -43 1087 -9
tri 1028 -55 1029 -54 se
rect 1029 -55 1087 -43
tri 711 -79 735 -55 sw
tri 1004 -79 1028 -55 se
rect 1028 -79 1087 -55
rect 1029 -137 1087 -79
use DFL1_CDNS_524688791851160  DFL1_CDNS_524688791851160_0
timestamp 1704896540
transform -1 0 591 0 -1 109
box 0 0 1 1
use DFL1_CDNS_524688791851160  DFL1_CDNS_524688791851160_1
timestamp 1704896540
transform -1 0 591 0 -1 373
box 0 0 1 1
use DFL1_CDNS_524688791851160  DFL1_CDNS_524688791851160_2
timestamp 1704896540
transform 1 0 61 0 -1 373
box 0 0 1 1
use DFL1_CDNS_524688791851160  DFL1_CDNS_524688791851160_3
timestamp 1704896540
transform 1 0 61 0 -1 109
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1704896540
transform -1 0 1096 0 1 843
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1704896540
transform 1 0 -121 0 1 843
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1704896540
transform 0 -1 343 -1 0 1101
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_1
timestamp 1704896540
transform 0 -1 31 -1 0 1101
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_2
timestamp 1704896540
transform 0 -1 655 -1 0 1101
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_3
timestamp 1704896540
transform 0 -1 795 -1 0 1101
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_4
timestamp 1704896540
transform 0 -1 979 -1 0 1101
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_0
timestamp 1704896540
transform 1 0 69 0 1 173
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_1
timestamp 1704896540
transform 1 0 549 0 1 73
box 0 0 1 1
use L1M1_CDNS_52468879185306  L1M1_CDNS_52468879185306_0
timestamp 1704896540
transform 1 0 1041 0 -1 351
box 0 0 1 1
use L1M1_CDNS_52468879185306  L1M1_CDNS_52468879185306_1
timestamp 1704896540
transform 1 0 -47 0 -1 351
box 0 0 1 1
use L1M1_CDNS_52468879185306  L1M1_CDNS_52468879185306_2
timestamp 1704896540
transform 1 0 665 0 -1 351
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_0
timestamp 1704896540
transform 1 0 1062 0 -1 1187
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_1
timestamp 1704896540
transform 1 0 -120 0 -1 1187
box 0 0 1 1
use L1M1_CDNS_524688791851055  L1M1_CDNS_524688791851055_0
timestamp 1704896540
transform 0 1 -43 1 0 -125
box -12 -6 46 1120
use L1M1_CDNS_524688791851057  L1M1_CDNS_524688791851057_0
timestamp 1704896540
transform 1 0 761 0 -1 351
box 0 0 1 1
use L1M1_CDNS_524688791851057  L1M1_CDNS_524688791851057_1
timestamp 1704896540
transform 1 0 945 0 -1 351
box 0 0 1 1
use nfet_CDNS_524688791851161  nfet_CDNS_524688791851161_0
timestamp 1704896540
transform 1 0 42 0 -1 1135
box -79 -26 335 226
use nfet_CDNS_524688791851161  nfet_CDNS_524688791851161_1
timestamp 1704896540
transform 1 0 354 0 -1 1135
box -79 -26 335 226
use nfet_CDNS_524688791851162  nfet_CDNS_524688791851162_0
timestamp 1704896540
transform 1 0 806 0 -1 1135
box -79 -26 207 226
use pfet_CDNS_524688791851163  pfet_CDNS_524688791851163_0
timestamp 1704896540
transform -1 0 526 0 -1 441
box -89 -36 489 146
use pfet_CDNS_524688791851163  pfet_CDNS_524688791851163_1
timestamp 1704896540
transform 1 0 126 0 1 -17
box -89 -36 489 146
use pfet_CDNS_524688791851165  pfet_CDNS_524688791851165_0
timestamp 1704896540
transform -1 0 934 0 1 -17
box -89 -36 217 636
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_0
timestamp 1704896540
transform 0 -1 119 -1 0 800
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_1
timestamp 1704896540
transform 0 1 533 -1 0 800
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_0
timestamp 1704896540
transform 0 -1 819 -1 0 868
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_0
timestamp 1704896540
transform 0 1 153 1 0 233
box 0 0 1 1
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_1
timestamp 1704896540
transform 0 -1 499 1 0 125
box 0 0 1 1
<< labels >>
flabel metal1 s -133 837 -103 883 3 FreeSans 200 0 0 0 vnb
port 1 nsew
flabel metal1 s -133 911 -103 1113 3 FreeSans 200 0 0 0 vgnd
port 2 nsew
flabel metal1 s -83 67 -66 357 0 FreeSans 200 0 0 0 vpwr_ka
port 3 nsew
flabel locali s 853 587 887 911 3 FreeSans 200 0 0 0 out_n
port 5 nsew
flabel locali s 53 682 119 784 0 FreeSans 200 0 0 0 in_h
port 6 nsew
flabel locali s 533 682 599 784 0 FreeSans 200 0 0 0 in_h_n
port 7 nsew
<< properties >>
string GDS_END 79605024
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 79593472
string path 17.050 -2.525 17.050 15.225 
<< end >>
