magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< poly >>
rect -50 131 0 160
rect -50 97 -34 131
rect -50 63 0 97
rect -50 29 -34 63
rect -50 0 0 29
rect -50 -125 0 -96
rect -50 -159 -34 -125
rect -50 -193 0 -159
rect -50 -227 -34 -193
rect -50 -256 0 -227
<< polycont >>
rect -34 97 0 131
rect -34 29 0 63
rect -34 -159 0 -125
rect -34 -227 0 -193
<< npolyres >>
rect 0 0 1232 160
rect 1072 -96 1232 0
rect 0 -256 1232 -96
<< locali >>
rect -34 131 0 147
rect -34 63 0 97
rect -34 13 0 29
rect -34 -125 0 -109
rect -34 -193 0 -159
rect -34 -243 0 -227
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_0
timestamp 1704896540
transform 1 0 -50 0 1 -243
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_1
timestamp 1704896540
transform 1 0 -50 0 1 13
box 0 0 1 1
<< properties >>
string GDS_END 90829736
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 90828996
<< end >>
