magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -36 -36 89 636
<< pdiff >>
rect 0 522 53 600
rect 0 488 11 522
rect 45 488 53 522
rect 0 454 53 488
rect 0 420 11 454
rect 45 420 53 454
rect 0 386 53 420
rect 0 352 11 386
rect 45 352 53 386
rect 0 318 53 352
rect 0 284 11 318
rect 45 284 53 318
rect 0 250 53 284
rect 0 216 11 250
rect 45 216 53 250
rect 0 182 53 216
rect 0 148 11 182
rect 45 148 53 182
rect 0 114 53 148
rect 0 80 11 114
rect 45 80 53 114
rect 0 46 53 80
rect 0 12 11 46
rect 45 12 53 46
rect 0 0 53 12
<< pdiffc >>
rect 11 488 45 522
rect 11 420 45 454
rect 11 352 45 386
rect 11 284 45 318
rect 11 216 45 250
rect 11 148 45 182
rect 11 80 45 114
rect 11 12 45 46
<< locali >>
rect 11 522 45 538
rect 11 454 45 488
rect 11 386 45 420
rect 11 318 45 352
rect 11 250 45 284
rect 11 182 45 216
rect 11 114 45 148
rect 11 46 45 80
rect 11 -4 45 12
<< properties >>
string GDS_END 7602338
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 7601566
<< end >>
