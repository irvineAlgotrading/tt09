magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -38 261 406 582
<< pwell >>
rect 1 21 367 157
rect 29 -17 63 21
<< locali >>
rect 212 406 249 487
rect 212 371 345 406
rect 85 149 157 265
rect 277 165 345 371
rect 208 131 345 165
rect 208 51 249 131
<< obsli1 >>
rect 0 527 368 561
rect 17 333 71 487
rect 105 371 171 527
rect 283 442 350 527
rect 17 299 243 333
rect 17 117 51 299
rect 193 199 243 299
rect 17 51 69 117
rect 111 17 166 113
rect 283 17 350 97
rect 0 -17 368 17
<< metal1 >>
rect 0 496 368 592
rect 0 -48 368 48
<< labels >>
rlabel locali s 85 149 157 265 6 A
port 1 nsew signal input
rlabel metal1 s 0 -48 368 48 8 VGND
port 2 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 3 nsew ground bidirectional
rlabel pwell s 1 21 367 157 6 VNB
port 3 nsew ground bidirectional
rlabel nwell s -38 261 406 582 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 496 368 592 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 208 51 249 131 6 X
port 6 nsew signal output
rlabel locali s 208 131 345 165 6 X
port 6 nsew signal output
rlabel locali s 277 165 345 371 6 X
port 6 nsew signal output
rlabel locali s 212 371 345 406 6 X
port 6 nsew signal output
rlabel locali s 212 406 249 487 6 X
port 6 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 368 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3193860
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3189314
<< end >>
