magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -89 -36 205 636
<< pmos >>
rect 0 0 30 600
rect 86 0 116 600
<< pdiff >>
rect -50 0 0 600
rect 116 0 166 600
<< poly >>
rect 0 600 30 626
rect 0 -26 30 0
rect 86 600 116 626
rect 86 -26 116 0
<< locali >>
rect -45 -4 -11 538
rect 41 -4 75 538
rect 127 -4 161 538
use hvDFL1sd2_CDNS_52468879185138  hvDFL1sd2_CDNS_52468879185138_0
timestamp 1704896540
transform 1 0 30 0 1 0
box -36 -36 92 636
use hvDFL1sd_CDNS_52468879185135  hvDFL1sd_CDNS_52468879185135_0
timestamp 1704896540
transform -1 0 0 0 1 0
box -36 -36 89 636
use hvDFL1sd_CDNS_52468879185135  hvDFL1sd_CDNS_52468879185135_1
timestamp 1704896540
transform 1 0 116 0 1 0
box -36 -36 89 636
<< labels >>
flabel comment s -28 267 -28 267 0 FreeSans 300 0 0 0 S
flabel comment s 58 267 58 267 0 FreeSans 300 0 0 0 D
flabel comment s 144 267 144 267 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 97511368
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 97509978
<< end >>
