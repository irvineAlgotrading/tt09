magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< pwell >>
rect -68 -26 668 92
<< ndiff >>
rect -42 50 0 66
rect -42 16 -34 50
rect -42 0 0 16
rect 600 50 642 66
rect 634 16 642 50
rect 600 0 642 16
<< ndiffc >>
rect -34 16 0 50
rect 600 16 634 50
<< ndiffres >>
rect 0 0 600 66
<< locali >>
rect -34 50 0 66
rect -34 0 0 16
rect 600 50 634 66
rect 600 0 634 16
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_0
timestamp 1704896540
transform -1 0 8 0 1 4
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_1
timestamp 1704896540
transform 1 0 592 0 1 4
box 0 0 1 1
<< properties >>
string GDS_END 86205306
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86204804
<< end >>
