magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect 8943 0 12298 701
<< pwell >>
rect 9013 1020 12249 1106
rect 9024 806 12224 1020
<< mvnmos >>
rect 9103 832 9223 972
rect 9279 832 9399 972
rect 9455 832 9575 972
rect 9744 832 9864 972
rect 9920 832 10040 972
rect 10096 832 10216 972
rect 10272 832 10392 972
rect 10573 832 10693 972
rect 10749 832 10869 972
rect 10925 832 11045 972
rect 11211 832 11331 972
rect 11387 832 11507 972
rect 11563 832 11683 972
rect 11849 832 11969 972
rect 12025 832 12145 972
<< mvpmos >>
rect 9103 434 9223 634
rect 9279 434 9399 634
rect 9455 434 9575 634
rect 9744 434 9864 634
rect 9920 434 10040 634
rect 10096 434 10216 634
rect 10272 434 10392 634
rect 10573 434 10693 634
rect 10749 434 10869 634
rect 10925 434 11045 634
rect 11211 434 11331 634
rect 11387 434 11507 634
rect 11563 434 11683 634
rect 11849 434 11969 634
rect 12025 434 12145 634
rect 9103 166 9223 366
rect 9279 166 9399 366
rect 9455 166 9575 366
rect 9744 166 9864 366
rect 9920 166 10040 366
rect 10096 166 10216 366
rect 10272 166 10392 366
rect 10573 166 10693 366
rect 10749 166 10869 366
rect 10925 166 11045 366
rect 11211 166 11331 366
rect 11387 166 11507 366
rect 11563 166 11683 366
rect 11849 166 11969 366
rect 12025 166 12145 366
<< mvndiff >>
rect 9050 946 9103 972
rect 9050 912 9058 946
rect 9092 912 9103 946
rect 9050 878 9103 912
rect 9050 844 9058 878
rect 9092 844 9103 878
rect 9050 832 9103 844
rect 9223 946 9279 972
rect 9223 912 9234 946
rect 9268 912 9279 946
rect 9223 878 9279 912
rect 9223 844 9234 878
rect 9268 844 9279 878
rect 9223 832 9279 844
rect 9399 946 9455 972
rect 9399 912 9410 946
rect 9444 912 9455 946
rect 9399 878 9455 912
rect 9399 844 9410 878
rect 9444 844 9455 878
rect 9399 832 9455 844
rect 9575 946 9631 972
rect 9575 912 9586 946
rect 9620 912 9631 946
rect 9575 878 9631 912
rect 9575 844 9586 878
rect 9620 844 9631 878
rect 9575 832 9631 844
rect 9691 946 9744 972
rect 9691 912 9699 946
rect 9733 912 9744 946
rect 9691 878 9744 912
rect 9691 844 9699 878
rect 9733 844 9744 878
rect 9691 832 9744 844
rect 9864 832 9920 972
rect 10040 946 10096 972
rect 10040 912 10051 946
rect 10085 912 10096 946
rect 10040 878 10096 912
rect 10040 844 10051 878
rect 10085 844 10096 878
rect 10040 832 10096 844
rect 10216 832 10272 972
rect 10392 946 10445 972
rect 10392 912 10403 946
rect 10437 912 10445 946
rect 10392 878 10445 912
rect 10392 844 10403 878
rect 10437 844 10445 878
rect 10392 832 10445 844
rect 10520 946 10573 972
rect 10520 912 10528 946
rect 10562 912 10573 946
rect 10520 878 10573 912
rect 10520 844 10528 878
rect 10562 844 10573 878
rect 10520 832 10573 844
rect 10693 946 10749 972
rect 10693 912 10704 946
rect 10738 912 10749 946
rect 10693 878 10749 912
rect 10693 844 10704 878
rect 10738 844 10749 878
rect 10693 832 10749 844
rect 10869 832 10925 972
rect 11045 946 11098 972
rect 11045 912 11056 946
rect 11090 912 11098 946
rect 11045 878 11098 912
rect 11045 844 11056 878
rect 11090 844 11098 878
rect 11045 832 11098 844
rect 11158 946 11211 972
rect 11158 912 11166 946
rect 11200 912 11211 946
rect 11158 878 11211 912
rect 11158 844 11166 878
rect 11200 844 11211 878
rect 11158 832 11211 844
rect 11331 832 11387 972
rect 11507 946 11563 972
rect 11507 912 11518 946
rect 11552 912 11563 946
rect 11507 878 11563 912
rect 11507 844 11518 878
rect 11552 844 11563 878
rect 11507 832 11563 844
rect 11683 946 11736 972
rect 11683 912 11694 946
rect 11728 912 11736 946
rect 11683 878 11736 912
rect 11683 844 11694 878
rect 11728 844 11736 878
rect 11683 832 11736 844
rect 11796 946 11849 972
rect 11796 912 11804 946
rect 11838 912 11849 946
rect 11796 878 11849 912
rect 11796 844 11804 878
rect 11838 844 11849 878
rect 11796 832 11849 844
rect 11969 832 12025 972
rect 12145 946 12198 972
rect 12145 912 12156 946
rect 12190 912 12198 946
rect 12145 878 12198 912
rect 12145 844 12156 878
rect 12190 844 12198 878
rect 12145 832 12198 844
<< mvpdiff >>
rect 9050 616 9103 634
rect 9050 582 9058 616
rect 9092 582 9103 616
rect 9050 548 9103 582
rect 9050 514 9058 548
rect 9092 514 9103 548
rect 9050 480 9103 514
rect 9050 446 9058 480
rect 9092 446 9103 480
rect 9050 434 9103 446
rect 9223 616 9279 634
rect 9223 582 9234 616
rect 9268 582 9279 616
rect 9223 548 9279 582
rect 9223 514 9234 548
rect 9268 514 9279 548
rect 9223 480 9279 514
rect 9223 446 9234 480
rect 9268 446 9279 480
rect 9223 434 9279 446
rect 9399 548 9455 634
rect 9399 514 9410 548
rect 9444 514 9455 548
rect 9399 480 9455 514
rect 9399 446 9410 480
rect 9444 446 9455 480
rect 9399 434 9455 446
rect 9575 616 9628 634
rect 9575 582 9586 616
rect 9620 582 9628 616
rect 9575 548 9628 582
rect 9575 514 9586 548
rect 9620 514 9628 548
rect 9575 480 9628 514
rect 9575 446 9586 480
rect 9620 446 9628 480
rect 9575 434 9628 446
rect 9691 616 9744 634
rect 9691 582 9699 616
rect 9733 582 9744 616
rect 9691 548 9744 582
rect 9691 514 9699 548
rect 9733 514 9744 548
rect 9691 480 9744 514
rect 9691 446 9699 480
rect 9733 446 9744 480
rect 9691 434 9744 446
rect 9864 616 9920 634
rect 9864 582 9875 616
rect 9909 582 9920 616
rect 9864 548 9920 582
rect 9864 514 9875 548
rect 9909 514 9920 548
rect 9864 480 9920 514
rect 9864 446 9875 480
rect 9909 446 9920 480
rect 9864 434 9920 446
rect 10040 616 10096 634
rect 10040 582 10051 616
rect 10085 582 10096 616
rect 10040 548 10096 582
rect 10040 514 10051 548
rect 10085 514 10096 548
rect 10040 480 10096 514
rect 10040 446 10051 480
rect 10085 446 10096 480
rect 10040 434 10096 446
rect 10216 616 10272 634
rect 10216 582 10227 616
rect 10261 582 10272 616
rect 10216 548 10272 582
rect 10216 514 10227 548
rect 10261 514 10272 548
rect 10216 480 10272 514
rect 10216 446 10227 480
rect 10261 446 10272 480
rect 10216 434 10272 446
rect 10392 616 10445 634
rect 10392 582 10403 616
rect 10437 582 10445 616
rect 10392 548 10445 582
rect 10392 514 10403 548
rect 10437 514 10445 548
rect 10392 480 10445 514
rect 10392 446 10403 480
rect 10437 446 10445 480
rect 10392 434 10445 446
rect 10520 616 10573 634
rect 10520 582 10528 616
rect 10562 582 10573 616
rect 10520 548 10573 582
rect 10520 514 10528 548
rect 10562 514 10573 548
rect 10520 480 10573 514
rect 10520 446 10528 480
rect 10562 446 10573 480
rect 10520 434 10573 446
rect 10693 616 10749 634
rect 10693 582 10704 616
rect 10738 582 10749 616
rect 10693 548 10749 582
rect 10693 514 10704 548
rect 10738 514 10749 548
rect 10693 480 10749 514
rect 10693 446 10704 480
rect 10738 446 10749 480
rect 10693 434 10749 446
rect 10869 616 10925 634
rect 10869 582 10880 616
rect 10914 582 10925 616
rect 10869 548 10925 582
rect 10869 514 10880 548
rect 10914 514 10925 548
rect 10869 480 10925 514
rect 10869 446 10880 480
rect 10914 446 10925 480
rect 10869 434 10925 446
rect 11045 616 11098 634
rect 11045 582 11056 616
rect 11090 582 11098 616
rect 11045 548 11098 582
rect 11045 514 11056 548
rect 11090 514 11098 548
rect 11045 480 11098 514
rect 11045 446 11056 480
rect 11090 446 11098 480
rect 11045 434 11098 446
rect 11158 616 11211 634
rect 11158 582 11166 616
rect 11200 582 11211 616
rect 11158 548 11211 582
rect 11158 514 11166 548
rect 11200 514 11211 548
rect 11158 480 11211 514
rect 11158 446 11166 480
rect 11200 446 11211 480
rect 11158 434 11211 446
rect 11331 616 11387 634
rect 11331 582 11342 616
rect 11376 582 11387 616
rect 11331 548 11387 582
rect 11331 514 11342 548
rect 11376 514 11387 548
rect 11331 480 11387 514
rect 11331 446 11342 480
rect 11376 446 11387 480
rect 11331 434 11387 446
rect 11507 616 11563 634
rect 11507 582 11518 616
rect 11552 582 11563 616
rect 11507 548 11563 582
rect 11507 514 11518 548
rect 11552 514 11563 548
rect 11507 480 11563 514
rect 11507 446 11518 480
rect 11552 446 11563 480
rect 11507 434 11563 446
rect 11683 616 11736 634
rect 11683 582 11694 616
rect 11728 582 11736 616
rect 11683 548 11736 582
rect 11683 514 11694 548
rect 11728 514 11736 548
rect 11683 480 11736 514
rect 11683 446 11694 480
rect 11728 446 11736 480
rect 11683 434 11736 446
rect 11796 616 11849 634
rect 11796 582 11804 616
rect 11838 582 11849 616
rect 11796 548 11849 582
rect 11796 514 11804 548
rect 11838 514 11849 548
rect 11796 480 11849 514
rect 11796 446 11804 480
rect 11838 446 11849 480
rect 11796 434 11849 446
rect 11969 616 12025 634
rect 11969 582 11980 616
rect 12014 582 12025 616
rect 11969 548 12025 582
rect 11969 514 11980 548
rect 12014 514 12025 548
rect 11969 480 12025 514
rect 11969 446 11980 480
rect 12014 446 12025 480
rect 11969 434 12025 446
rect 12145 616 12198 634
rect 12145 582 12156 616
rect 12190 582 12198 616
rect 12145 548 12198 582
rect 12145 514 12156 548
rect 12190 514 12198 548
rect 12145 480 12198 514
rect 12145 446 12156 480
rect 12190 446 12198 480
rect 12145 434 12198 446
rect 9050 354 9103 366
rect 9050 320 9058 354
rect 9092 320 9103 354
rect 9050 286 9103 320
rect 9050 252 9058 286
rect 9092 252 9103 286
rect 9050 218 9103 252
rect 9050 184 9058 218
rect 9092 184 9103 218
rect 9050 166 9103 184
rect 9223 354 9279 366
rect 9223 320 9234 354
rect 9268 320 9279 354
rect 9223 286 9279 320
rect 9223 252 9234 286
rect 9268 252 9279 286
rect 9223 218 9279 252
rect 9223 184 9234 218
rect 9268 184 9279 218
rect 9223 166 9279 184
rect 9399 354 9455 366
rect 9399 320 9410 354
rect 9444 320 9455 354
rect 9399 286 9455 320
rect 9399 252 9410 286
rect 9444 252 9455 286
rect 9399 218 9455 252
rect 9399 184 9410 218
rect 9444 184 9455 218
rect 9399 166 9455 184
rect 9575 354 9628 366
rect 9575 320 9586 354
rect 9620 320 9628 354
rect 9575 286 9628 320
rect 9575 252 9586 286
rect 9620 252 9628 286
rect 9575 218 9628 252
rect 9575 184 9586 218
rect 9620 184 9628 218
rect 9575 166 9628 184
rect 9691 354 9744 366
rect 9691 320 9699 354
rect 9733 320 9744 354
rect 9691 286 9744 320
rect 9691 252 9699 286
rect 9733 252 9744 286
rect 9691 218 9744 252
rect 9691 184 9699 218
rect 9733 184 9744 218
rect 9691 166 9744 184
rect 9864 354 9920 366
rect 9864 320 9875 354
rect 9909 320 9920 354
rect 9864 286 9920 320
rect 9864 252 9875 286
rect 9909 252 9920 286
rect 9864 218 9920 252
rect 9864 184 9875 218
rect 9909 184 9920 218
rect 9864 166 9920 184
rect 10040 354 10096 366
rect 10040 320 10051 354
rect 10085 320 10096 354
rect 10040 286 10096 320
rect 10040 252 10051 286
rect 10085 252 10096 286
rect 10040 218 10096 252
rect 10040 184 10051 218
rect 10085 184 10096 218
rect 10040 166 10096 184
rect 10216 354 10272 366
rect 10216 320 10227 354
rect 10261 320 10272 354
rect 10216 286 10272 320
rect 10216 252 10227 286
rect 10261 252 10272 286
rect 10216 218 10272 252
rect 10216 184 10227 218
rect 10261 184 10272 218
rect 10216 166 10272 184
rect 10392 354 10445 366
rect 10392 320 10403 354
rect 10437 320 10445 354
rect 10392 286 10445 320
rect 10392 252 10403 286
rect 10437 252 10445 286
rect 10392 218 10445 252
rect 10392 184 10403 218
rect 10437 184 10445 218
rect 10392 166 10445 184
rect 10520 354 10573 366
rect 10520 320 10528 354
rect 10562 320 10573 354
rect 10520 286 10573 320
rect 10520 252 10528 286
rect 10562 252 10573 286
rect 10520 218 10573 252
rect 10520 184 10528 218
rect 10562 184 10573 218
rect 10520 166 10573 184
rect 10693 354 10749 366
rect 10693 320 10704 354
rect 10738 320 10749 354
rect 10693 286 10749 320
rect 10693 252 10704 286
rect 10738 252 10749 286
rect 10693 218 10749 252
rect 10693 184 10704 218
rect 10738 184 10749 218
rect 10693 166 10749 184
rect 10869 354 10925 366
rect 10869 320 10880 354
rect 10914 320 10925 354
rect 10869 286 10925 320
rect 10869 252 10880 286
rect 10914 252 10925 286
rect 10869 218 10925 252
rect 10869 184 10880 218
rect 10914 184 10925 218
rect 10869 166 10925 184
rect 11045 354 11098 366
rect 11045 320 11056 354
rect 11090 320 11098 354
rect 11045 286 11098 320
rect 11045 252 11056 286
rect 11090 252 11098 286
rect 11045 218 11098 252
rect 11045 184 11056 218
rect 11090 184 11098 218
rect 11045 166 11098 184
rect 11158 354 11211 366
rect 11158 320 11166 354
rect 11200 320 11211 354
rect 11158 286 11211 320
rect 11158 252 11166 286
rect 11200 252 11211 286
rect 11158 218 11211 252
rect 11158 184 11166 218
rect 11200 184 11211 218
rect 11158 166 11211 184
rect 11331 354 11387 366
rect 11331 320 11342 354
rect 11376 320 11387 354
rect 11331 286 11387 320
rect 11331 252 11342 286
rect 11376 252 11387 286
rect 11331 218 11387 252
rect 11331 184 11342 218
rect 11376 184 11387 218
rect 11331 166 11387 184
rect 11507 354 11563 366
rect 11507 320 11518 354
rect 11552 320 11563 354
rect 11507 286 11563 320
rect 11507 252 11518 286
rect 11552 252 11563 286
rect 11507 218 11563 252
rect 11507 184 11518 218
rect 11552 184 11563 218
rect 11507 166 11563 184
rect 11683 354 11736 366
rect 11683 320 11694 354
rect 11728 320 11736 354
rect 11683 286 11736 320
rect 11683 252 11694 286
rect 11728 252 11736 286
rect 11683 218 11736 252
rect 11683 184 11694 218
rect 11728 184 11736 218
rect 11683 166 11736 184
rect 11796 354 11849 366
rect 11796 320 11804 354
rect 11838 320 11849 354
rect 11796 286 11849 320
rect 11796 252 11804 286
rect 11838 252 11849 286
rect 11796 218 11849 252
rect 11796 184 11804 218
rect 11838 184 11849 218
rect 11796 166 11849 184
rect 11969 354 12025 366
rect 11969 320 11980 354
rect 12014 320 12025 354
rect 11969 286 12025 320
rect 11969 252 11980 286
rect 12014 252 12025 286
rect 11969 218 12025 252
rect 11969 184 11980 218
rect 12014 184 12025 218
rect 11969 166 12025 184
rect 12145 354 12198 366
rect 12145 320 12156 354
rect 12190 320 12198 354
rect 12145 286 12198 320
rect 12145 252 12156 286
rect 12190 252 12198 286
rect 12145 218 12198 252
rect 12145 184 12156 218
rect 12190 184 12198 218
rect 12145 166 12198 184
<< mvndiffc >>
rect 9058 912 9092 946
rect 9058 844 9092 878
rect 9234 912 9268 946
rect 9234 844 9268 878
rect 9410 912 9444 946
rect 9410 844 9444 878
rect 9586 912 9620 946
rect 9586 844 9620 878
rect 9699 912 9733 946
rect 9699 844 9733 878
rect 10051 912 10085 946
rect 10051 844 10085 878
rect 10403 912 10437 946
rect 10403 844 10437 878
rect 10528 912 10562 946
rect 10528 844 10562 878
rect 10704 912 10738 946
rect 10704 844 10738 878
rect 11056 912 11090 946
rect 11056 844 11090 878
rect 11166 912 11200 946
rect 11166 844 11200 878
rect 11518 912 11552 946
rect 11518 844 11552 878
rect 11694 912 11728 946
rect 11694 844 11728 878
rect 11804 912 11838 946
rect 11804 844 11838 878
rect 12156 912 12190 946
rect 12156 844 12190 878
<< mvpdiffc >>
rect 9058 582 9092 616
rect 9058 514 9092 548
rect 9058 446 9092 480
rect 9234 582 9268 616
rect 9234 514 9268 548
rect 9234 446 9268 480
rect 9410 514 9444 548
rect 9410 446 9444 480
rect 9586 582 9620 616
rect 9586 514 9620 548
rect 9586 446 9620 480
rect 9699 582 9733 616
rect 9699 514 9733 548
rect 9699 446 9733 480
rect 9875 582 9909 616
rect 9875 514 9909 548
rect 9875 446 9909 480
rect 10051 582 10085 616
rect 10051 514 10085 548
rect 10051 446 10085 480
rect 10227 582 10261 616
rect 10227 514 10261 548
rect 10227 446 10261 480
rect 10403 582 10437 616
rect 10403 514 10437 548
rect 10403 446 10437 480
rect 10528 582 10562 616
rect 10528 514 10562 548
rect 10528 446 10562 480
rect 10704 582 10738 616
rect 10704 514 10738 548
rect 10704 446 10738 480
rect 10880 582 10914 616
rect 10880 514 10914 548
rect 10880 446 10914 480
rect 11056 582 11090 616
rect 11056 514 11090 548
rect 11056 446 11090 480
rect 11166 582 11200 616
rect 11166 514 11200 548
rect 11166 446 11200 480
rect 11342 582 11376 616
rect 11342 514 11376 548
rect 11342 446 11376 480
rect 11518 582 11552 616
rect 11518 514 11552 548
rect 11518 446 11552 480
rect 11694 582 11728 616
rect 11694 514 11728 548
rect 11694 446 11728 480
rect 11804 582 11838 616
rect 11804 514 11838 548
rect 11804 446 11838 480
rect 11980 582 12014 616
rect 11980 514 12014 548
rect 11980 446 12014 480
rect 12156 582 12190 616
rect 12156 514 12190 548
rect 12156 446 12190 480
rect 9058 320 9092 354
rect 9058 252 9092 286
rect 9058 184 9092 218
rect 9234 320 9268 354
rect 9234 252 9268 286
rect 9234 184 9268 218
rect 9410 320 9444 354
rect 9410 252 9444 286
rect 9410 184 9444 218
rect 9586 320 9620 354
rect 9586 252 9620 286
rect 9586 184 9620 218
rect 9699 320 9733 354
rect 9699 252 9733 286
rect 9699 184 9733 218
rect 9875 320 9909 354
rect 9875 252 9909 286
rect 9875 184 9909 218
rect 10051 320 10085 354
rect 10051 252 10085 286
rect 10051 184 10085 218
rect 10227 320 10261 354
rect 10227 252 10261 286
rect 10227 184 10261 218
rect 10403 320 10437 354
rect 10403 252 10437 286
rect 10403 184 10437 218
rect 10528 320 10562 354
rect 10528 252 10562 286
rect 10528 184 10562 218
rect 10704 320 10738 354
rect 10704 252 10738 286
rect 10704 184 10738 218
rect 10880 320 10914 354
rect 10880 252 10914 286
rect 10880 184 10914 218
rect 11056 320 11090 354
rect 11056 252 11090 286
rect 11056 184 11090 218
rect 11166 320 11200 354
rect 11166 252 11200 286
rect 11166 184 11200 218
rect 11342 320 11376 354
rect 11342 252 11376 286
rect 11342 184 11376 218
rect 11518 320 11552 354
rect 11518 252 11552 286
rect 11518 184 11552 218
rect 11694 320 11728 354
rect 11694 252 11728 286
rect 11694 184 11728 218
rect 11804 320 11838 354
rect 11804 252 11838 286
rect 11804 184 11838 218
rect 11980 320 12014 354
rect 11980 252 12014 286
rect 11980 184 12014 218
rect 12156 320 12190 354
rect 12156 252 12190 286
rect 12156 184 12190 218
<< mvpsubdiff >>
rect 9039 1046 9063 1080
rect 9097 1046 9131 1080
rect 9165 1046 9199 1080
rect 9233 1046 9267 1080
rect 9301 1046 9335 1080
rect 9369 1046 9403 1080
rect 9437 1046 9471 1080
rect 9505 1046 9539 1080
rect 9573 1046 9607 1080
rect 9641 1046 9675 1080
rect 9709 1046 9743 1080
rect 9777 1046 9811 1080
rect 9845 1046 9879 1080
rect 9913 1046 9947 1080
rect 9981 1046 10015 1080
rect 10049 1046 10083 1080
rect 10117 1046 10151 1080
rect 10185 1046 10219 1080
rect 10253 1046 10287 1080
rect 10321 1046 10355 1080
rect 10389 1046 10423 1080
rect 10457 1046 10491 1080
rect 10525 1046 10559 1080
rect 10593 1046 10627 1080
rect 10661 1046 10695 1080
rect 10729 1046 10763 1080
rect 10797 1046 10831 1080
rect 10865 1046 10899 1080
rect 10933 1046 10967 1080
rect 11001 1046 11035 1080
rect 11069 1046 11103 1080
rect 11137 1046 11171 1080
rect 11205 1046 11239 1080
rect 11273 1046 11307 1080
rect 11341 1046 11375 1080
rect 11409 1046 11443 1080
rect 11477 1046 11511 1080
rect 11545 1046 11579 1080
rect 11613 1046 11647 1080
rect 11681 1046 11715 1080
rect 11749 1046 11783 1080
rect 11817 1046 11851 1080
rect 11885 1046 11919 1080
rect 11953 1046 11987 1080
rect 12021 1046 12055 1080
rect 12089 1046 12123 1080
rect 12157 1046 12223 1080
<< mvnsubdiff >>
rect 9053 66 9077 100
rect 9111 66 9145 100
rect 9179 66 9213 100
rect 9247 66 9281 100
rect 9315 66 9349 100
rect 9383 66 9417 100
rect 9451 66 9485 100
rect 9519 66 9553 100
rect 9587 66 9621 100
rect 9655 66 9689 100
rect 9723 66 9757 100
rect 9791 66 9825 100
rect 9859 66 9893 100
rect 9927 66 9961 100
rect 9995 66 10029 100
rect 10063 66 10097 100
rect 10131 66 10165 100
rect 10199 66 10233 100
rect 10267 66 10301 100
rect 10335 66 10369 100
rect 10403 66 10437 100
rect 10471 66 10505 100
rect 10539 66 10573 100
rect 10607 66 10641 100
rect 10675 66 10709 100
rect 10743 66 10777 100
rect 10811 66 10845 100
rect 10879 66 10913 100
rect 10947 66 10981 100
rect 11015 66 11049 100
rect 11083 66 11117 100
rect 11151 66 11185 100
rect 11219 66 11253 100
rect 11287 66 11321 100
rect 11355 66 11389 100
rect 11423 66 11457 100
rect 11491 66 11525 100
rect 11559 66 11593 100
rect 11627 66 11661 100
rect 11695 66 11729 100
rect 11763 66 11797 100
rect 11831 66 11865 100
rect 11899 66 11933 100
rect 11967 66 12001 100
rect 12035 66 12069 100
rect 12103 66 12137 100
rect 12171 66 12198 100
<< mvpsubdiffcont >>
rect 9063 1046 9097 1080
rect 9131 1046 9165 1080
rect 9199 1046 9233 1080
rect 9267 1046 9301 1080
rect 9335 1046 9369 1080
rect 9403 1046 9437 1080
rect 9471 1046 9505 1080
rect 9539 1046 9573 1080
rect 9607 1046 9641 1080
rect 9675 1046 9709 1080
rect 9743 1046 9777 1080
rect 9811 1046 9845 1080
rect 9879 1046 9913 1080
rect 9947 1046 9981 1080
rect 10015 1046 10049 1080
rect 10083 1046 10117 1080
rect 10151 1046 10185 1080
rect 10219 1046 10253 1080
rect 10287 1046 10321 1080
rect 10355 1046 10389 1080
rect 10423 1046 10457 1080
rect 10491 1046 10525 1080
rect 10559 1046 10593 1080
rect 10627 1046 10661 1080
rect 10695 1046 10729 1080
rect 10763 1046 10797 1080
rect 10831 1046 10865 1080
rect 10899 1046 10933 1080
rect 10967 1046 11001 1080
rect 11035 1046 11069 1080
rect 11103 1046 11137 1080
rect 11171 1046 11205 1080
rect 11239 1046 11273 1080
rect 11307 1046 11341 1080
rect 11375 1046 11409 1080
rect 11443 1046 11477 1080
rect 11511 1046 11545 1080
rect 11579 1046 11613 1080
rect 11647 1046 11681 1080
rect 11715 1046 11749 1080
rect 11783 1046 11817 1080
rect 11851 1046 11885 1080
rect 11919 1046 11953 1080
rect 11987 1046 12021 1080
rect 12055 1046 12089 1080
rect 12123 1046 12157 1080
<< mvnsubdiffcont >>
rect 9077 66 9111 100
rect 9145 66 9179 100
rect 9213 66 9247 100
rect 9281 66 9315 100
rect 9349 66 9383 100
rect 9417 66 9451 100
rect 9485 66 9519 100
rect 9553 66 9587 100
rect 9621 66 9655 100
rect 9689 66 9723 100
rect 9757 66 9791 100
rect 9825 66 9859 100
rect 9893 66 9927 100
rect 9961 66 9995 100
rect 10029 66 10063 100
rect 10097 66 10131 100
rect 10165 66 10199 100
rect 10233 66 10267 100
rect 10301 66 10335 100
rect 10369 66 10403 100
rect 10437 66 10471 100
rect 10505 66 10539 100
rect 10573 66 10607 100
rect 10641 66 10675 100
rect 10709 66 10743 100
rect 10777 66 10811 100
rect 10845 66 10879 100
rect 10913 66 10947 100
rect 10981 66 11015 100
rect 11049 66 11083 100
rect 11117 66 11151 100
rect 11185 66 11219 100
rect 11253 66 11287 100
rect 11321 66 11355 100
rect 11389 66 11423 100
rect 11457 66 11491 100
rect 11525 66 11559 100
rect 11593 66 11627 100
rect 11661 66 11695 100
rect 11729 66 11763 100
rect 11797 66 11831 100
rect 11865 66 11899 100
rect 11933 66 11967 100
rect 12001 66 12035 100
rect 12069 66 12103 100
rect 12137 66 12171 100
<< poly >>
rect 9103 972 9223 998
rect 9279 972 9399 998
rect 9455 972 9575 998
rect 9744 972 9864 998
rect 9920 972 10040 998
rect 10096 972 10216 998
rect 10272 972 10392 998
rect 10573 972 10693 998
rect 10749 972 10869 998
rect 10925 972 11045 998
rect 11211 972 11331 998
rect 11387 972 11507 998
rect 11563 972 11683 998
rect 11849 972 11969 998
rect 12025 972 12145 998
rect 9103 784 9223 832
rect 9103 750 9145 784
rect 9179 750 9223 784
rect 9103 716 9223 750
rect 9103 682 9145 716
rect 9179 682 9223 716
rect 9103 634 9223 682
rect 9279 784 9399 832
rect 9279 750 9322 784
rect 9356 750 9399 784
rect 9279 716 9399 750
rect 9279 682 9322 716
rect 9356 682 9399 716
rect 9279 634 9399 682
rect 9455 784 9575 832
rect 9455 750 9500 784
rect 9534 750 9575 784
rect 9455 716 9575 750
rect 9455 682 9500 716
rect 9534 682 9575 716
rect 9455 634 9575 682
rect 9744 784 9864 832
rect 9744 750 9789 784
rect 9823 750 9864 784
rect 9744 716 9864 750
rect 9744 682 9789 716
rect 9823 682 9864 716
rect 9744 634 9864 682
rect 9920 784 10040 832
rect 9920 750 9960 784
rect 9994 750 10040 784
rect 9920 716 10040 750
rect 9920 682 9960 716
rect 9994 682 10040 716
rect 9920 634 10040 682
rect 10096 784 10216 832
rect 10096 750 10142 784
rect 10176 750 10216 784
rect 10096 716 10216 750
rect 10096 682 10142 716
rect 10176 682 10216 716
rect 10096 634 10216 682
rect 10272 784 10392 832
rect 10272 750 10313 784
rect 10347 750 10392 784
rect 10272 716 10392 750
rect 10272 682 10313 716
rect 10347 682 10392 716
rect 10272 634 10392 682
rect 10573 784 10693 832
rect 10573 750 10615 784
rect 10649 750 10693 784
rect 10573 716 10693 750
rect 10573 682 10615 716
rect 10649 682 10693 716
rect 10573 634 10693 682
rect 10749 784 10869 832
rect 10749 750 10795 784
rect 10829 750 10869 784
rect 10749 716 10869 750
rect 10749 682 10795 716
rect 10829 682 10869 716
rect 10749 634 10869 682
rect 10925 784 11045 832
rect 10925 750 10966 784
rect 11000 750 11045 784
rect 10925 716 11045 750
rect 10925 682 10966 716
rect 11000 682 11045 716
rect 10925 634 11045 682
rect 11211 784 11331 832
rect 11211 750 11256 784
rect 11290 750 11331 784
rect 11211 716 11331 750
rect 11211 682 11256 716
rect 11290 682 11331 716
rect 11211 634 11331 682
rect 11387 784 11507 832
rect 11387 750 11427 784
rect 11461 750 11507 784
rect 11387 716 11507 750
rect 11387 682 11427 716
rect 11461 682 11507 716
rect 11387 634 11507 682
rect 11563 784 11683 832
rect 11563 750 11607 784
rect 11641 750 11683 784
rect 11563 716 11683 750
rect 11563 682 11607 716
rect 11641 682 11683 716
rect 11563 634 11683 682
rect 11849 784 11969 832
rect 11849 750 11894 784
rect 11928 750 11969 784
rect 11849 716 11969 750
rect 11849 682 11894 716
rect 11928 682 11969 716
rect 11849 634 11969 682
rect 12025 784 12145 832
rect 12025 750 12065 784
rect 12099 750 12145 784
rect 12025 716 12145 750
rect 12025 682 12065 716
rect 12099 682 12145 716
rect 12025 634 12145 682
rect 9103 366 9223 434
rect 9279 366 9399 434
rect 9455 366 9575 434
rect 9744 366 9864 434
rect 9920 366 10040 434
rect 10096 366 10216 434
rect 10272 366 10392 434
rect 10573 366 10693 434
rect 10749 366 10869 434
rect 10925 366 11045 434
rect 11211 366 11331 434
rect 11387 366 11507 434
rect 11563 366 11683 434
rect 11849 366 11969 434
rect 12025 366 12145 434
rect 9103 140 9223 166
rect 9279 140 9399 166
rect 9455 140 9575 166
rect 9744 140 9864 166
rect 9920 140 10040 166
rect 10096 140 10216 166
rect 10272 140 10392 166
rect 10573 140 10693 166
rect 10749 140 10869 166
rect 10925 140 11045 166
rect 11211 140 11331 166
rect 11387 140 11507 166
rect 11563 140 11683 166
rect 11849 140 11969 166
rect 12025 140 12145 166
<< polycont >>
rect 9145 750 9179 784
rect 9145 682 9179 716
rect 9322 750 9356 784
rect 9322 682 9356 716
rect 9500 750 9534 784
rect 9500 682 9534 716
rect 9789 750 9823 784
rect 9789 682 9823 716
rect 9960 750 9994 784
rect 9960 682 9994 716
rect 10142 750 10176 784
rect 10142 682 10176 716
rect 10313 750 10347 784
rect 10313 682 10347 716
rect 10615 750 10649 784
rect 10615 682 10649 716
rect 10795 750 10829 784
rect 10795 682 10829 716
rect 10966 750 11000 784
rect 10966 682 11000 716
rect 11256 750 11290 784
rect 11256 682 11290 716
rect 11427 750 11461 784
rect 11427 682 11461 716
rect 11607 750 11641 784
rect 11607 682 11641 716
rect 11894 750 11928 784
rect 11894 682 11928 716
rect 12065 750 12099 784
rect 12065 682 12099 716
<< locali >>
rect 9039 1046 9051 1080
rect 9097 1046 9123 1080
rect 9165 1046 9195 1080
rect 9233 1046 9267 1080
rect 9301 1046 9335 1080
rect 9373 1046 9403 1080
rect 9445 1046 9471 1080
rect 9517 1046 9539 1080
rect 9589 1046 9607 1080
rect 9661 1046 9675 1080
rect 9733 1046 9743 1080
rect 9805 1046 9811 1080
rect 9877 1046 9879 1080
rect 9913 1046 9915 1080
rect 9981 1046 9987 1080
rect 10049 1046 10059 1080
rect 10117 1046 10131 1080
rect 10185 1046 10203 1080
rect 10253 1046 10275 1080
rect 10321 1046 10347 1080
rect 10389 1046 10419 1080
rect 10457 1046 10491 1080
rect 10525 1046 10559 1080
rect 10597 1046 10627 1080
rect 10669 1046 10695 1080
rect 10741 1046 10763 1080
rect 10813 1046 10831 1080
rect 10885 1046 10899 1080
rect 10957 1046 10967 1080
rect 11029 1046 11035 1080
rect 11101 1046 11103 1080
rect 11137 1046 11139 1080
rect 11205 1046 11211 1080
rect 11273 1046 11283 1080
rect 11341 1046 11355 1080
rect 11409 1046 11427 1080
rect 11477 1046 11499 1080
rect 11545 1046 11571 1080
rect 11613 1046 11643 1080
rect 11681 1046 11715 1080
rect 11749 1046 11783 1080
rect 11821 1046 11851 1080
rect 11893 1046 11919 1080
rect 11965 1046 11987 1080
rect 12037 1046 12055 1080
rect 12109 1046 12123 1080
rect 12181 1046 12223 1080
rect 9058 946 9092 962
rect 9058 878 9092 912
rect 9058 616 9092 844
rect 9234 946 9268 961
rect 9234 878 9268 889
rect 9234 828 9268 844
rect 9410 946 9444 962
rect 9410 878 9444 912
rect 9129 750 9145 784
rect 9179 750 9195 784
rect 9129 725 9195 750
rect 9129 716 9149 725
rect 9129 682 9145 716
rect 9183 691 9195 725
rect 9179 682 9195 691
rect 9306 750 9322 784
rect 9365 753 9372 784
rect 9356 750 9372 753
rect 9306 716 9372 750
rect 9306 682 9322 716
rect 9356 715 9372 716
rect 9365 682 9372 715
rect 9129 653 9195 682
rect 9129 619 9149 653
rect 9183 619 9195 653
rect 9410 632 9444 844
rect 9586 946 9620 961
rect 9586 878 9620 889
rect 9586 828 9620 844
rect 9657 962 9733 965
rect 9657 946 9738 962
rect 9657 912 9699 946
rect 9733 912 9738 946
rect 9657 889 9738 912
rect 10051 946 10085 961
rect 10398 946 10437 962
rect 10398 912 10403 946
rect 10398 889 10437 912
rect 9657 878 9909 889
rect 9657 844 9699 878
rect 9733 855 9909 878
rect 9657 794 9733 844
rect 9484 787 9733 794
rect 9484 784 9611 787
rect 9484 750 9500 784
rect 9534 753 9611 784
rect 9645 753 9733 787
rect 9534 750 9733 753
rect 9484 716 9733 750
rect 9484 682 9500 716
rect 9534 715 9733 716
rect 9534 682 9611 715
rect 9645 682 9733 715
rect 9773 753 9785 784
rect 9773 750 9789 753
rect 9823 750 9839 784
rect 9773 716 9839 750
rect 9773 715 9789 716
rect 9773 682 9785 715
rect 9823 682 9839 716
rect 9058 548 9092 582
rect 9058 480 9092 514
rect 9058 354 9092 446
rect 9056 320 9058 325
rect 9234 616 9268 632
rect 9437 598 9475 632
rect 9509 616 9620 632
rect 9509 598 9586 616
rect 9234 548 9268 582
rect 9234 480 9268 514
rect 9234 354 9268 446
rect 9092 320 9094 325
rect 9056 291 9094 320
rect 9058 286 9092 291
rect 9058 218 9092 252
rect 9058 166 9092 184
rect 9234 286 9268 320
rect 9234 244 9268 252
rect 9234 172 9268 184
rect 9410 548 9444 564
rect 9410 480 9444 514
rect 9410 354 9444 446
rect 9410 286 9444 320
rect 9410 218 9444 252
rect 9410 168 9444 184
rect 9586 548 9620 582
rect 9586 480 9620 514
rect 9586 354 9620 446
rect 9586 286 9620 320
rect 9586 218 9620 252
rect 9586 138 9620 184
rect 9699 616 9733 632
rect 9699 548 9733 582
rect 9699 480 9733 514
rect 9699 354 9733 446
rect 9699 286 9733 320
rect 9699 244 9733 252
rect 9699 172 9733 184
rect 9875 616 9909 855
rect 10051 878 10085 889
rect 10051 828 10085 844
rect 10227 878 10437 889
rect 10227 855 10403 878
rect 9944 750 9960 784
rect 9994 753 10051 784
rect 10085 753 10142 784
rect 9994 750 10142 753
rect 10176 750 10192 784
rect 9944 716 10192 750
rect 9944 682 9960 716
rect 9994 715 10142 716
rect 9994 682 10051 715
rect 10085 682 10142 715
rect 10176 682 10192 716
rect 10227 752 10261 855
rect 10403 828 10437 844
rect 10528 946 10562 962
rect 10528 878 10562 912
rect 10528 787 10562 844
rect 10704 946 10738 961
rect 11051 946 11090 962
rect 11051 912 11056 946
rect 11051 889 11090 912
rect 10704 878 10738 889
rect 10704 828 10738 844
rect 10880 878 11090 889
rect 10880 855 11056 878
rect 10227 718 10228 752
rect 10227 680 10262 718
rect 10297 750 10313 784
rect 10347 752 10363 784
rect 10297 718 10315 750
rect 10349 718 10363 752
rect 10297 716 10363 718
rect 10297 682 10313 716
rect 10347 682 10363 716
rect 10528 715 10562 753
rect 10227 646 10228 680
rect 10315 680 10349 682
rect 10599 750 10615 784
rect 10649 758 10665 784
rect 10779 760 10795 784
rect 10829 760 10845 784
rect 10599 724 10621 750
rect 10655 724 10665 758
rect 10722 726 10727 760
rect 10761 750 10795 760
rect 10761 726 10799 750
rect 10833 726 10845 760
rect 10599 716 10665 724
rect 10599 682 10615 716
rect 10649 686 10665 716
rect 10655 682 10665 686
rect 10779 716 10845 726
rect 10779 682 10795 716
rect 10829 682 10845 716
rect 9875 548 9909 582
rect 9875 480 9909 514
rect 9875 354 9909 446
rect 9875 286 9909 320
rect 9875 218 9909 252
rect 9875 166 9909 184
rect 10051 616 10085 632
rect 10051 548 10085 582
rect 10051 480 10085 514
rect 10051 354 10085 446
rect 10051 286 10085 320
rect 10051 244 10085 252
rect 10051 172 10085 184
rect 10227 616 10261 646
rect 10227 548 10261 582
rect 10227 480 10261 514
rect 10227 354 10261 446
rect 10227 286 10261 320
rect 10227 218 10261 252
rect 10227 166 10261 184
rect 10403 616 10437 632
rect 10403 548 10437 582
rect 10403 480 10437 514
rect 10403 354 10437 446
rect 10403 286 10437 320
rect 10403 244 10437 252
rect 10403 172 10437 184
rect 10528 616 10562 681
rect 10621 647 10655 652
rect 10528 567 10562 582
rect 10528 495 10562 514
rect 10528 354 10562 446
rect 10528 286 10562 320
rect 10528 218 10562 252
rect 10528 166 10562 184
rect 10704 616 10738 632
rect 10704 548 10738 582
rect 10704 480 10738 514
rect 10704 354 10738 446
rect 10704 286 10738 320
rect 10704 244 10738 252
rect 10704 172 10738 184
rect 10880 616 10914 855
rect 11056 828 11090 844
rect 11166 946 11205 962
rect 11200 912 11205 946
rect 11166 889 11205 912
rect 11518 946 11552 961
rect 11166 878 11376 889
rect 11200 855 11376 878
rect 11166 828 11200 844
rect 10880 548 10914 582
rect 10880 480 10914 505
rect 10880 354 10914 433
rect 10950 750 10966 784
rect 11000 750 11016 784
rect 10950 716 11016 750
rect 10950 682 10966 716
rect 11000 682 11016 716
rect 11185 760 11256 784
rect 11290 760 11306 784
rect 11185 726 11190 760
rect 11224 750 11256 760
rect 11224 726 11262 750
rect 11296 726 11306 760
rect 11185 716 11306 726
rect 11185 682 11256 716
rect 11290 682 11306 716
rect 10950 475 11016 682
rect 10950 441 10968 475
rect 11002 441 11016 475
rect 10950 403 11016 441
rect 10950 369 10968 403
rect 11002 369 11016 403
rect 10950 364 11016 369
rect 11056 616 11090 632
rect 11056 548 11090 582
rect 11056 480 11090 514
rect 10880 286 10914 320
rect 10880 218 10914 252
rect 10880 166 10914 184
rect 11056 354 11090 446
rect 11056 286 11090 320
rect 11056 244 11090 252
rect 11056 172 11090 184
rect 11166 616 11200 632
rect 11166 548 11200 582
rect 11166 480 11200 514
rect 11166 354 11200 446
rect 11166 286 11200 320
rect 11166 244 11200 252
rect 11166 172 11200 184
rect 11342 616 11376 855
rect 11518 878 11552 889
rect 11518 828 11552 844
rect 11694 946 11728 962
rect 11694 878 11728 912
rect 11411 726 11427 784
rect 11461 760 11477 784
rect 11461 726 11499 760
rect 11591 750 11607 784
rect 11641 750 11657 784
rect 11411 716 11477 726
rect 11411 682 11427 716
rect 11461 682 11477 716
rect 11591 720 11657 750
rect 11591 682 11607 720
rect 11641 682 11657 720
rect 11607 681 11641 682
rect 11342 548 11376 582
rect 11342 501 11376 514
rect 11342 429 11376 446
rect 11342 354 11376 395
rect 11342 286 11376 320
rect 11342 218 11376 252
rect 11342 166 11376 184
rect 11518 616 11552 632
rect 11518 548 11552 582
rect 11518 480 11552 514
rect 11518 354 11552 446
rect 11518 286 11552 320
rect 11518 244 11552 252
rect 11518 172 11552 184
rect 11694 616 11728 844
rect 11804 946 11843 962
rect 11838 912 11843 946
rect 11804 889 11843 912
rect 12156 946 12190 961
rect 11804 878 12014 889
rect 11838 855 12014 878
rect 11804 828 11838 844
rect 11872 760 11894 784
rect 11928 760 11944 784
rect 11818 726 11827 760
rect 11861 750 11894 760
rect 11861 726 11899 750
rect 11933 726 11944 760
rect 11872 716 11944 726
rect 11872 682 11894 716
rect 11928 682 11944 716
rect 11980 659 12014 855
rect 12156 878 12190 889
rect 12156 828 12190 844
rect 12049 726 12065 784
rect 12099 760 12115 784
rect 12099 726 12137 760
rect 12049 716 12115 726
rect 12049 682 12065 716
rect 12099 682 12115 716
rect 11694 548 11728 560
rect 11694 480 11728 488
rect 11694 354 11728 446
rect 11694 286 11728 320
rect 11694 218 11728 252
rect 11694 166 11728 184
rect 11804 616 11838 632
rect 11804 548 11838 582
rect 11804 480 11838 514
rect 11804 354 11838 446
rect 11804 286 11838 320
rect 11804 244 11838 252
rect 11804 172 11838 184
rect 11980 616 12014 625
rect 11980 548 12014 553
rect 11980 480 12014 514
rect 11980 354 12014 446
rect 11980 286 12014 320
rect 11980 218 12014 252
rect 11980 166 12014 184
rect 12156 616 12190 632
rect 12156 548 12190 582
rect 12156 480 12190 514
rect 12156 354 12190 446
rect 12156 286 12190 320
rect 12156 244 12190 252
rect 12156 172 12190 184
rect 9053 66 9065 100
rect 9111 66 9137 100
rect 9179 66 9209 100
rect 9247 66 9281 100
rect 9315 66 9349 100
rect 9387 66 9417 100
rect 9459 66 9485 100
rect 9531 66 9553 100
rect 9603 66 9621 100
rect 9675 66 9689 100
rect 9747 66 9757 100
rect 9819 66 9825 100
rect 9891 66 9893 100
rect 9927 66 9929 100
rect 9995 66 10001 100
rect 10063 66 10073 100
rect 10131 66 10145 100
rect 10199 66 10217 100
rect 10267 66 10289 100
rect 10335 66 10361 100
rect 10403 66 10433 100
rect 10471 66 10505 100
rect 10539 66 10573 100
rect 10611 66 10641 100
rect 10683 66 10709 100
rect 10755 66 10777 100
rect 10827 66 10845 100
rect 10899 66 10913 100
rect 10971 66 10981 100
rect 11043 66 11049 100
rect 11115 66 11117 100
rect 11151 66 11153 100
rect 11219 66 11225 100
rect 11287 66 11297 100
rect 11355 66 11369 100
rect 11423 66 11441 100
rect 11491 66 11513 100
rect 11559 66 11585 100
rect 11627 66 11657 100
rect 11695 66 11729 100
rect 11763 66 11797 100
rect 11835 66 11865 100
rect 11907 66 11933 100
rect 11979 66 12001 100
rect 12051 66 12069 100
rect 12123 66 12137 100
rect 12171 66 12198 100
<< viali >>
rect 9051 1046 9063 1080
rect 9063 1046 9085 1080
rect 9123 1046 9131 1080
rect 9131 1046 9157 1080
rect 9195 1046 9199 1080
rect 9199 1046 9229 1080
rect 9267 1046 9301 1080
rect 9339 1046 9369 1080
rect 9369 1046 9373 1080
rect 9411 1046 9437 1080
rect 9437 1046 9445 1080
rect 9483 1046 9505 1080
rect 9505 1046 9517 1080
rect 9555 1046 9573 1080
rect 9573 1046 9589 1080
rect 9627 1046 9641 1080
rect 9641 1046 9661 1080
rect 9699 1046 9709 1080
rect 9709 1046 9733 1080
rect 9771 1046 9777 1080
rect 9777 1046 9805 1080
rect 9843 1046 9845 1080
rect 9845 1046 9877 1080
rect 9915 1046 9947 1080
rect 9947 1046 9949 1080
rect 9987 1046 10015 1080
rect 10015 1046 10021 1080
rect 10059 1046 10083 1080
rect 10083 1046 10093 1080
rect 10131 1046 10151 1080
rect 10151 1046 10165 1080
rect 10203 1046 10219 1080
rect 10219 1046 10237 1080
rect 10275 1046 10287 1080
rect 10287 1046 10309 1080
rect 10347 1046 10355 1080
rect 10355 1046 10381 1080
rect 10419 1046 10423 1080
rect 10423 1046 10453 1080
rect 10491 1046 10525 1080
rect 10563 1046 10593 1080
rect 10593 1046 10597 1080
rect 10635 1046 10661 1080
rect 10661 1046 10669 1080
rect 10707 1046 10729 1080
rect 10729 1046 10741 1080
rect 10779 1046 10797 1080
rect 10797 1046 10813 1080
rect 10851 1046 10865 1080
rect 10865 1046 10885 1080
rect 10923 1046 10933 1080
rect 10933 1046 10957 1080
rect 10995 1046 11001 1080
rect 11001 1046 11029 1080
rect 11067 1046 11069 1080
rect 11069 1046 11101 1080
rect 11139 1046 11171 1080
rect 11171 1046 11173 1080
rect 11211 1046 11239 1080
rect 11239 1046 11245 1080
rect 11283 1046 11307 1080
rect 11307 1046 11317 1080
rect 11355 1046 11375 1080
rect 11375 1046 11389 1080
rect 11427 1046 11443 1080
rect 11443 1046 11461 1080
rect 11499 1046 11511 1080
rect 11511 1046 11533 1080
rect 11571 1046 11579 1080
rect 11579 1046 11605 1080
rect 11643 1046 11647 1080
rect 11647 1046 11677 1080
rect 11715 1046 11749 1080
rect 11787 1046 11817 1080
rect 11817 1046 11821 1080
rect 11859 1046 11885 1080
rect 11885 1046 11893 1080
rect 11931 1046 11953 1080
rect 11953 1046 11965 1080
rect 12003 1046 12021 1080
rect 12021 1046 12037 1080
rect 12075 1046 12089 1080
rect 12089 1046 12109 1080
rect 12147 1046 12157 1080
rect 12157 1046 12181 1080
rect 9234 961 9268 995
rect 9234 912 9268 923
rect 9234 889 9268 912
rect 9331 784 9365 787
rect 9149 716 9183 725
rect 9149 691 9179 716
rect 9179 691 9183 716
rect 9331 753 9356 784
rect 9356 753 9365 784
rect 9331 682 9356 715
rect 9356 682 9365 715
rect 9331 681 9365 682
rect 9149 619 9183 653
rect 9586 961 9620 995
rect 9586 912 9620 923
rect 9586 889 9620 912
rect 10051 961 10085 995
rect 10051 912 10085 923
rect 10051 889 10085 912
rect 9611 753 9645 787
rect 9785 784 9819 787
rect 9611 681 9645 715
rect 9785 753 9789 784
rect 9789 753 9819 784
rect 9785 682 9789 715
rect 9789 682 9819 715
rect 9785 681 9819 682
rect 9022 291 9056 325
rect 9403 598 9437 632
rect 9475 598 9509 632
rect 9094 291 9128 325
rect 9234 218 9268 244
rect 9234 210 9268 218
rect 9234 138 9268 172
rect 9699 218 9733 244
rect 9699 210 9733 218
rect 9699 138 9733 172
rect 10051 753 10085 787
rect 10051 681 10085 715
rect 10704 961 10738 995
rect 10704 912 10738 923
rect 10704 889 10738 912
rect 10228 718 10262 752
rect 10315 750 10347 752
rect 10347 750 10349 752
rect 10315 718 10349 750
rect 10528 753 10562 787
rect 10228 646 10262 680
rect 10315 646 10349 680
rect 10528 681 10562 715
rect 10621 750 10649 758
rect 10649 750 10655 758
rect 10621 724 10655 750
rect 10727 726 10761 760
rect 10799 750 10829 760
rect 10829 750 10833 760
rect 10799 726 10833 750
rect 10621 682 10649 686
rect 10649 682 10655 686
rect 10051 218 10085 244
rect 10051 210 10085 218
rect 10051 138 10085 172
rect 10403 218 10437 244
rect 10403 210 10437 218
rect 10403 138 10437 172
rect 10621 652 10655 682
rect 10528 548 10562 567
rect 10528 533 10562 548
rect 10528 480 10562 495
rect 10528 461 10562 480
rect 10704 218 10738 244
rect 10704 210 10738 218
rect 10704 138 10738 172
rect 11518 961 11552 995
rect 11518 912 11552 923
rect 11518 889 11552 912
rect 10880 514 10914 539
rect 10880 505 10914 514
rect 10880 446 10914 467
rect 10880 433 10914 446
rect 11190 726 11224 760
rect 11262 750 11290 760
rect 11290 750 11296 760
rect 11262 726 11296 750
rect 10968 441 11002 475
rect 10968 369 11002 403
rect 11056 218 11090 244
rect 11056 210 11090 218
rect 11056 138 11090 172
rect 11166 218 11200 244
rect 11166 210 11200 218
rect 11166 138 11200 172
rect 11607 784 11641 792
rect 11427 750 11461 760
rect 11427 726 11461 750
rect 11499 726 11533 760
rect 11607 758 11641 784
rect 11607 716 11641 720
rect 11607 686 11641 716
rect 11342 480 11376 501
rect 11342 467 11376 480
rect 11342 395 11376 429
rect 11518 218 11552 244
rect 11518 210 11552 218
rect 11518 138 11552 172
rect 12156 961 12190 995
rect 12156 912 12190 923
rect 12156 889 12190 912
rect 11827 726 11861 760
rect 11899 750 11928 760
rect 11928 750 11933 760
rect 11899 726 11933 750
rect 12065 750 12099 760
rect 12065 726 12099 750
rect 12137 726 12171 760
rect 11694 582 11728 594
rect 11694 560 11728 582
rect 11694 514 11728 522
rect 11694 488 11728 514
rect 11804 218 11838 244
rect 11804 210 11838 218
rect 11804 138 11838 172
rect 11980 625 12014 659
rect 11980 582 12014 587
rect 11980 553 12014 582
rect 12156 218 12190 244
rect 12156 210 12190 218
rect 12156 138 12190 172
rect 9065 66 9077 100
rect 9077 66 9099 100
rect 9137 66 9145 100
rect 9145 66 9171 100
rect 9209 66 9213 100
rect 9213 66 9243 100
rect 9281 66 9315 100
rect 9353 66 9383 100
rect 9383 66 9387 100
rect 9425 66 9451 100
rect 9451 66 9459 100
rect 9497 66 9519 100
rect 9519 66 9531 100
rect 9569 66 9587 100
rect 9587 66 9603 100
rect 9641 66 9655 100
rect 9655 66 9675 100
rect 9713 66 9723 100
rect 9723 66 9747 100
rect 9785 66 9791 100
rect 9791 66 9819 100
rect 9857 66 9859 100
rect 9859 66 9891 100
rect 9929 66 9961 100
rect 9961 66 9963 100
rect 10001 66 10029 100
rect 10029 66 10035 100
rect 10073 66 10097 100
rect 10097 66 10107 100
rect 10145 66 10165 100
rect 10165 66 10179 100
rect 10217 66 10233 100
rect 10233 66 10251 100
rect 10289 66 10301 100
rect 10301 66 10323 100
rect 10361 66 10369 100
rect 10369 66 10395 100
rect 10433 66 10437 100
rect 10437 66 10467 100
rect 10505 66 10539 100
rect 10577 66 10607 100
rect 10607 66 10611 100
rect 10649 66 10675 100
rect 10675 66 10683 100
rect 10721 66 10743 100
rect 10743 66 10755 100
rect 10793 66 10811 100
rect 10811 66 10827 100
rect 10865 66 10879 100
rect 10879 66 10899 100
rect 10937 66 10947 100
rect 10947 66 10971 100
rect 11009 66 11015 100
rect 11015 66 11043 100
rect 11081 66 11083 100
rect 11083 66 11115 100
rect 11153 66 11185 100
rect 11185 66 11187 100
rect 11225 66 11253 100
rect 11253 66 11259 100
rect 11297 66 11321 100
rect 11321 66 11331 100
rect 11369 66 11389 100
rect 11389 66 11403 100
rect 11441 66 11457 100
rect 11457 66 11475 100
rect 11513 66 11525 100
rect 11525 66 11547 100
rect 11585 66 11593 100
rect 11593 66 11619 100
rect 11657 66 11661 100
rect 11661 66 11691 100
rect 11729 66 11763 100
rect 11801 66 11831 100
rect 11831 66 11835 100
rect 11873 66 11899 100
rect 11899 66 11907 100
rect 11945 66 11967 100
rect 11967 66 11979 100
rect 12017 66 12035 100
rect 12035 66 12051 100
rect 12089 66 12103 100
rect 12103 66 12123 100
<< metal1 >>
tri 3115 39968 3147 40000 se
rect 2697 39916 2703 39968
rect 2755 39916 2793 39968
rect 2845 39916 2883 39968
rect 2935 39916 2973 39968
rect 3025 39916 3063 39968
rect 3115 39916 3158 39968
rect 2697 39876 3158 39916
rect 2697 39824 2703 39876
rect 2755 39824 2793 39876
rect 2845 39824 2883 39876
rect 2935 39824 2973 39876
rect 3025 39824 3063 39876
rect 3115 39824 3158 39876
rect 2697 39784 3158 39824
rect 2697 39732 2703 39784
rect 2755 39732 2793 39784
rect 2845 39732 2883 39784
rect 2935 39732 2973 39784
rect 3025 39732 3063 39784
rect 3115 39732 3158 39784
rect 3342 39782 3799 39961
rect 15429 39770 15848 39986
tri 3115 39700 3147 39732 ne
rect 954 38664 960 38716
rect 1012 38664 1024 38716
rect 1076 38664 2546 38716
tri 2460 38630 2494 38664 ne
rect 1014 38387 1020 38439
rect 1072 38387 1084 38439
rect 1136 38387 2466 38439
tri 2380 38353 2414 38387 ne
rect 2414 38204 2466 38387
rect 2494 38322 2546 38664
rect 3449 38545 3455 38597
rect 3507 38545 3519 38597
rect 3571 38545 3577 38597
tri 2546 38322 2580 38356 sw
rect 2494 38270 3455 38322
rect 3507 38270 3519 38322
rect 3571 38270 3577 38322
tri 2466 38204 2500 38238 sw
rect 2414 38152 3210 38204
rect 3262 38152 3274 38204
rect 3326 38152 3332 38204
rect 2470 38107 3333 38113
rect 2522 38061 3333 38107
rect 2470 38043 2522 38055
tri 2522 38027 2556 38061 nw
rect 15862 38051 15914 38057
tri 15846 38027 15862 38043 se
tri 15828 38009 15846 38027 se
rect 15846 38009 15862 38027
rect 2470 37985 2522 37991
rect 2774 37907 2780 37959
rect 2832 37907 2844 37959
rect 2896 37958 2902 37959
tri 2902 37958 2903 37959 sw
rect 2896 37907 8463 37958
rect 13588 37929 13594 37981
rect 13646 37929 13660 37981
rect 13712 37929 13718 37981
rect 15473 37934 15595 38006
rect 15818 37999 15862 38009
rect 15818 37987 15914 37999
rect 15818 37935 15862 37987
rect 15818 37929 15914 37935
rect 2774 37894 8463 37907
rect 2774 37891 8341 37894
rect 2774 37839 2780 37891
rect 2832 37839 2844 37891
rect 2896 37842 8341 37891
rect 8393 37842 8405 37894
rect 8457 37842 8463 37894
rect 2896 37839 8463 37842
tri 8463 37839 8530 37906 nw
rect 2550 37664 2556 37716
rect 2608 37664 2620 37716
rect 2672 37664 4271 37716
rect 4323 37664 4335 37716
rect 4387 37664 4395 37716
rect 2390 37407 2442 37413
rect 3301 37377 3307 37429
rect 3359 37377 3371 37429
rect 3423 37377 3429 37429
rect 2390 37343 2442 37355
tri 2442 37337 2476 37371 sw
rect 2442 37291 3333 37337
rect 2390 37285 3333 37291
tri 15426 37210 15460 37244 ne
rect 2435 37101 2902 37124
rect 2435 37049 2780 37101
rect 2832 37049 2844 37101
rect 2896 37049 2902 37101
rect 2435 37028 2902 37049
rect 13866 37101 13918 37107
rect 15723 37101 15775 37107
rect 13866 37037 13918 37049
rect 1284 36946 2058 36998
rect 2162 36482 2259 36998
rect 2131 36459 2137 36482
tri 2024 36354 2129 36459 ne
rect 2129 36430 2137 36459
rect 2189 36430 2201 36482
rect 2253 36430 2259 36482
rect 2129 36406 2259 36430
rect 2129 36354 2137 36406
rect 2189 36354 2201 36406
rect 2253 36354 2259 36406
tri 2401 36222 2435 36256 se
rect 2435 36222 2517 37028
tri 2517 36994 2551 37028 nw
tri 13918 37031 13952 37065 sw
tri 15689 37031 15723 37065 se
rect 15723 37037 15775 37049
rect 13918 36985 15723 37031
rect 13866 36979 15775 36985
rect 794 36203 2517 36222
rect 794 36151 800 36203
rect 852 36151 864 36203
rect 916 36151 2517 36203
rect 2612 36202 3014 36319
rect 794 36140 2517 36151
rect 0 36079 3141 36080
rect 0 36074 397 36079
rect 0 36022 157 36074
rect 209 36022 269 36074
rect 321 36027 397 36074
rect 449 36027 489 36079
rect 541 36027 581 36079
rect 633 36027 673 36079
rect 725 36074 3141 36079
rect 725 36027 2131 36074
rect 321 36022 2131 36027
rect 2183 36022 2207 36074
rect 2259 36022 3141 36074
rect 0 35997 3141 36022
rect 0 35996 397 35997
rect 0 35944 157 35996
rect 209 35944 269 35996
rect 321 35945 397 35996
rect 449 35945 489 35997
rect 541 35945 581 35997
rect 633 35945 673 35997
rect 725 35996 3141 35997
rect 725 35945 2131 35996
rect 321 35944 2131 35945
rect 2183 35944 2207 35996
rect 2259 35944 3141 35996
rect 0 35917 3141 35944
rect 0 35865 157 35917
rect 209 35865 269 35917
rect 321 35915 2131 35917
rect 321 35865 397 35915
rect 0 35863 397 35865
rect 449 35863 489 35915
rect 541 35863 581 35915
rect 633 35863 673 35915
rect 725 35865 2131 35915
rect 2183 35865 2207 35917
rect 2259 35865 3141 35917
rect 725 35863 3141 35865
rect 0 35838 3141 35863
rect 0 35786 157 35838
rect 209 35786 269 35838
rect 321 35833 2131 35838
rect 321 35786 397 35833
rect 0 35781 397 35786
rect 449 35781 489 35833
rect 541 35781 581 35833
rect 633 35781 673 35833
rect 725 35786 2131 35833
rect 2183 35786 2207 35838
rect 2259 35786 3141 35838
rect 725 35781 3141 35786
rect 0 35780 3141 35781
tri 2058 35701 2064 35707 se
rect 2064 35655 2070 35707
rect 2122 35655 2149 35707
rect 2201 35655 2227 35707
rect 2279 35655 2305 35707
rect 2357 35655 2363 35707
tri 2363 35701 2369 35707 sw
tri 5489 3800 5496 3807 se
rect 5496 3800 8566 3807
rect 1090 3770 1142 3776
tri 1142 3731 1185 3774 sw
tri 1844 3731 1878 3765 se
rect 1878 3760 2175 3800
tri 5453 3764 5489 3800 se
rect 5489 3767 8566 3800
rect 5489 3764 5496 3767
rect 1878 3731 1918 3760
rect 1142 3718 1918 3731
tri 1918 3726 1952 3760 nw
tri 2101 3726 2135 3760 ne
rect 2135 3730 2175 3760
tri 2175 3730 2209 3764 sw
tri 5438 3749 5453 3764 se
rect 5453 3749 5496 3764
tri 5496 3749 5514 3767 nw
tri 8548 3749 8566 3767 ne
tri 8566 3751 8622 3807 sw
rect 8566 3749 8764 3751
tri 5419 3730 5438 3749 se
rect 5438 3730 5477 3749
tri 5477 3730 5496 3749 nw
tri 8566 3730 8585 3749 ne
rect 8585 3730 8764 3749
rect 1090 3706 1918 3718
rect 1142 3691 1918 3706
rect 1090 3648 1142 3654
tri 1142 3648 1185 3691 nw
rect 2135 3690 5437 3730
tri 5437 3690 5477 3730 nw
tri 8585 3699 8616 3730 ne
rect 8616 3699 8764 3730
rect 8816 3699 8828 3751
rect 8880 3699 8886 3751
rect 1134 3460 1140 3512
rect 1192 3460 1204 3512
rect 1256 3509 1262 3512
tri 1262 3509 1265 3512 sw
tri 9503 3509 9505 3511 se
rect 9505 3509 9511 3511
rect 1256 3469 9511 3509
rect 1256 3460 1262 3469
tri 1262 3460 1271 3469 nw
tri 9500 3464 9505 3469 ne
rect 9505 3459 9511 3469
rect 9563 3459 9575 3511
rect 9627 3459 9633 3511
tri 1340 3432 1344 3436 se
rect 1344 3432 9298 3436
rect 1073 3380 1079 3432
rect 1131 3380 1143 3432
rect 1195 3431 9298 3432
tri 9298 3431 9303 3436 sw
rect 1195 3396 9434 3431
rect 1195 3392 1384 3396
tri 1384 3392 1388 3396 nw
tri 9253 3392 9257 3396 ne
rect 9257 3392 9434 3396
rect 1195 3380 1201 3392
tri 1201 3380 1213 3392 nw
tri 9257 3391 9258 3392 ne
rect 9258 3391 9434 3392
tri 9421 3384 9428 3391 ne
rect 9428 3379 9434 3391
rect 9486 3379 9498 3431
rect 9550 3379 9556 3431
rect 9003 1080 12240 1092
rect 9003 1046 9051 1080
rect 9085 1046 9123 1080
rect 9157 1046 9195 1080
rect 9229 1046 9267 1080
rect 9301 1046 9339 1080
rect 9373 1046 9411 1080
rect 9445 1046 9483 1080
rect 9517 1046 9555 1080
rect 9589 1046 9627 1080
rect 9661 1046 9699 1080
rect 9733 1046 9771 1080
rect 9805 1046 9843 1080
rect 9877 1046 9915 1080
rect 9949 1046 9987 1080
rect 10021 1046 10059 1080
rect 10093 1046 10131 1080
rect 10165 1046 10203 1080
rect 10237 1046 10275 1080
rect 10309 1046 10347 1080
rect 10381 1046 10419 1080
rect 10453 1046 10491 1080
rect 10525 1046 10563 1080
rect 10597 1046 10635 1080
rect 10669 1046 10707 1080
rect 10741 1046 10779 1080
rect 10813 1046 10851 1080
rect 10885 1046 10923 1080
rect 10957 1046 10995 1080
rect 11029 1046 11067 1080
rect 11101 1046 11139 1080
rect 11173 1046 11211 1080
rect 11245 1046 11283 1080
rect 11317 1046 11355 1080
rect 11389 1046 11427 1080
rect 11461 1046 11499 1080
rect 11533 1046 11571 1080
rect 11605 1046 11643 1080
rect 11677 1046 11715 1080
rect 11749 1046 11787 1080
rect 11821 1046 11859 1080
rect 11893 1046 11931 1080
rect 11965 1046 12003 1080
rect 12037 1046 12075 1080
rect 12109 1046 12147 1080
rect 12181 1046 12240 1080
rect 9003 995 12240 1046
rect 9003 961 9234 995
rect 9268 961 9586 995
rect 9620 961 10051 995
rect 10085 961 10704 995
rect 10738 961 11518 995
rect 11552 961 12156 995
rect 12190 961 12240 995
rect 9003 923 12240 961
rect 9003 889 9234 923
rect 9268 889 9586 923
rect 9620 889 10051 923
rect 10085 889 10704 923
rect 10738 889 11518 923
rect 11552 889 12156 923
rect 12190 889 12240 923
rect 9003 877 12240 889
rect 10045 803 10568 849
rect 9325 787 9371 799
rect 9325 753 9331 787
rect 9365 753 9371 787
rect 9143 725 9195 737
rect 9143 710 9149 725
rect 9183 710 9195 725
rect 9325 715 9371 753
rect 9325 681 9331 715
rect 9365 681 9371 715
tri 9195 669 9198 672 sw
rect 9325 669 9371 681
rect 9602 789 9654 799
rect 9602 725 9654 737
rect 9195 667 9198 669
tri 9198 667 9200 669 sw
rect 9602 667 9654 673
rect 9779 787 9825 799
rect 9779 753 9785 787
rect 9819 753 9825 787
rect 9779 715 9825 753
rect 9779 681 9785 715
rect 9819 681 9825 715
rect 9779 669 9825 681
rect 10045 795 10117 803
tri 10117 795 10125 803 nw
tri 10488 795 10496 803 ne
rect 10496 795 10568 803
rect 10045 792 10114 795
tri 10114 792 10117 795 nw
tri 10496 792 10499 795 ne
rect 10499 792 10568 795
rect 10045 787 10109 792
tri 10109 787 10114 792 nw
tri 10499 787 10504 792 ne
rect 10504 787 10568 792
rect 10045 753 10051 787
rect 10085 753 10091 787
tri 10091 769 10109 787 nw
tri 10504 769 10522 787 ne
rect 10045 715 10091 753
rect 10045 681 10051 715
rect 10085 681 10091 715
rect 10045 669 10091 681
rect 10222 752 10268 764
rect 10222 718 10228 752
rect 10262 718 10268 752
rect 10222 680 10268 718
rect 9195 658 9200 667
rect 9143 653 9200 658
rect 9143 646 9149 653
rect 9183 646 9200 653
tri 9200 646 9221 667 sw
rect 10222 646 10228 680
rect 10262 646 10268 680
rect 9195 638 9221 646
tri 9221 638 9229 646 sw
rect 9195 632 9521 638
rect 10222 634 10268 646
rect 10309 752 10355 764
rect 10309 718 10315 752
rect 10349 718 10355 752
rect 10309 680 10355 718
rect 10309 646 10315 680
rect 10349 646 10355 680
rect 10522 753 10528 787
rect 10562 753 10568 787
rect 11601 792 11647 804
rect 10522 715 10568 753
rect 10522 681 10528 715
rect 10562 681 10568 715
rect 10522 664 10568 681
rect 10615 758 10661 770
rect 10615 724 10621 758
rect 10655 724 10661 758
rect 10615 686 10661 724
rect 10710 760 10853 766
tri 10853 760 10859 766 sw
rect 11173 760 11309 766
tri 11309 760 11315 766 sw
rect 11410 760 11545 766
rect 10710 726 10727 760
rect 10761 726 10799 760
rect 10833 726 10859 760
tri 10859 726 10893 760 sw
rect 11173 726 11190 760
rect 11224 726 11262 760
rect 11296 736 11315 760
tri 11315 736 11339 760 sw
rect 11296 726 11339 736
tri 11339 726 11349 736 sw
rect 11410 726 11427 760
rect 11461 726 11499 760
rect 11533 726 11545 760
rect 10710 720 10893 726
tri 10893 720 10899 726 sw
rect 11173 720 11349 726
tri 11349 720 11355 726 sw
rect 11410 720 11545 726
rect 11601 758 11607 792
rect 11641 758 11647 792
rect 11601 726 11647 758
rect 11806 760 11945 766
tri 11647 726 11668 747 sw
rect 11806 726 11827 760
rect 11861 726 11899 760
rect 11933 726 11945 760
rect 11601 720 11668 726
tri 11668 720 11674 726 sw
rect 11806 720 11945 726
rect 12048 760 12183 766
rect 12048 726 12065 760
rect 12099 726 12137 760
rect 12171 726 12183 760
rect 12048 720 12183 726
tri 10833 715 10838 720 ne
rect 10838 715 10899 720
tri 10661 686 10690 715 sw
tri 10838 686 10867 715 ne
rect 10867 692 10899 715
tri 10899 692 10927 720 sw
tri 11289 692 11317 720 ne
rect 11317 692 11355 720
tri 11355 692 11383 720 sw
rect 10867 686 10927 692
tri 10927 686 10933 692 sw
tri 11317 686 11323 692 ne
rect 11323 691 11383 692
tri 11383 691 11384 692 sw
rect 11323 690 11384 691
tri 11384 690 11385 691 sw
rect 11323 689 11385 690
tri 11385 689 11386 690 sw
rect 11323 688 11386 689
tri 11386 688 11387 689 sw
rect 11323 687 11387 688
tri 11387 687 11388 688 sw
rect 11323 686 11388 687
tri 11388 686 11389 687 sw
rect 11601 686 11607 720
rect 11641 713 11674 720
tri 11674 713 11681 720 sw
rect 11641 686 11761 713
rect 10309 634 10355 646
rect 10615 652 10621 686
rect 10655 681 10690 686
tri 10690 681 10695 686 sw
tri 10867 681 10872 686 ne
rect 10872 681 10933 686
rect 10655 667 10757 681
tri 10757 667 10771 681 sw
tri 10872 667 10886 681 ne
rect 10886 667 10933 681
tri 10933 667 10952 686 sw
tri 11323 667 11342 686 ne
rect 11342 685 11389 686
tri 11389 685 11390 686 sw
rect 11342 684 11390 685
tri 11390 684 11391 685 sw
rect 11342 683 11391 684
tri 11391 683 11392 684 sw
rect 11342 682 11392 683
tri 11392 682 11393 683 sw
rect 11342 681 11393 682
tri 11393 681 11394 682 sw
rect 11342 680 11394 681
tri 11394 680 11395 681 sw
rect 11342 679 11395 680
tri 11395 679 11396 680 sw
rect 11342 678 11396 679
tri 11396 678 11397 679 sw
rect 11342 677 11397 678
tri 11397 677 11398 678 sw
rect 11342 676 11398 677
tri 11398 676 11399 677 sw
rect 11342 675 11399 676
tri 11399 675 11400 676 sw
rect 11342 674 11400 675
tri 11400 674 11401 675 sw
rect 11342 673 11401 674
tri 11401 673 11402 674 sw
rect 11342 672 11402 673
tri 11402 672 11403 673 sw
rect 11342 671 11403 672
tri 11403 671 11404 672 sw
rect 11601 671 11761 686
tri 11761 671 11803 713 sw
rect 11342 669 11404 671
tri 11404 669 11406 671 sw
rect 11601 669 12020 671
rect 11342 667 11406 669
tri 11406 667 11408 669 sw
tri 11742 667 11744 669 ne
rect 11744 667 12020 669
rect 10655 665 10771 667
tri 10771 665 10773 667 sw
tri 10886 665 10888 667 ne
rect 10888 665 10952 667
tri 10952 665 10954 667 sw
tri 11342 665 11344 667 ne
rect 11344 665 11408 667
rect 10655 659 10773 665
tri 10773 659 10779 665 sw
tri 10888 659 10894 665 ne
rect 10894 659 10954 665
tri 10954 659 10960 665 sw
tri 11344 659 11350 665 ne
rect 11350 659 11408 665
tri 11408 659 11416 667 sw
tri 11744 659 11752 667 ne
rect 11752 659 12020 667
rect 10655 652 10779 659
rect 10615 635 10779 652
tri 10779 635 10803 659 sw
tri 10894 635 10918 659 ne
rect 10918 635 10960 659
tri 10735 634 10736 635 ne
rect 10736 634 10803 635
rect 9195 598 9403 632
rect 9437 598 9475 632
rect 9509 598 9521 632
tri 10736 625 10745 634 ne
rect 10745 625 10803 634
tri 10803 625 10813 635 sw
tri 10918 625 10928 635 ne
rect 10928 626 10960 635
tri 10960 626 10993 659 sw
tri 11350 626 11383 659 ne
rect 11383 626 11416 659
tri 11416 626 11449 659 sw
tri 11752 626 11785 659 ne
rect 11785 626 11980 659
rect 10928 625 10993 626
tri 10993 625 10994 626 sw
tri 11383 625 11384 626 ne
rect 11384 625 11449 626
tri 11449 625 11450 626 sw
tri 11785 625 11786 626 ne
rect 11786 625 11980 626
rect 12014 625 12020 659
rect 9195 594 9521 598
tri 10745 594 10776 625 ne
rect 10776 599 10813 625
tri 10813 599 10839 625 sw
tri 10928 599 10954 625 ne
rect 10954 599 10994 625
tri 10994 599 11020 625 sw
tri 11384 599 11410 625 ne
rect 11410 624 11450 625
tri 11450 624 11451 625 sw
tri 11940 624 11941 625 ne
rect 11941 624 12020 625
rect 11410 623 11451 624
tri 11451 623 11452 624 sw
tri 11941 623 11942 624 ne
rect 11942 623 12020 624
rect 11410 622 11452 623
tri 11452 622 11453 623 sw
tri 11942 622 11943 623 ne
rect 11943 622 12020 623
rect 11410 621 11453 622
tri 11453 621 11454 622 sw
tri 11943 621 11944 622 ne
rect 11944 621 12020 622
rect 11410 620 11454 621
tri 11454 620 11455 621 sw
tri 11944 620 11945 621 ne
rect 11945 620 12020 621
rect 11410 619 11455 620
tri 11455 619 11456 620 sw
tri 11945 619 11946 620 ne
rect 11946 619 12020 620
rect 11410 618 11456 619
tri 11456 618 11457 619 sw
tri 11946 618 11947 619 ne
rect 11947 618 12020 619
rect 11410 617 11457 618
tri 11457 617 11458 618 sw
tri 11947 617 11948 618 ne
rect 11948 617 12020 618
rect 11410 616 11458 617
tri 11458 616 11459 617 sw
tri 11948 616 11949 617 ne
rect 11949 616 12020 617
rect 11410 615 11459 616
tri 11459 615 11460 616 sw
tri 11949 615 11950 616 ne
rect 11950 615 12020 616
rect 11410 614 11460 615
tri 11460 614 11461 615 sw
tri 11950 614 11951 615 ne
rect 11951 614 12020 615
rect 11410 613 11461 614
tri 11461 613 11462 614 sw
tri 11951 613 11952 614 ne
rect 11952 613 12020 614
rect 11410 612 11462 613
tri 11462 612 11463 613 sw
tri 11952 612 11953 613 ne
rect 11953 612 12020 613
rect 11410 611 11463 612
tri 11463 611 11464 612 sw
tri 11953 611 11954 612 ne
rect 11954 611 12020 612
rect 11410 610 11464 611
tri 11464 610 11465 611 sw
tri 11954 610 11955 611 ne
rect 11955 610 12020 611
rect 11410 609 11465 610
tri 11465 609 11466 610 sw
tri 11955 609 11956 610 ne
rect 11956 609 12020 610
rect 11410 608 11466 609
tri 11466 608 11467 609 sw
tri 11956 608 11957 609 ne
rect 11957 608 12020 609
rect 11410 607 11467 608
tri 11467 607 11468 608 sw
tri 11957 607 11958 608 ne
rect 11958 607 12020 608
rect 11410 606 11468 607
tri 11468 606 11469 607 sw
tri 11958 606 11959 607 ne
rect 11959 606 12020 607
rect 11410 599 11734 606
rect 10776 594 10839 599
tri 10839 594 10844 599 sw
tri 10954 594 10959 599 ne
rect 10959 594 11020 599
tri 11020 594 11025 599 sw
tri 11410 594 11415 599 ne
rect 11415 594 11734 599
rect 9143 592 9521 594
tri 10776 592 10778 594 ne
rect 10778 592 10844 594
rect 9143 588 9195 592
tri 9195 588 9199 592 nw
tri 10778 588 10782 592 ne
rect 10782 588 10844 592
tri 10844 588 10850 594 sw
tri 10959 588 10965 594 ne
rect 10965 588 11025 594
tri 11025 588 11031 594 sw
tri 11415 588 11421 594 ne
rect 11421 588 11694 594
tri 10782 579 10791 588 ne
rect 10791 579 10850 588
rect 10522 567 10568 579
tri 10791 567 10803 579 ne
rect 10803 567 10850 579
tri 10850 567 10871 588 sw
tri 10965 567 10986 588 ne
rect 10986 567 11031 588
rect 10522 533 10528 567
rect 10562 533 10568 567
tri 10803 560 10810 567 ne
rect 10810 560 10871 567
tri 10871 560 10878 567 sw
tri 10986 560 10993 567 ne
rect 10993 560 11031 567
tri 11031 560 11059 588 sw
tri 11421 560 11449 588 ne
rect 11449 560 11694 588
rect 11728 560 11734 594
tri 11959 591 11974 606 ne
tri 10810 553 10817 560 ne
rect 10817 553 10878 560
tri 10878 553 10885 560 sw
tri 10993 553 11000 560 ne
rect 11000 553 11059 560
tri 11059 553 11066 560 sw
tri 11654 553 11661 560 ne
rect 11661 553 11734 560
tri 10817 539 10831 553 ne
rect 10831 551 10885 553
tri 10885 551 10887 553 sw
tri 11000 551 11002 553 ne
rect 11002 551 11066 553
rect 10831 539 10920 551
rect 10522 495 10568 533
tri 10831 505 10865 539 ne
rect 10865 505 10880 539
rect 10914 505 10920 539
tri 11002 533 11020 551 ne
rect 11020 533 11066 551
tri 11066 533 11086 553 sw
tri 11661 533 11681 553 ne
rect 11681 533 11734 553
rect 11974 587 12020 606
rect 11974 553 11980 587
rect 12014 553 12020 587
rect 11974 536 12020 553
tri 11020 522 11031 533 ne
rect 11031 526 11086 533
tri 11086 526 11093 533 sw
tri 11681 526 11688 533 ne
rect 11031 522 11093 526
tri 11093 522 11097 526 sw
rect 11688 522 11734 533
tri 10865 501 10869 505 ne
rect 10869 501 10920 505
tri 11031 501 11052 522 ne
rect 11052 513 11097 522
tri 11097 513 11106 522 sw
rect 11052 501 11382 513
tri 10869 499 10871 501 ne
rect 10871 499 10920 501
tri 10871 496 10874 499 ne
rect 10522 461 10528 495
rect 10562 461 10568 495
rect 10522 444 10568 461
rect 10874 467 10920 499
tri 11052 487 11066 501 ne
rect 11066 487 11342 501
rect 10874 433 10880 467
rect 10914 433 10920 467
rect 10874 416 10920 433
rect 10962 475 11008 487
rect 10962 441 10968 475
rect 11002 441 11008 475
tri 11066 467 11086 487 ne
rect 11086 467 11342 487
rect 11376 467 11382 501
rect 11688 488 11694 522
rect 11728 488 11734 522
rect 11688 471 11734 488
rect 10962 403 11008 441
tri 11302 433 11336 467 ne
rect 10962 369 10968 403
rect 11002 369 11008 403
rect 11336 429 11382 467
rect 11336 395 11342 429
rect 11376 395 11382 429
rect 11336 378 11382 395
rect 10962 352 11008 369
rect 9008 325 9360 337
rect 9008 291 9022 325
rect 9056 291 9094 325
rect 9128 291 9360 325
rect 9008 285 9360 291
rect 9412 285 9445 337
rect 9497 285 9503 337
rect 9003 244 12239 257
rect 9003 210 9234 244
rect 9268 210 9699 244
rect 9733 210 10051 244
rect 10085 210 10403 244
rect 10437 210 10704 244
rect 10738 210 11056 244
rect 11090 210 11166 244
rect 11200 210 11518 244
rect 11552 210 11804 244
rect 11838 210 12156 244
rect 12190 210 12239 244
rect 9003 172 12239 210
rect 9003 138 9234 172
rect 9268 138 9699 172
rect 9733 138 10051 172
rect 10085 138 10403 172
rect 10437 138 10704 172
rect 10738 138 11056 172
rect 11090 138 11166 172
rect 11200 138 11518 172
rect 11552 138 11804 172
rect 11838 138 12156 172
rect 12190 138 12239 172
rect 9003 100 12239 138
rect 9003 66 9065 100
rect 9099 66 9137 100
rect 9171 66 9209 100
rect 9243 66 9281 100
rect 9315 66 9353 100
rect 9387 66 9425 100
rect 9459 66 9497 100
rect 9531 66 9569 100
rect 9603 66 9641 100
rect 9675 66 9713 100
rect 9747 66 9785 100
rect 9819 66 9857 100
rect 9891 66 9929 100
rect 9963 66 10001 100
rect 10035 66 10073 100
rect 10107 66 10145 100
rect 10179 66 10217 100
rect 10251 66 10289 100
rect 10323 66 10361 100
rect 10395 66 10433 100
rect 10467 66 10505 100
rect 10539 66 10577 100
rect 10611 66 10649 100
rect 10683 66 10721 100
rect 10755 66 10793 100
rect 10827 66 10865 100
rect 10899 66 10937 100
rect 10971 66 11009 100
rect 11043 66 11081 100
rect 11115 66 11153 100
rect 11187 66 11225 100
rect 11259 66 11297 100
rect 11331 66 11369 100
rect 11403 66 11441 100
rect 11475 66 11513 100
rect 11547 66 11585 100
rect 11619 66 11657 100
rect 11691 66 11729 100
rect 11763 66 11801 100
rect 11835 66 11873 100
rect 11907 66 11945 100
rect 11979 66 12017 100
rect 12051 66 12089 100
rect 12123 66 12239 100
rect 9003 54 12239 66
<< via1 >>
rect 2703 39916 2755 39968
rect 2793 39916 2845 39968
rect 2883 39916 2935 39968
rect 2973 39916 3025 39968
rect 3063 39916 3115 39968
rect 2703 39824 2755 39876
rect 2793 39824 2845 39876
rect 2883 39824 2935 39876
rect 2973 39824 3025 39876
rect 3063 39824 3115 39876
rect 2703 39732 2755 39784
rect 2793 39732 2845 39784
rect 2883 39732 2935 39784
rect 2973 39732 3025 39784
rect 3063 39732 3115 39784
rect 960 38664 1012 38716
rect 1024 38664 1076 38716
rect 1020 38387 1072 38439
rect 1084 38387 1136 38439
rect 3455 38545 3507 38597
rect 3519 38545 3571 38597
rect 3455 38270 3507 38322
rect 3519 38270 3571 38322
rect 3210 38152 3262 38204
rect 3274 38152 3326 38204
rect 2470 38055 2522 38107
rect 2470 37991 2522 38043
rect 2780 37907 2832 37959
rect 2844 37907 2896 37959
rect 13594 37929 13646 37981
rect 13660 37929 13712 37981
rect 15862 37999 15914 38051
rect 15862 37935 15914 37987
rect 2780 37839 2832 37891
rect 2844 37839 2896 37891
rect 8341 37842 8393 37894
rect 8405 37842 8457 37894
rect 2556 37664 2608 37716
rect 2620 37664 2672 37716
rect 4271 37664 4323 37716
rect 4335 37664 4387 37716
rect 2390 37355 2442 37407
rect 3307 37377 3359 37429
rect 3371 37377 3423 37429
rect 2390 37291 2442 37343
rect 2780 37049 2832 37101
rect 2844 37049 2896 37101
rect 13866 37049 13918 37101
rect 2137 36430 2189 36482
rect 2201 36430 2253 36482
rect 2137 36354 2189 36406
rect 2201 36354 2253 36406
rect 13866 36985 13918 37037
rect 15723 37049 15775 37101
rect 15723 36985 15775 37037
rect 800 36151 852 36203
rect 864 36151 916 36203
rect 157 36022 209 36074
rect 269 36022 321 36074
rect 397 36027 449 36079
rect 489 36027 541 36079
rect 581 36027 633 36079
rect 673 36027 725 36079
rect 2131 36022 2183 36074
rect 2207 36022 2259 36074
rect 157 35944 209 35996
rect 269 35944 321 35996
rect 397 35945 449 35997
rect 489 35945 541 35997
rect 581 35945 633 35997
rect 673 35945 725 35997
rect 2131 35944 2183 35996
rect 2207 35944 2259 35996
rect 157 35865 209 35917
rect 269 35865 321 35917
rect 397 35863 449 35915
rect 489 35863 541 35915
rect 581 35863 633 35915
rect 673 35863 725 35915
rect 2131 35865 2183 35917
rect 2207 35865 2259 35917
rect 157 35786 209 35838
rect 269 35786 321 35838
rect 397 35781 449 35833
rect 489 35781 541 35833
rect 581 35781 633 35833
rect 673 35781 725 35833
rect 2131 35786 2183 35838
rect 2207 35786 2259 35838
rect 2070 35655 2122 35707
rect 2149 35655 2201 35707
rect 2227 35655 2279 35707
rect 2305 35655 2357 35707
rect 1090 3718 1142 3770
rect 1090 3654 1142 3706
rect 8764 3699 8816 3751
rect 8828 3699 8880 3751
rect 1140 3460 1192 3512
rect 1204 3460 1256 3512
rect 9511 3459 9563 3511
rect 9575 3459 9627 3511
rect 1079 3380 1131 3432
rect 1143 3380 1195 3432
rect 9434 3379 9486 3431
rect 9498 3379 9550 3431
rect 9143 691 9149 710
rect 9149 691 9183 710
rect 9183 691 9195 710
rect 9143 658 9195 691
rect 9602 787 9654 789
rect 9602 753 9611 787
rect 9611 753 9645 787
rect 9645 753 9654 787
rect 9602 737 9654 753
rect 9602 715 9654 725
rect 9602 681 9611 715
rect 9611 681 9645 715
rect 9645 681 9654 715
rect 9602 673 9654 681
rect 9143 619 9149 646
rect 9149 619 9183 646
rect 9183 619 9195 646
rect 9143 594 9195 619
rect 9360 285 9412 337
rect 9445 285 9497 337
<< metal2 >>
rect 1351 39916 2703 39968
rect 2755 39916 2793 39968
rect 2845 39916 2883 39968
rect 2935 39916 2973 39968
rect 3025 39916 3063 39968
rect 3115 39916 3121 39968
rect 1351 39876 3121 39916
rect 1351 39824 2703 39876
rect 2755 39824 2793 39876
rect 2845 39824 2883 39876
rect 2935 39824 2973 39876
rect 3025 39824 3063 39876
rect 3115 39824 3121 39876
rect 1351 39784 3121 39824
rect 1351 39732 2703 39784
rect 2755 39732 2793 39784
rect 2845 39732 2883 39784
rect 2935 39732 2973 39784
rect 3025 39732 3063 39784
rect 3115 39732 3121 39784
tri 1752 39524 1960 39732 nw
rect 954 38664 960 38716
rect 1012 38664 1024 38716
rect 1076 38664 1082 38716
rect 8392 38683 8418 38696
tri 225 37101 359 37235 se
rect 359 37101 457 37152
tri 457 37101 508 37152 nw
tri 173 37049 225 37101 se
rect 225 37049 405 37101
tri 405 37049 457 37101 nw
tri 549 37049 580 37080 se
rect 580 37049 921 37050
tri 161 37037 173 37049 se
rect 173 37037 393 37049
tri 393 37037 405 37049 nw
tri 537 37037 549 37049 se
rect 549 37037 921 37049
tri 157 37033 161 37037 se
rect 161 37033 389 37037
tri 389 37033 393 37037 nw
tri 533 37033 537 37037 se
rect 537 37033 921 37037
rect 157 36985 341 37033
tri 341 36985 389 37033 nw
tri 485 36985 533 37033 se
rect 533 36985 921 37033
rect 157 36074 321 36985
tri 321 36965 341 36985 nw
tri 465 36965 485 36985 se
rect 485 36965 921 36985
rect 209 36022 269 36074
rect 157 35996 321 36022
rect 209 35944 269 35996
rect 157 35917 321 35944
rect 209 35865 269 35917
rect 157 35838 321 35865
rect 209 35786 269 35838
rect 157 35780 321 35786
tri 391 36891 465 36965 se
rect 465 36891 921 36965
rect 391 36528 921 36891
rect 391 36482 875 36528
tri 875 36482 921 36528 nw
rect 391 36430 823 36482
tri 823 36430 875 36482 nw
rect 391 36406 799 36430
tri 799 36406 823 36430 nw
rect 391 36354 747 36406
tri 747 36354 799 36406 nw
rect 391 36079 731 36354
tri 731 36338 747 36354 nw
rect 794 36151 800 36203
rect 852 36151 864 36203
rect 916 36151 922 36203
tri 794 36123 822 36151 ne
rect 391 36027 397 36079
rect 449 36027 489 36079
rect 541 36027 581 36079
rect 633 36027 673 36079
rect 725 36027 731 36079
rect 391 35997 731 36027
rect 391 35945 397 35997
rect 449 35945 489 35997
rect 541 35945 581 35997
rect 633 35945 673 35997
rect 725 35945 731 35997
rect 391 35915 731 35945
rect 391 35863 397 35915
rect 449 35863 489 35915
rect 541 35863 581 35915
rect 633 35863 673 35915
rect 725 35863 731 35915
rect 391 35833 731 35863
rect 391 35781 397 35833
rect 449 35781 489 35833
rect 541 35781 581 35833
rect 633 35781 673 35833
rect 725 35781 731 35833
rect 391 35780 731 35781
rect 822 35669 922 36151
rect 954 7453 986 38664
tri 986 38630 1020 38664 nw
rect 1014 38387 1020 38439
rect 1072 38387 1084 38439
rect 1136 38387 1142 38439
rect 1014 7499 1046 38387
tri 1046 38353 1080 38387 nw
rect 3204 38204 3332 38639
rect 3449 38545 3455 38597
rect 3507 38545 3519 38597
rect 3571 38545 3577 38597
rect 3449 38322 3577 38545
rect 3449 38270 3455 38322
rect 3507 38270 3519 38322
rect 3571 38270 3577 38322
rect 3204 38152 3210 38204
rect 3262 38152 3274 38204
rect 3326 38152 3332 38204
rect 2470 38107 2522 38113
rect 2470 38043 2522 38055
rect 2390 37407 2442 37413
rect 2390 37343 2442 37355
tri 2356 36879 2390 36913 se
rect 2390 36831 2442 37291
tri 2454 36793 2470 36809 se
rect 2470 36793 2522 37991
rect 15848 38051 15914 38057
rect 15848 38048 15862 38051
rect 15848 37992 15853 38048
rect 15909 37992 15914 37999
rect 15848 37987 15914 37992
rect 2774 37907 2780 37959
rect 2832 37907 2844 37959
rect 2896 37907 2902 37959
rect 13588 37929 13594 37981
rect 13646 37929 13660 37981
rect 13712 37929 13718 37981
tri 13632 37916 13645 37929 ne
rect 13645 37916 13718 37929
rect 2774 37891 2902 37907
rect 2774 37839 2780 37891
rect 2832 37839 2844 37891
rect 2896 37839 2902 37891
rect 8335 37894 8463 37916
tri 13645 37895 13666 37916 ne
rect 8335 37842 8341 37894
rect 8393 37842 8405 37894
rect 8457 37842 8463 37894
rect 8335 37839 8463 37842
tri 2017 36779 2031 36793 se
tri 2440 36779 2454 36793 se
rect 2454 36779 2522 36793
rect 1621 36711 2048 36779
tri 2436 36775 2440 36779 se
rect 2440 36775 2522 36779
rect 2470 36728 2522 36775
rect 2550 37664 2556 37716
rect 2608 37664 2620 37716
rect 2672 37664 2678 37716
tri 1587 36207 1621 36241 se
rect 1621 36207 1653 36711
tri 1653 36677 1687 36711 nw
tri 1997 36677 2031 36711 ne
tri 2516 36623 2550 36657 se
rect 2550 36575 2602 37664
tri 2602 37630 2636 37664 nw
rect 2774 37101 2902 37839
rect 4265 37664 4271 37716
rect 4323 37664 4335 37716
rect 4387 37664 4393 37716
rect 3301 37377 3307 37429
rect 3359 37377 3371 37429
rect 3423 37377 3429 37429
tri 3363 37343 3397 37377 ne
rect 2774 37049 2780 37101
rect 2832 37049 2844 37101
rect 2896 37049 2902 37101
rect 2774 37028 2902 37049
tri 3395 36575 3397 36577 se
rect 3397 36575 3429 37377
rect 13666 37317 13718 37916
rect 15848 37968 15862 37987
rect 15848 37912 15853 37968
rect 15909 37912 15914 37935
rect 15848 37903 15914 37912
tri 13666 37265 13718 37317 ne
tri 13718 37287 13770 37339 sw
rect 13718 37265 13770 37287
tri 13718 37213 13770 37265 ne
tri 13770 37213 13844 37287 sw
rect 15184 37213 15187 37244
tri 15187 37213 15218 37244 nw
tri 13770 37139 13844 37213 ne
tri 13844 37139 13918 37213 sw
tri 15184 37210 15187 37213 nw
tri 13844 37117 13866 37139 ne
rect 13866 37101 13918 37139
rect 13866 37037 13918 37049
rect 13866 36979 13918 36985
rect 15721 37101 15777 37107
rect 15721 37091 15723 37101
rect 15775 37091 15777 37101
rect 15721 37011 15723 37035
rect 15775 37011 15777 37035
rect 15721 36946 15777 36955
tri 15184 36845 15218 36879 sw
tri 3363 36543 3395 36575 se
rect 3395 36543 3429 36575
tri 2017 36497 2063 36543 se
rect 2063 36511 3429 36543
tri 2063 36497 2077 36511 nw
tri 2002 36482 2017 36497 se
rect 2017 36482 2048 36497
tri 2048 36482 2063 36497 nw
tri 1971 36451 2002 36482 se
rect 2002 36451 2017 36482
tri 2017 36451 2048 36482 nw
tri 1950 36430 1971 36451 se
rect 1971 36430 1996 36451
tri 1996 36430 2017 36451 nw
rect 2131 36430 2137 36482
rect 2189 36430 2201 36482
rect 2253 36430 2259 36482
tri 1926 36406 1950 36430 se
rect 1950 36406 1972 36430
tri 1972 36406 1996 36430 nw
rect 2131 36406 2259 36430
tri 1925 36405 1926 36406 se
rect 1926 36405 1971 36406
tri 1971 36405 1972 36406 nw
tri 1879 36359 1925 36405 se
tri 1925 36359 1971 36405 nw
tri 1874 36354 1879 36359 se
rect 1879 36354 1920 36359
tri 1920 36354 1925 36359 nw
rect 2131 36354 2137 36406
rect 2189 36354 2201 36406
rect 2253 36354 2259 36406
tri 1833 36313 1874 36354 se
rect 1874 36313 1879 36354
tri 1879 36313 1920 36354 nw
tri 1787 36267 1833 36313 se
tri 1833 36267 1879 36313 nw
tri 1741 36221 1787 36267 se
tri 1787 36221 1833 36267 nw
rect 1074 36175 1653 36207
tri 1695 36175 1741 36221 se
tri 1741 36175 1787 36221 nw
rect 1074 7537 1104 36175
tri 1104 36141 1138 36175 nw
tri 1661 36141 1695 36175 se
rect 1695 36141 1707 36175
tri 1707 36141 1741 36175 nw
tri 1142 36095 1188 36141 se
rect 1188 36109 1675 36141
tri 1675 36109 1707 36141 nw
tri 1188 36095 1202 36109 nw
tri 1133 36086 1142 36095 se
rect 1142 36086 1167 36095
rect 1133 36074 1167 36086
tri 1167 36074 1188 36095 nw
rect 2131 36074 2259 36354
rect 1133 7603 1165 36074
tri 1165 36072 1167 36074 nw
rect 2183 36022 2207 36074
rect 2131 35996 2259 36022
rect 2183 35944 2207 35996
rect 2131 35917 2259 35944
rect 2183 35865 2207 35917
rect 2131 35838 2259 35865
rect 2183 35786 2207 35838
rect 2131 35780 2259 35786
rect 2064 35655 2070 35707
rect 2122 35655 2149 35707
rect 2201 35655 2227 35707
rect 2279 35655 2305 35707
rect 2357 35655 2363 35707
tri 1165 7603 1179 7617 sw
tri 1133 7557 1179 7603 ne
tri 1179 7557 1225 7603 sw
tri 1179 7549 1187 7557 ne
rect 1187 7549 1225 7557
tri 1104 7537 1116 7549 sw
tri 1187 7537 1199 7549 ne
rect 1199 7537 1225 7549
tri 1074 7503 1108 7537 ne
rect 1108 7503 1116 7537
tri 1046 7499 1050 7503 sw
tri 1108 7499 1112 7503 ne
rect 1112 7499 1116 7503
rect 1014 7495 1050 7499
tri 1050 7495 1054 7499 sw
tri 1112 7495 1116 7499 ne
tri 1116 7495 1158 7537 sw
tri 1199 7511 1225 7537 ne
tri 1225 7520 1262 7557 sw
rect 1225 7511 1262 7520
tri 1225 7506 1230 7511 ne
rect 1014 7489 1054 7495
tri 1014 7459 1044 7489 ne
rect 1044 7459 1054 7489
tri 986 7453 992 7459 sw
tri 1044 7453 1050 7459 ne
rect 1050 7453 1054 7459
tri 1054 7453 1096 7495 sw
tri 1116 7453 1158 7495 ne
tri 1158 7482 1171 7495 sw
rect 1158 7453 1171 7482
rect 954 7445 992 7453
tri 954 7413 986 7445 ne
rect 986 7429 992 7445
tri 992 7429 1016 7453 sw
tri 1050 7429 1074 7453 ne
rect 1074 7429 1096 7453
rect 986 7413 1016 7429
tri 986 7383 1016 7413 ne
tri 1016 7407 1038 7429 sw
tri 1074 7407 1096 7429 ne
tri 1096 7407 1142 7453 sw
tri 1158 7440 1171 7453 ne
tri 1171 7452 1201 7482 sw
rect 1016 7383 1038 7407
tri 1038 7383 1062 7407 sw
tri 1096 7393 1110 7407 ne
tri 1016 7369 1030 7383 ne
rect 1030 4044 1062 7383
rect 1110 4285 1142 7407
rect 1171 4377 1201 7452
rect 1230 4518 1262 7511
tri 1262 4518 1287 4543 sw
rect 1230 4486 1287 4518
tri 1230 4461 1255 4486 ne
tri 1201 4377 1226 4402 sw
rect 1171 4363 1226 4377
tri 1171 4338 1196 4363 ne
tri 1142 4285 1167 4310 sw
rect 1110 4253 1167 4285
tri 1110 4228 1135 4253 ne
tri 1110 3943 1135 3968 se
rect 1135 3943 1167 4253
rect 1110 3911 1167 3943
tri 1090 3776 1110 3796 se
rect 1110 3776 1142 3911
tri 1142 3886 1167 3911 nw
rect 1090 3770 1142 3776
rect 1090 3706 1142 3718
rect 1090 3648 1142 3654
tri 1171 3854 1196 3879 se
rect 1196 3854 1226 4363
rect 1171 3824 1226 3854
tri 1129 3595 1171 3637 se
rect 1171 3625 1201 3824
tri 1201 3799 1226 3824 nw
tri 1251 3799 1255 3803 se
rect 1255 3799 1287 4486
tri 1171 3595 1201 3625 nw
tri 1230 3778 1251 3799 se
rect 1251 3778 1287 3799
rect 1230 3746 1287 3778
tri 1087 3553 1129 3595 se
tri 1129 3553 1171 3595 nw
tri 1051 3517 1087 3553 se
rect 1087 3517 1093 3553
tri 1093 3517 1129 3553 nw
tri 1208 3517 1230 3539 se
rect 1230 3517 1262 3746
tri 1262 3721 1287 3746 nw
rect 8758 3699 8764 3751
rect 8816 3699 8828 3751
rect 8880 3699 9689 3751
tri 9606 3644 9661 3699 ne
rect 1051 3512 1088 3517
tri 1088 3512 1093 3517 nw
tri 1203 3512 1208 3517 se
rect 1208 3512 1262 3517
rect 1051 3460 1081 3512
tri 1081 3505 1088 3512 nw
tri 1081 3460 1084 3463 sw
rect 1134 3460 1140 3512
rect 1192 3460 1204 3512
rect 1256 3460 1262 3512
rect 1051 3459 1084 3460
tri 1084 3459 1085 3460 sw
rect 9505 3459 9511 3511
rect 9563 3459 9575 3511
rect 9627 3459 9633 3511
rect 1051 3432 1085 3459
tri 1085 3432 1112 3459 sw
tri 9578 3432 9605 3459 ne
rect 1051 3380 1079 3432
rect 1131 3380 1143 3432
rect 1195 3380 1201 3432
rect 9428 3379 9434 3431
rect 9486 3379 9498 3431
rect 9550 3384 9556 3431
tri 9556 3384 9571 3399 sw
rect 9550 3379 9571 3384
tri 9510 3346 9543 3379 ne
tri 9513 973 9543 1003 se
rect 9543 973 9571 3379
rect 9143 945 9571 973
rect 9143 710 9195 945
tri 9195 911 9229 945 nw
tri 9581 911 9605 935 se
rect 9605 911 9633 3459
tri 9575 905 9581 911 se
rect 9581 905 9633 911
rect 9143 646 9195 658
rect 9143 588 9195 594
rect 9475 877 9633 905
tri 9441 337 9475 371 se
rect 9475 337 9503 877
tri 9503 843 9537 877 nw
tri 9643 843 9661 861 se
rect 9661 843 9689 3699
tri 9627 827 9643 843 se
rect 9643 827 9689 843
rect 9602 795 9689 827
rect 9602 789 9654 795
tri 9654 761 9688 795 nw
rect 9602 725 9654 737
rect 9602 667 9654 673
rect 9354 285 9360 337
rect 9412 285 9445 337
rect 9497 285 9503 337
<< via2 >>
rect 15853 37999 15862 38048
rect 15862 37999 15909 38048
rect 15853 37992 15909 37999
rect 15853 37935 15862 37968
rect 15862 37935 15909 37968
rect 15853 37912 15909 37935
rect 15721 37049 15723 37091
rect 15723 37049 15775 37091
rect 15775 37049 15777 37091
rect 15721 37037 15777 37049
rect 15721 37035 15723 37037
rect 15723 37035 15775 37037
rect 15775 37035 15777 37037
rect 15721 36985 15723 37011
rect 15723 36985 15775 37011
rect 15775 36985 15777 37011
rect 15721 36955 15777 36985
<< metal3 >>
rect 15848 38048 15914 38053
rect 15848 37992 15853 38048
rect 15909 37992 15914 38048
rect 15848 37968 15914 37992
rect 15848 37912 15853 37968
rect 15909 37912 15914 37968
rect 15716 37091 15782 37107
rect 15716 37035 15721 37091
rect 15777 37035 15782 37091
rect 15716 37011 15782 37035
rect 15716 36955 15721 37011
rect 15777 36955 15782 37011
rect 15716 35292 15782 36955
rect 15848 35292 15914 37912
use sky130_fd_io__gpiov2_buf_localesd  sky130_fd_io__gpiov2_buf_localesd_0
timestamp 1704896540
transform -1 0 3161 0 1 36196
box 146 0 3161 3800
use sky130_fd_io__gpiov2_ibuf_se  sky130_fd_io__gpiov2_ibuf_se_0
timestamp 1704896540
transform 1 0 3079 0 1 36000
box -467 -220 12925 4000
use sky130_fd_io__gpiov2_ictl_logic  sky130_fd_io__gpiov2_ictl_logic_0
timestamp 1704896540
transform -1 0 12264 0 -1 1116
box 107 226 3162 873
<< labels >>
flabel metal3 s 15726 35819 15775 36078 3 FreeSans 200 0 0 0 ENABLE_VDDIO_LV
port 1 nsew
flabel metal2 s 824 35975 904 36127 3 FreeSans 400 180 0 0 OUT_H
port 2 nsew
flabel metal2 s 1042 4136 1042 4136 0 FreeSans 200 90 0 0 MODE_VCCHIB_N
flabel metal1 s 10245 704 10245 704 0 FreeSans 200 90 0 0 MODE_VCCHIB_N
flabel metal1 s 15429 39770 15848 39986 3 FreeSans 400 180 0 0 VCCHIB
port 4 nsew
flabel metal1 s 3342 39782 3799 39961 3 FreeSans 400 180 0 0 VDDIO_Q
port 5 nsew
flabel metal1 s 911 35817 1231 36038 3 FreeSans 400 180 0 0 VSSD
port 6 nsew
flabel metal1 s 2702 36238 2938 36301 3 FreeSans 400 180 0 0 PAD
port 7 nsew
flabel metal1 s 15473 37934 15595 38006 3 FreeSans 400 180 0 0 OUT
port 8 nsew
flabel metal1 s 12069 729 12160 763 3 FreeSans 200 0 0 0 DM_H_N[1]
port 9 nsew
flabel metal1 s 11816 725 11876 762 3 FreeSans 200 0 0 0 DM_H_N[0]
port 10 nsew
flabel metal1 s 11416 728 11524 760 3 FreeSans 200 0 0 0 DM_H_N[2]
port 11 nsew
flabel metal1 s 10972 361 11001 477 3 FreeSans 200 0 0 0 INP_DIS_H_N
port 12 nsew
flabel metal1 s 10320 642 10351 759 3 FreeSans 200 0 0 0 IB_MODE_SEL_H
port 13 nsew
flabel metal1 s 9786 678 9818 789 3 FreeSans 200 0 0 0 IB_MODE_SEL_H_N
port 14 nsew
flabel metal1 s 9330 687 9363 788 3 FreeSans 200 0 0 0 VTRIP_SEL_H_N
port 15 nsew
flabel metal1 s 9334 910 9654 1086 3 FreeSans 400 180 0 0 VSSD
port 6 nsew
flabel metal1 s 10366 69 10823 248 3 FreeSans 400 180 0 0 VDDIO_Q
port 5 nsew
flabel comment s 13712 38624 13712 38624 0 FreeSans 440 0 0 0 LV_NET
flabel comment s 1148 35565 1148 35565 0 FreeSans 200 90 0 0 TRIPSEL_I_H_N
flabel comment s 1084 35565 1084 35565 0 FreeSans 200 90 0 0 VTRIP_SEL_H
flabel comment s 1026 35565 1026 35565 0 FreeSans 200 90 0 0 MODE_NORMAL_N
flabel comment s 967 35565 967 35565 0 FreeSans 200 90 0 0 MODE_VCCHIB_N
flabel comment s 15882 35630 15882 35630 0 FreeSans 400 0 0 0 OUT
flabel comment s 15740 35546 15740 35546 0 FreeSans 400 90 0 0 ENABLE_VDDIO_LV
flabel comment s 870 35708 870 35708 0 FreeSans 400 0 0 0 OUT_H
<< properties >>
string GDS_END 17302498
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 17281300
<< end >>
