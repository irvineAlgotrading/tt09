magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -89 -36 189 1036
<< pmos >>
rect 0 0 100 1000
<< pdiff >>
rect -50 0 0 1000
rect 100 0 150 1000
<< poly >>
rect 0 1000 100 1026
rect 0 -26 100 0
<< metal1 >>
rect -51 -16 -5 978
rect 105 -16 151 978
use DFM1sd_CDNS_52468879185574  DFM1sd_CDNS_52468879185574_0
timestamp 1704896540
transform -1 0 0 0 1 0
box -36 -36 89 1036
use DFM1sd_CDNS_52468879185574  DFM1sd_CDNS_52468879185574_1
timestamp 1704896540
transform 1 0 100 0 1 0
box -36 -36 89 1036
<< labels >>
flabel comment s -28 481 -28 481 0 FreeSans 300 0 0 0 S
flabel comment s 128 481 128 481 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 86595954
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86595068
<< end >>
