magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect 1450 -561 1618 347
rect 2656 -561 2824 347
rect 1450 -729 2824 -561
<< pwell >>
rect 1678 -13 2596 73
rect 1678 -415 1764 -13
rect 2510 -415 2596 -13
rect 1678 -501 2596 -415
<< psubdiff >>
rect 1704 31 1822 47
rect 1856 31 1890 47
rect 1924 31 1958 47
rect 1992 31 2026 47
rect 2060 31 2094 47
rect 2128 31 2162 47
rect 2196 31 2230 47
rect 2264 31 2298 47
rect 2332 31 2366 47
rect 2400 31 2434 47
rect 2468 31 2502 47
rect 2536 31 2570 47
<< nsubdiff >>
rect 1518 110 1552 138
rect 1518 39 1552 76
rect 2722 109 2756 138
rect 2722 38 2756 75
<< mvpsubdiff >>
rect 1704 13 1822 31
rect 1856 13 1890 31
rect 1924 13 1958 31
rect 1992 13 2026 31
rect 2060 13 2094 31
rect 2128 13 2162 31
rect 2196 13 2230 31
rect 2264 13 2298 31
rect 2332 13 2366 31
rect 2400 13 2434 31
rect 2468 13 2502 31
rect 1704 -55 1738 -21
rect 1704 -123 1738 -89
rect 2536 -67 2570 31
rect 1704 -191 1738 -157
rect 1704 -259 1738 -225
rect 1704 -327 1738 -293
rect 2536 -135 2570 -101
rect 2536 -203 2570 -169
rect 2536 -271 2570 -237
rect 1704 -475 1738 -361
rect 2536 -339 2570 -305
rect 2536 -407 2570 -373
rect 1772 -475 1890 -441
rect 1924 -475 1958 -441
rect 1992 -475 2026 -441
rect 2060 -475 2094 -441
rect 2128 -475 2162 -441
rect 2196 -475 2230 -441
rect 2264 -475 2298 -441
rect 2332 -475 2366 -441
rect 2400 -475 2434 -441
rect 2468 -475 2570 -441
<< mvnsubdiff >>
rect 1518 181 1552 205
rect 1518 138 1552 147
rect 2722 180 2756 204
rect 2722 138 2756 146
rect 1518 -32 1552 5
rect 1518 -103 1552 -66
rect 1518 -174 1552 -137
rect 1518 -245 1552 -208
rect 1518 -316 1552 -279
rect 1518 -387 1552 -350
rect 1518 -458 1552 -421
rect 2722 -33 2756 4
rect 2722 -104 2756 -67
rect 2722 -175 2756 -138
rect 2722 -246 2756 -209
rect 2722 -317 2756 -280
rect 2722 -388 2756 -351
rect 2722 -459 2756 -422
rect 1518 -529 1552 -492
rect 1518 -627 1552 -563
rect 2722 -531 2756 -493
rect 2722 -603 2756 -565
rect 1518 -661 1542 -627
rect 1576 -661 1610 -627
rect 1644 -661 1678 -627
rect 1712 -661 1746 -627
rect 1780 -661 1814 -627
rect 1848 -661 1882 -627
rect 1916 -661 1950 -627
rect 1984 -661 2018 -627
rect 2052 -661 2086 -627
rect 2120 -661 2154 -627
rect 2188 -661 2222 -627
rect 2256 -661 2290 -627
rect 2324 -661 2358 -627
rect 2392 -661 2426 -627
rect 2460 -661 2494 -627
rect 2528 -661 2562 -627
rect 2596 -661 2630 -627
rect 2664 -637 2722 -627
rect 2664 -661 2756 -637
<< psubdiffcont >>
rect 1822 31 1856 47
rect 1890 31 1924 47
rect 1958 31 1992 47
rect 2026 31 2060 47
rect 2094 31 2128 47
rect 2162 31 2196 47
rect 2230 31 2264 47
rect 2298 31 2332 47
rect 2366 31 2400 47
rect 2434 31 2468 47
rect 2502 31 2536 47
<< nsubdiffcont >>
rect 1518 76 1552 110
rect 2722 75 2756 109
rect 1518 31 1552 39
rect 2722 31 2756 38
<< mvpsubdiffcont >>
rect 1822 13 1856 31
rect 1890 13 1924 31
rect 1958 13 1992 31
rect 2026 13 2060 31
rect 2094 13 2128 31
rect 2162 13 2196 31
rect 2230 13 2264 31
rect 2298 13 2332 31
rect 2366 13 2400 31
rect 2434 13 2468 31
rect 2502 13 2536 31
rect 1704 -21 1738 13
rect 1704 -89 1738 -55
rect 2536 -101 2570 -67
rect 1704 -157 1738 -123
rect 1704 -225 1738 -191
rect 1704 -293 1738 -259
rect 2536 -169 2570 -135
rect 2536 -237 2570 -203
rect 2536 -305 2570 -271
rect 1704 -361 1738 -327
rect 2536 -373 2570 -339
rect 2536 -441 2570 -407
rect 1738 -475 1772 -441
rect 1890 -475 1924 -441
rect 1958 -475 1992 -441
rect 2026 -475 2060 -441
rect 2094 -475 2128 -441
rect 2162 -475 2196 -441
rect 2230 -475 2264 -441
rect 2298 -475 2332 -441
rect 2366 -475 2400 -441
rect 2434 -475 2468 -441
<< mvnsubdiffcont >>
rect 1518 147 1552 181
rect 2722 146 2756 180
rect 1518 5 1552 31
rect 1518 -66 1552 -32
rect 1518 -137 1552 -103
rect 1518 -208 1552 -174
rect 1518 -279 1552 -245
rect 1518 -350 1552 -316
rect 1518 -421 1552 -387
rect 1518 -492 1552 -458
rect 2722 4 2756 31
rect 2722 -67 2756 -33
rect 2722 -138 2756 -104
rect 2722 -209 2756 -175
rect 2722 -280 2756 -246
rect 2722 -351 2756 -317
rect 2722 -422 2756 -388
rect 1518 -563 1552 -529
rect 2722 -493 2756 -459
rect 2722 -565 2756 -531
rect 1542 -661 1576 -627
rect 1610 -661 1644 -627
rect 1678 -661 1712 -627
rect 1746 -661 1780 -627
rect 1814 -661 1848 -627
rect 1882 -661 1916 -627
rect 1950 -661 1984 -627
rect 2018 -661 2052 -627
rect 2086 -661 2120 -627
rect 2154 -661 2188 -627
rect 2222 -661 2256 -627
rect 2290 -661 2324 -627
rect 2358 -661 2392 -627
rect 2426 -661 2460 -627
rect 2494 -661 2528 -627
rect 2562 -661 2596 -627
rect 2630 -661 2664 -627
rect 2722 -637 2756 -603
<< poly >>
rect 1770 -130 1836 -114
rect 1770 -164 1786 -130
rect 1820 -164 1836 -130
rect 1770 -198 1836 -164
rect 1770 -232 1786 -198
rect 1820 -232 1836 -198
rect 1770 -266 1836 -232
rect 1770 -300 1786 -266
rect 1820 -300 1836 -266
rect 1770 -316 1836 -300
<< polycont >>
rect 1786 -164 1820 -130
rect 1786 -232 1820 -198
rect 1786 -300 1820 -266
<< locali >>
rect 2272 4572 2310 4606
rect 2344 4572 2382 4606
rect 2272 246 2310 280
rect 2344 246 2382 280
rect 1518 192 1552 205
rect 1518 118 1552 147
rect 1518 44 1552 76
rect 2722 192 2756 204
rect 2722 117 2756 146
rect 1518 -30 1552 5
rect 1518 -103 1552 -66
rect 1518 -174 1552 -139
rect 1518 -245 1552 -214
rect 1518 -316 1552 -289
rect 1518 -387 1552 -364
rect 1518 -458 1552 -439
rect 1704 13 1822 47
rect 1856 13 1890 47
rect 1924 13 1958 47
rect 1992 13 2026 47
rect 2060 13 2094 47
rect 2128 13 2162 47
rect 2196 13 2230 47
rect 2264 13 2298 47
rect 2332 13 2366 47
rect 2400 13 2434 47
rect 2468 13 2502 47
rect 1704 -43 1738 -21
rect 1704 -123 1738 -89
rect 2536 -48 2570 47
rect 1704 -191 1738 -159
rect 1704 -259 1738 -241
rect 1786 -130 1820 -114
rect 1786 -198 1820 -196
rect 1786 -234 1820 -232
rect 1786 -316 1820 -300
rect 2536 -120 2570 -101
rect 2536 -192 2570 -169
rect 2536 -264 2570 -237
rect 1704 -327 1738 -322
rect 1981 -359 2019 -325
rect 2053 -359 2091 -325
rect 2125 -359 2163 -325
rect 2404 -359 2442 -325
rect 2536 -336 2570 -305
rect 1704 -369 1738 -361
rect 1704 -475 1738 -403
rect 2536 -407 2570 -373
rect 1776 -475 1814 -441
rect 1848 -475 1886 -441
rect 1924 -475 1958 -441
rect 1992 -475 2026 -441
rect 2128 -475 2132 -441
rect 2196 -475 2204 -441
rect 2264 -475 2298 -441
rect 2332 -475 2366 -441
rect 2426 -475 2434 -441
rect 2498 -475 2536 -441
rect 2722 42 2756 75
rect 2722 -33 2756 4
rect 2722 -104 2756 -67
rect 2722 -175 2756 -142
rect 2722 -246 2756 -217
rect 2722 -317 2756 -291
rect 2722 -388 2756 -365
rect 2722 -459 2756 -439
rect 1518 -529 1552 -514
rect 1518 -627 1552 -589
rect 2722 -531 2756 -513
rect 2722 -603 2756 -587
rect 1518 -661 1542 -627
rect 1576 -661 1593 -627
rect 1644 -661 1668 -627
rect 1712 -661 1743 -627
rect 1780 -661 1814 -627
rect 1852 -661 1882 -627
rect 1927 -661 1950 -627
rect 2002 -661 2018 -627
rect 2077 -661 2086 -627
rect 2152 -661 2154 -627
rect 2188 -661 2194 -627
rect 2256 -661 2270 -627
rect 2324 -661 2346 -627
rect 2392 -661 2422 -627
rect 2460 -661 2494 -627
rect 2532 -661 2562 -627
rect 2608 -661 2630 -627
rect 2684 -637 2722 -627
rect 2684 -661 2756 -637
<< viali >>
rect 2238 4572 2272 4606
rect 2310 4572 2344 4606
rect 2382 4572 2416 4606
rect 2238 246 2272 280
rect 2310 246 2344 280
rect 2382 246 2416 280
rect 1518 181 1552 192
rect 1518 158 1552 181
rect 1518 110 1552 118
rect 1518 84 1552 110
rect 2722 180 2756 192
rect 2722 158 2756 180
rect 2722 109 2756 117
rect 2722 83 2756 109
rect 1518 39 1552 44
rect 1518 31 1552 39
rect 1518 10 1552 31
rect 1518 -32 1552 -30
rect 1518 -64 1552 -32
rect 1518 -137 1552 -105
rect 1518 -139 1552 -137
rect 1518 -208 1552 -180
rect 1518 -214 1552 -208
rect 1518 -279 1552 -255
rect 1518 -289 1552 -279
rect 1518 -350 1552 -330
rect 1518 -364 1552 -350
rect 1518 -421 1552 -405
rect 1518 -439 1552 -421
rect 1704 -55 1738 -43
rect 1704 -77 1738 -55
rect 2536 -67 2570 -48
rect 2536 -82 2570 -67
rect 1704 -157 1738 -125
rect 1704 -159 1738 -157
rect 1704 -225 1738 -207
rect 1704 -241 1738 -225
rect 1704 -293 1738 -288
rect 1704 -322 1738 -293
rect 1786 -164 1820 -162
rect 1786 -196 1820 -164
rect 1786 -266 1820 -234
rect 1786 -268 1820 -266
rect 2536 -135 2570 -120
rect 2536 -154 2570 -135
rect 2536 -203 2570 -192
rect 2536 -226 2570 -203
rect 2536 -271 2570 -264
rect 2536 -298 2570 -271
rect 1947 -359 1981 -325
rect 2019 -359 2053 -325
rect 2091 -359 2125 -325
rect 2163 -359 2197 -325
rect 2370 -359 2404 -325
rect 2442 -359 2476 -325
rect 2536 -339 2570 -336
rect 1704 -403 1738 -369
rect 2536 -370 2570 -339
rect 1742 -475 1772 -441
rect 1772 -475 1776 -441
rect 1814 -475 1848 -441
rect 1886 -475 1890 -441
rect 1890 -475 1920 -441
rect 2060 -475 2094 -441
rect 2132 -475 2162 -441
rect 2162 -475 2166 -441
rect 2204 -475 2230 -441
rect 2230 -475 2238 -441
rect 2392 -475 2400 -441
rect 2400 -475 2426 -441
rect 2464 -475 2468 -441
rect 2468 -475 2498 -441
rect 2536 -475 2570 -441
rect 2722 38 2756 42
rect 2722 31 2756 38
rect 2722 8 2756 31
rect 2722 -67 2756 -33
rect 2722 -138 2756 -108
rect 2722 -142 2756 -138
rect 2722 -209 2756 -183
rect 2722 -217 2756 -209
rect 2722 -280 2756 -257
rect 2722 -291 2756 -280
rect 2722 -351 2756 -331
rect 2722 -365 2756 -351
rect 2722 -422 2756 -405
rect 2722 -439 2756 -422
rect 1518 -492 1552 -480
rect 1518 -514 1552 -492
rect 1518 -563 1552 -555
rect 1518 -589 1552 -563
rect 2722 -493 2756 -479
rect 2722 -513 2756 -493
rect 2722 -565 2756 -553
rect 2722 -587 2756 -565
rect 1593 -661 1610 -627
rect 1610 -661 1627 -627
rect 1668 -661 1678 -627
rect 1678 -661 1702 -627
rect 1743 -661 1746 -627
rect 1746 -661 1777 -627
rect 1818 -661 1848 -627
rect 1848 -661 1852 -627
rect 1893 -661 1916 -627
rect 1916 -661 1927 -627
rect 1968 -661 1984 -627
rect 1984 -661 2002 -627
rect 2043 -661 2052 -627
rect 2052 -661 2077 -627
rect 2118 -661 2120 -627
rect 2120 -661 2152 -627
rect 2194 -661 2222 -627
rect 2222 -661 2228 -627
rect 2270 -661 2290 -627
rect 2290 -661 2304 -627
rect 2346 -661 2358 -627
rect 2358 -661 2380 -627
rect 2422 -661 2426 -627
rect 2426 -661 2456 -627
rect 2498 -661 2528 -627
rect 2528 -661 2532 -627
rect 2574 -661 2596 -627
rect 2596 -661 2608 -627
rect 2650 -661 2664 -627
rect 2664 -661 2684 -627
<< metal1 >>
rect 1468 4510 1474 4626
rect 1590 4510 1596 4626
rect 2230 4510 2236 4626
rect 2416 4510 2422 4626
rect 440 4066 446 4182
rect 562 4066 568 4182
rect 1158 4066 1164 4182
rect 1280 4066 1286 4182
rect 1780 4066 1786 4182
rect 1902 4066 1908 4182
rect 2495 4066 2501 4182
rect 2617 4066 2623 4182
rect 2948 4066 2954 4182
rect 3070 4066 3076 4182
rect 645 4032 825 4038
rect 645 3910 825 3916
rect 1977 4032 2157 4038
rect 1977 3910 2157 3916
rect 440 3766 446 3882
rect 562 3766 568 3882
rect 1159 3766 1165 3882
rect 1281 3766 1287 3882
rect 1775 3766 1781 3882
rect 1897 3766 1903 3882
rect 2495 3766 2501 3882
rect 2617 3766 2623 3882
rect 1131 3610 1309 3616
rect 1131 3110 1162 3610
rect 1278 3110 1309 3610
rect 1131 3097 1309 3110
rect 1131 3045 1162 3097
rect 1214 3045 1226 3097
rect 1278 3045 1309 3097
rect 1131 3032 1309 3045
tri 838 2923 895 2980 se
rect 895 2950 1095 3005
rect 895 2876 1021 2950
tri 1021 2876 1095 2950 nw
rect 1131 2980 1162 3032
rect 1214 2980 1226 3032
rect 1278 2980 1309 3032
rect 1131 2967 1309 2980
rect 1131 2915 1162 2967
rect 1214 2915 1226 2967
rect 1278 2915 1309 2967
rect 1131 2902 1309 2915
tri 964 2819 1021 2876 nw
rect 1131 2850 1162 2902
rect 1214 2850 1226 2902
rect 1278 2850 1309 2902
rect 1131 2837 1309 2850
rect 1131 2785 1162 2837
rect 1214 2785 1226 2837
rect 1278 2785 1309 2837
rect 1131 2772 1309 2785
rect 1131 2720 1162 2772
rect 1214 2720 1226 2772
rect 1278 2720 1309 2772
rect 1131 2714 1309 2720
rect 1753 3610 1931 3616
rect 1753 3110 1784 3610
rect 1900 3110 1931 3610
rect 1753 3097 1931 3110
rect 1753 3045 1784 3097
rect 1836 3045 1848 3097
rect 1900 3045 1931 3097
rect 1753 3032 1931 3045
rect 1753 2980 1784 3032
rect 1836 2980 1848 3032
rect 1900 2980 1931 3032
rect 1753 2967 1931 2980
rect 1753 2915 1784 2967
rect 1836 2915 1848 2967
rect 1900 2915 1931 2967
rect 1753 2902 1931 2915
rect 1753 2850 1784 2902
rect 1836 2850 1848 2902
rect 1900 2850 1931 2902
rect 1753 2837 1931 2850
rect 1753 2785 1784 2837
rect 1836 2785 1848 2837
rect 1900 2785 1931 2837
rect 1753 2772 1931 2785
rect 1753 2720 1784 2772
rect 1836 2720 1848 2772
rect 1900 2720 1931 2772
rect 1753 2714 1931 2720
rect 2948 3010 3076 4066
rect 2948 2894 2954 3010
rect 3070 2894 3076 3010
rect 2948 2861 3076 2894
tri 3076 2861 3110 2895 sw
rect 2948 2855 3287 2861
rect 2948 2675 2954 2855
rect 3070 2675 3084 2855
rect 3200 2809 3287 2855
rect 3339 2809 3377 2861
rect 3429 2809 3467 2861
rect 3519 2809 3525 2861
rect 3200 2791 3525 2809
rect 3200 2739 3287 2791
rect 3339 2739 3377 2791
rect 3429 2739 3467 2791
rect 3519 2739 3525 2791
rect 3200 2721 3525 2739
rect 3200 2675 3287 2721
rect 2948 2669 3287 2675
rect 3339 2669 3377 2721
rect 3429 2669 3467 2721
rect 3519 2669 3525 2721
rect 197 2403 223 2452
rect 1518 2415 1544 2437
rect 2839 2404 2865 2453
rect 998 2198 1130 2204
rect 998 2146 1006 2198
rect 1058 2146 1070 2198
rect 1122 2146 1130 2198
rect 998 2099 1130 2146
rect 1932 2198 2064 2204
rect 1932 2146 1940 2198
rect 1992 2146 2004 2198
rect 2056 2146 2064 2198
rect 998 2047 1006 2099
rect 1058 2047 1070 2099
rect 1122 2047 1130 2099
rect 998 2041 1130 2047
rect 1131 2132 1309 2138
rect 1131 2080 1162 2132
rect 1214 2080 1226 2132
rect 1278 2080 1309 2132
rect 1131 2067 1309 2080
tri 964 1976 1021 2033 sw
rect 1131 2015 1162 2067
rect 1214 2015 1226 2067
rect 1278 2015 1309 2067
rect 1131 2002 1309 2015
tri 838 1872 895 1929 ne
rect 895 1902 1021 1976
tri 1021 1902 1095 1976 sw
rect 1131 1950 1162 2002
rect 1214 1950 1226 2002
rect 1278 1950 1309 2002
rect 1131 1944 1309 1950
rect 1753 2132 1931 2138
rect 1753 2080 1784 2132
rect 1836 2080 1848 2132
rect 1900 2080 1931 2132
rect 1753 2067 1931 2080
rect 1753 2015 1784 2067
rect 1836 2015 1848 2067
rect 1900 2015 1931 2067
rect 1932 2099 2064 2146
rect 1932 2047 1940 2099
rect 1992 2047 2004 2099
rect 2056 2047 2064 2099
rect 1932 2041 2064 2047
rect 2281 2179 2483 2203
rect 2281 2127 2287 2179
rect 2339 2127 2356 2179
rect 2408 2127 2425 2179
rect 2477 2127 2483 2179
rect 2281 2115 2483 2127
rect 2281 2063 2287 2115
rect 2339 2063 2356 2115
rect 2408 2063 2425 2115
rect 2477 2063 2483 2115
rect 2281 2039 2483 2063
rect 2488 2132 2628 2138
rect 2488 2080 2500 2132
rect 2552 2080 2564 2132
rect 2616 2080 2628 2132
rect 2488 2067 2628 2080
rect 1753 2002 1931 2015
rect 1753 1950 1784 2002
rect 1836 1950 1848 2002
rect 1900 1950 1931 2002
rect 1753 1944 1931 1950
rect 2488 2015 2500 2067
rect 2552 2015 2564 2067
rect 2616 2015 2628 2067
rect 2488 2002 2628 2015
rect 2488 1950 2500 2002
rect 2552 1950 2564 2002
rect 2616 1950 2628 2002
rect 2488 1944 2628 1950
rect 895 1847 1095 1902
rect 647 1503 827 1509
rect 647 1381 827 1387
rect 1977 1503 2157 1509
rect 1977 1381 2157 1387
rect 2948 1353 3076 2669
tri 3076 2642 3103 2669 nw
rect 3106 2405 3508 2411
rect 3106 2353 3122 2405
rect 3174 2353 3186 2405
rect 3238 2353 3250 2405
rect 3302 2353 3314 2405
rect 3366 2353 3508 2405
rect 3106 2291 3508 2353
rect 3106 2239 3122 2291
rect 3174 2239 3186 2291
rect 3238 2239 3250 2291
rect 3302 2239 3314 2291
rect 3366 2239 3508 2291
rect 3106 2233 3508 2239
rect 3524 1537 3962 1739
rect 439 1237 445 1353
rect 561 1237 567 1353
rect 1167 1237 1173 1353
rect 1289 1237 1295 1353
rect 1780 1237 1786 1353
rect 1902 1237 1908 1353
rect 2499 1237 2505 1353
rect 2621 1237 2627 1353
rect 2948 1237 2954 1353
rect 3070 1237 3076 1353
rect 3524 741 4014 923
rect 1468 227 1474 343
rect 1590 227 1596 343
rect 2230 227 2236 343
rect 2416 227 2422 343
tri 1461 192 1473 204 ne
rect 1473 192 1589 204
tri 1589 192 1601 204 nw
tri 1473 158 1507 192 ne
rect 1507 158 1518 192
rect 1552 158 1558 192
tri 1558 161 1589 192 nw
tri 1507 153 1512 158 ne
rect 1512 118 1558 158
rect 1512 84 1518 118
rect 1552 84 1558 118
rect 1512 44 1558 84
rect 1967 146 2167 204
tri 2652 192 2664 204 ne
rect 2664 192 2762 204
tri 2664 158 2698 192 ne
rect 2698 158 2722 192
rect 2756 158 2762 192
tri 2762 188 2778 204 nw
rect 1967 94 1973 146
rect 2025 94 2041 146
rect 2093 94 2109 146
rect 2161 94 2167 146
tri 2698 140 2716 158 ne
rect 1967 81 2167 94
rect 2716 117 2762 158
rect 2716 83 2722 117
rect 2756 83 2762 117
tri 2296 53 2302 59 se
rect 1512 10 1518 44
rect 1552 10 1558 44
rect 1512 -30 1558 10
rect 1512 -64 1518 -30
rect 1552 -64 1558 -30
rect 1512 -105 1558 -64
rect 1512 -139 1518 -105
rect 1552 -139 1558 -105
rect 1512 -180 1558 -139
rect 1512 -214 1518 -180
rect 1552 -214 1558 -180
rect 1512 -255 1558 -214
rect 1512 -289 1518 -255
rect 1552 -289 1558 -255
rect 1512 -330 1558 -289
rect 1512 -364 1518 -330
rect 1552 -364 1558 -330
rect 1512 -405 1558 -364
rect 1512 -439 1518 -405
rect 1552 -439 1558 -405
rect 1512 -480 1558 -439
rect 1512 -514 1518 -480
rect 1552 -514 1558 -480
rect 1698 45 1714 53
rect 1698 -43 1744 45
rect 2302 7 2308 59
rect 2360 7 2380 59
rect 2432 7 2452 59
rect 2504 7 2524 59
rect 2576 7 2582 59
tri 1744 -31 1782 7 nw
tri 2492 -31 2530 7 ne
rect 1698 -77 1704 -43
rect 1738 -77 1744 -43
rect 2530 -48 2582 7
rect 1698 -125 1744 -77
rect 1913 -112 2228 -60
rect 2280 -112 2292 -60
rect 2344 -112 2356 -60
rect 2408 -112 2420 -60
rect 2472 -112 2478 -60
rect 2530 -82 2536 -48
rect 2570 -82 2582 -48
rect 1698 -159 1704 -125
rect 1738 -159 1744 -125
rect 2530 -120 2582 -82
rect 1698 -207 1744 -159
rect 1698 -241 1704 -207
rect 1738 -241 1744 -207
rect 1698 -288 1744 -241
rect 1777 -157 2424 -150
rect 1777 -162 2369 -157
rect 1777 -196 1786 -162
rect 1820 -196 2369 -162
rect 1777 -209 2369 -196
rect 2421 -209 2424 -157
rect 1777 -221 2424 -209
rect 1777 -234 2369 -221
rect 1777 -268 1786 -234
rect 1820 -268 2369 -234
rect 1777 -273 2369 -268
rect 2421 -273 2424 -221
rect 1777 -280 2424 -273
rect 2530 -154 2536 -120
rect 2570 -154 2582 -120
rect 2530 -192 2582 -154
rect 2530 -226 2536 -192
rect 2570 -226 2582 -192
rect 2530 -264 2582 -226
rect 1698 -322 1704 -288
rect 1738 -322 1744 -288
rect 2530 -298 2536 -264
rect 2570 -298 2582 -264
rect 1698 -369 1744 -322
rect 1897 -368 1903 -316
rect 1955 -325 1967 -316
rect 2019 -325 2031 -316
rect 2083 -325 2095 -316
rect 2083 -359 2091 -325
rect 1955 -368 1967 -359
rect 2019 -368 2031 -359
rect 2083 -368 2095 -359
rect 2147 -368 2159 -316
rect 2211 -368 2217 -316
rect 2358 -368 2364 -316
rect 2416 -368 2428 -316
rect 2480 -368 2488 -316
rect 2530 -336 2582 -298
rect 1698 -403 1704 -369
rect 1738 -403 1744 -369
rect 2530 -370 2536 -336
rect 2570 -370 2582 -336
rect 1698 -405 1744 -403
tri 1744 -405 1752 -397 sw
tri 2522 -405 2530 -397 se
rect 2530 -405 2582 -370
rect 1698 -435 1752 -405
tri 1752 -435 1782 -405 sw
tri 2492 -435 2522 -405 se
rect 2522 -435 2582 -405
rect 1698 -441 1753 -435
rect 1805 -441 1817 -435
rect 1698 -475 1742 -441
rect 1805 -475 1814 -441
rect 1698 -487 1753 -475
rect 1805 -487 1817 -475
rect 1869 -487 1881 -435
rect 1933 -487 1940 -435
rect 2048 -487 2058 -435
rect 2110 -487 2122 -435
rect 2174 -487 2186 -435
rect 2238 -487 2250 -435
rect 2358 -487 2364 -435
rect 2416 -441 2428 -435
rect 2480 -441 2582 -435
rect 2426 -475 2428 -441
rect 2498 -475 2536 -441
rect 2570 -475 2582 -441
rect 2416 -487 2428 -475
rect 2480 -487 2582 -475
rect 2716 42 2762 83
rect 2716 8 2722 42
rect 2756 8 2762 42
rect 2716 -33 2762 8
rect 2716 -67 2722 -33
rect 2756 -67 2762 -33
rect 2716 -108 2762 -67
rect 2716 -142 2722 -108
rect 2756 -142 2762 -108
rect 2716 -183 2762 -142
rect 2716 -217 2722 -183
rect 2756 -217 2762 -183
rect 2716 -257 2762 -217
rect 2716 -291 2722 -257
rect 2756 -291 2762 -257
rect 2716 -331 2762 -291
rect 2716 -365 2722 -331
rect 2756 -365 2762 -331
rect 2716 -405 2762 -365
rect 2716 -439 2722 -405
rect 2756 -439 2762 -405
rect 2716 -479 2762 -439
rect 1512 -555 1558 -514
rect 2716 -513 2722 -479
rect 2756 -513 2762 -479
tri 2685 -553 2716 -522 se
rect 2716 -553 2762 -513
tri 2684 -554 2685 -553 se
rect 2685 -554 2722 -553
rect 1512 -589 1518 -555
rect 1552 -587 1558 -555
tri 1558 -587 1591 -554 sw
tri 2651 -587 2684 -554 se
rect 2684 -587 2722 -554
rect 2756 -587 2762 -553
rect 1552 -589 1591 -587
rect 1512 -621 1591 -589
tri 1591 -621 1625 -587 sw
tri 2617 -621 2651 -587 se
rect 2651 -621 2762 -587
rect 1512 -627 2762 -621
rect 1512 -661 1593 -627
rect 1627 -661 1668 -627
rect 1702 -661 1743 -627
rect 1777 -661 1818 -627
rect 1852 -661 1893 -627
rect 1927 -661 1968 -627
rect 2002 -661 2043 -627
rect 2077 -661 2118 -627
rect 2152 -661 2194 -627
rect 2228 -661 2270 -627
rect 2304 -661 2346 -627
rect 2380 -661 2422 -627
rect 2456 -661 2498 -627
rect 2532 -661 2574 -627
rect 2608 -661 2650 -627
rect 2684 -661 2762 -627
rect 1512 -667 2762 -661
rect 3106 -589 3508 -37
rect 3106 -641 3112 -589
rect 3164 -641 3197 -589
rect 3249 -641 3282 -589
rect 3334 -641 3366 -589
rect 3418 -641 3450 -589
rect 3502 -641 3508 -589
rect 3106 -657 3508 -641
rect 3106 -709 3112 -657
rect 3164 -709 3197 -657
rect 3249 -709 3282 -657
rect 3334 -709 3366 -657
rect 3418 -709 3450 -657
rect 3502 -709 3508 -657
rect 3106 -713 3508 -709
<< via1 >>
rect 1474 4510 1590 4626
rect 2236 4606 2416 4626
rect 2236 4572 2238 4606
rect 2238 4572 2272 4606
rect 2272 4572 2310 4606
rect 2310 4572 2344 4606
rect 2344 4572 2382 4606
rect 2382 4572 2416 4606
rect 2236 4510 2416 4572
rect 446 4066 562 4182
rect 1164 4066 1280 4182
rect 1786 4066 1902 4182
rect 2501 4066 2617 4182
rect 2954 4066 3070 4182
rect 645 3916 825 4032
rect 1977 3916 2157 4032
rect 446 3766 562 3882
rect 1165 3766 1281 3882
rect 1781 3766 1897 3882
rect 2501 3766 2617 3882
rect 1162 3110 1278 3610
rect 1162 3045 1214 3097
rect 1226 3045 1278 3097
rect 1162 2980 1214 3032
rect 1226 2980 1278 3032
rect 1162 2915 1214 2967
rect 1226 2915 1278 2967
rect 1162 2850 1214 2902
rect 1226 2850 1278 2902
rect 1162 2785 1214 2837
rect 1226 2785 1278 2837
rect 1162 2720 1214 2772
rect 1226 2720 1278 2772
rect 1784 3110 1900 3610
rect 1784 3045 1836 3097
rect 1848 3045 1900 3097
rect 1784 2980 1836 3032
rect 1848 2980 1900 3032
rect 1784 2915 1836 2967
rect 1848 2915 1900 2967
rect 1784 2850 1836 2902
rect 1848 2850 1900 2902
rect 1784 2785 1836 2837
rect 1848 2785 1900 2837
rect 1784 2720 1836 2772
rect 1848 2720 1900 2772
rect 2954 2894 3070 3010
rect 2954 2675 3070 2855
rect 3084 2675 3200 2855
rect 3287 2809 3339 2861
rect 3377 2809 3429 2861
rect 3467 2809 3519 2861
rect 3287 2739 3339 2791
rect 3377 2739 3429 2791
rect 3467 2739 3519 2791
rect 3287 2669 3339 2721
rect 3377 2669 3429 2721
rect 3467 2669 3519 2721
rect 1006 2146 1058 2198
rect 1070 2146 1122 2198
rect 1940 2146 1992 2198
rect 2004 2146 2056 2198
rect 1006 2047 1058 2099
rect 1070 2047 1122 2099
rect 1162 2080 1214 2132
rect 1226 2080 1278 2132
rect 1162 2015 1214 2067
rect 1226 2015 1278 2067
rect 1162 1950 1214 2002
rect 1226 1950 1278 2002
rect 1784 2080 1836 2132
rect 1848 2080 1900 2132
rect 1784 2015 1836 2067
rect 1848 2015 1900 2067
rect 1940 2047 1992 2099
rect 2004 2047 2056 2099
rect 2287 2127 2339 2179
rect 2356 2127 2408 2179
rect 2425 2127 2477 2179
rect 2287 2063 2339 2115
rect 2356 2063 2408 2115
rect 2425 2063 2477 2115
rect 2500 2080 2552 2132
rect 2564 2080 2616 2132
rect 1784 1950 1836 2002
rect 1848 1950 1900 2002
rect 2500 2015 2552 2067
rect 2564 2015 2616 2067
rect 2500 1950 2552 2002
rect 2564 1950 2616 2002
rect 647 1387 827 1503
rect 1977 1387 2157 1503
rect 3122 2353 3174 2405
rect 3186 2353 3238 2405
rect 3250 2353 3302 2405
rect 3314 2353 3366 2405
rect 3122 2239 3174 2291
rect 3186 2239 3238 2291
rect 3250 2239 3302 2291
rect 3314 2239 3366 2291
rect 445 1237 561 1353
rect 1173 1237 1289 1353
rect 1786 1237 1902 1353
rect 2505 1237 2621 1353
rect 2954 1237 3070 1353
rect 1474 227 1590 343
rect 2236 280 2416 343
rect 2236 246 2238 280
rect 2238 246 2272 280
rect 2272 246 2310 280
rect 2310 246 2344 280
rect 2344 246 2382 280
rect 2382 246 2416 280
rect 2236 227 2416 246
rect 1973 94 2025 146
rect 2041 94 2093 146
rect 2109 94 2161 146
rect 2308 7 2360 59
rect 2380 7 2432 59
rect 2452 7 2504 59
rect 2524 7 2576 59
rect 2228 -112 2280 -60
rect 2292 -112 2344 -60
rect 2356 -112 2408 -60
rect 2420 -112 2472 -60
rect 2369 -209 2421 -157
rect 2369 -273 2421 -221
rect 1903 -325 1955 -316
rect 1967 -325 2019 -316
rect 2031 -325 2083 -316
rect 2095 -325 2147 -316
rect 1903 -359 1947 -325
rect 1947 -359 1955 -325
rect 1967 -359 1981 -325
rect 1981 -359 2019 -325
rect 2031 -359 2053 -325
rect 2053 -359 2083 -325
rect 2095 -359 2125 -325
rect 2125 -359 2147 -325
rect 1903 -368 1955 -359
rect 1967 -368 2019 -359
rect 2031 -368 2083 -359
rect 2095 -368 2147 -359
rect 2159 -325 2211 -316
rect 2159 -359 2163 -325
rect 2163 -359 2197 -325
rect 2197 -359 2211 -325
rect 2159 -368 2211 -359
rect 2364 -325 2416 -316
rect 2364 -359 2370 -325
rect 2370 -359 2404 -325
rect 2404 -359 2416 -325
rect 2364 -368 2416 -359
rect 2428 -325 2480 -316
rect 2428 -359 2442 -325
rect 2442 -359 2476 -325
rect 2476 -359 2480 -325
rect 2428 -368 2480 -359
rect 1753 -441 1805 -435
rect 1817 -441 1869 -435
rect 1753 -475 1776 -441
rect 1776 -475 1805 -441
rect 1817 -475 1848 -441
rect 1848 -475 1869 -441
rect 1753 -487 1805 -475
rect 1817 -487 1869 -475
rect 1881 -441 1933 -435
rect 1881 -475 1886 -441
rect 1886 -475 1920 -441
rect 1920 -475 1933 -441
rect 1881 -487 1933 -475
rect 2058 -441 2110 -435
rect 2058 -475 2060 -441
rect 2060 -475 2094 -441
rect 2094 -475 2110 -441
rect 2058 -487 2110 -475
rect 2122 -441 2174 -435
rect 2122 -475 2132 -441
rect 2132 -475 2166 -441
rect 2166 -475 2174 -441
rect 2122 -487 2174 -475
rect 2186 -441 2238 -435
rect 2186 -475 2204 -441
rect 2204 -475 2238 -441
rect 2186 -487 2238 -475
rect 2364 -441 2416 -435
rect 2428 -441 2480 -435
rect 2364 -475 2392 -441
rect 2392 -475 2416 -441
rect 2428 -475 2464 -441
rect 2464 -475 2480 -441
rect 2364 -487 2416 -475
rect 2428 -487 2480 -475
rect 3112 -641 3164 -589
rect 3197 -641 3249 -589
rect 3282 -641 3334 -589
rect 3366 -641 3418 -589
rect 3450 -641 3502 -589
rect 3112 -709 3164 -657
rect 3197 -709 3249 -657
rect 3282 -709 3334 -657
rect 3366 -709 3418 -657
rect 3450 -709 3502 -657
<< metal2 >>
rect 0 -221 120 4667
rect 596 4510 1474 4626
rect 1590 4510 2236 4626
rect 2416 4510 2541 4626
rect 440 4066 446 4182
rect 562 4066 1164 4182
rect 1280 4066 1786 4182
rect 1902 4066 2501 4182
rect 2617 4066 2954 4182
rect 3070 4066 3076 4182
rect 148 4032 3233 4038
rect 148 3916 645 4032
rect 825 3916 1977 4032
rect 2157 3916 3233 4032
rect 148 3910 3233 3916
rect 148 2015 403 3910
tri 403 3885 428 3910 nw
rect 440 3766 446 3882
rect 562 3766 1165 3882
rect 1281 3766 1781 3882
rect 1897 3766 2501 3882
rect 2617 3766 3076 3882
tri 2922 3740 2948 3766 ne
rect 826 3610 2667 3616
rect 826 3110 1162 3610
rect 1278 3110 1784 3610
rect 1900 3110 2667 3610
rect 826 3097 2667 3110
rect 826 3045 1162 3097
rect 1214 3045 1226 3097
rect 1278 3045 1784 3097
rect 1836 3045 1848 3097
rect 1900 3045 2667 3097
rect 826 3032 2667 3045
rect 826 2980 1162 3032
rect 1214 2980 1226 3032
rect 1278 2980 1784 3032
rect 1836 2980 1848 3032
rect 1900 2980 2667 3032
rect 826 2967 2667 2980
rect 826 2915 1162 2967
rect 1214 2915 1226 2967
rect 1278 2915 1784 2967
rect 1836 2915 1848 2967
rect 1900 2915 2667 2967
rect 826 2902 2667 2915
rect 826 2850 1162 2902
rect 1214 2850 1226 2902
rect 1278 2850 1784 2902
rect 1836 2850 1848 2902
rect 1900 2850 2667 2902
rect 826 2837 2667 2850
rect 826 2785 1162 2837
rect 1214 2785 1226 2837
rect 1278 2785 1784 2837
rect 1836 2785 1848 2837
rect 1900 2785 2667 2837
rect 826 2772 2667 2785
rect 826 2720 1162 2772
rect 1214 2720 1226 2772
rect 1278 2720 1784 2772
rect 1836 2720 1848 2772
rect 1900 2720 2667 2772
rect 826 2291 2667 2720
rect 2948 3010 3076 3766
rect 2948 2894 2954 3010
rect 3070 2894 3076 3010
rect 2948 2861 3076 2894
tri 3076 2861 3285 3070 sw
rect 2948 2855 3287 2861
rect 2948 2675 2954 2855
rect 3070 2675 3084 2855
rect 3200 2809 3287 2855
rect 3339 2809 3377 2861
rect 3429 2809 3467 2861
rect 3519 2809 3525 2861
rect 3200 2791 3525 2809
rect 3200 2739 3287 2791
rect 3339 2739 3377 2791
rect 3429 2739 3467 2791
rect 3519 2739 3525 2791
rect 3200 2721 3525 2739
rect 3200 2675 3287 2721
rect 2948 2669 3287 2675
rect 3339 2669 3377 2721
rect 3429 2669 3467 2721
rect 3519 2669 3525 2721
rect 2948 2556 3525 2669
tri 2667 2291 2704 2328 sw
tri 2932 2291 2948 2307 se
rect 2948 2291 3066 2556
tri 3066 2456 3166 2556 nw
tri 3309 2456 3409 2556 ne
rect 3409 2456 3525 2556
tri 3409 2411 3454 2456 ne
rect 3454 2411 3525 2456
rect 826 2252 2704 2291
tri 2704 2252 2743 2291 sw
tri 2893 2252 2932 2291 se
rect 2932 2252 3066 2291
rect 3106 2405 3412 2411
rect 3106 2353 3122 2405
rect 3174 2353 3186 2405
rect 3238 2353 3250 2405
rect 3302 2353 3314 2405
rect 3366 2353 3412 2405
rect 3106 2291 3412 2353
tri 3454 2341 3524 2411 ne
rect 3524 2383 3525 2411
tri 3525 2383 3768 2626 sw
rect 826 2198 3066 2252
tri 3066 2246 3076 2256 sw
rect 826 2146 1006 2198
rect 1058 2146 1070 2198
rect 1122 2146 1940 2198
rect 1992 2146 2004 2198
rect 2056 2179 3066 2198
rect 2056 2146 2287 2179
rect 826 2132 2287 2146
rect 826 2099 1162 2132
rect 826 2047 1006 2099
rect 1058 2047 1070 2099
rect 1122 2080 1162 2099
rect 1214 2080 1226 2132
rect 1278 2080 1784 2132
rect 1836 2080 1848 2132
rect 1900 2127 2287 2132
rect 2339 2127 2356 2179
rect 2408 2127 2425 2179
rect 2477 2132 3066 2179
rect 2477 2127 2500 2132
rect 1900 2115 2500 2127
rect 1900 2099 2287 2115
rect 1900 2080 1940 2099
rect 1122 2067 1940 2080
rect 1122 2047 1162 2067
tri 403 2015 425 2037 sw
rect 826 2015 1162 2047
rect 1214 2015 1226 2067
rect 1278 2015 1784 2067
rect 1836 2015 1848 2067
rect 1900 2047 1940 2067
rect 1992 2047 2004 2099
rect 2056 2063 2287 2099
rect 2339 2063 2356 2115
rect 2408 2063 2425 2115
rect 2477 2080 2500 2115
rect 2552 2080 2564 2132
rect 2616 2080 3066 2132
rect 2477 2067 3066 2080
rect 2477 2063 2500 2067
rect 2056 2047 2500 2063
rect 1900 2015 2500 2047
rect 2552 2015 2564 2067
rect 2616 2066 3066 2067
rect 3106 2239 3122 2291
rect 3174 2239 3186 2291
rect 3238 2239 3250 2291
rect 3302 2239 3314 2291
rect 3366 2239 3412 2291
rect 2616 2015 2976 2066
rect 148 2002 425 2015
tri 425 2002 438 2015 sw
rect 826 2002 2976 2015
rect 148 1950 438 2002
tri 438 1950 490 2002 sw
rect 826 1950 1162 2002
rect 1214 1950 1226 2002
rect 1278 1950 1784 2002
rect 1836 1950 1848 2002
rect 1900 1950 2500 2002
rect 2552 1950 2564 2002
rect 2616 1985 2976 2002
tri 2976 1985 3057 2066 nw
tri 3057 1985 3106 2034 se
rect 3106 1985 3412 2239
rect 2616 1950 2935 1985
rect 148 1888 490 1950
tri 490 1888 552 1950 sw
rect 826 1944 2935 1950
tri 2935 1944 2976 1985 nw
tri 3016 1944 3057 1985 se
rect 3057 1944 3412 1985
tri 2960 1888 3016 1944 se
rect 3016 1888 3412 1944
rect 148 1571 3412 1888
rect 148 1537 3378 1571
tri 3378 1537 3412 1571 nw
rect 647 1503 2375 1509
rect 827 1387 1977 1503
rect 2157 1387 2375 1503
rect 647 1381 2375 1387
rect 437 1237 445 1353
rect 561 1237 1173 1353
rect 1289 1237 1786 1353
rect 1902 1237 2505 1353
rect 2621 1237 2954 1353
rect 3070 1237 3076 1353
rect 3524 900 3768 2383
tri 3068 343 3157 432 ne
rect 3157 393 3189 432
rect 3157 343 3299 393
rect 596 227 1474 343
rect 1590 227 2236 343
rect 2416 227 2541 343
tri 3157 313 3187 343 ne
tri 3183 159 3187 163 se
rect 3187 159 3299 343
tri 3299 271 3420 392 nw
rect 1967 146 2167 159
rect 1967 94 1973 146
rect 2025 94 2041 146
rect 2093 94 2109 146
rect 2161 94 2167 146
tri 3139 115 3183 159 se
rect 3183 115 3299 159
rect 1967 -209 2167 94
rect 2302 59 3299 115
rect 2302 7 2308 59
rect 2360 7 2380 59
rect 2432 7 2452 59
rect 2504 7 2524 59
rect 2576 7 3299 59
rect 2302 3 3299 7
tri 3575 3 3591 19 se
tri 3512 -60 3575 3 se
rect 3575 -60 3591 3
rect 2222 -112 2228 -60
rect 2280 -112 2292 -60
rect 2344 -112 2356 -60
rect 2408 -112 2420 -60
rect 2472 -63 3591 -60
rect 2472 -112 3643 -63
rect 2369 -157 3643 -151
tri 2167 -209 2179 -197 sw
rect 2421 -209 3643 -157
tri 120 -221 130 -211 sw
rect 1967 -221 2179 -209
tri 2179 -221 2191 -209 sw
rect 2369 -221 3643 -209
rect 0 -261 130 -221
tri 130 -261 170 -221 sw
tri 1952 -261 1967 -246 se
rect 1967 -261 2191 -221
tri 0 -273 12 -261 ne
rect 12 -273 170 -261
tri 170 -273 182 -261 sw
tri 1940 -273 1952 -261 se
rect 1952 -273 2191 -261
tri 2191 -273 2243 -221 sw
rect 2421 -273 3643 -221
tri 12 -316 55 -273 ne
rect 55 -316 182 -273
tri 182 -316 225 -273 sw
tri 1897 -316 1940 -273 se
rect 1940 -316 2243 -273
tri 2243 -316 2286 -273 sw
rect 2369 -279 3643 -273
tri 55 -368 107 -316 ne
rect 107 -368 225 -316
tri 225 -368 277 -316 sw
rect 1897 -368 1903 -316
rect 1955 -368 1967 -316
rect 2019 -368 2031 -316
rect 2083 -368 2095 -316
rect 2147 -368 2159 -316
rect 2211 -368 2364 -316
rect 2416 -368 2428 -316
rect 2480 -368 3643 -316
tri 107 -431 170 -368 ne
rect 170 -431 277 -368
tri 277 -431 340 -368 sw
tri 3515 -431 3578 -368 ne
rect 3578 -431 3591 -368
tri 170 -435 174 -431 ne
rect 174 -435 340 -431
tri 340 -435 344 -431 sw
tri 3578 -435 3582 -431 ne
rect 3582 -435 3591 -431
tri 174 -487 226 -435 ne
rect 226 -487 344 -435
tri 344 -487 396 -435 sw
rect 1747 -487 1753 -435
rect 1805 -487 1817 -435
rect 1869 -487 1881 -435
rect 1933 -487 2058 -435
rect 2110 -487 2122 -435
rect 2174 -487 2186 -435
rect 2238 -487 2364 -435
rect 2416 -487 2428 -435
rect 2480 -487 2486 -435
tri 3582 -444 3591 -435 ne
tri 226 -589 328 -487 ne
rect 328 -589 396 -487
tri 396 -589 498 -487 sw
tri 328 -601 340 -589 ne
rect 340 -601 3112 -589
tri 340 -641 380 -601 ne
rect 380 -641 3112 -601
rect 3164 -641 3197 -589
rect 3249 -641 3282 -589
rect 3334 -641 3366 -589
rect 3418 -641 3450 -589
rect 3502 -641 3508 -589
tri 380 -657 396 -641 ne
rect 396 -657 3508 -641
tri 396 -709 448 -657 ne
rect 448 -709 3112 -657
rect 3164 -709 3197 -657
rect 3249 -709 3282 -657
rect 3334 -709 3366 -657
rect 3418 -709 3450 -657
rect 3502 -709 3508 -657
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1704896540
transform 0 -1 1820 -1 0 -162
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1704896540
transform -1 0 2476 0 -1 -325
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1704896540
transform -1 0 2570 0 1 -475
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_1
timestamp 1704896540
transform 1 0 1742 0 1 -475
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_2
timestamp 1704896540
transform 1 0 2060 0 1 -475
box 0 0 1 1
use L1M1_CDNS_52468879185191  L1M1_CDNS_52468879185191_0
timestamp 1704896540
transform 1 0 1726 0 1 13
box -12 -6 838 40
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_0
timestamp 1704896540
transform 0 1 2238 -1 0 4606
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_1
timestamp 1704896540
transform 0 1 2238 -1 0 280
box 0 0 1 1
use L1M1_CDNS_52468879185193  L1M1_CDNS_52468879185193_0
timestamp 1704896540
transform 0 -1 2570 -1 0 -48
box 0 0 1 1
use L1M1_CDNS_52468879185195  L1M1_CDNS_52468879185195_0
timestamp 1704896540
transform 1 0 1925 0 -1 -69
box -12 -6 550 40
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_0
timestamp 1704896540
transform 1 0 1947 0 -1 -325
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1704896540
transform -1 0 2486 0 -1 -435
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_1
timestamp 1704896540
transform -1 0 2486 0 -1 -316
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_2
timestamp 1704896540
transform 0 1 2369 1 0 -279
box 0 0 1 1
use M1M2_CDNS_52468879185197  M1M2_CDNS_52468879185197_0
timestamp 1704896540
transform -1 0 2721 0 1 4510
box 0 0 256 116
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_0
timestamp 1704896540
transform 0 1 3084 -1 0 2861
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_1
timestamp 1704896540
transform 1 0 2230 0 1 227
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_2
timestamp 1704896540
transform 1 0 2230 0 1 4510
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_0
timestamp 1704896540
transform -1 0 1295 0 -1 1353
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_1
timestamp 1704896540
transform -1 0 2627 0 -1 1353
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_2
timestamp 1704896540
transform 1 0 1775 0 -1 3882
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_3
timestamp 1704896540
transform 1 0 2948 0 -1 1353
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_4
timestamp 1704896540
transform 1 0 1159 0 -1 3882
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_5
timestamp 1704896540
transform 1 0 1780 0 -1 1353
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_6
timestamp 1704896540
transform 1 0 440 0 -1 3882
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_7
timestamp 1704896540
transform 1 0 2495 0 -1 3882
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_8
timestamp 1704896540
transform 1 0 1780 0 -1 4182
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_9
timestamp 1704896540
transform 1 0 1158 0 -1 4182
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_10
timestamp 1704896540
transform 1 0 440 0 -1 4182
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_11
timestamp 1704896540
transform 1 0 439 0 -1 1353
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_12
timestamp 1704896540
transform 1 0 2948 0 -1 3010
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_13
timestamp 1704896540
transform 1 0 2948 0 1 4066
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_14
timestamp 1704896540
transform 1 0 2495 0 1 4066
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_15
timestamp 1704896540
transform 1 0 1468 0 1 4510
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_16
timestamp 1704896540
transform 1 0 1468 0 1 227
box 0 0 1 1
use M1M2_CDNS_52468879185200  M1M2_CDNS_52468879185200_0
timestamp 1704896540
transform 0 1 1977 1 0 3910
box 0 0 1 1
use M1M2_CDNS_52468879185200  M1M2_CDNS_52468879185200_1
timestamp 1704896540
transform 0 1 1977 1 0 1381
box 0 0 1 1
use M1M2_CDNS_52468879185200  M1M2_CDNS_52468879185200_2
timestamp 1704896540
transform 0 1 645 1 0 3910
box 0 0 1 1
use M1M2_CDNS_52468879185200  M1M2_CDNS_52468879185200_3
timestamp 1704896540
transform 0 1 647 1 0 1381
box 0 0 1 1
use M1M2_CDNS_52468879185201  M1M2_CDNS_52468879185201_0
timestamp 1704896540
transform -1 0 596 0 1 4510
box 0 0 320 116
use M1M2_CDNS_52468879185201  M1M2_CDNS_52468879185201_1
timestamp 1704896540
transform -1 0 596 0 1 227
box 0 0 320 116
use M1M2_CDNS_52468879185201  M1M2_CDNS_52468879185201_2
timestamp 1704896540
transform -1 0 2787 0 1 227
box 0 0 320 116
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_0
timestamp 1704896540
transform 1 0 1897 0 -1 -316
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_0
timestamp 1704896540
transform -1 0 2244 0 -1 -435
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_1
timestamp 1704896540
transform -1 0 1939 0 -1 -435
box 0 0 1 1
use M1M2_CDNS_52468879185205  M1M2_CDNS_52468879185205_0
timestamp 1704896540
transform 1 0 2948 0 1 3247
box 0 0 128 628
use M1M2_CDNS_52468879185206  M1M2_CDNS_52468879185206_0
timestamp 1704896540
transform 1 0 826 0 1 1944
box 0 0 128 948
use M1M2_CDNS_52468879185206  M1M2_CDNS_52468879185206_1
timestamp 1704896540
transform 1 0 2108 0 1 1944
box 0 0 128 948
use M1M2_CDNS_52468879185207  M1M2_CDNS_52468879185207_0
timestamp 1704896540
transform 1 0 899 0 -1 3616
box 0 0 192 692
use M1M2_CDNS_52468879185208  M1M2_CDNS_52468879185208_0
timestamp 1704896540
transform 0 1 3524 -1 0 1733
box 0 0 192 244
use M1M2_CDNS_52468879185209  M1M2_CDNS_52468879185209_0
timestamp 1704896540
transform 0 1 3524 -1 0 900
box 0 0 128 244
use M1M2_CDNS_52468879185297  M1M2_CDNS_52468879185297_0
timestamp 1704896540
transform -1 0 2478 0 -1 -60
box 0 0 1 1
use nfet_CDNS_52468879185210  nfet_CDNS_52468879185210_0
timestamp 1704896540
transform 0 -1 2462 1 0 -314
box -79 -26 279 626
use PYL1_CDNS_52468879185136  PYL1_CDNS_52468879185136_0
timestamp 1704896540
transform -1 0 1836 0 -1 -114
box 0 0 1 1
use s8_esd_res250only_small  s8_esd_res250only_small_0
timestamp 1704896540
transform 0 -1 3509 1 0 -37
box 0 0 2270 404
use s8_esd_signal_5_sym_hv_local_5term  s8_esd_signal_5_sym_hv_local_5term_0
timestamp 1704896540
transform -1 0 1667 0 1 138
box 0 0 1591 2424
use s8_esd_signal_5_sym_hv_local_5term  s8_esd_signal_5_sym_hv_local_5term_1
timestamp 1704896540
transform -1 0 1667 0 -1 4714
box 0 0 1591 2424
use s8_esd_signal_5_sym_hv_local_5term  s8_esd_signal_5_sym_hv_local_5term_2
timestamp 1704896540
transform 1 0 1395 0 -1 4714
box 0 0 1591 2424
use s8_esd_signal_5_sym_hv_local_5term  s8_esd_signal_5_sym_hv_local_5term_3
timestamp 1704896540
transform 1 0 1395 0 1 138
box 0 0 1591 2424
<< labels >>
flabel comment s 59 4554 59 4554 0 FreeSans 200 0 0 0 Pad
flabel metal1 s 3106 -149 3508 -129 3 FreeSans 520 0 0 0 in_h
port 2 nsew
flabel metal1 s 3952 1537 3962 1739 7 FreeSans 200 0 0 0 vgnd
port 3 nsew
flabel metal2 s 3592 -368 3643 -316 3 FreeSans 520 180 0 0 out_vt
port 4 nsew
flabel metal2 s 3592 -109 3643 -63 3 FreeSans 520 180 0 0 out_h
port 5 nsew
flabel metal2 s 1424 4525 1635 4597 0 FreeSans 200 0 0 0 vcc_io
port 6 nsew
flabel metal2 s 3592 -279 3643 -151 0 FreeSans 200 270 0 0 vtrip_sel_h
port 7 nsew
<< properties >>
string GDS_END 85875670
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85848746
string path 49.175 3.000 54.175 3.000 
<< end >>
