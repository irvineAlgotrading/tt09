magic
tech sky130A
timestamp 1704896540
<< properties >>
string GDS_END 89696170
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 89695910
<< end >>
