magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< obsli1 >>
rect 80 719 214 735
rect 80 685 94 719
rect 128 685 166 719
rect 200 685 214 719
rect 80 667 214 685
rect 44 605 78 621
rect 44 533 78 571
rect 44 461 78 499
rect 44 389 78 427
rect 44 317 78 355
rect 44 245 78 283
rect 44 173 78 211
rect 44 101 78 139
rect 44 47 78 67
rect 130 51 164 621
rect 216 605 250 621
rect 216 533 250 571
rect 216 461 250 499
rect 216 389 250 427
rect 216 317 250 355
rect 216 245 250 283
rect 216 173 250 211
rect 216 101 250 139
rect 216 51 250 67
<< obsli1c >>
rect 94 685 128 719
rect 166 685 200 719
rect 44 571 78 605
rect 44 499 78 533
rect 44 427 78 461
rect 44 355 78 389
rect 44 283 78 317
rect 44 211 78 245
rect 44 139 78 173
rect 44 67 78 101
rect 216 571 250 605
rect 216 499 250 533
rect 216 427 250 461
rect 216 355 250 389
rect 216 283 250 317
rect 216 211 250 245
rect 216 139 250 173
rect 216 67 250 101
<< metal1 >>
rect 82 719 212 731
rect 82 685 94 719
rect 128 685 166 719
rect 200 685 212 719
rect 82 673 212 685
rect 38 605 84 621
rect 38 571 44 605
rect 78 571 84 605
rect 38 533 84 571
rect 38 499 44 533
rect 78 499 84 533
rect 38 461 84 499
rect 38 427 44 461
rect 78 427 84 461
rect 38 389 84 427
rect 38 355 44 389
rect 78 355 84 389
rect 38 317 84 355
rect 38 283 44 317
rect 78 283 84 317
rect 38 245 84 283
rect 38 211 44 245
rect 78 211 84 245
rect 38 173 84 211
rect 38 139 44 173
rect 78 139 84 173
rect 38 101 84 139
rect 38 67 44 101
rect 78 67 84 101
rect 38 -29 84 67
rect 210 605 256 621
rect 210 571 216 605
rect 250 571 256 605
rect 210 533 256 571
rect 210 499 216 533
rect 250 499 256 533
rect 210 461 256 499
rect 210 427 216 461
rect 250 427 256 461
rect 210 389 256 427
rect 210 355 216 389
rect 250 355 256 389
rect 210 317 256 355
rect 210 283 216 317
rect 250 283 256 317
rect 210 245 256 283
rect 210 211 216 245
rect 250 211 256 245
rect 210 173 256 211
rect 210 139 216 173
rect 250 139 256 173
rect 210 101 256 139
rect 210 67 216 101
rect 250 67 256 101
rect 210 -29 256 67
rect 38 -89 256 -29
<< obsm1 >>
rect 121 51 173 621
<< metal2 >>
rect 121 488 173 616
<< labels >>
rlabel metal2 s 121 488 173 616 6 DRAIN
port 1 nsew
rlabel metal1 s 82 673 212 731 6 GATE
port 2 nsew
rlabel metal1 s 210 -29 256 621 6 SOURCE
port 3 nsew
rlabel metal1 s 38 -29 84 621 6 SOURCE
port 3 nsew
rlabel metal1 s 38 -89 256 -29 8 SOURCE
port 3 nsew
<< properties >>
string FIXED_BBOX 0 -89 294 735
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 10417414
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 10411090
string device primitive
<< end >>
