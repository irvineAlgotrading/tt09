magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -89 -36 217 1036
<< pmos >>
rect 0 0 36 1000
rect 92 0 128 1000
<< pdiff >>
rect -50 0 0 1000
rect 128 0 178 1000
<< poly >>
rect 0 1000 36 1026
rect 0 -26 36 0
rect 92 1000 128 1026
rect 92 -26 128 0
<< locali >>
rect -45 -4 -11 946
rect 47 -4 81 946
rect 139 -4 173 946
use DFL1sd2_CDNS_52468879185113  DFL1sd2_CDNS_52468879185113_0
timestamp 1704896540
transform 1 0 36 0 1 0
box -36 -36 92 1036
use DFL1sd_CDNS_52468879185122  DFL1sd_CDNS_52468879185122_0
timestamp 1704896540
transform -1 0 0 0 1 0
box -36 -36 89 1036
use DFL1sd_CDNS_52468879185122  DFL1sd_CDNS_52468879185122_1
timestamp 1704896540
transform 1 0 128 0 1 0
box -36 -36 89 1036
<< labels >>
flabel comment s -28 471 -28 471 0 FreeSans 300 0 0 0 S
flabel comment s 64 471 64 471 0 FreeSans 300 0 0 0 D
flabel comment s 156 471 156 471 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 85794410
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85793026
<< end >>
