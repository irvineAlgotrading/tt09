magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< pwell >>
rect -76 -26 724 1026
<< mvnmos >>
rect 0 0 120 1000
rect 176 0 296 1000
rect 352 0 472 1000
rect 528 0 648 1000
<< mvndiff >>
rect -50 0 0 1000
rect 648 0 698 1000
<< poly >>
rect 0 1000 120 1026
rect 0 -26 120 0
rect 176 1000 296 1026
rect 176 -26 296 0
rect 352 1000 472 1026
rect 352 -26 472 0
rect 528 1000 648 1026
rect 528 -26 648 0
<< locali >>
rect -45 -4 -11 946
rect 131 -4 165 946
rect 307 -4 341 946
rect 483 -4 517 946
rect 659 -4 693 946
use hvDFL1sd2_CDNS_524688791858  hvDFL1sd2_CDNS_524688791858_0
timestamp 1704896540
transform 1 0 472 0 1 0
box -26 -26 82 1026
use hvDFL1sd2_CDNS_524688791858  hvDFL1sd2_CDNS_524688791858_1
timestamp 1704896540
transform 1 0 296 0 1 0
box -26 -26 82 1026
use hvDFL1sd2_CDNS_524688791858  hvDFL1sd2_CDNS_524688791858_2
timestamp 1704896540
transform 1 0 120 0 1 0
box -26 -26 82 1026
use hvDFL1sd_CDNS_5246887918592  hvDFL1sd_CDNS_5246887918592_0
timestamp 1704896540
transform -1 0 0 0 1 0
box -26 -26 79 1026
use hvDFL1sd_CDNS_5246887918592  hvDFL1sd_CDNS_5246887918592_1
timestamp 1704896540
transform 1 0 648 0 1 0
box -26 -26 79 1026
<< labels >>
flabel comment s -28 471 -28 471 0 FreeSans 300 0 0 0 S
flabel comment s 148 471 148 471 0 FreeSans 300 0 0 0 D
flabel comment s 324 471 324 471 0 FreeSans 300 0 0 0 S
flabel comment s 500 471 500 471 0 FreeSans 300 0 0 0 D
flabel comment s 676 471 676 471 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 87828158
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 87825774
<< end >>
