magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 1 21 643 203
rect 27 -17 61 21
<< locali >>
rect 18 337 71 491
rect 18 53 85 337
rect 205 199 261 265
rect 297 199 412 265
rect 448 199 535 265
rect 571 199 625 265
<< obsli1 >>
rect 0 527 644 561
rect 105 383 171 527
rect 209 419 261 491
rect 295 453 361 527
rect 395 419 447 491
rect 209 373 447 419
rect 561 337 619 491
rect 120 301 619 337
rect 120 163 165 301
rect 120 125 617 163
rect 121 17 270 91
rect 383 53 434 125
rect 470 17 536 91
rect 572 53 617 125
rect 0 -17 644 17
<< metal1 >>
rect 0 496 644 592
rect 0 -48 644 48
<< labels >>
rlabel locali s 297 199 412 265 6 A1
port 1 nsew signal input
rlabel locali s 205 199 261 265 6 A2
port 2 nsew signal input
rlabel locali s 448 199 535 265 6 B1
port 3 nsew signal input
rlabel locali s 571 199 625 265 6 C1
port 4 nsew signal input
rlabel metal1 s 0 -48 644 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 27 -17 61 21 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1 21 643 203 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 682 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 644 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 18 53 85 337 6 X
port 9 nsew signal output
rlabel locali s 18 337 71 491 6 X
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 644 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3627924
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3621578
<< end >>
