magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< locali >>
rect 11923 32808 11954 32846
rect 18056 32815 18086 32844
rect 18234 32813 18269 32838
rect 18234 32803 18242 32813
rect 16799 32751 16831 32795
rect 16965 32758 16996 32798
rect 18216 32779 18242 32781
rect 18420 32797 18456 32833
rect 18276 32779 18282 32781
rect 18216 32741 18282 32779
rect 19211 32744 19267 32788
rect 18216 32707 18242 32741
rect 18276 32707 18282 32741
<< viali >>
rect 18242 32779 18276 32813
rect 18242 32707 18276 32741
<< metal1 >>
rect 18522 33471 19108 33673
rect 17266 33331 17272 33383
rect 17324 33331 17336 33383
rect 17388 33331 17394 33383
rect 17875 33269 18003 33399
tri 27460 33067 27488 33095 ne
rect 18228 32814 18282 32825
rect 18280 32762 18282 32814
rect 18228 32750 18282 32762
rect 18280 32698 18282 32750
rect 18228 32692 18282 32698
rect 11513 32365 11551 32404
rect 18581 32317 19176 32472
tri 27665 32197 27695 32227 ne
rect 27695 32197 27698 32227
rect 27140 32164 27192 32197
tri 27695 32194 27698 32197 ne
tri 27750 32194 27783 32227 nw
rect 19853 31506 19905 31512
rect 19853 31442 19905 31454
rect 19853 31384 19905 31390
rect 24432 30637 24634 30679
rect 25923 30641 26053 30683
rect 26335 30641 26537 30683
rect 26861 30641 27063 30683
rect 27575 30646 27721 30683
rect 27321 30418 27352 30562
tri 26781 29926 26787 29932 se
rect 26787 29926 26833 30165
rect 26781 29920 26833 29926
tri 27359 29893 27365 29899 nw
rect 26781 29856 26833 29868
rect 26781 29798 26833 29804
rect 24184 29706 24386 29748
rect 27091 24877 27137 24917
rect 27091 24740 27137 24781
rect 26721 23039 26752 23133
rect 27171 22975 27217 23015
rect 27289 22777 27335 22823
rect 26650 22321 26674 22407
rect 27289 21535 27335 21581
rect 25465 20856 25511 20902
rect 27247 20545 27293 20585
rect 25923 17881 26053 17923
rect 26335 17905 26537 17947
rect 24184 17775 24386 17817
rect 24710 17775 24912 17817
rect 25307 17775 25437 17817
rect 26861 17775 27063 17817
rect 27575 17775 27721 17812
<< via1 >>
rect 17272 33331 17324 33383
rect 17336 33331 17388 33383
rect 18228 32813 18280 32814
rect 18228 32779 18242 32813
rect 18242 32779 18276 32813
rect 18276 32779 18280 32813
rect 18228 32762 18280 32779
rect 18228 32741 18280 32750
rect 18228 32707 18242 32741
rect 18242 32707 18276 32741
rect 18276 32707 18280 32741
rect 18228 32698 18280 32707
rect 19853 31454 19905 31506
rect 19853 31390 19905 31442
rect 26781 29868 26833 29920
rect 26781 29804 26833 29856
<< metal2 >>
rect 11274 33500 11643 33685
rect 17260 33453 17269 33509
rect 17325 33453 17349 33509
rect 17405 33453 17414 33509
rect 17266 33383 17394 33453
tri 17394 33433 17414 33453 nw
rect 17266 33331 17272 33383
rect 17324 33331 17336 33383
rect 17388 33331 17394 33383
rect 20036 33327 20045 33383
rect 20101 33327 20125 33383
rect 20181 33327 20190 33383
tri 20037 33322 20042 33327 ne
tri 15704 33201 15760 33257 se
rect 15760 33201 16206 33257
rect 16262 33201 16307 33257
rect 16363 33201 16408 33257
rect 16464 33201 16473 33257
tri 15658 33155 15704 33201 se
rect 15704 33155 15736 33201
tri 15736 33155 15782 33201 nw
tri 15580 33077 15658 33155 se
tri 15658 33077 15736 33155 nw
tri 15811 33077 15865 33131 se
rect 15865 33077 16206 33131
tri 15502 32999 15580 33077 se
tri 15580 32999 15658 33077 nw
tri 15787 33053 15811 33077 se
rect 15811 33075 16206 33077
rect 16262 33075 16307 33131
rect 16363 33075 16408 33131
rect 16464 33075 16473 33131
rect 15811 33053 15865 33075
tri 15865 33053 15887 33075 nw
tri 15733 32999 15787 33053 se
tri 15424 32921 15502 32999 se
tri 15502 32921 15580 32999 nw
tri 15709 32975 15733 32999 se
rect 15733 32975 15787 32999
tri 15787 32975 15865 33053 nw
tri 15655 32921 15709 32975 se
tri 15402 32899 15424 32921 se
rect 14766 32843 14775 32899
rect 14831 32843 14876 32899
rect 14932 32843 14977 32899
rect 15033 32843 15424 32899
tri 15424 32843 15502 32921 nw
tri 15631 32897 15655 32921 se
rect 15655 32897 15709 32921
tri 15709 32897 15787 32975 nw
tri 15577 32843 15631 32897 se
tri 15553 32819 15577 32843 se
rect 15577 32819 15631 32843
tri 15631 32819 15709 32897 nw
rect 16933 32823 16942 32879
rect 16998 32823 17022 32879
rect 17078 32823 17087 32879
tri 15548 32814 15553 32819 se
rect 15553 32814 15626 32819
tri 15626 32814 15631 32819 nw
tri 15507 32773 15548 32814 se
rect 15548 32773 15585 32814
tri 15585 32773 15626 32814 nw
rect 16951 32805 17003 32823
rect 18228 32814 18280 32820
rect 14766 32717 14775 32773
rect 14831 32717 14876 32773
rect 14932 32717 14977 32773
rect 15033 32762 15574 32773
tri 15574 32762 15585 32773 nw
rect 15033 32750 15562 32762
tri 15562 32750 15574 32762 nw
rect 18228 32753 18280 32762
rect 15033 32717 15529 32750
tri 15529 32717 15562 32750 nw
rect 18129 32697 18138 32753
rect 18194 32697 18218 32753
rect 18274 32750 18283 32753
rect 18280 32698 18283 32750
rect 18274 32697 18283 32698
rect 18228 32692 18280 32697
tri 19968 31516 20042 31590 se
rect 20042 31516 20097 33327
tri 20097 33292 20132 33327 nw
rect 19853 31506 20097 31516
rect 19905 31454 20097 31506
rect 19853 31442 20097 31454
rect 19905 31390 20097 31442
rect 19853 31384 20097 31390
rect 24402 29926 24458 29929
tri 24458 29926 24461 29929 sw
rect 24402 29920 26833 29926
tri 23413 29868 23418 29873 sw
rect 23413 29856 23418 29868
tri 23418 29856 23430 29868 sw
rect 24458 29868 26781 29920
rect 24458 29864 26833 29868
rect 24402 29856 26833 29864
rect 23413 29842 23430 29856
tri 23430 29842 23444 29856 sw
rect 24402 29840 26781 29856
tri 23409 29751 23443 29785 ne
rect 24458 29804 26781 29840
rect 24458 29798 26833 29804
rect 24402 29775 24458 29784
tri 24458 29775 24481 29798 nw
rect 2214 29431 2333 29489
rect 5497 29432 5506 29488
rect 5562 29432 5586 29488
rect 5642 29432 5651 29488
rect 2028 29282 2200 29364
rect 5291 29332 5300 29388
rect 5356 29332 5380 29388
rect 5436 29332 5445 29388
rect 4839 28595 4994 28884
rect 18919 27043 19027 27411
rect 22701 27039 22809 27407
rect 26693 23756 26745 23808
rect 25722 23272 25873 23315
rect 25032 21231 25088 21240
rect 25032 21151 25088 21175
rect 25032 21086 25088 21095
rect 25159 21137 25465 21146
rect 25215 21081 25465 21137
rect 25159 21057 25465 21081
rect 25215 21018 25465 21057
rect 25159 20992 25215 21001
rect 24780 20822 24836 20831
rect 25098 20781 25150 20828
rect 24780 20742 24836 20766
rect 24780 20677 24836 20686
rect 26781 20301 26833 20359
tri 27553 20199 27585 20231 ne
rect 24906 20105 24962 20114
tri 24962 20081 24995 20114 sw
rect 24962 20064 26751 20081
tri 26751 20064 26768 20081 sw
tri 27573 20064 27585 20076 se
rect 27585 20064 27671 20231
tri 27671 20199 27703 20231 nw
rect 24962 20049 26768 20064
rect 24906 20025 26768 20049
rect 24962 19995 26768 20025
rect 24906 19960 24962 19969
tri 24962 19961 24996 19995 nw
tri 26715 19961 26749 19995 ne
rect 26749 19961 26768 19995
tri 26749 19960 26750 19961 ne
rect 26750 19960 26768 19961
tri 26750 19942 26768 19960 ne
tri 26768 19942 26890 20064 sw
tri 27463 19954 27573 20064 se
rect 27573 20040 27671 20064
rect 27573 19954 27585 20040
tri 27585 19954 27671 20040 nw
tri 27451 19942 27463 19954 se
rect 27463 19942 27487 19954
tri 26768 19856 26854 19942 ne
rect 26854 19856 27487 19942
tri 27487 19856 27585 19954 nw
tri 24644 18588 24654 18598 se
rect 24654 18589 24710 18598
tri 24710 18588 24720 18598 sw
tri 25406 18588 25410 18592 se
rect 25410 18588 25468 18592
tri 25468 18588 25472 18592 sw
rect 24654 18509 24710 18533
tri 24638 18444 24654 18460 ne
tri 25376 18460 25388 18472 ne
rect 25388 18460 25410 18472
rect 24654 18444 24710 18453
tri 24710 18444 24726 18460 nw
tri 25388 18444 25404 18460 ne
rect 25404 18444 25410 18460
tri 25404 18438 25410 18444 ne
tri 25466 18438 25500 18472 nw
rect 26621 17940 26673 17987
<< via2 >>
rect 17269 33453 17325 33509
rect 17349 33453 17405 33509
rect 20045 33327 20101 33383
rect 20125 33327 20181 33383
rect 16206 33201 16262 33257
rect 16307 33201 16363 33257
rect 16408 33201 16464 33257
rect 16206 33075 16262 33131
rect 16307 33075 16363 33131
rect 16408 33075 16464 33131
rect 14775 32843 14831 32899
rect 14876 32843 14932 32899
rect 14977 32843 15033 32899
rect 16942 32823 16998 32879
rect 17022 32823 17078 32879
rect 14775 32717 14831 32773
rect 14876 32717 14932 32773
rect 14977 32717 15033 32773
rect 18138 32697 18194 32753
rect 18218 32750 18274 32753
rect 18218 32698 18228 32750
rect 18228 32698 18274 32750
rect 18218 32697 18274 32698
rect 24402 29864 24458 29920
rect 24402 29784 24458 29840
rect 5506 29432 5562 29488
rect 5586 29432 5642 29488
rect 5300 29332 5356 29388
rect 5380 29332 5436 29388
rect 25032 21175 25088 21231
rect 25032 21095 25088 21151
rect 25159 21081 25215 21137
rect 25159 21001 25215 21057
rect 24780 20766 24836 20822
rect 24780 20686 24836 20742
rect 24906 20049 24962 20105
rect 24906 19969 24962 20025
rect 24654 18533 24710 18589
rect 24654 18453 24710 18509
<< metal3 >>
rect 17264 33509 23690 33514
rect 17264 33453 17269 33509
rect 17325 33453 17349 33509
rect 17405 33488 23690 33509
tri 23690 33488 23716 33514 sw
rect 17405 33453 23716 33488
rect 17264 33448 23716 33453
tri 23662 33394 23716 33448 ne
tri 23716 33394 23810 33488 sw
tri 23716 33388 23722 33394 ne
rect 23722 33388 23810 33394
rect 20040 33383 23635 33388
rect 20040 33327 20045 33383
rect 20101 33327 20125 33383
rect 20181 33340 23635 33383
tri 23635 33340 23683 33388 sw
tri 23722 33340 23770 33388 ne
rect 23770 33340 23810 33388
rect 20181 33327 23683 33340
rect 20040 33322 23683 33327
tri 23607 33262 23667 33322 ne
rect 23667 33307 23683 33322
tri 23683 33307 23716 33340 sw
tri 23770 33307 23803 33340 ne
rect 23803 33307 23810 33340
rect 23667 33262 23716 33307
rect 16183 33257 23581 33262
rect 16183 33201 16206 33257
rect 16262 33201 16307 33257
rect 16363 33201 16408 33257
rect 16464 33246 23581 33257
tri 23581 33246 23597 33262 sw
tri 23667 33246 23683 33262 ne
rect 23683 33246 23716 33262
tri 23716 33246 23777 33307 sw
tri 23803 33300 23810 33307 ne
tri 23810 33300 23904 33394 sw
tri 23810 33246 23864 33300 ne
rect 23864 33246 23904 33300
rect 16464 33201 23597 33246
rect 16183 33196 23597 33201
tri 23553 33168 23581 33196 ne
rect 23581 33192 23597 33196
tri 23597 33192 23651 33246 sw
tri 23683 33192 23737 33246 ne
rect 23737 33213 23777 33246
tri 23777 33213 23810 33246 sw
tri 23864 33213 23897 33246 ne
rect 23897 33213 23904 33246
rect 23737 33192 23810 33213
rect 23581 33184 23651 33192
tri 23651 33184 23659 33192 sw
tri 23737 33184 23745 33192 ne
rect 23745 33184 23810 33192
rect 23581 33168 23659 33184
tri 23581 33136 23613 33168 ne
rect 23613 33136 23659 33168
rect 16183 33131 23527 33136
rect 16183 33075 16206 33131
rect 16262 33075 16307 33131
rect 16363 33075 16408 33131
rect 16464 33130 23527 33131
tri 23527 33130 23533 33136 sw
tri 23613 33130 23619 33136 ne
rect 23619 33130 23659 33136
rect 16464 33098 23533 33130
tri 23533 33098 23565 33130 sw
tri 23619 33098 23651 33130 ne
rect 23651 33098 23659 33130
tri 23659 33098 23745 33184 sw
tri 23745 33152 23777 33184 ne
rect 23777 33152 23810 33184
tri 23810 33152 23871 33213 sw
tri 23897 33206 23904 33213 ne
tri 23904 33206 23998 33300 sw
tri 23904 33152 23958 33206 ne
rect 23958 33152 23998 33206
tri 23777 33098 23831 33152 ne
rect 23831 33119 23871 33152
tri 23871 33119 23904 33152 sw
tri 23958 33119 23991 33152 ne
rect 23991 33119 23998 33152
rect 23831 33098 23904 33119
rect 16464 33075 23565 33098
rect 16183 33070 23565 33075
tri 23499 33042 23527 33070 ne
rect 23527 33044 23565 33070
tri 23565 33044 23619 33098 sw
tri 23651 33044 23705 33098 ne
rect 23705 33090 23745 33098
tri 23745 33090 23753 33098 sw
tri 23831 33090 23839 33098 ne
rect 23839 33090 23904 33098
rect 23705 33044 23753 33090
rect 23527 33042 23619 33044
tri 23527 33010 23559 33042 ne
rect 23559 33036 23619 33042
tri 23619 33036 23627 33044 sw
tri 23705 33036 23713 33044 ne
rect 23713 33036 23753 33044
rect 23559 33010 23627 33036
rect 16649 32990 23473 33010
tri 23473 32990 23493 33010 sw
tri 23559 32990 23579 33010 ne
rect 23579 32990 23627 33010
rect 16649 32956 23493 32990
tri 23493 32956 23527 32990 sw
tri 23579 32956 23613 32990 ne
rect 23613 32956 23627 32990
rect 16649 32944 23527 32956
tri 23445 32904 23485 32944 ne
rect 23485 32904 23527 32944
tri 5608 32899 5613 32904 se
rect 5613 32899 15041 32904
tri 5552 32843 5608 32899 se
rect 5608 32843 14775 32899
rect 14831 32843 14876 32899
rect 14932 32843 14977 32899
rect 15033 32843 15041 32899
tri 23485 32896 23493 32904 ne
rect 23493 32896 23527 32904
tri 23527 32896 23587 32956 sw
tri 23613 32950 23619 32956 ne
rect 23619 32950 23627 32956
tri 23627 32950 23713 33036 sw
tri 23713 33004 23745 33036 ne
rect 23745 33004 23753 33036
tri 23753 33004 23839 33090 sw
tri 23839 33058 23871 33090 ne
rect 23871 33058 23904 33090
tri 23904 33058 23965 33119 sw
tri 23991 33112 23998 33119 ne
tri 23998 33112 24092 33206 sw
tri 23998 33058 24052 33112 ne
rect 24052 33058 24092 33112
tri 23871 33004 23925 33058 ne
rect 23925 33025 23965 33058
tri 23965 33025 23998 33058 sw
tri 24052 33025 24085 33058 ne
rect 24085 33025 24092 33058
rect 23925 33004 23998 33025
tri 23745 32950 23799 33004 ne
rect 23799 32996 23839 33004
tri 23839 32996 23847 33004 sw
tri 23925 32996 23933 33004 ne
rect 23933 32996 23998 33004
rect 23799 32950 23847 32996
tri 23619 32896 23673 32950 ne
rect 23673 32942 23713 32950
tri 23713 32942 23721 32950 sw
tri 23799 32942 23807 32950 ne
rect 23807 32942 23847 32950
rect 23673 32896 23721 32942
tri 23493 32884 23505 32896 ne
rect 23505 32884 23587 32896
tri 5532 32823 5552 32843 se
rect 5552 32838 15041 32843
rect 16937 32879 23419 32884
rect 5552 32823 5660 32838
tri 5660 32823 5675 32838 nw
rect 16937 32823 16942 32879
rect 16998 32823 17022 32879
rect 17078 32842 23419 32879
tri 23419 32842 23461 32884 sw
tri 23505 32842 23547 32884 ne
rect 23547 32864 23587 32884
tri 23587 32864 23619 32896 sw
tri 23673 32864 23705 32896 ne
rect 23705 32864 23721 32896
rect 23547 32842 23619 32864
rect 17078 32823 23461 32842
tri 5485 32776 5532 32823 se
rect 5532 32776 5613 32823
tri 5613 32776 5660 32823 nw
rect 16937 32818 23461 32823
tri 23391 32778 23431 32818 ne
rect 23431 32810 23461 32818
tri 23461 32810 23493 32842 sw
tri 23547 32810 23579 32842 ne
rect 23579 32810 23619 32842
rect 23431 32778 23493 32810
tri 5747 32776 5749 32778 se
rect 5749 32776 15041 32778
tri 5482 32773 5485 32776 se
rect 5485 32773 5610 32776
tri 5610 32773 5613 32776 nw
tri 5744 32773 5747 32776 se
rect 5747 32773 15041 32776
tri 5426 32717 5482 32773 se
rect 5482 32761 5598 32773
tri 5598 32761 5610 32773 nw
tri 5732 32761 5744 32773 se
rect 5744 32761 14775 32773
rect 5482 32717 5554 32761
tri 5554 32717 5598 32761 nw
tri 5688 32717 5732 32761 se
rect 5732 32717 14775 32761
rect 14831 32717 14876 32773
rect 14932 32717 14977 32773
rect 15033 32717 15041 32773
tri 23431 32758 23451 32778 ne
rect 23451 32758 23493 32778
tri 5406 32697 5426 32717 se
rect 5426 32697 5534 32717
tri 5534 32697 5554 32717 nw
tri 5683 32712 5688 32717 se
rect 5688 32712 15041 32717
rect 18133 32753 23365 32758
tri 5668 32697 5683 32712 se
rect 5683 32697 5819 32712
tri 5819 32697 5834 32712 nw
rect 18133 32697 18138 32753
rect 18194 32697 18218 32753
rect 18274 32748 23365 32753
tri 23365 32748 23375 32758 sw
tri 23451 32748 23461 32758 ne
rect 23461 32748 23493 32758
tri 23493 32748 23555 32810 sw
tri 23579 32802 23587 32810 ne
rect 23587 32802 23619 32810
tri 23619 32802 23681 32864 sw
tri 23705 32856 23713 32864 ne
rect 23713 32856 23721 32864
tri 23721 32856 23807 32942 sw
tri 23807 32910 23839 32942 ne
rect 23839 32910 23847 32942
tri 23847 32910 23933 32996 sw
tri 23933 32964 23965 32996 ne
rect 23965 32964 23998 32996
tri 23998 32964 24059 33025 sw
tri 24085 33018 24092 33025 ne
tri 24092 33018 24186 33112 sw
tri 24092 32964 24146 33018 ne
rect 24146 32964 24186 33018
tri 23965 32910 24019 32964 ne
rect 24019 32931 24059 32964
tri 24059 32931 24092 32964 sw
tri 24146 32931 24179 32964 ne
rect 24179 32931 24186 32964
rect 24019 32910 24092 32931
tri 23839 32856 23893 32910 ne
rect 23893 32902 23933 32910
tri 23933 32902 23941 32910 sw
tri 24019 32902 24027 32910 ne
rect 24027 32902 24092 32910
rect 23893 32856 23941 32902
tri 23713 32802 23767 32856 ne
rect 23767 32848 23807 32856
tri 23807 32848 23815 32856 sw
tri 23893 32848 23901 32856 ne
rect 23901 32848 23941 32856
rect 23767 32802 23815 32848
tri 23587 32748 23641 32802 ne
rect 23641 32770 23681 32802
tri 23681 32770 23713 32802 sw
tri 23767 32770 23799 32802 ne
rect 23799 32770 23815 32802
rect 23641 32748 23713 32770
rect 18274 32697 23375 32748
tri 5375 32666 5406 32697 se
rect 5406 32666 5503 32697
tri 5503 32666 5534 32697 nw
tri 5637 32666 5668 32697 se
rect 5668 32666 5749 32697
tri 5334 29432 5375 29473 se
rect 5375 29432 5441 32666
tri 5441 32604 5503 32666 nw
tri 5598 32627 5637 32666 se
rect 5637 32627 5749 32666
tri 5749 32627 5819 32697 nw
rect 18133 32694 23375 32697
tri 23375 32694 23429 32748 sw
tri 23461 32694 23515 32748 ne
rect 23515 32716 23555 32748
tri 23555 32716 23587 32748 sw
tri 23641 32716 23673 32748 ne
rect 23673 32716 23713 32748
rect 23515 32694 23587 32716
rect 18133 32692 23429 32694
tri 23337 32627 23402 32692 ne
rect 23402 32662 23429 32692
tri 23429 32662 23461 32694 sw
tri 23515 32662 23547 32694 ne
rect 23547 32662 23587 32694
rect 23402 32627 23461 32662
tri 5575 32604 5598 32627 se
rect 5598 32604 5652 32627
tri 5571 32600 5575 32604 se
rect 5575 32600 5652 32604
tri 5295 29393 5334 29432 se
rect 5334 29393 5441 29432
tri 5501 32530 5571 32600 se
rect 5571 32530 5652 32600
tri 5652 32530 5749 32627 nw
tri 23402 32600 23429 32627 ne
rect 23429 32600 23461 32627
tri 23461 32600 23523 32662 sw
tri 23547 32654 23555 32662 ne
rect 23555 32654 23587 32662
tri 23587 32654 23649 32716 sw
tri 23673 32708 23681 32716 ne
rect 23681 32708 23713 32716
tri 23713 32708 23775 32770 sw
tri 23799 32762 23807 32770 ne
rect 23807 32762 23815 32770
tri 23815 32762 23901 32848 sw
tri 23901 32816 23933 32848 ne
rect 23933 32816 23941 32848
tri 23941 32816 24027 32902 sw
tri 24027 32870 24059 32902 ne
rect 24059 32870 24092 32902
tri 24092 32870 24153 32931 sw
tri 24179 32924 24186 32931 ne
tri 24186 32924 24280 33018 sw
tri 24186 32870 24240 32924 ne
rect 24240 32870 24280 32924
tri 24059 32816 24113 32870 ne
rect 24113 32837 24153 32870
tri 24153 32837 24186 32870 sw
tri 24240 32837 24273 32870 ne
rect 24273 32837 24280 32870
rect 24113 32816 24186 32837
tri 23933 32762 23987 32816 ne
rect 23987 32808 24027 32816
tri 24027 32808 24035 32816 sw
tri 24113 32808 24121 32816 ne
rect 24121 32808 24186 32816
rect 23987 32762 24035 32808
tri 23807 32708 23861 32762 ne
rect 23861 32754 23901 32762
tri 23901 32754 23909 32762 sw
tri 23987 32754 23995 32762 ne
rect 23995 32754 24035 32762
rect 23861 32708 23909 32754
tri 23681 32654 23735 32708 ne
rect 23735 32676 23775 32708
tri 23775 32676 23807 32708 sw
tri 23861 32676 23893 32708 ne
rect 23893 32676 23909 32708
rect 23735 32654 23807 32676
tri 23555 32600 23609 32654 ne
rect 23609 32622 23649 32654
tri 23649 32622 23681 32654 sw
tri 23735 32622 23767 32654 ne
rect 23767 32622 23807 32654
rect 23609 32600 23681 32622
tri 23429 32530 23499 32600 ne
rect 23499 32568 23523 32600
tri 23523 32568 23555 32600 sw
tri 23609 32568 23641 32600 ne
rect 23641 32568 23681 32600
rect 23499 32530 23555 32568
rect 5501 29493 5567 32530
tri 5567 32445 5652 32530 nw
tri 23499 32506 23523 32530 ne
rect 23523 32506 23555 32530
tri 23555 32506 23617 32568 sw
tri 23641 32560 23649 32568 ne
rect 23649 32560 23681 32568
tri 23681 32560 23743 32622 sw
tri 23767 32614 23775 32622 ne
rect 23775 32614 23807 32622
tri 23807 32614 23869 32676 sw
tri 23893 32668 23901 32676 ne
rect 23901 32668 23909 32676
tri 23909 32668 23995 32754 sw
tri 23995 32722 24027 32754 ne
rect 24027 32722 24035 32754
tri 24035 32722 24121 32808 sw
tri 24121 32776 24153 32808 ne
rect 24153 32776 24186 32808
tri 24186 32776 24247 32837 sw
tri 24273 32830 24280 32837 ne
tri 24280 32830 24374 32924 sw
tri 24280 32776 24334 32830 ne
rect 24334 32776 24374 32830
tri 24153 32722 24207 32776 ne
rect 24207 32743 24247 32776
tri 24247 32743 24280 32776 sw
tri 24334 32743 24367 32776 ne
rect 24367 32743 24374 32776
rect 24207 32722 24280 32743
tri 24027 32668 24081 32722 ne
rect 24081 32714 24121 32722
tri 24121 32714 24129 32722 sw
tri 24207 32714 24215 32722 ne
rect 24215 32714 24280 32722
rect 24081 32668 24129 32714
tri 23901 32614 23955 32668 ne
rect 23955 32660 23995 32668
tri 23995 32660 24003 32668 sw
tri 24081 32660 24089 32668 ne
rect 24089 32660 24129 32668
rect 23955 32614 24003 32660
tri 23775 32560 23829 32614 ne
rect 23829 32582 23869 32614
tri 23869 32582 23901 32614 sw
tri 23955 32582 23987 32614 ne
rect 23987 32582 24003 32614
rect 23829 32560 23901 32582
tri 23649 32506 23703 32560 ne
rect 23703 32528 23743 32560
tri 23743 32528 23775 32560 sw
tri 23829 32528 23861 32560 ne
rect 23861 32528 23901 32560
rect 23703 32506 23775 32528
tri 23523 32445 23584 32506 ne
rect 23584 32474 23617 32506
tri 23617 32474 23649 32506 sw
tri 23703 32474 23735 32506 ne
rect 23735 32474 23775 32506
rect 23584 32445 23649 32474
tri 23584 32412 23617 32445 ne
rect 23617 32412 23649 32445
tri 23649 32412 23711 32474 sw
tri 23735 32466 23743 32474 ne
rect 23743 32466 23775 32474
tri 23775 32466 23837 32528 sw
tri 23861 32520 23869 32528 ne
rect 23869 32520 23901 32528
tri 23901 32520 23963 32582 sw
tri 23987 32574 23995 32582 ne
rect 23995 32574 24003 32582
tri 24003 32574 24089 32660 sw
tri 24089 32628 24121 32660 ne
rect 24121 32628 24129 32660
tri 24129 32628 24215 32714 sw
tri 24215 32682 24247 32714 ne
rect 24247 32682 24280 32714
tri 24280 32682 24341 32743 sw
tri 24367 32736 24374 32743 ne
tri 24374 32736 24468 32830 sw
tri 24374 32682 24428 32736 ne
rect 24428 32682 24468 32736
tri 24247 32628 24301 32682 ne
rect 24301 32649 24341 32682
tri 24341 32649 24374 32682 sw
tri 24428 32649 24461 32682 ne
rect 24461 32649 24468 32682
rect 24301 32628 24374 32649
tri 24121 32574 24175 32628 ne
rect 24175 32620 24215 32628
tri 24215 32620 24223 32628 sw
tri 24301 32620 24309 32628 ne
rect 24309 32620 24374 32628
rect 24175 32574 24223 32620
tri 23995 32520 24049 32574 ne
rect 24049 32566 24089 32574
tri 24089 32566 24097 32574 sw
tri 24175 32566 24183 32574 ne
rect 24183 32566 24223 32574
rect 24049 32520 24097 32566
tri 23869 32466 23923 32520 ne
rect 23923 32488 23963 32520
tri 23963 32488 23995 32520 sw
tri 24049 32488 24081 32520 ne
rect 24081 32488 24097 32520
rect 23923 32466 23995 32488
tri 23743 32412 23797 32466 ne
rect 23797 32434 23837 32466
tri 23837 32434 23869 32466 sw
tri 23923 32434 23955 32466 ne
rect 23955 32434 23995 32466
rect 23797 32412 23869 32434
tri 23617 32318 23711 32412 ne
tri 23711 32380 23743 32412 sw
tri 23797 32380 23829 32412 ne
rect 23829 32380 23869 32412
rect 23711 32318 23743 32380
tri 23743 32318 23805 32380 sw
tri 23829 32372 23837 32380 ne
rect 23837 32372 23869 32380
tri 23869 32372 23931 32434 sw
tri 23955 32426 23963 32434 ne
rect 23963 32426 23995 32434
tri 23995 32426 24057 32488 sw
tri 24081 32480 24089 32488 ne
rect 24089 32480 24097 32488
tri 24097 32480 24183 32566 sw
tri 24183 32534 24215 32566 ne
rect 24215 32534 24223 32566
tri 24223 32534 24309 32620 sw
tri 24309 32588 24341 32620 ne
rect 24341 32588 24374 32620
tri 24374 32588 24435 32649 sw
tri 24461 32642 24468 32649 ne
tri 24468 32642 24562 32736 sw
tri 24468 32588 24522 32642 ne
rect 24522 32588 24562 32642
tri 24341 32534 24395 32588 ne
rect 24395 32555 24435 32588
tri 24435 32555 24468 32588 sw
tri 24522 32555 24555 32588 ne
rect 24555 32555 24562 32588
rect 24395 32534 24468 32555
tri 24215 32480 24269 32534 ne
rect 24269 32526 24309 32534
tri 24309 32526 24317 32534 sw
tri 24395 32526 24403 32534 ne
rect 24403 32526 24468 32534
rect 24269 32480 24317 32526
tri 24089 32426 24143 32480 ne
rect 24143 32472 24183 32480
tri 24183 32472 24191 32480 sw
tri 24269 32472 24277 32480 ne
rect 24277 32472 24317 32480
rect 24143 32426 24191 32472
tri 23963 32372 24017 32426 ne
rect 24017 32394 24057 32426
tri 24057 32394 24089 32426 sw
tri 24143 32394 24175 32426 ne
rect 24175 32394 24191 32426
rect 24017 32372 24089 32394
tri 23837 32318 23891 32372 ne
rect 23891 32340 23931 32372
tri 23931 32340 23963 32372 sw
tri 24017 32340 24049 32372 ne
rect 24049 32340 24089 32372
rect 23891 32318 23963 32340
tri 23711 32224 23805 32318 ne
tri 23805 32286 23837 32318 sw
tri 23891 32286 23923 32318 ne
rect 23923 32286 23963 32318
rect 23805 32224 23837 32286
tri 23837 32224 23899 32286 sw
tri 23923 32278 23931 32286 ne
rect 23931 32278 23963 32286
tri 23963 32278 24025 32340 sw
tri 24049 32332 24057 32340 ne
rect 24057 32332 24089 32340
tri 24089 32332 24151 32394 sw
tri 24175 32386 24183 32394 ne
rect 24183 32386 24191 32394
tri 24191 32386 24277 32472 sw
tri 24277 32440 24309 32472 ne
rect 24309 32440 24317 32472
tri 24317 32440 24403 32526 sw
tri 24403 32494 24435 32526 ne
rect 24435 32494 24468 32526
tri 24468 32494 24529 32555 sw
tri 24555 32548 24562 32555 ne
tri 24562 32548 24656 32642 sw
tri 24562 32494 24616 32548 ne
rect 24616 32494 24656 32548
tri 24435 32440 24489 32494 ne
rect 24489 32461 24529 32494
tri 24529 32461 24562 32494 sw
tri 24616 32461 24649 32494 ne
rect 24649 32461 24656 32494
rect 24489 32440 24562 32461
tri 24309 32386 24363 32440 ne
rect 24363 32432 24403 32440
tri 24403 32432 24411 32440 sw
tri 24489 32432 24497 32440 ne
rect 24497 32432 24562 32440
rect 24363 32386 24411 32432
tri 24183 32332 24237 32386 ne
rect 24237 32378 24277 32386
tri 24277 32378 24285 32386 sw
tri 24363 32378 24371 32386 ne
rect 24371 32378 24411 32386
rect 24237 32332 24285 32378
tri 24057 32278 24111 32332 ne
rect 24111 32300 24151 32332
tri 24151 32300 24183 32332 sw
tri 24237 32300 24269 32332 ne
rect 24269 32300 24285 32332
rect 24111 32278 24183 32300
tri 23931 32224 23985 32278 ne
rect 23985 32246 24025 32278
tri 24025 32246 24057 32278 sw
tri 24111 32246 24143 32278 ne
rect 24143 32246 24183 32278
rect 23985 32224 24057 32246
tri 23805 32130 23899 32224 ne
tri 23899 32192 23931 32224 sw
tri 23985 32192 24017 32224 ne
rect 24017 32192 24057 32224
rect 23899 32130 23931 32192
tri 23931 32130 23993 32192 sw
tri 24017 32184 24025 32192 ne
rect 24025 32184 24057 32192
tri 24057 32184 24119 32246 sw
tri 24143 32238 24151 32246 ne
rect 24151 32238 24183 32246
tri 24183 32238 24245 32300 sw
tri 24269 32292 24277 32300 ne
rect 24277 32292 24285 32300
tri 24285 32292 24371 32378 sw
tri 24371 32346 24403 32378 ne
rect 24403 32346 24411 32378
tri 24411 32346 24497 32432 sw
tri 24497 32400 24529 32432 ne
rect 24529 32400 24562 32432
tri 24562 32400 24623 32461 sw
tri 24649 32454 24656 32461 ne
tri 24656 32454 24750 32548 sw
tri 24656 32400 24710 32454 ne
rect 24710 32400 24750 32454
tri 24529 32346 24583 32400 ne
rect 24583 32367 24623 32400
tri 24623 32367 24656 32400 sw
tri 24710 32367 24743 32400 ne
rect 24743 32367 24750 32400
rect 24583 32346 24656 32367
tri 24403 32292 24457 32346 ne
rect 24457 32338 24497 32346
tri 24497 32338 24505 32346 sw
tri 24583 32338 24591 32346 ne
rect 24591 32338 24656 32346
rect 24457 32292 24505 32338
tri 24277 32238 24331 32292 ne
rect 24331 32284 24371 32292
tri 24371 32284 24379 32292 sw
tri 24457 32284 24465 32292 ne
rect 24465 32284 24505 32292
rect 24331 32238 24379 32284
tri 24151 32184 24205 32238 ne
rect 24205 32206 24245 32238
tri 24245 32206 24277 32238 sw
tri 24331 32206 24363 32238 ne
rect 24363 32206 24379 32238
rect 24205 32184 24277 32206
tri 24025 32130 24079 32184 ne
rect 24079 32152 24119 32184
tri 24119 32152 24151 32184 sw
tri 24205 32152 24237 32184 ne
rect 24237 32152 24277 32184
rect 24079 32130 24151 32152
tri 23899 32036 23993 32130 ne
tri 23993 32098 24025 32130 sw
tri 24079 32098 24111 32130 ne
rect 24111 32098 24151 32130
rect 23993 32036 24025 32098
tri 24025 32036 24087 32098 sw
tri 24111 32090 24119 32098 ne
rect 24119 32090 24151 32098
tri 24151 32090 24213 32152 sw
tri 24237 32144 24245 32152 ne
rect 24245 32144 24277 32152
tri 24277 32144 24339 32206 sw
tri 24363 32198 24371 32206 ne
rect 24371 32198 24379 32206
tri 24379 32198 24465 32284 sw
tri 24465 32252 24497 32284 ne
rect 24497 32252 24505 32284
tri 24505 32252 24591 32338 sw
tri 24591 32306 24623 32338 ne
rect 24623 32306 24656 32338
tri 24656 32306 24717 32367 sw
tri 24743 32360 24750 32367 ne
tri 24750 32360 24844 32454 sw
tri 24750 32306 24804 32360 ne
rect 24804 32306 24844 32360
tri 24623 32252 24677 32306 ne
rect 24677 32273 24717 32306
tri 24717 32273 24750 32306 sw
tri 24804 32273 24837 32306 ne
rect 24837 32273 24844 32306
rect 24677 32252 24750 32273
tri 24497 32198 24551 32252 ne
rect 24551 32244 24591 32252
tri 24591 32244 24599 32252 sw
tri 24677 32244 24685 32252 ne
rect 24685 32244 24750 32252
rect 24551 32198 24599 32244
tri 24371 32144 24425 32198 ne
rect 24425 32190 24465 32198
tri 24465 32190 24473 32198 sw
tri 24551 32190 24559 32198 ne
rect 24559 32190 24599 32198
rect 24425 32144 24473 32190
tri 24245 32090 24299 32144 ne
rect 24299 32112 24339 32144
tri 24339 32112 24371 32144 sw
tri 24425 32112 24457 32144 ne
rect 24457 32112 24473 32144
rect 24299 32090 24371 32112
tri 24119 32036 24173 32090 ne
rect 24173 32058 24213 32090
tri 24213 32058 24245 32090 sw
tri 24299 32058 24331 32090 ne
rect 24331 32058 24371 32090
rect 24173 32036 24245 32058
tri 23993 31942 24087 32036 ne
tri 24087 32004 24119 32036 sw
tri 24173 32004 24205 32036 ne
rect 24205 32004 24245 32036
rect 24087 31942 24119 32004
tri 24119 31942 24181 32004 sw
tri 24205 31996 24213 32004 ne
rect 24213 31996 24245 32004
tri 24245 31996 24307 32058 sw
tri 24331 32050 24339 32058 ne
rect 24339 32050 24371 32058
tri 24371 32050 24433 32112 sw
tri 24457 32104 24465 32112 ne
rect 24465 32104 24473 32112
tri 24473 32104 24559 32190 sw
tri 24559 32158 24591 32190 ne
rect 24591 32158 24599 32190
tri 24599 32158 24685 32244 sw
tri 24685 32212 24717 32244 ne
rect 24717 32212 24750 32244
tri 24750 32212 24811 32273 sw
tri 24837 32266 24844 32273 ne
tri 24844 32266 24938 32360 sw
tri 24844 32212 24898 32266 ne
rect 24898 32212 24938 32266
tri 24717 32158 24771 32212 ne
rect 24771 32179 24811 32212
tri 24811 32179 24844 32212 sw
tri 24898 32179 24931 32212 ne
rect 24931 32179 24938 32212
rect 24771 32158 24844 32179
tri 24591 32104 24645 32158 ne
rect 24645 32150 24685 32158
tri 24685 32150 24693 32158 sw
tri 24771 32150 24779 32158 ne
rect 24779 32150 24844 32158
rect 24645 32104 24693 32150
tri 24465 32050 24519 32104 ne
rect 24519 32096 24559 32104
tri 24559 32096 24567 32104 sw
tri 24645 32096 24653 32104 ne
rect 24653 32096 24693 32104
rect 24519 32050 24567 32096
tri 24339 31996 24393 32050 ne
rect 24393 32018 24433 32050
tri 24433 32018 24465 32050 sw
tri 24519 32018 24551 32050 ne
rect 24551 32018 24567 32050
rect 24393 31996 24465 32018
tri 24213 31942 24267 31996 ne
rect 24267 31964 24307 31996
tri 24307 31964 24339 31996 sw
tri 24393 31964 24425 31996 ne
rect 24425 31964 24465 31996
rect 24267 31942 24339 31964
tri 24087 31848 24181 31942 ne
tri 24181 31910 24213 31942 sw
tri 24267 31910 24299 31942 ne
rect 24299 31910 24339 31942
rect 24181 31848 24213 31910
tri 24213 31848 24275 31910 sw
tri 24299 31902 24307 31910 ne
rect 24307 31902 24339 31910
tri 24339 31902 24401 31964 sw
tri 24425 31956 24433 31964 ne
rect 24433 31956 24465 31964
tri 24465 31956 24527 32018 sw
tri 24551 32010 24559 32018 ne
rect 24559 32010 24567 32018
tri 24567 32010 24653 32096 sw
tri 24653 32064 24685 32096 ne
rect 24685 32064 24693 32096
tri 24693 32064 24779 32150 sw
tri 24779 32118 24811 32150 ne
rect 24811 32118 24844 32150
tri 24844 32118 24905 32179 sw
tri 24931 32172 24938 32179 ne
tri 24938 32172 25032 32266 sw
tri 24938 32118 24992 32172 ne
rect 24992 32118 25032 32172
tri 24811 32064 24865 32118 ne
rect 24865 32085 24905 32118
tri 24905 32085 24938 32118 sw
tri 24992 32085 25025 32118 ne
rect 25025 32085 25032 32118
rect 24865 32064 24938 32085
tri 24685 32010 24739 32064 ne
rect 24739 32056 24779 32064
tri 24779 32056 24787 32064 sw
tri 24865 32056 24873 32064 ne
rect 24873 32056 24938 32064
rect 24739 32010 24787 32056
tri 24559 31956 24613 32010 ne
rect 24613 32002 24653 32010
tri 24653 32002 24661 32010 sw
tri 24739 32002 24747 32010 ne
rect 24747 32002 24787 32010
rect 24613 31956 24661 32002
tri 24433 31902 24487 31956 ne
rect 24487 31924 24527 31956
tri 24527 31924 24559 31956 sw
tri 24613 31924 24645 31956 ne
rect 24645 31924 24661 31956
rect 24487 31902 24559 31924
tri 24307 31848 24361 31902 ne
rect 24361 31870 24401 31902
tri 24401 31870 24433 31902 sw
tri 24487 31870 24519 31902 ne
rect 24519 31870 24559 31902
rect 24361 31848 24433 31870
tri 24181 31754 24275 31848 ne
tri 24275 31816 24307 31848 sw
tri 24361 31816 24393 31848 ne
rect 24393 31816 24433 31848
rect 24275 31754 24307 31816
tri 24307 31754 24369 31816 sw
tri 24393 31808 24401 31816 ne
rect 24401 31808 24433 31816
tri 24433 31808 24495 31870 sw
tri 24519 31862 24527 31870 ne
rect 24527 31862 24559 31870
tri 24559 31862 24621 31924 sw
tri 24645 31916 24653 31924 ne
rect 24653 31916 24661 31924
tri 24661 31916 24747 32002 sw
tri 24747 31970 24779 32002 ne
rect 24779 31970 24787 32002
tri 24787 31970 24873 32056 sw
tri 24873 32024 24905 32056 ne
rect 24905 32024 24938 32056
tri 24938 32024 24999 32085 sw
tri 25025 32078 25032 32085 ne
tri 25032 32078 25126 32172 sw
tri 25032 32024 25086 32078 ne
rect 25086 32024 25126 32078
tri 24905 31970 24959 32024 ne
rect 24959 31991 24999 32024
tri 24999 31991 25032 32024 sw
tri 25086 31991 25119 32024 ne
rect 25119 31991 25126 32024
rect 24959 31970 25032 31991
tri 24779 31916 24833 31970 ne
rect 24833 31962 24873 31970
tri 24873 31962 24881 31970 sw
tri 24959 31962 24967 31970 ne
rect 24967 31962 25032 31970
rect 24833 31916 24881 31962
tri 24653 31862 24707 31916 ne
rect 24707 31908 24747 31916
tri 24747 31908 24755 31916 sw
tri 24833 31908 24841 31916 ne
rect 24841 31908 24881 31916
rect 24707 31862 24755 31908
tri 24527 31808 24581 31862 ne
rect 24581 31830 24621 31862
tri 24621 31830 24653 31862 sw
tri 24707 31830 24739 31862 ne
rect 24739 31830 24755 31862
rect 24581 31808 24653 31830
tri 24401 31754 24455 31808 ne
rect 24455 31776 24495 31808
tri 24495 31776 24527 31808 sw
tri 24581 31776 24613 31808 ne
rect 24613 31776 24653 31808
rect 24455 31754 24527 31776
tri 24275 31660 24369 31754 ne
tri 24369 31722 24401 31754 sw
tri 24455 31722 24487 31754 ne
rect 24487 31722 24527 31754
rect 24369 31660 24401 31722
tri 24401 31660 24463 31722 sw
tri 24487 31714 24495 31722 ne
rect 24495 31714 24527 31722
tri 24527 31714 24589 31776 sw
tri 24613 31768 24621 31776 ne
rect 24621 31768 24653 31776
tri 24653 31768 24715 31830 sw
tri 24739 31822 24747 31830 ne
rect 24747 31822 24755 31830
tri 24755 31822 24841 31908 sw
tri 24841 31876 24873 31908 ne
rect 24873 31876 24881 31908
tri 24881 31876 24967 31962 sw
tri 24967 31902 25027 31962 ne
rect 25027 31930 25032 31962
tri 25032 31930 25093 31991 sw
tri 25119 31984 25126 31991 ne
tri 25126 31984 25220 32078 sw
tri 25126 31956 25154 31984 ne
tri 24873 31848 24901 31876 ne
tri 24747 31794 24775 31822 ne
tri 24621 31740 24649 31768 ne
tri 24495 31686 24523 31714 ne
tri 24369 31632 24397 31660 ne
rect 24397 29920 24463 31660
rect 24397 29864 24402 29920
rect 24458 29864 24463 29920
rect 24397 29840 24463 29864
rect 24397 29784 24402 29840
rect 24458 29784 24463 29840
rect 24397 29767 24463 29784
tri 5567 29493 5647 29573 sw
rect 5501 29488 5647 29493
rect 5501 29432 5506 29488
rect 5562 29432 5586 29488
rect 5642 29432 5647 29488
rect 5501 29427 5647 29432
rect 5295 29388 5441 29393
rect 5295 29332 5300 29388
rect 5356 29332 5380 29388
rect 5436 29332 5441 29388
rect 5295 29327 5441 29332
rect 21299 27345 21892 27790
rect 24523 21096 24589 31714
rect 24649 18589 24715 31768
rect 24775 20822 24841 31822
rect 24775 20766 24780 20822
rect 24836 20766 24841 20822
rect 24775 20742 24841 20766
rect 24775 20686 24780 20742
rect 24836 20686 24841 20742
rect 24775 20677 24841 20686
rect 24901 20105 24967 31876
rect 25027 21231 25093 31930
rect 25027 21175 25032 21231
rect 25088 21175 25093 21231
rect 25027 21151 25093 21175
rect 25027 21095 25032 21151
rect 25088 21095 25093 21151
rect 25027 21090 25093 21095
rect 25154 21137 25220 31984
rect 25154 21081 25159 21137
rect 25215 21081 25220 21137
rect 25154 21057 25220 21081
rect 25154 21001 25159 21057
rect 25215 21001 25220 21057
rect 25154 20996 25220 21001
rect 24901 20049 24906 20105
rect 24962 20049 24967 20105
rect 24901 20025 24967 20049
rect 24901 19969 24906 20025
rect 24962 19969 24967 20025
rect 24901 19960 24967 19969
rect 24649 18533 24654 18589
rect 24710 18533 24715 18589
rect 24649 18509 24715 18533
rect 2646 18462 2686 18491
rect 24649 18453 24654 18509
rect 24710 18453 24715 18509
rect 24649 18444 24715 18453
use sky130_fd_io__gpio_ovtv2_obpredrvr_new_i2c_fix_leak_fix  sky130_fd_io__gpio_ovtv2_obpredrvr_new_i2c_fix_leak_fix_0
timestamp 1704896540
transform 1 0 -49 0 1 28727
box 255 -19630 28132 5180
use sky130_fd_io__gpio_ovtv2_obpredrvr_old  sky130_fd_io__gpio_ovtv2_obpredrvr_old_0
timestamp 1704896540
transform 0 1 23158 -1 0 30683
box -255 631 13433 4925
<< labels >>
flabel metal3 s 2646 18462 2686 18491 0 FreeSans 200 0 0 0 NGHS_H
port 2 nsew
flabel metal3 s 21299 27345 21892 27790 3 FreeSans 520 270 0 0 VGND_IO
port 3 nsew
flabel metal3 s 21595 27567 21595 27567 3 FreeSans 520 270 0 0 VGND_IO
flabel metal1 s 11513 32365 11551 32404 3 FreeSans 520 90 0 0 OE_I_H_N
port 5 nsew
flabel metal1 s 26335 17905 26537 17947 7 FreeSans 300 270 0 0 VGND_IO
port 3 nsew
flabel metal1 s 25923 17881 26053 17923 7 FreeSans 300 270 0 0 VGND_IO
port 3 nsew
flabel metal1 s 25307 17775 25437 17817 7 FreeSans 300 270 0 0 VGND_IO
port 3 nsew
flabel metal1 s 24184 17775 24386 17817 7 FreeSans 300 270 0 0 VGND_IO
port 3 nsew
flabel metal1 s 24184 29706 24386 29748 3 FreeSans 300 270 0 0 VGND_IO
port 3 nsew
flabel metal1 s 25923 30641 26053 30683 3 FreeSans 300 270 0 0 VGND_IO
port 3 nsew
flabel metal1 s 26335 30641 26537 30683 3 FreeSans 300 270 0 0 VGND_IO
port 3 nsew
flabel metal1 s 26861 17775 27063 17817 7 FreeSans 300 270 0 0 VCC_IO
port 6 nsew
flabel metal1 s 27575 17775 27721 17812 7 FreeSans 300 270 0 0 VCC_IO
port 6 nsew
flabel metal1 s 24710 17775 24912 17817 7 FreeSans 300 270 0 0 VCC_IO
port 6 nsew
flabel metal1 s 24432 30637 24634 30679 3 FreeSans 300 270 0 0 VCC_IO
port 6 nsew
flabel metal1 s 27575 30646 27721 30683 3 FreeSans 300 270 0 0 VCC_IO
port 6 nsew
flabel metal1 s 26861 30641 27063 30683 3 FreeSans 300 270 0 0 VCC_IO
port 6 nsew
flabel metal1 s 25465 20856 25511 20902 3 FreeSans 300 270 0 0 SLOW_H
port 7 nsew
flabel metal1 s 27321 30418 27352 30562 3 FreeSans 520 270 0 0 PUEN_H[1]
port 8 nsew
flabel metal1 s 26721 23039 26752 23133 3 FreeSans 520 270 0 0 PUEN_H[0]
port 9 nsew
flabel metal1 s 27091 24740 27137 24781 3 FreeSans 300 270 0 0 PU_H_N[3]
port 10 nsew
flabel metal1 s 27091 24877 27137 24917 7 FreeSans 300 270 0 0 PU_H_N[2]
port 11 nsew
flabel metal1 s 27247 20545 27293 20585 3 FreeSans 300 270 0 0 PU_H_N[1]
port 12 nsew
flabel metal1 s 27171 22975 27217 23015 3 FreeSans 300 270 0 0 PU_H_N[0]
port 13 nsew
flabel metal1 s 27289 21535 27335 21581 3 FreeSans 300 270 0 0 PD_H[1]
port 14 nsew
flabel metal1 s 18581 32317 19176 32472 3 FreeSans 520 90 0 0 VGND_IO
port 3 nsew
flabel metal1 s 18522 33471 19108 33673 3 FreeSans 520 90 0 0 VCC_IO
port 6 nsew
flabel metal1 s 27289 22777 27335 22823 3 FreeSans 300 270 0 0 PD_H[0]
port 15 nsew
flabel metal1 s 26650 22321 26674 22407 3 FreeSans 520 270 0 0 PDEN_H_N[0]
port 16 nsew
flabel metal2 s 4839 28595 4994 28884 3 FreeSans 520 180 0 0 VGND_IO
port 3 nsew
flabel metal2 s 4916 28739 4916 28739 3 FreeSans 520 180 0 0 VGND_IO
flabel metal2 s 11274 33500 11643 33685 3 FreeSans 520 90 0 0 VCC_IO
port 6 nsew
flabel metal2 s 2028 29282 2200 29364 3 FreeSans 520 0 0 0 PD_H[3]
port 18 nsew
flabel metal2 s 2114 29323 2114 29323 3 FreeSans 520 0 0 0 PD_H[3]
flabel metal2 s 2214 29431 2333 29489 3 FreeSans 520 0 0 0 PD_H[2]
port 19 nsew
flabel metal2 s 18919 27043 19027 27411 3 FreeSans 520 180 0 0 PAD
port 20 nsew
flabel metal2 s 22701 27039 22809 27407 3 FreeSans 520 0 0 0 PAD
port 20 nsew
flabel metal2 s 22755 27223 22755 27223 3 FreeSans 520 0 0 0 PAD
flabel metal2 s 25722 23272 25873 23315 3 FreeSans 520 270 0 0 PDEN_H_N[1]
port 21 nsew
flabel metal2 s 26781 20301 26833 20359 3 FreeSans 300 270 0 0 PD_H[3]
port 18 nsew
flabel metal2 s 25098 20781 25150 20828 3 FreeSans 300 270 0 0 PD_H[2]
port 19 nsew
flabel metal2 s 26621 17940 26673 17987 7 FreeSans 300 270 0 0 DRVLO_H_N
port 22 nsew
flabel metal2 s 26693 23756 26745 23808 3 FreeSans 300 270 0 0 DRVHI_H
port 23 nsew
flabel locali s 18234 32803 18269 32838 3 FreeSans 520 90 0 0 SLOW_H_N
port 24 nsew
flabel locali s 19211 32744 19267 32788 3 FreeSans 520 90 0 0 SLEW_CTL_H_N[0]
port 25 nsew
flabel locali s 18420 32797 18456 32833 3 FreeSans 520 90 0 0 SLEW_CTL_H[1]
port 26 nsew
flabel locali s 16965 32758 16996 32798 3 FreeSans 520 90 0 0 PDEN_H_N[1]
port 21 nsew
flabel locali s 11923 32808 11954 32846 3 FreeSans 520 90 0 0 PD_DIS_H
port 27 nsew
flabel locali s 18056 32815 18086 32844 3 FreeSans 520 90 0 0 I2C_MODE_H_N
port 28 nsew
flabel locali s 16799 32751 16831 32795 3 FreeSans 520 90 0 0 DRVLO_H_N
port 22 nsew
<< properties >>
string GDS_END 69053838
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 69037980
<< end >>
