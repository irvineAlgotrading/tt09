magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -119 -66 687 366
<< mvpmos >>
rect 0 0 100 300
rect 156 0 256 300
rect 312 0 412 300
rect 468 0 568 300
<< mvpdiff >>
rect -53 250 0 300
rect -53 216 -45 250
rect -11 216 0 250
rect -53 182 0 216
rect -53 148 -45 182
rect -11 148 0 182
rect -53 114 0 148
rect -53 80 -45 114
rect -11 80 0 114
rect -53 46 0 80
rect -53 12 -45 46
rect -11 12 0 46
rect -53 0 0 12
rect 100 250 156 300
rect 100 216 111 250
rect 145 216 156 250
rect 100 182 156 216
rect 100 148 111 182
rect 145 148 156 182
rect 100 114 156 148
rect 100 80 111 114
rect 145 80 156 114
rect 100 46 156 80
rect 100 12 111 46
rect 145 12 156 46
rect 100 0 156 12
rect 256 250 312 300
rect 256 216 267 250
rect 301 216 312 250
rect 256 182 312 216
rect 256 148 267 182
rect 301 148 312 182
rect 256 114 312 148
rect 256 80 267 114
rect 301 80 312 114
rect 256 46 312 80
rect 256 12 267 46
rect 301 12 312 46
rect 256 0 312 12
rect 412 250 468 300
rect 412 216 423 250
rect 457 216 468 250
rect 412 182 468 216
rect 412 148 423 182
rect 457 148 468 182
rect 412 114 468 148
rect 412 80 423 114
rect 457 80 468 114
rect 412 46 468 80
rect 412 12 423 46
rect 457 12 468 46
rect 412 0 468 12
rect 568 250 621 300
rect 568 216 579 250
rect 613 216 621 250
rect 568 182 621 216
rect 568 148 579 182
rect 613 148 621 182
rect 568 114 621 148
rect 568 80 579 114
rect 613 80 621 114
rect 568 46 621 80
rect 568 12 579 46
rect 613 12 621 46
rect 568 0 621 12
<< mvpdiffc >>
rect -45 216 -11 250
rect -45 148 -11 182
rect -45 80 -11 114
rect -45 12 -11 46
rect 111 216 145 250
rect 111 148 145 182
rect 111 80 145 114
rect 111 12 145 46
rect 267 216 301 250
rect 267 148 301 182
rect 267 80 301 114
rect 267 12 301 46
rect 423 216 457 250
rect 423 148 457 182
rect 423 80 457 114
rect 423 12 457 46
rect 579 216 613 250
rect 579 148 613 182
rect 579 80 613 114
rect 579 12 613 46
<< poly >>
rect 0 300 100 332
rect 156 300 256 332
rect 312 300 412 332
rect 468 300 568 332
rect 0 -32 100 0
rect 156 -32 256 0
rect 312 -32 412 0
rect 468 -32 568 0
<< locali >>
rect -45 250 -11 266
rect -45 182 -11 216
rect -45 114 -11 148
rect -45 46 -11 80
rect -45 -4 -11 12
rect 111 250 145 266
rect 111 182 145 216
rect 111 114 145 148
rect 111 46 145 80
rect 111 -4 145 12
rect 267 250 301 266
rect 267 182 301 216
rect 267 114 301 148
rect 267 46 301 80
rect 267 -4 301 12
rect 423 250 457 266
rect 423 182 457 216
rect 423 114 457 148
rect 423 46 457 80
rect 423 -4 457 12
rect 579 250 613 266
rect 579 182 613 216
rect 579 114 613 148
rect 579 46 613 80
rect 579 -4 613 12
use DFL1sd2_CDNS_52468879185253  DFL1sd2_CDNS_52468879185253_0
timestamp 1704896540
transform 1 0 412 0 1 0
box 0 0 1 1
use DFL1sd2_CDNS_52468879185253  DFL1sd2_CDNS_52468879185253_1
timestamp 1704896540
transform 1 0 256 0 1 0
box 0 0 1 1
use DFL1sd2_CDNS_52468879185253  DFL1sd2_CDNS_52468879185253_2
timestamp 1704896540
transform 1 0 100 0 1 0
box 0 0 1 1
use DFL1sd_CDNS_52468879185252  DFL1sd_CDNS_52468879185252_0
timestamp 1704896540
transform -1 0 0 0 1 0
box 0 0 1 1
use DFL1sd_CDNS_52468879185252  DFL1sd_CDNS_52468879185252_1
timestamp 1704896540
transform 1 0 568 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s -28 131 -28 131 0 FreeSans 300 0 0 0 S
flabel comment s 128 131 128 131 0 FreeSans 300 0 0 0 D
flabel comment s 284 131 284 131 0 FreeSans 300 0 0 0 S
flabel comment s 440 131 440 131 0 FreeSans 300 0 0 0 D
flabel comment s 596 131 596 131 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 6083018
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 6080510
<< end >>
