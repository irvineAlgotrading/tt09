magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< pwell >>
rect -105 -26 607 4026
rect 815 -26 1527 4026
rect 1735 -26 2447 4026
rect 2655 -26 3367 4026
rect 3575 -26 4287 4026
rect 4495 -26 5207 4026
rect 5415 -26 6127 4026
rect 6335 -26 7047 4026
rect 7255 -26 7967 4026
rect 8175 -26 8887 4026
rect 9095 -26 9807 4026
<< mvnmos >>
rect 0 0 100 4000
rect 402 0 502 4000
rect 920 0 1020 4000
rect 1322 0 1422 4000
rect 1840 0 1940 4000
rect 2242 0 2342 4000
rect 2760 0 2860 4000
rect 3162 0 3262 4000
rect 3680 0 3780 4000
rect 4082 0 4182 4000
rect 4600 0 4700 4000
rect 5002 0 5102 4000
rect 5520 0 5620 4000
rect 5922 0 6022 4000
rect 6440 0 6540 4000
rect 6842 0 6942 4000
rect 7360 0 7460 4000
rect 7762 0 7862 4000
rect 8280 0 8380 4000
rect 8682 0 8782 4000
rect 9200 0 9300 4000
rect 9602 0 9702 4000
<< mvndiff >>
rect -79 0 0 4000
rect 100 0 402 4000
rect 502 0 581 4000
rect 841 0 920 4000
rect 1020 0 1322 4000
rect 1422 0 1501 4000
rect 1761 0 1840 4000
rect 1940 0 2242 4000
rect 2342 0 2421 4000
rect 2681 0 2760 4000
rect 2860 0 3162 4000
rect 3262 0 3341 4000
rect 3601 0 3680 4000
rect 3780 0 4082 4000
rect 4182 0 4261 4000
rect 4521 0 4600 4000
rect 4700 0 5002 4000
rect 5102 0 5181 4000
rect 5441 0 5520 4000
rect 5620 0 5922 4000
rect 6022 0 6101 4000
rect 6361 0 6440 4000
rect 6540 0 6842 4000
rect 6942 0 7021 4000
rect 7281 0 7360 4000
rect 7460 0 7762 4000
rect 7862 0 7941 4000
rect 8201 0 8280 4000
rect 8380 0 8682 4000
rect 8782 0 8861 4000
rect 9121 0 9200 4000
rect 9300 0 9602 4000
rect 9702 0 9781 4000
<< poly >>
rect 0 4000 100 4032
rect 402 4000 502 4032
rect 920 4000 1020 4032
rect 1322 4000 1422 4032
rect 1840 4000 1940 4032
rect 2242 4000 2342 4032
rect 2760 4000 2860 4032
rect 3162 4000 3262 4032
rect 3680 4000 3780 4032
rect 4082 4000 4182 4032
rect 4600 4000 4700 4032
rect 5002 4000 5102 4032
rect 5520 4000 5620 4032
rect 5922 4000 6022 4032
rect 6440 4000 6540 4032
rect 6842 4000 6942 4032
rect 7360 4000 7460 4032
rect 7762 4000 7862 4032
rect 8280 4000 8380 4032
rect 8682 4000 8782 4032
rect 9200 4000 9300 4032
rect 9602 4000 9702 4032
rect 0 -32 100 0
rect 402 -32 502 0
rect 920 -32 1020 0
rect 1322 -32 1422 0
rect 1840 -32 1940 0
rect 2242 -32 2342 0
rect 2760 -32 2860 0
rect 3162 -32 3262 0
rect 3680 -32 3780 0
rect 4082 -32 4182 0
rect 4600 -32 4700 0
rect 5002 -32 5102 0
rect 5520 -32 5620 0
rect 5922 -32 6022 0
rect 6440 -32 6540 0
rect 6842 -32 6942 0
rect 7360 -32 7460 0
rect 7762 -32 7862 0
rect 8280 -32 8380 0
rect 8682 -32 8782 0
rect 9200 -32 9300 0
rect 9602 -32 9702 0
<< locali >>
rect -192 -4 -90 3950
rect 592 -4 830 3938
rect 1512 -4 1750 3938
rect 2432 -4 2670 3938
rect 3352 -4 3590 3938
rect 4272 -4 4510 3938
rect 5192 -4 5430 3938
rect 6112 -4 6350 3938
rect 7032 -4 7270 3938
rect 7952 -4 8190 3938
rect 8872 -4 9110 3938
rect 9792 -4 9894 3950
use hvDFTPL1s2_CDNS_52468879185832  hvDFTPL1s2_CDNS_52468879185832_0
timestamp 1704896540
transform 1 0 8861 0 1 0
box -26 -26 286 4026
use hvDFTPL1s2_CDNS_52468879185832  hvDFTPL1s2_CDNS_52468879185832_1
timestamp 1704896540
transform 1 0 7941 0 1 0
box -26 -26 286 4026
use hvDFTPL1s2_CDNS_52468879185832  hvDFTPL1s2_CDNS_52468879185832_2
timestamp 1704896540
transform 1 0 7021 0 1 0
box -26 -26 286 4026
use hvDFTPL1s2_CDNS_52468879185832  hvDFTPL1s2_CDNS_52468879185832_3
timestamp 1704896540
transform 1 0 6101 0 1 0
box -26 -26 286 4026
use hvDFTPL1s2_CDNS_52468879185832  hvDFTPL1s2_CDNS_52468879185832_4
timestamp 1704896540
transform 1 0 5181 0 1 0
box -26 -26 286 4026
use hvDFTPL1s2_CDNS_52468879185832  hvDFTPL1s2_CDNS_52468879185832_5
timestamp 1704896540
transform 1 0 4261 0 1 0
box -26 -26 286 4026
use hvDFTPL1s2_CDNS_52468879185832  hvDFTPL1s2_CDNS_52468879185832_6
timestamp 1704896540
transform 1 0 3341 0 1 0
box -26 -26 286 4026
use hvDFTPL1s2_CDNS_52468879185832  hvDFTPL1s2_CDNS_52468879185832_7
timestamp 1704896540
transform 1 0 2421 0 1 0
box -26 -26 286 4026
use hvDFTPL1s2_CDNS_52468879185832  hvDFTPL1s2_CDNS_52468879185832_8
timestamp 1704896540
transform 1 0 1501 0 1 0
box -26 -26 286 4026
use hvDFTPL1s2_CDNS_52468879185832  hvDFTPL1s2_CDNS_52468879185832_9
timestamp 1704896540
transform 1 0 581 0 1 0
box -26 -26 286 4026
use hvDFTPL1s_CDNS_52468879185831  hvDFTPL1s_CDNS_52468879185831_0
timestamp 1704896540
transform -1 0 -79 0 1 0
box -26 -26 226 4026
use hvDFTPL1s_CDNS_52468879185831  hvDFTPL1s_CDNS_52468879185831_1
timestamp 1704896540
transform 1 0 9781 0 1 0
box -26 -26 226 4026
<< labels >>
flabel comment s -141 1973 -141 1973 0 FreeSans 300 0 0 0 S
flabel comment s 251 2000 251 2000 0 FreeSans 300 0 0 0 D
flabel comment s 711 1967 711 1967 0 FreeSans 300 0 0 0 S
flabel comment s 1171 2000 1171 2000 0 FreeSans 300 0 0 0 D
flabel comment s 1631 1967 1631 1967 0 FreeSans 300 0 0 0 S
flabel comment s 2091 2000 2091 2000 0 FreeSans 300 0 0 0 D
flabel comment s 2551 1967 2551 1967 0 FreeSans 300 0 0 0 S
flabel comment s 3011 2000 3011 2000 0 FreeSans 300 0 0 0 D
flabel comment s 3471 1967 3471 1967 0 FreeSans 300 0 0 0 S
flabel comment s 3931 2000 3931 2000 0 FreeSans 300 0 0 0 D
flabel comment s 4391 1967 4391 1967 0 FreeSans 300 0 0 0 S
flabel comment s 4851 2000 4851 2000 0 FreeSans 300 0 0 0 D
flabel comment s 5311 1967 5311 1967 0 FreeSans 300 0 0 0 S
flabel comment s 5771 2000 5771 2000 0 FreeSans 300 0 0 0 D
flabel comment s 6231 1967 6231 1967 0 FreeSans 300 0 0 0 S
flabel comment s 6691 2000 6691 2000 0 FreeSans 300 0 0 0 D
flabel comment s 7151 1967 7151 1967 0 FreeSans 300 0 0 0 S
flabel comment s 7611 2000 7611 2000 0 FreeSans 300 0 0 0 D
flabel comment s 8071 1967 8071 1967 0 FreeSans 300 0 0 0 S
flabel comment s 8531 2000 8531 2000 0 FreeSans 300 0 0 0 D
flabel comment s 8991 1967 8991 1967 0 FreeSans 300 0 0 0 S
flabel comment s 9451 2000 9451 2000 0 FreeSans 300 0 0 0 D
flabel comment s 9843 1973 9843 1973 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 34463156
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 34451652
<< end >>
