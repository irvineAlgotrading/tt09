magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -36 679 294 1471
<< poly >>
rect 114 702 144 1113
rect 48 686 144 702
rect 48 652 64 686
rect 98 652 144 686
rect 48 636 144 652
rect 114 149 144 636
<< polycont >>
rect 64 652 98 686
<< locali >>
rect 0 1397 258 1431
rect 62 1218 96 1397
rect 64 686 98 702
rect 64 636 98 652
rect 162 686 196 1284
rect 162 652 213 686
rect 162 54 196 652
rect 62 17 96 54
rect 0 -17 258 17
use contact_12  contact_12_0
timestamp 1704896540
transform 1 0 48 0 1 636
box 0 0 1 1
use nmos_m1_w0_360_sli_dli_da_p  nmos_m1_w0_360_sli_dli_da_p_0
timestamp 1704896540
transform 1 0 54 0 1 51
box -26 -26 176 98
use pmos_m1_w1_120_sli_dli_da_p  pmos_m1_w1_120_sli_dli_da_p_0
timestamp 1704896540
transform 1 0 54 0 1 1139
box -59 -54 209 278
<< labels >>
rlabel locali s 196 669 196 669 4 Z
port 2 nsew
rlabel locali s 81 669 81 669 4 A
port 1 nsew
rlabel locali s 129 1414 129 1414 4 vdd
port 3 nsew
rlabel locali s 129 0 129 0 4 gnd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 258 1414
string GDS_END 4172490
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 4171096
<< end >>
