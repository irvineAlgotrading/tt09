magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< pwell >>
rect -76 -26 372 226
<< mvnmos >>
rect 0 0 120 200
rect 176 0 296 200
<< mvndiff >>
rect -50 0 0 200
rect 120 182 176 200
rect 120 148 131 182
rect 165 148 176 182
rect 120 114 176 148
rect 120 80 131 114
rect 165 80 176 114
rect 120 46 176 80
rect 120 12 131 46
rect 165 12 176 46
rect 120 0 176 12
rect 296 0 346 200
<< mvndiffc >>
rect 131 148 165 182
rect 131 80 165 114
rect 131 12 165 46
<< poly >>
rect 0 200 120 226
rect 176 200 296 226
rect 0 -26 120 0
rect 176 -26 296 0
<< locali >>
rect 131 182 165 198
rect 131 114 165 148
rect 131 46 165 80
rect 131 -4 165 12
use hvDFL1sd2_CDNS_52468879185133  hvDFL1sd2_CDNS_52468879185133_0
timestamp 1704896540
transform 1 0 120 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s -25 100 -25 100 0 FreeSans 300 0 0 0 S
flabel comment s 148 97 148 97 0 FreeSans 300 0 0 0 D
flabel comment s 321 100 321 100 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 87661346
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 87660142
<< end >>
