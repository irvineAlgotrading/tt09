magic
tech sky130A
timestamp 1704896540
<< nwell >>
rect -18 -18 127 263
<< nsubdiff >>
rect 0 233 109 245
rect 0 12 12 233
rect 97 12 109 233
rect 0 0 109 12
<< nsubdiffcont >>
rect 12 12 97 233
<< locali >>
rect 12 233 97 241
rect 12 4 97 12
<< properties >>
string GDS_END 87769288
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 87767684
<< end >>
