magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< pwell >>
rect 15 163 787 545
<< nmoslvt >>
rect 171 189 201 519
rect 257 189 287 519
rect 343 189 373 519
rect 429 189 459 519
rect 515 189 545 519
rect 601 189 631 519
<< ndiff >>
rect 111 507 171 519
rect 111 473 126 507
rect 160 473 171 507
rect 111 439 171 473
rect 111 405 126 439
rect 160 405 171 439
rect 111 371 171 405
rect 111 337 126 371
rect 160 337 171 371
rect 111 303 171 337
rect 111 269 126 303
rect 160 269 171 303
rect 111 235 171 269
rect 111 201 126 235
rect 160 201 171 235
rect 111 189 171 201
rect 201 507 257 519
rect 201 473 212 507
rect 246 473 257 507
rect 201 439 257 473
rect 201 405 212 439
rect 246 405 257 439
rect 201 371 257 405
rect 201 337 212 371
rect 246 337 257 371
rect 201 303 257 337
rect 201 269 212 303
rect 246 269 257 303
rect 201 235 257 269
rect 201 201 212 235
rect 246 201 257 235
rect 201 189 257 201
rect 287 507 343 519
rect 287 473 298 507
rect 332 473 343 507
rect 287 439 343 473
rect 287 405 298 439
rect 332 405 343 439
rect 287 371 343 405
rect 287 337 298 371
rect 332 337 343 371
rect 287 303 343 337
rect 287 269 298 303
rect 332 269 343 303
rect 287 235 343 269
rect 287 201 298 235
rect 332 201 343 235
rect 287 189 343 201
rect 373 507 429 519
rect 373 473 384 507
rect 418 473 429 507
rect 373 439 429 473
rect 373 405 384 439
rect 418 405 429 439
rect 373 371 429 405
rect 373 337 384 371
rect 418 337 429 371
rect 373 303 429 337
rect 373 269 384 303
rect 418 269 429 303
rect 373 235 429 269
rect 373 201 384 235
rect 418 201 429 235
rect 373 189 429 201
rect 459 507 515 519
rect 459 473 470 507
rect 504 473 515 507
rect 459 439 515 473
rect 459 405 470 439
rect 504 405 515 439
rect 459 371 515 405
rect 459 337 470 371
rect 504 337 515 371
rect 459 303 515 337
rect 459 269 470 303
rect 504 269 515 303
rect 459 235 515 269
rect 459 201 470 235
rect 504 201 515 235
rect 459 189 515 201
rect 545 507 601 519
rect 545 473 556 507
rect 590 473 601 507
rect 545 439 601 473
rect 545 405 556 439
rect 590 405 601 439
rect 545 371 601 405
rect 545 337 556 371
rect 590 337 601 371
rect 545 303 601 337
rect 545 269 556 303
rect 590 269 601 303
rect 545 235 601 269
rect 545 201 556 235
rect 590 201 601 235
rect 545 189 601 201
rect 631 507 691 519
rect 631 473 642 507
rect 676 473 691 507
rect 631 439 691 473
rect 631 405 642 439
rect 676 405 691 439
rect 631 371 691 405
rect 631 337 642 371
rect 676 337 691 371
rect 631 303 691 337
rect 631 269 642 303
rect 676 269 691 303
rect 631 235 691 269
rect 631 201 642 235
rect 676 201 691 235
rect 631 189 691 201
<< ndiffc >>
rect 126 473 160 507
rect 126 405 160 439
rect 126 337 160 371
rect 126 269 160 303
rect 126 201 160 235
rect 212 473 246 507
rect 212 405 246 439
rect 212 337 246 371
rect 212 269 246 303
rect 212 201 246 235
rect 298 473 332 507
rect 298 405 332 439
rect 298 337 332 371
rect 298 269 332 303
rect 298 201 332 235
rect 384 473 418 507
rect 384 405 418 439
rect 384 337 418 371
rect 384 269 418 303
rect 384 201 418 235
rect 470 473 504 507
rect 470 405 504 439
rect 470 337 504 371
rect 470 269 504 303
rect 470 201 504 235
rect 556 473 590 507
rect 556 405 590 439
rect 556 337 590 371
rect 556 269 590 303
rect 556 201 590 235
rect 642 473 676 507
rect 642 405 676 439
rect 642 337 676 371
rect 642 269 676 303
rect 642 201 676 235
<< psubdiff >>
rect 41 507 111 519
rect 41 473 58 507
rect 92 473 111 507
rect 41 439 111 473
rect 41 405 58 439
rect 92 405 111 439
rect 41 371 111 405
rect 41 337 58 371
rect 92 337 111 371
rect 41 303 111 337
rect 41 269 58 303
rect 92 269 111 303
rect 41 235 111 269
rect 41 201 58 235
rect 92 201 111 235
rect 41 189 111 201
rect 691 507 761 519
rect 691 473 710 507
rect 744 473 761 507
rect 691 439 761 473
rect 691 405 710 439
rect 744 405 761 439
rect 691 371 761 405
rect 691 337 710 371
rect 744 337 761 371
rect 691 303 761 337
rect 691 269 710 303
rect 744 269 761 303
rect 691 235 761 269
rect 691 201 710 235
rect 744 201 761 235
rect 691 189 761 201
<< psubdiffcont >>
rect 58 473 92 507
rect 58 405 92 439
rect 58 337 92 371
rect 58 269 92 303
rect 58 201 92 235
rect 710 473 744 507
rect 710 405 744 439
rect 710 337 744 371
rect 710 269 744 303
rect 710 201 744 235
<< poly >>
rect 243 687 559 708
rect 243 653 264 687
rect 298 653 344 687
rect 378 653 424 687
rect 458 653 504 687
rect 538 653 559 687
rect 243 619 559 653
rect 120 595 201 611
rect 120 561 136 595
rect 170 561 201 595
rect 243 585 264 619
rect 298 585 344 619
rect 378 585 424 619
rect 458 585 504 619
rect 538 585 559 619
rect 243 569 559 585
rect 601 595 682 611
rect 120 545 201 561
rect 171 519 201 545
rect 257 519 287 569
rect 343 519 373 569
rect 429 519 459 569
rect 515 519 545 569
rect 601 561 632 595
rect 666 561 682 595
rect 601 545 682 561
rect 601 519 631 545
rect 171 163 201 189
rect 120 147 201 163
rect 120 113 136 147
rect 170 113 201 147
rect 257 139 287 189
rect 343 139 373 189
rect 429 139 459 189
rect 515 139 545 189
rect 601 163 631 189
rect 601 147 682 163
rect 120 97 201 113
rect 243 123 559 139
rect 243 89 264 123
rect 298 89 344 123
rect 378 89 424 123
rect 458 89 504 123
rect 538 89 559 123
rect 601 113 632 147
rect 666 113 682 147
rect 601 97 682 113
rect 243 55 559 89
rect 243 21 264 55
rect 298 21 344 55
rect 378 21 424 55
rect 458 21 504 55
rect 538 21 559 55
rect 243 0 559 21
<< polycont >>
rect 264 653 298 687
rect 344 653 378 687
rect 424 653 458 687
rect 504 653 538 687
rect 136 561 170 595
rect 264 585 298 619
rect 344 585 378 619
rect 424 585 458 619
rect 504 585 538 619
rect 632 561 666 595
rect 136 113 170 147
rect 264 89 298 123
rect 344 89 378 123
rect 424 89 458 123
rect 504 89 538 123
rect 632 113 666 147
rect 264 21 298 55
rect 344 21 378 55
rect 424 21 458 55
rect 504 21 538 55
<< locali >>
rect 243 689 559 708
rect 243 655 255 689
rect 289 687 337 689
rect 371 687 431 689
rect 465 687 513 689
rect 298 655 337 687
rect 243 653 264 655
rect 298 653 344 655
rect 378 653 424 687
rect 465 655 504 687
rect 547 655 559 689
rect 458 653 504 655
rect 538 653 559 655
rect 243 619 559 653
rect 243 617 264 619
rect 298 617 344 619
rect 120 595 186 611
rect 120 561 136 595
rect 170 561 186 595
rect 243 583 255 617
rect 298 585 337 617
rect 378 585 424 619
rect 458 617 504 619
rect 538 617 559 619
rect 465 585 504 617
rect 289 583 337 585
rect 371 583 431 585
rect 465 583 513 585
rect 547 583 559 617
rect 243 569 559 583
rect 616 595 682 611
rect 120 545 186 561
rect 616 561 632 595
rect 666 561 682 595
rect 616 545 682 561
rect 120 523 160 545
rect 642 523 682 545
rect 41 507 160 523
rect 41 473 58 507
rect 92 479 126 507
rect 94 473 126 479
rect 41 445 60 473
rect 94 445 160 473
rect 41 439 160 445
rect 41 405 58 439
rect 92 407 126 439
rect 94 405 126 407
rect 41 373 60 405
rect 94 373 160 405
rect 41 371 160 373
rect 41 337 58 371
rect 92 337 126 371
rect 41 335 160 337
rect 41 303 60 335
rect 94 303 160 335
rect 41 269 58 303
rect 94 301 126 303
rect 92 269 126 301
rect 41 263 160 269
rect 41 235 60 263
rect 94 235 160 263
rect 41 201 58 235
rect 94 229 126 235
rect 92 201 126 229
rect 41 185 160 201
rect 212 507 246 523
rect 212 439 246 445
rect 212 371 246 373
rect 212 335 246 337
rect 212 263 246 269
rect 212 185 246 201
rect 298 507 332 523
rect 298 439 332 445
rect 298 371 332 373
rect 298 335 332 337
rect 298 263 332 269
rect 298 185 332 201
rect 384 507 418 523
rect 384 439 418 445
rect 384 371 418 373
rect 384 335 418 337
rect 384 263 418 269
rect 384 185 418 201
rect 470 507 504 523
rect 470 439 504 445
rect 470 371 504 373
rect 470 335 504 337
rect 470 263 504 269
rect 470 185 504 201
rect 556 507 590 523
rect 556 439 590 445
rect 556 371 590 373
rect 556 335 590 337
rect 556 263 590 269
rect 556 185 590 201
rect 642 507 761 523
rect 676 479 710 507
rect 676 473 708 479
rect 744 473 761 507
rect 642 445 708 473
rect 742 445 761 473
rect 642 439 761 445
rect 676 407 710 439
rect 676 405 708 407
rect 744 405 761 439
rect 642 373 708 405
rect 742 373 761 405
rect 642 371 761 373
rect 676 337 710 371
rect 744 337 761 371
rect 642 335 761 337
rect 642 303 708 335
rect 742 303 761 335
rect 676 301 708 303
rect 676 269 710 301
rect 744 269 761 303
rect 642 263 761 269
rect 642 235 708 263
rect 742 235 761 263
rect 676 229 708 235
rect 676 201 710 229
rect 744 201 761 235
rect 642 185 761 201
rect 120 163 160 185
rect 642 163 682 185
rect 120 147 186 163
rect 120 113 136 147
rect 170 113 186 147
rect 616 147 682 163
rect 120 97 186 113
rect 243 125 559 139
rect 243 91 255 125
rect 289 123 337 125
rect 371 123 431 125
rect 465 123 513 125
rect 298 91 337 123
rect 243 89 264 91
rect 298 89 344 91
rect 378 89 424 123
rect 465 91 504 123
rect 547 91 559 125
rect 616 113 632 147
rect 666 113 682 147
rect 616 97 682 113
rect 458 89 504 91
rect 538 89 559 91
rect 243 55 559 89
rect 243 53 264 55
rect 298 53 344 55
rect 243 19 255 53
rect 298 21 337 53
rect 378 21 424 55
rect 458 53 504 55
rect 538 53 559 55
rect 465 21 504 53
rect 289 19 337 21
rect 371 19 431 21
rect 465 19 513 21
rect 547 19 559 53
rect 243 0 559 19
<< viali >>
rect 255 687 289 689
rect 337 687 371 689
rect 431 687 465 689
rect 513 687 547 689
rect 255 655 264 687
rect 264 655 289 687
rect 337 655 344 687
rect 344 655 371 687
rect 431 655 458 687
rect 458 655 465 687
rect 513 655 538 687
rect 538 655 547 687
rect 255 585 264 617
rect 264 585 289 617
rect 337 585 344 617
rect 344 585 371 617
rect 431 585 458 617
rect 458 585 465 617
rect 513 585 538 617
rect 538 585 547 617
rect 255 583 289 585
rect 337 583 371 585
rect 431 583 465 585
rect 513 583 547 585
rect 60 473 92 479
rect 92 473 94 479
rect 60 445 94 473
rect 60 405 92 407
rect 92 405 94 407
rect 60 373 94 405
rect 60 303 94 335
rect 60 301 92 303
rect 92 301 94 303
rect 60 235 94 263
rect 60 229 92 235
rect 92 229 94 235
rect 212 473 246 479
rect 212 445 246 473
rect 212 405 246 407
rect 212 373 246 405
rect 212 303 246 335
rect 212 301 246 303
rect 212 235 246 263
rect 212 229 246 235
rect 298 473 332 479
rect 298 445 332 473
rect 298 405 332 407
rect 298 373 332 405
rect 298 303 332 335
rect 298 301 332 303
rect 298 235 332 263
rect 298 229 332 235
rect 384 473 418 479
rect 384 445 418 473
rect 384 405 418 407
rect 384 373 418 405
rect 384 303 418 335
rect 384 301 418 303
rect 384 235 418 263
rect 384 229 418 235
rect 470 473 504 479
rect 470 445 504 473
rect 470 405 504 407
rect 470 373 504 405
rect 470 303 504 335
rect 470 301 504 303
rect 470 235 504 263
rect 470 229 504 235
rect 556 473 590 479
rect 556 445 590 473
rect 556 405 590 407
rect 556 373 590 405
rect 556 303 590 335
rect 556 301 590 303
rect 556 235 590 263
rect 556 229 590 235
rect 708 473 710 479
rect 710 473 742 479
rect 708 445 742 473
rect 708 405 710 407
rect 710 405 742 407
rect 708 373 742 405
rect 708 303 742 335
rect 708 301 710 303
rect 710 301 742 303
rect 708 235 742 263
rect 708 229 710 235
rect 710 229 742 235
rect 255 123 289 125
rect 337 123 371 125
rect 431 123 465 125
rect 513 123 547 125
rect 255 91 264 123
rect 264 91 289 123
rect 337 91 344 123
rect 344 91 371 123
rect 431 91 458 123
rect 458 91 465 123
rect 513 91 538 123
rect 538 91 547 123
rect 255 21 264 53
rect 264 21 289 53
rect 337 21 344 53
rect 344 21 371 53
rect 431 21 458 53
rect 458 21 465 53
rect 513 21 538 53
rect 538 21 547 53
rect 255 19 289 21
rect 337 19 371 21
rect 431 19 465 21
rect 513 19 547 21
<< metal1 >>
rect 243 689 559 708
rect 243 655 255 689
rect 289 655 337 689
rect 371 655 431 689
rect 465 655 513 689
rect 547 655 559 689
rect 243 617 559 655
rect 243 583 255 617
rect 289 583 337 617
rect 371 583 431 617
rect 465 583 513 617
rect 547 583 559 617
rect 243 571 559 583
rect 41 479 100 507
rect 41 445 60 479
rect 94 445 100 479
rect 41 407 100 445
rect 41 373 60 407
rect 94 373 100 407
rect 41 335 100 373
rect 41 301 60 335
rect 94 301 100 335
rect 41 263 100 301
rect 41 229 60 263
rect 94 229 100 263
rect 41 201 100 229
rect 203 479 255 507
rect 203 445 212 479
rect 246 445 255 479
rect 203 407 255 445
rect 203 373 212 407
rect 246 373 255 407
rect 203 335 255 373
rect 203 323 212 335
rect 246 323 255 335
rect 203 263 255 271
rect 203 259 212 263
rect 246 259 255 263
rect 203 201 255 207
rect 289 501 341 507
rect 289 445 298 449
rect 332 445 341 449
rect 289 437 341 445
rect 289 373 298 385
rect 332 373 341 385
rect 289 335 341 373
rect 289 301 298 335
rect 332 301 341 335
rect 289 263 341 301
rect 289 229 298 263
rect 332 229 341 263
rect 289 201 341 229
rect 375 479 427 507
rect 375 445 384 479
rect 418 445 427 479
rect 375 407 427 445
rect 375 373 384 407
rect 418 373 427 407
rect 375 335 427 373
rect 375 323 384 335
rect 418 323 427 335
rect 375 263 427 271
rect 375 259 384 263
rect 418 259 427 263
rect 375 201 427 207
rect 461 501 513 507
rect 461 445 470 449
rect 504 445 513 449
rect 461 437 513 445
rect 461 373 470 385
rect 504 373 513 385
rect 461 335 513 373
rect 461 301 470 335
rect 504 301 513 335
rect 461 263 513 301
rect 461 229 470 263
rect 504 229 513 263
rect 461 201 513 229
rect 547 479 599 507
rect 547 445 556 479
rect 590 445 599 479
rect 547 407 599 445
rect 547 373 556 407
rect 590 373 599 407
rect 547 335 599 373
rect 547 323 556 335
rect 590 323 599 335
rect 547 263 599 271
rect 547 259 556 263
rect 590 259 599 263
rect 547 201 599 207
rect 702 479 761 507
rect 702 445 708 479
rect 742 445 761 479
rect 702 407 761 445
rect 702 373 708 407
rect 742 373 761 407
rect 702 335 761 373
rect 702 301 708 335
rect 742 301 761 335
rect 702 263 761 301
rect 702 229 708 263
rect 742 229 761 263
rect 702 201 761 229
rect 243 125 559 137
rect 243 91 255 125
rect 289 91 337 125
rect 371 91 431 125
rect 465 91 513 125
rect 547 91 559 125
rect 243 53 559 91
rect 243 19 255 53
rect 289 19 337 53
rect 371 19 431 53
rect 465 19 513 53
rect 547 19 559 53
rect 243 0 559 19
<< via1 >>
rect 203 301 212 323
rect 212 301 246 323
rect 246 301 255 323
rect 203 271 255 301
rect 203 229 212 259
rect 212 229 246 259
rect 246 229 255 259
rect 203 207 255 229
rect 289 479 341 501
rect 289 449 298 479
rect 298 449 332 479
rect 332 449 341 479
rect 289 407 341 437
rect 289 385 298 407
rect 298 385 332 407
rect 332 385 341 407
rect 375 301 384 323
rect 384 301 418 323
rect 418 301 427 323
rect 375 271 427 301
rect 375 229 384 259
rect 384 229 418 259
rect 418 229 427 259
rect 375 207 427 229
rect 461 479 513 501
rect 461 449 470 479
rect 470 449 504 479
rect 504 449 513 479
rect 461 407 513 437
rect 461 385 470 407
rect 470 385 504 407
rect 504 385 513 407
rect 547 301 556 323
rect 556 301 590 323
rect 590 301 599 323
rect 547 271 599 301
rect 547 229 556 259
rect 556 229 590 259
rect 590 229 599 259
rect 547 207 599 229
<< metal2 >>
rect 14 501 788 507
rect 14 449 289 501
rect 341 449 461 501
rect 513 449 788 501
rect 14 437 788 449
rect 14 385 289 437
rect 341 385 461 437
rect 513 385 788 437
rect 14 379 788 385
rect 14 323 788 329
rect 14 271 203 323
rect 255 271 375 323
rect 427 271 547 323
rect 599 271 788 323
rect 14 259 788 271
rect 14 207 203 259
rect 255 207 375 259
rect 427 207 547 259
rect 599 207 788 259
rect 14 201 788 207
<< labels >>
flabel comment s 184 356 184 356 0 FreeSans 180 90 0 0 dummy_poly
flabel comment s 612 355 612 355 0 FreeSans 180 90 0 0 dummy_poly
flabel metal1 s 301 606 511 656 0 FreeSans 200 0 0 0 GATE
port 3 nsew
flabel metal1 s 301 42 511 92 0 FreeSans 200 0 0 0 GATE
port 3 nsew
flabel metal1 s 715 339 761 369 0 FreeSans 200 90 0 0 SUBSTRATE
port 2 nsew
flabel metal1 s 41 339 87 369 0 FreeSans 200 90 0 0 SUBSTRATE
port 2 nsew
flabel metal2 s 14 201 35 329 7 FreeSans 300 180 0 0 SOURCE
port 4 nsew
flabel metal2 s 14 379 35 507 7 FreeSans 300 180 0 0 DRAIN
port 5 nsew
<< properties >>
string GDS_END 6251654
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 6236730
<< end >>
