magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 1 21 779 203
rect 30 -17 64 21
<< locali >>
rect 459 349 493 425
rect 627 349 661 425
rect 459 289 811 349
rect 28 215 360 255
rect 424 215 697 255
rect 731 181 811 289
rect 107 145 811 181
rect 107 51 173 145
rect 275 51 341 145
rect 443 51 509 145
rect 611 51 677 145
<< obsli1 >>
rect 0 527 828 561
rect 18 333 73 493
rect 107 367 173 527
rect 207 333 241 493
rect 275 367 325 527
rect 359 459 778 493
rect 359 333 425 459
rect 18 291 425 333
rect 527 387 593 459
rect 695 383 778 459
rect 18 17 73 181
rect 207 17 241 111
rect 375 17 409 111
rect 543 17 577 111
rect 711 17 768 111
rect 0 -17 828 17
<< metal1 >>
rect 0 496 828 592
rect 0 -48 828 48
<< labels >>
rlabel locali s 28 215 360 255 6 A
port 1 nsew signal input
rlabel locali s 424 215 697 255 6 B
port 2 nsew signal input
rlabel metal1 s 0 -48 828 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 1 21 779 203 6 VNB
port 4 nsew ground bidirectional
rlabel nwell s -38 261 866 582 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 496 828 592 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 611 51 677 145 6 Y
port 7 nsew signal output
rlabel locali s 443 51 509 145 6 Y
port 7 nsew signal output
rlabel locali s 275 51 341 145 6 Y
port 7 nsew signal output
rlabel locali s 107 51 173 145 6 Y
port 7 nsew signal output
rlabel locali s 107 145 811 181 6 Y
port 7 nsew signal output
rlabel locali s 731 181 811 289 6 Y
port 7 nsew signal output
rlabel locali s 459 289 811 349 6 Y
port 7 nsew signal output
rlabel locali s 627 349 661 425 6 Y
port 7 nsew signal output
rlabel locali s 459 349 493 425 6 Y
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 828 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1964744
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1957698
<< end >>
