magic
tech sky130A
timestamp 1704896540
<< metal1 >>
rect 0 0 3 90
rect 93 0 96 90
<< via1 >>
rect 3 0 93 90
<< metal2 >>
rect 0 0 3 90
rect 93 0 96 90
<< properties >>
string GDS_END 78447090
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 78446382
<< end >>
