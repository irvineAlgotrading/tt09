magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -38 261 2890 582
<< pwell >>
rect 2382 201 2851 203
rect 1240 157 1694 201
rect 2015 157 2851 201
rect 1 21 2851 157
rect 29 -17 63 21
<< locali >>
rect 17 195 87 325
rect 288 205 344 337
rect 392 203 436 339
rect 765 265 805 475
rect 392 169 483 203
rect 392 69 436 169
rect 2500 326 2557 493
rect 2307 219 2398 265
rect 2521 143 2557 326
rect 2500 51 2557 143
rect 2783 321 2835 493
rect 2793 165 2835 321
rect 2783 51 2835 165
<< obsli1 >>
rect 0 527 2852 561
rect 34 393 69 493
rect 103 427 169 527
rect 34 359 167 393
rect 121 161 167 359
rect 34 127 167 161
rect 34 69 69 127
rect 103 17 169 93
rect 203 69 248 493
rect 291 377 357 527
rect 447 375 513 477
rect 579 381 613 493
rect 662 443 728 527
rect 470 273 513 375
rect 549 349 613 381
rect 549 315 729 349
rect 470 237 615 273
rect 517 215 615 237
rect 695 219 729 315
rect 291 17 341 127
rect 517 119 551 215
rect 695 159 754 219
rect 470 53 551 119
rect 585 153 754 159
rect 585 125 729 153
rect 585 61 625 125
rect 674 17 740 89
rect 846 61 891 493
rect 927 450 1093 484
rect 925 315 1025 391
rect 925 141 969 315
rect 1059 281 1093 450
rect 1141 441 1217 527
rect 1277 407 1311 475
rect 1127 357 1397 407
rect 1435 383 1501 527
rect 1710 450 1876 484
rect 1924 451 2000 527
rect 1127 315 1177 357
rect 1279 281 1329 297
rect 1059 247 1329 281
rect 1059 239 1143 247
rect 1005 129 1075 203
rect 1109 93 1143 239
rect 1285 231 1329 247
rect 1363 213 1397 357
rect 1431 283 1632 331
rect 1672 315 1719 397
rect 1431 247 1497 283
rect 1767 261 1808 381
rect 1559 213 1625 247
rect 1177 193 1243 213
rect 1177 147 1259 193
rect 1363 179 1625 213
rect 1684 225 1808 261
rect 1842 281 1876 450
rect 2048 417 2082 475
rect 2188 451 2466 527
rect 1910 383 2466 417
rect 1910 315 1960 383
rect 1842 247 2112 281
rect 1363 153 1406 179
rect 1340 119 1406 153
rect 940 53 1143 93
rect 1177 17 1211 105
rect 1245 85 1311 93
rect 1440 85 1479 143
rect 1684 141 1741 225
rect 1842 93 1876 247
rect 2068 215 2112 247
rect 1951 147 2026 213
rect 2146 163 2181 383
rect 2115 129 2181 163
rect 2216 315 2371 349
rect 2216 185 2271 315
rect 2432 265 2466 383
rect 2432 199 2485 265
rect 2216 151 2353 185
rect 1245 51 1479 85
rect 1528 17 1595 93
rect 1723 53 1876 93
rect 1912 17 1964 105
rect 2016 85 2086 93
rect 2215 85 2250 117
rect 2016 51 2250 85
rect 2313 53 2353 151
rect 2400 17 2466 161
rect 2592 265 2655 483
rect 2690 353 2749 527
rect 2592 199 2759 265
rect 2592 51 2655 199
rect 2691 17 2749 109
rect 0 -17 2852 17
<< metal1 >>
rect 0 496 2852 592
rect 1213 184 1271 193
rect 1949 184 2007 193
rect 1213 156 2007 184
rect 1213 147 1271 156
rect 1949 147 2007 156
rect 0 -48 2852 48
<< obsm1 >>
rect 109 388 167 397
rect 937 388 995 397
rect 1673 388 1731 397
rect 109 360 1731 388
rect 109 351 167 360
rect 937 351 995 360
rect 1673 351 1731 360
rect 1581 320 1639 329
rect 2225 320 2283 329
rect 1581 292 2283 320
rect 1581 283 1639 292
rect 2225 283 2283 292
rect 569 252 627 261
rect 845 252 903 261
rect 1673 252 1731 261
rect 569 224 903 252
rect 569 215 627 224
rect 845 215 903 224
rect 1044 224 1731 252
rect 1044 193 1087 224
rect 1673 215 1731 224
rect 201 184 259 193
rect 1029 184 1087 193
rect 201 156 1087 184
rect 201 147 259 156
rect 1029 147 1087 156
<< labels >>
rlabel locali s 17 195 87 325 6 CLK
port 1 nsew clock input
rlabel locali s 765 265 805 475 6 D
port 2 nsew signal input
rlabel locali s 2307 219 2398 265 6 RESET_B
port 3 nsew signal input
rlabel locali s 288 205 344 337 6 SCD
port 4 nsew signal input
rlabel locali s 392 69 436 169 6 SCE
port 5 nsew signal input
rlabel locali s 392 169 483 203 6 SCE
port 5 nsew signal input
rlabel locali s 392 203 436 339 6 SCE
port 5 nsew signal input
rlabel metal1 s 1949 147 2007 156 6 SET_B
port 6 nsew signal input
rlabel metal1 s 1213 147 1271 156 6 SET_B
port 6 nsew signal input
rlabel metal1 s 1213 156 2007 184 6 SET_B
port 6 nsew signal input
rlabel metal1 s 1949 184 2007 193 6 SET_B
port 6 nsew signal input
rlabel metal1 s 1213 184 1271 193 6 SET_B
port 6 nsew signal input
rlabel metal1 s 0 -48 2852 48 8 VGND
port 7 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 8 nsew ground bidirectional
rlabel pwell s 1 21 2851 157 6 VNB
port 8 nsew ground bidirectional
rlabel pwell s 2015 157 2851 201 6 VNB
port 8 nsew ground bidirectional
rlabel pwell s 1240 157 1694 201 6 VNB
port 8 nsew ground bidirectional
rlabel pwell s 2382 201 2851 203 6 VNB
port 8 nsew ground bidirectional
rlabel nwell s -38 261 2890 582 6 VPB
port 9 nsew power bidirectional
rlabel metal1 s 0 496 2852 592 6 VPWR
port 10 nsew power bidirectional abutment
rlabel locali s 2783 51 2835 165 6 Q
port 11 nsew signal output
rlabel locali s 2793 165 2835 321 6 Q
port 11 nsew signal output
rlabel locali s 2783 321 2835 493 6 Q
port 11 nsew signal output
rlabel locali s 2500 51 2557 143 6 Q_N
port 12 nsew signal output
rlabel locali s 2521 143 2557 326 6 Q_N
port 12 nsew signal output
rlabel locali s 2500 326 2557 493 6 Q_N
port 12 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2852 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 240892
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 218578
<< end >>
