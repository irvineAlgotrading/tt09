magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -42 415 569 1122
<< poly >>
rect 119 790 239 799
rect 105 774 239 790
rect 105 740 121 774
rect 155 740 189 774
rect 223 740 239 774
rect 105 724 239 740
rect 119 708 239 724
rect 295 790 415 798
rect 295 774 429 790
rect 295 740 311 774
rect 345 740 379 774
rect 413 740 429 774
rect 295 724 429 740
rect 295 708 415 724
rect 119 434 239 496
rect 119 400 165 434
rect 199 400 239 434
rect 119 366 239 400
rect 119 332 165 366
rect 199 332 239 366
rect 119 306 239 332
rect 295 434 415 496
rect 295 400 336 434
rect 370 400 415 434
rect 295 366 415 400
rect 295 332 336 366
rect 370 332 415 366
rect 295 310 415 332
<< polycont >>
rect 121 740 155 774
rect 189 740 223 774
rect 311 740 345 774
rect 379 740 413 774
rect 165 400 199 434
rect 165 332 199 366
rect 336 400 370 434
rect 336 332 370 366
<< locali >>
rect 74 1042 108 1043
rect 74 970 108 1008
rect 74 924 108 936
rect 426 971 460 1009
rect 426 920 460 937
rect 247 834 285 868
rect 105 740 121 774
rect 155 740 189 774
rect 223 740 239 774
rect 295 740 311 774
rect 345 740 379 774
rect 413 740 429 774
rect 74 628 108 666
rect 149 434 215 740
rect 250 554 284 592
rect 149 400 165 434
rect 199 400 215 434
rect 149 366 215 400
rect 149 332 165 366
rect 199 332 215 366
rect 320 434 386 740
rect 426 598 460 636
rect 320 400 336 434
rect 370 400 386 434
rect 320 366 386 400
rect 320 332 336 366
rect 370 332 386 366
rect 423 254 461 288
rect 74 136 108 174
<< viali >>
rect 74 1008 108 1042
rect 74 936 108 970
rect 426 1009 460 1043
rect 426 937 460 971
rect 213 834 247 868
rect 285 834 319 868
rect 74 666 108 700
rect 74 594 108 628
rect 250 592 284 626
rect 250 520 284 554
rect 426 636 460 670
rect 426 564 460 598
rect 389 254 423 288
rect 461 254 495 288
rect 74 174 108 208
rect 74 102 108 136
<< metal1 >>
rect 25 1043 503 1127
rect 25 1042 426 1043
rect 25 1008 74 1042
rect 108 1009 426 1042
rect 460 1009 503 1043
rect 108 1008 503 1009
rect 25 971 503 1008
rect 25 970 426 971
rect 25 936 74 970
rect 108 937 426 970
rect 460 937 503 971
rect 108 936 503 937
rect 25 924 503 936
rect 68 700 114 924
rect 201 868 331 874
rect 201 834 213 868
rect 247 834 285 868
rect 319 834 331 868
rect 201 828 331 834
rect 68 666 74 700
rect 108 666 114 700
rect 68 628 114 666
rect 68 594 74 628
rect 108 594 114 628
rect 68 582 114 594
rect 244 626 290 828
rect 244 592 250 626
rect 284 592 290 626
rect 244 554 290 592
rect 244 520 250 554
rect 284 520 290 554
rect 420 670 466 924
rect 420 636 426 670
rect 460 636 466 670
rect 420 598 466 636
rect 420 564 426 598
rect 460 564 466 598
rect 420 552 466 564
rect 244 294 290 520
rect 244 288 507 294
rect 244 254 389 288
rect 423 254 461 288
rect 495 254 507 288
rect 244 248 507 254
rect 24 208 503 220
rect 24 174 74 208
rect 108 174 503 208
rect 24 136 503 174
rect 24 102 74 136
rect 108 102 503 136
rect 24 24 503 102
use L1M1_CDNS_559591418084  L1M1_CDNS_559591418084_0
timestamp 1704896540
transform 0 -1 460 1 0 937
box 0 0 1 1
use L1M1_CDNS_559591418084  L1M1_CDNS_559591418084_1
timestamp 1704896540
transform 0 -1 108 -1 0 208
box 0 0 1 1
use nfet_CDNS_559591418087  nfet_CDNS_559591418087_0
timestamp 1704896540
transform 1 0 295 0 -1 284
box -76 -26 199 166
use nfet_CDNS_559591418089  nfet_CDNS_559591418089_0
timestamp 1704896540
transform 1 0 119 0 -1 284
box -79 -26 196 166
use pfet_CDNS_559591418085  pfet_CDNS_559591418085_0
timestamp 1704896540
transform 1 0 119 0 -1 1022
box -119 -66 239 266
use pfet_CDNS_559591418085  pfet_CDNS_559591418085_1
timestamp 1704896540
transform 1 0 295 0 -1 1022
box -119 -66 239 266
use pfet_CDNS_559591418085  pfet_CDNS_559591418085_2
timestamp 1704896540
transform 1 0 119 0 -1 682
box -119 -66 239 266
use pfet_CDNS_559591418085  pfet_CDNS_559591418085_3
timestamp 1704896540
transform 1 0 295 0 -1 682
box -119 -66 239 266
use PYL1_CDNS_559591418083  PYL1_CDNS_559591418083_0
timestamp 1704896540
transform 0 -1 386 1 0 316
box 0 0 1 1
use PYL1_CDNS_559591418083  PYL1_CDNS_559591418083_1
timestamp 1704896540
transform 0 -1 215 1 0 316
box 0 0 1 1
<< labels >>
flabel metal1 s 24 24 107 220 0 FreeSans 320 0 0 0 vgnd
port 2 nsew
flabel metal1 s 420 924 503 1127 0 FreeSans 320 0 0 0 vpwr
port 3 nsew
flabel locali s 156 353 207 394 0 FreeSans 400 0 0 0 in0
port 4 nsew
<< properties >>
string GDS_END 804178
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 799830
<< end >>
