magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -66 377 1698 897
<< pwell >>
rect 1191 217 1628 283
rect 45 43 1628 217
rect -26 -43 1658 43
<< mvnmos >>
rect 128 107 228 191
rect 284 107 384 191
rect 550 107 650 191
rect 706 107 806 191
rect 862 107 962 191
rect 1004 107 1104 191
rect 1270 173 1370 257
rect 1449 107 1549 257
<< mvpmos >>
rect 83 443 183 593
rect 297 443 397 593
rect 564 587 664 737
rect 735 587 835 737
rect 914 587 1014 671
rect 1056 587 1156 671
rect 1266 443 1366 527
rect 1445 443 1545 743
<< mvndiff >>
rect 1217 232 1270 257
rect 1217 198 1225 232
rect 1259 198 1270 232
rect 71 166 128 191
rect 71 132 83 166
rect 117 132 128 166
rect 71 107 128 132
rect 228 166 284 191
rect 228 132 239 166
rect 273 132 284 166
rect 228 107 284 132
rect 384 166 437 191
rect 384 132 395 166
rect 429 132 437 166
rect 384 107 437 132
rect 497 166 550 191
rect 497 132 505 166
rect 539 132 550 166
rect 497 107 550 132
rect 650 166 706 191
rect 650 132 661 166
rect 695 132 706 166
rect 650 107 706 132
rect 806 166 862 191
rect 806 132 817 166
rect 851 132 862 166
rect 806 107 862 132
rect 962 107 1004 191
rect 1104 166 1157 191
rect 1217 173 1270 198
rect 1370 249 1449 257
rect 1370 215 1404 249
rect 1438 215 1449 249
rect 1370 173 1449 215
rect 1104 132 1115 166
rect 1149 132 1157 166
rect 1392 149 1449 173
rect 1104 107 1157 132
rect 1392 115 1404 149
rect 1438 115 1449 149
rect 1392 107 1449 115
rect 1549 245 1602 257
rect 1549 211 1560 245
rect 1594 211 1602 245
rect 1549 153 1602 211
rect 1549 119 1560 153
rect 1594 119 1602 153
rect 1549 107 1602 119
<< mvpdiff >>
rect 510 725 564 737
rect 510 691 518 725
rect 552 691 564 725
rect 510 633 564 691
rect 510 599 518 633
rect 552 599 564 633
rect 30 581 83 593
rect 30 547 38 581
rect 72 547 83 581
rect 30 489 83 547
rect 30 455 38 489
rect 72 455 83 489
rect 30 443 83 455
rect 183 585 297 593
rect 183 551 194 585
rect 228 551 297 585
rect 183 485 297 551
rect 183 451 194 485
rect 228 451 297 485
rect 183 443 297 451
rect 397 491 450 593
rect 510 587 564 599
rect 664 660 735 737
rect 664 626 690 660
rect 724 626 735 660
rect 664 587 735 626
rect 835 729 892 737
rect 835 695 846 729
rect 880 695 892 729
rect 1388 735 1445 743
rect 1388 701 1400 735
rect 1434 701 1445 735
rect 835 671 892 695
rect 835 629 914 671
rect 835 595 846 629
rect 880 595 914 629
rect 835 587 914 595
rect 1014 587 1056 671
rect 1156 646 1213 671
rect 1156 612 1167 646
rect 1201 612 1213 646
rect 1156 587 1213 612
rect 1388 638 1445 701
rect 1388 604 1400 638
rect 1434 604 1445 638
rect 397 457 408 491
rect 442 457 450 491
rect 397 443 450 457
rect 1388 541 1445 604
rect 1388 527 1400 541
rect 1209 502 1266 527
rect 1209 468 1221 502
rect 1255 468 1266 502
rect 1209 443 1266 468
rect 1366 507 1400 527
rect 1434 507 1445 541
rect 1366 443 1445 507
rect 1545 735 1602 743
rect 1545 701 1556 735
rect 1590 701 1602 735
rect 1545 652 1602 701
rect 1545 618 1556 652
rect 1590 618 1602 652
rect 1545 568 1602 618
rect 1545 534 1556 568
rect 1590 534 1602 568
rect 1545 485 1602 534
rect 1545 451 1556 485
rect 1590 451 1602 485
rect 1545 443 1602 451
<< mvndiffc >>
rect 1225 198 1259 232
rect 83 132 117 166
rect 239 132 273 166
rect 395 132 429 166
rect 505 132 539 166
rect 661 132 695 166
rect 817 132 851 166
rect 1404 215 1438 249
rect 1115 132 1149 166
rect 1404 115 1438 149
rect 1560 211 1594 245
rect 1560 119 1594 153
<< mvpdiffc >>
rect 518 691 552 725
rect 518 599 552 633
rect 38 547 72 581
rect 38 455 72 489
rect 194 551 228 585
rect 194 451 228 485
rect 690 626 724 660
rect 846 695 880 729
rect 1400 701 1434 735
rect 846 595 880 629
rect 1167 612 1201 646
rect 1400 604 1434 638
rect 408 457 442 491
rect 1221 468 1255 502
rect 1400 507 1434 541
rect 1556 701 1590 735
rect 1556 618 1590 652
rect 1556 534 1590 568
rect 1556 451 1590 485
<< mvpsubdiff >>
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1632 831
<< mvpsubdiffcont >>
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
<< poly >>
rect 564 737 664 763
rect 735 737 835 763
rect 1445 743 1545 769
rect 83 593 183 619
rect 297 593 397 619
rect 914 671 1014 697
rect 1056 671 1156 697
rect 564 561 664 587
rect 550 477 664 561
rect 735 539 835 587
rect 914 561 1014 587
rect 735 505 760 539
rect 794 505 835 539
rect 735 485 835 505
rect 550 443 570 477
rect 604 443 664 477
rect 908 443 1014 561
rect 83 361 183 443
rect 297 417 397 443
rect 284 387 397 417
rect 83 341 228 361
rect 83 307 124 341
rect 158 307 228 341
rect 83 273 228 307
rect 83 239 124 273
rect 158 239 228 273
rect 83 217 228 239
rect 128 191 228 217
rect 284 353 324 387
rect 358 353 397 387
rect 284 319 397 353
rect 284 285 324 319
rect 358 285 397 319
rect 284 265 397 285
rect 550 409 664 443
rect 550 375 570 409
rect 604 375 664 409
rect 550 355 664 375
rect 706 397 1008 443
rect 706 394 812 397
rect 706 360 726 394
rect 760 360 812 394
rect 284 191 384 265
rect 550 191 650 355
rect 706 326 812 360
rect 706 292 726 326
rect 760 292 812 326
rect 706 272 812 292
rect 862 335 962 355
rect 862 301 898 335
rect 932 301 962 335
rect 1056 331 1156 587
rect 1266 527 1366 553
rect 1056 313 1102 331
rect 706 191 806 272
rect 862 267 962 301
rect 862 233 898 267
rect 932 233 962 267
rect 862 191 962 233
rect 1004 297 1102 313
rect 1136 297 1156 331
rect 1004 263 1156 297
rect 1266 417 1366 443
rect 1445 417 1545 443
rect 1266 395 1549 417
rect 1266 361 1286 395
rect 1320 361 1549 395
rect 1266 317 1549 361
rect 1266 283 1370 317
rect 1004 229 1102 263
rect 1136 229 1156 263
rect 1270 257 1370 283
rect 1449 257 1549 317
rect 1004 213 1156 229
rect 1004 191 1104 213
rect 1270 147 1370 173
rect 128 81 228 107
rect 284 81 384 107
rect 550 81 650 107
rect 706 81 806 107
rect 862 81 962 107
rect 1004 81 1104 107
rect 1449 81 1549 107
<< polycont >>
rect 760 505 794 539
rect 570 443 604 477
rect 124 307 158 341
rect 124 239 158 273
rect 324 353 358 387
rect 324 285 358 319
rect 570 375 604 409
rect 726 360 760 394
rect 726 292 760 326
rect 898 301 932 335
rect 898 233 932 267
rect 1102 297 1136 331
rect 1286 361 1320 395
rect 1102 229 1136 263
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1632 831
rect 108 735 286 741
rect 142 701 180 735
rect 214 701 252 735
rect 22 581 72 597
rect 22 547 38 581
rect 22 489 72 547
rect 22 455 38 489
rect 22 415 72 455
rect 108 585 286 701
rect 378 735 568 741
rect 378 701 384 735
rect 418 701 456 735
rect 490 725 528 735
rect 490 701 518 725
rect 562 701 568 735
rect 378 691 518 701
rect 552 691 568 701
rect 378 633 568 691
rect 378 599 518 633
rect 552 599 568 633
rect 604 727 810 761
rect 108 551 194 585
rect 228 551 286 585
rect 604 563 638 727
rect 108 485 286 551
rect 108 451 194 485
rect 228 451 286 485
rect 322 529 638 563
rect 674 660 740 691
rect 674 626 690 660
rect 724 626 740 660
rect 674 579 740 626
rect 322 415 356 529
rect 392 491 458 493
rect 392 457 408 491
rect 442 457 458 491
rect 392 439 458 457
rect 22 403 356 415
rect 22 387 359 403
rect 22 381 324 387
rect 22 199 72 381
rect 308 353 324 381
rect 358 353 359 387
rect 108 341 174 345
rect 108 307 124 341
rect 158 307 174 341
rect 108 273 174 307
rect 108 239 124 273
rect 158 239 174 273
rect 308 319 359 353
rect 308 285 324 319
rect 358 285 359 319
rect 308 269 359 285
rect 395 323 458 439
rect 505 477 620 493
rect 505 443 570 477
rect 604 443 620 477
rect 505 409 620 443
rect 674 467 708 579
rect 776 543 810 727
rect 846 729 896 745
rect 880 695 896 729
rect 846 629 896 695
rect 880 613 896 629
rect 1054 735 1244 741
rect 1054 701 1060 735
rect 1094 701 1132 735
rect 1166 701 1204 735
rect 1238 701 1244 735
rect 1054 646 1244 701
rect 880 595 1018 613
rect 846 579 1018 595
rect 1054 612 1167 646
rect 1201 612 1244 646
rect 1054 579 1244 612
rect 1307 735 1497 751
rect 1307 701 1313 735
rect 1347 701 1385 735
rect 1434 701 1457 735
rect 1491 701 1497 735
rect 1307 638 1497 701
rect 1307 604 1400 638
rect 1434 604 1497 638
rect 744 539 948 543
rect 744 505 760 539
rect 794 505 948 539
rect 744 503 948 505
rect 674 433 846 467
rect 505 375 570 409
rect 604 375 620 409
rect 505 359 620 375
rect 710 394 776 397
rect 710 360 726 394
rect 760 360 776 394
rect 710 326 776 360
rect 710 323 726 326
rect 395 292 726 323
rect 760 292 776 326
rect 395 289 776 292
rect 108 235 174 239
rect 22 166 133 199
rect 22 132 83 166
rect 117 132 133 166
rect 22 99 133 132
rect 169 166 359 199
rect 169 132 239 166
rect 273 132 359 166
rect 169 113 359 132
rect 169 79 175 113
rect 209 79 247 113
rect 281 79 319 113
rect 353 79 359 113
rect 395 166 445 289
rect 812 253 846 433
rect 677 219 846 253
rect 882 335 948 503
rect 882 301 898 335
rect 932 301 948 335
rect 882 267 948 301
rect 882 233 898 267
rect 932 233 948 267
rect 882 219 948 233
rect 984 401 1018 579
rect 1307 541 1497 604
rect 1205 502 1271 535
rect 1307 507 1400 541
rect 1434 507 1497 541
rect 1540 735 1610 751
rect 1540 701 1556 735
rect 1590 701 1610 735
rect 1540 652 1610 701
rect 1540 618 1556 652
rect 1590 618 1610 652
rect 1540 568 1610 618
rect 1540 534 1556 568
rect 1590 534 1610 568
rect 1205 468 1221 502
rect 1255 471 1271 502
rect 1540 485 1610 534
rect 1255 468 1406 471
rect 1205 437 1406 468
rect 984 395 1336 401
rect 984 367 1286 395
rect 677 199 711 219
rect 429 132 445 166
rect 395 103 445 132
rect 481 166 599 195
rect 481 132 505 166
rect 539 132 599 166
rect 481 113 599 132
rect 169 73 359 79
rect 481 79 487 113
rect 521 79 559 113
rect 593 79 599 113
rect 645 166 711 199
rect 984 183 1018 367
rect 1270 361 1286 367
rect 1320 361 1336 395
rect 1270 355 1336 361
rect 1086 297 1102 331
rect 1136 319 1152 331
rect 1372 319 1406 437
rect 1136 297 1406 319
rect 1086 285 1406 297
rect 1540 451 1556 485
rect 1590 451 1610 485
rect 1086 263 1152 285
rect 1086 229 1102 263
rect 1136 229 1152 263
rect 1086 215 1152 229
rect 1209 232 1275 285
rect 645 132 661 166
rect 695 132 711 166
rect 645 99 711 132
rect 801 166 1018 183
rect 1209 198 1225 232
rect 1259 198 1275 232
rect 801 132 817 166
rect 851 149 1018 166
rect 1054 166 1172 179
rect 1209 169 1275 198
rect 1311 215 1404 249
rect 1438 215 1501 249
rect 851 132 867 149
rect 801 99 867 132
rect 1054 132 1115 166
rect 1149 132 1172 166
rect 1054 113 1172 132
rect 481 73 599 79
rect 1054 79 1060 113
rect 1094 79 1132 113
rect 1166 79 1172 113
rect 1054 73 1172 79
rect 1311 149 1501 215
rect 1311 115 1404 149
rect 1438 115 1501 149
rect 1311 113 1501 115
rect 1311 79 1317 113
rect 1351 79 1389 113
rect 1423 79 1461 113
rect 1495 79 1501 113
rect 1540 245 1610 451
rect 1540 211 1560 245
rect 1594 211 1610 245
rect 1540 153 1610 211
rect 1540 119 1560 153
rect 1594 119 1610 153
rect 1540 103 1610 119
rect 1311 73 1501 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 1087 797 1121 831
rect 1183 797 1217 831
rect 1279 797 1313 831
rect 1375 797 1409 831
rect 1471 797 1505 831
rect 1567 797 1601 831
rect 108 701 142 735
rect 180 701 214 735
rect 252 701 286 735
rect 384 701 418 735
rect 456 701 490 735
rect 528 725 562 735
rect 528 701 552 725
rect 552 701 562 725
rect 1060 701 1094 735
rect 1132 701 1166 735
rect 1204 701 1238 735
rect 1313 701 1347 735
rect 1385 701 1400 735
rect 1400 701 1419 735
rect 1457 701 1491 735
rect 175 79 209 113
rect 247 79 281 113
rect 319 79 353 113
rect 487 79 521 113
rect 559 79 593 113
rect 1060 79 1094 113
rect 1132 79 1166 113
rect 1317 79 1351 113
rect 1389 79 1423 113
rect 1461 79 1495 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
rect 1087 -17 1121 17
rect 1183 -17 1217 17
rect 1279 -17 1313 17
rect 1375 -17 1409 17
rect 1471 -17 1505 17
rect 1567 -17 1601 17
<< metal1 >>
rect 0 831 1632 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1087 831
rect 1121 797 1183 831
rect 1217 797 1279 831
rect 1313 797 1375 831
rect 1409 797 1471 831
rect 1505 797 1567 831
rect 1601 797 1632 831
rect 0 791 1632 797
rect 0 735 1632 763
rect 0 701 108 735
rect 142 701 180 735
rect 214 701 252 735
rect 286 701 384 735
rect 418 701 456 735
rect 490 701 528 735
rect 562 701 1060 735
rect 1094 701 1132 735
rect 1166 701 1204 735
rect 1238 701 1313 735
rect 1347 701 1385 735
rect 1419 701 1457 735
rect 1491 701 1632 735
rect 0 689 1632 701
rect 0 113 1632 125
rect 0 79 175 113
rect 209 79 247 113
rect 281 79 319 113
rect 353 79 487 113
rect 521 79 559 113
rect 593 79 1060 113
rect 1094 79 1132 113
rect 1166 79 1317 113
rect 1351 79 1389 113
rect 1423 79 1461 113
rect 1495 79 1632 113
rect 0 51 1632 79
rect 0 17 1632 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1087 17
rect 1121 -17 1183 17
rect 1217 -17 1279 17
rect 1313 -17 1375 17
rect 1409 -17 1471 17
rect 1505 -17 1567 17
rect 1601 -17 1632 17
rect 0 -23 1632 -17
<< labels >>
rlabel comment s 0 0 0 0 4 dlxtp_1
flabel metal1 s 0 51 1632 125 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel metal1 s 0 0 1632 23 0 FreeSans 340 0 0 0 VNB
port 4 nsew ground bidirectional
flabel metal1 s 0 689 1632 763 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 791 1632 814 0 FreeSans 340 0 0 0 VPB
port 5 nsew power bidirectional
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 D
port 1 nsew signal input
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 GATE
port 2 nsew clock input
flabel locali s 1567 316 1601 350 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
flabel locali s 1567 390 1601 424 0 FreeSans 340 0 0 0 Q
port 7 nsew signal output
rlabel locali s 481 73 599 195 1 VGND
port 3 nsew ground bidirectional
rlabel locali s 1054 73 1172 179 1 VGND
port 3 nsew ground bidirectional
rlabel locali s 1311 73 1501 249 1 VGND
port 3 nsew ground bidirectional
rlabel metal1 s 0 51 1632 125 1 VGND
port 3 nsew ground bidirectional
rlabel metal1 s 0 -23 1632 23 1 VNB
port 4 nsew ground bidirectional
rlabel metal1 s 0 791 1632 837 1 VPB
port 5 nsew power bidirectional
rlabel locali s 378 599 568 741 1 VPWR
port 6 nsew power bidirectional
rlabel locali s 1054 579 1244 741 1 VPWR
port 6 nsew power bidirectional
rlabel locali s 1307 507 1497 751 1 VPWR
port 6 nsew power bidirectional
rlabel metal1 s 0 689 1632 763 1 VPWR
port 6 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 1632 814
string GDS_END 1220156
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 1203716
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
<< end >>
