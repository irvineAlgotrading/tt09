magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect 0 0 294 408
<< pmos >>
rect 89 36 119 372
rect 175 36 205 372
<< pdiff >>
rect 36 329 89 372
rect 36 295 44 329
rect 78 295 89 329
rect 36 257 89 295
rect 36 223 44 257
rect 78 223 89 257
rect 36 185 89 223
rect 36 151 44 185
rect 78 151 89 185
rect 36 113 89 151
rect 36 79 44 113
rect 78 79 89 113
rect 36 36 89 79
rect 119 329 175 372
rect 119 295 130 329
rect 164 295 175 329
rect 119 257 175 295
rect 119 223 130 257
rect 164 223 175 257
rect 119 185 175 223
rect 119 151 130 185
rect 164 151 175 185
rect 119 113 175 151
rect 119 79 130 113
rect 164 79 175 113
rect 119 36 175 79
rect 205 329 258 372
rect 205 295 216 329
rect 250 295 258 329
rect 205 257 258 295
rect 205 223 216 257
rect 250 223 258 257
rect 205 185 258 223
rect 205 151 216 185
rect 250 151 258 185
rect 205 113 258 151
rect 205 79 216 113
rect 250 79 258 113
rect 205 36 258 79
<< pdiffc >>
rect 44 295 78 329
rect 44 223 78 257
rect 44 151 78 185
rect 44 79 78 113
rect 130 295 164 329
rect 130 223 164 257
rect 130 151 164 185
rect 130 79 164 113
rect 216 295 250 329
rect 216 223 250 257
rect 216 151 250 185
rect 216 79 250 113
<< poly >>
rect 80 459 214 475
rect 80 425 96 459
rect 130 425 164 459
rect 198 425 214 459
rect 80 409 214 425
rect 89 398 205 409
rect 89 372 119 398
rect 175 372 205 398
rect 89 10 119 36
rect 175 10 205 36
<< polycont >>
rect 96 425 130 459
rect 164 425 198 459
<< locali >>
rect 80 459 214 475
rect 80 425 94 459
rect 130 425 164 459
rect 200 425 214 459
rect 80 409 214 425
rect 44 329 78 370
rect 44 257 78 295
rect 44 185 78 223
rect 44 113 78 151
rect 44 36 78 79
rect 130 329 164 370
rect 130 257 164 295
rect 130 185 164 223
rect 130 113 164 151
rect 130 36 164 79
rect 216 329 250 370
rect 216 257 250 295
rect 216 185 250 223
rect 216 113 250 151
rect 216 36 250 79
<< viali >>
rect 94 425 96 459
rect 96 425 128 459
rect 166 425 198 459
rect 198 425 200 459
rect 44 295 78 329
rect 44 223 78 257
rect 44 151 78 185
rect 44 79 78 113
rect 130 295 164 329
rect 130 223 164 257
rect 130 151 164 185
rect 130 79 164 113
rect 216 295 250 329
rect 216 223 250 257
rect 216 151 250 185
rect 216 79 250 113
<< metal1 >>
rect 82 459 212 471
rect 82 425 94 459
rect 128 425 166 459
rect 200 425 212 459
rect 82 413 212 425
rect 38 329 84 370
rect 38 295 44 329
rect 78 295 84 329
rect 38 257 84 295
rect 38 223 44 257
rect 78 223 84 257
rect 38 185 84 223
rect 38 151 44 185
rect 78 151 84 185
rect 38 113 84 151
rect 38 79 44 113
rect 78 79 84 113
rect 38 -29 84 79
rect 121 363 173 370
rect 121 299 130 311
rect 164 299 173 311
rect 121 223 130 247
rect 164 223 173 247
rect 121 185 173 223
rect 121 151 130 185
rect 164 151 173 185
rect 121 113 173 151
rect 121 79 130 113
rect 164 79 173 113
rect 121 36 173 79
rect 210 329 256 370
rect 210 295 216 329
rect 250 295 256 329
rect 210 257 256 295
rect 210 223 216 257
rect 250 223 256 257
rect 210 185 256 223
rect 210 151 216 185
rect 250 151 256 185
rect 210 113 256 151
rect 210 79 216 113
rect 250 79 256 113
rect 210 -29 256 79
rect 38 -89 256 -29
<< via1 >>
rect 121 329 173 363
rect 121 311 130 329
rect 130 311 164 329
rect 164 311 173 329
rect 121 295 130 299
rect 130 295 164 299
rect 164 295 173 299
rect 121 257 173 295
rect 121 247 130 257
rect 130 247 164 257
rect 164 247 173 257
<< metal2 >>
rect 121 363 173 369
rect 121 299 173 311
rect 121 241 173 247
<< labels >>
flabel metal2 s 121 241 173 369 0 FreeSans 400 0 0 0 DRAIN
port 1 nsew
flabel metal1 s 38 -89 256 -29 0 FreeSans 400 0 0 0 SOURCE
port 3 nsew
flabel metal1 s 82 413 212 471 0 FreeSans 400 0 0 0 GATE
port 2 nsew
flabel nwell s 74 399 81 405 0 FreeSans 400 0 0 0 BULK
port 4 nsew
<< properties >>
string GDS_END 10482564
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 10477520
string path 0.950 -1.475 6.400 -1.475 
string device primitive
<< end >>
