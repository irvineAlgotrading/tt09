magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect 8827 2833 9559 2999
rect -181 1296 1108 1462
rect 2297 1422 3774 1527
rect 2297 1421 4153 1422
rect -181 -128 -15 1296
rect 935 1128 1108 1296
rect 935 962 2205 1128
rect 979 -128 1002 962
rect 3708 721 4153 1421
rect -181 -187 1681 -128
rect 2192 -132 2358 358
rect 2192 -134 2380 -132
rect 2192 -146 2358 -134
rect -167 -975 1681 -187
rect 1458 -978 1466 -975
<< pwell >>
rect 5989 1512 6149 1516
rect 5989 1426 10151 1512
rect 5989 1242 6296 1426
rect 4994 1156 6296 1242
rect 4994 1068 5080 1156
rect 2567 -3 3761 83
rect 4236 -48 4322 934
rect 5011 -88 8147 -2
rect 10065 -20 10151 1426
<< ndiff >>
rect 6051 1290 6123 1490
<< mvndiff >>
rect 6041 1290 6051 1490
<< psubdiff >>
rect 4262 884 4296 908
rect 4262 814 4296 850
rect 4262 744 4296 780
rect 4262 674 4296 710
rect 4262 604 4296 640
rect 4262 533 4296 570
rect 4262 462 4296 499
rect 4262 391 4296 428
rect 4262 320 4296 357
rect 4262 249 4296 286
rect 4262 178 4296 215
rect 4262 107 4296 144
rect 2593 23 2657 57
rect 2691 23 2725 57
rect 2759 23 2793 57
rect 2827 23 2861 57
rect 2895 23 2929 57
rect 2963 23 2997 57
rect 3031 23 3065 57
rect 3099 23 3133 57
rect 3167 23 3201 57
rect 3235 23 3269 57
rect 3303 23 3337 57
rect 3371 23 3405 57
rect 3439 23 3473 57
rect 3507 23 3541 57
rect 3575 23 3609 57
rect 3643 23 3677 57
rect 3711 23 3735 57
rect 4262 36 4296 73
rect 4262 -22 4296 2
<< nsubdiff >>
rect 2333 1457 2357 1491
rect 2391 1457 2425 1491
rect 2459 1457 2493 1491
rect 2527 1457 2561 1491
rect 2595 1457 2629 1491
rect 2663 1457 2697 1491
rect 2731 1457 2765 1491
rect 2799 1457 2833 1491
rect 2867 1457 2901 1491
rect 2935 1457 2969 1491
rect 3003 1457 3037 1491
rect 3071 1457 3105 1491
rect 3139 1457 3173 1491
rect 3207 1457 3241 1491
rect 3275 1457 3309 1491
rect 3343 1457 3377 1491
rect 3411 1457 3445 1491
rect 3479 1457 3513 1491
rect 3547 1457 3581 1491
rect 3615 1457 3649 1491
rect 3683 1457 3738 1491
<< mvpsubdiff >>
rect 6236 1452 6304 1486
rect 6338 1452 6372 1486
rect 6406 1452 6440 1486
rect 6474 1452 6508 1486
rect 6542 1452 6576 1486
rect 6610 1452 6644 1486
rect 6678 1452 6712 1486
rect 6746 1452 6780 1486
rect 6814 1452 6848 1486
rect 6882 1452 6916 1486
rect 6950 1452 6984 1486
rect 7018 1452 7052 1486
rect 7086 1452 7120 1486
rect 7154 1452 7188 1486
rect 7222 1452 7256 1486
rect 7290 1452 7324 1486
rect 7358 1452 7392 1486
rect 7426 1452 7460 1486
rect 7494 1452 7528 1486
rect 7562 1452 7596 1486
rect 7630 1452 7664 1486
rect 7698 1452 7732 1486
rect 7766 1452 7800 1486
rect 7834 1452 7868 1486
rect 7902 1452 7936 1486
rect 7970 1452 8004 1486
rect 8038 1452 8072 1486
rect 8106 1452 8140 1486
rect 8174 1452 8208 1486
rect 8242 1452 8276 1486
rect 8310 1452 8344 1486
rect 8378 1452 8412 1486
rect 8446 1452 8480 1486
rect 8514 1452 8548 1486
rect 8582 1452 8616 1486
rect 8650 1452 8684 1486
rect 8718 1452 8752 1486
rect 8786 1452 8820 1486
rect 8854 1452 8888 1486
rect 8922 1452 8956 1486
rect 8990 1452 9024 1486
rect 9058 1452 9092 1486
rect 9126 1452 9160 1486
rect 9194 1452 9228 1486
rect 9262 1452 9296 1486
rect 9330 1452 9364 1486
rect 9398 1452 9432 1486
rect 9466 1452 9500 1486
rect 9534 1452 9568 1486
rect 9602 1452 9636 1486
rect 9670 1452 9704 1486
rect 9738 1452 9772 1486
rect 9806 1452 9840 1486
rect 9874 1452 9908 1486
rect 9942 1452 9976 1486
rect 10010 1452 10125 1486
rect 6236 1352 6270 1452
rect 6236 1284 6270 1318
rect 6236 1216 6270 1250
rect 5020 1182 5159 1216
rect 5193 1182 5227 1216
rect 5261 1182 5295 1216
rect 5329 1182 5363 1216
rect 5397 1182 5431 1216
rect 5465 1182 5499 1216
rect 5533 1182 5567 1216
rect 5601 1182 5635 1216
rect 5669 1182 5703 1216
rect 5737 1182 5771 1216
rect 5805 1182 5839 1216
rect 5873 1182 5907 1216
rect 5941 1182 5975 1216
rect 6009 1182 6043 1216
rect 6077 1182 6165 1216
rect 6199 1182 6270 1216
rect 10091 1418 10125 1452
rect 10091 1350 10125 1384
rect 10091 1282 10125 1316
rect 10091 1214 10125 1248
rect 5020 1094 5054 1182
rect 10091 1146 10125 1180
rect 10091 1078 10125 1112
rect 10091 1010 10125 1044
rect 10091 942 10125 976
rect 10091 874 10125 908
rect 10091 806 10125 840
rect 10091 738 10125 772
rect 10091 670 10125 704
rect 10091 602 10125 636
rect 10091 534 10125 568
rect 10091 466 10125 500
rect 10091 398 10125 432
rect 10091 330 10125 364
rect 10091 262 10125 296
rect 10091 194 10125 228
rect 10091 126 10125 160
rect 10091 6 10125 92
rect 5037 -62 5071 -28
rect 5105 -62 5139 -28
rect 5173 -62 5207 -28
rect 5241 -62 5275 -28
rect 5309 -62 5343 -28
rect 5377 -62 5411 -28
rect 5445 -62 5479 -28
rect 5513 -62 5547 -28
rect 5581 -62 5615 -28
rect 5649 -62 5683 -28
rect 5717 -62 5751 -28
rect 5785 -62 5819 -28
rect 5853 -62 5887 -28
rect 5921 -62 5955 -28
rect 5989 -62 6023 -28
rect 6057 -62 6091 -28
rect 6125 -62 6159 -28
rect 6193 -62 6285 -28
rect 6319 -62 6353 -28
rect 6387 -62 6421 -28
rect 6455 -62 6489 -28
rect 6523 -62 6557 -28
rect 6591 -62 6625 -28
rect 6659 -62 6693 -28
rect 6727 -62 6761 -28
rect 6795 -62 6829 -28
rect 6863 -62 6897 -28
rect 6931 -62 6965 -28
rect 6999 -62 7033 -28
rect 7067 -62 7101 -28
rect 7135 -62 7169 -28
rect 7203 -62 7237 -28
rect 7271 -62 7305 -28
rect 7339 -62 7373 -28
rect 7407 -62 7441 -28
rect 7475 -62 7509 -28
rect 7543 -62 7577 -28
rect 7611 -62 7645 -28
rect 7679 -62 7713 -28
rect 7747 -62 7781 -28
rect 7815 -62 7849 -28
rect 7883 -62 7917 -28
rect 7951 -62 7985 -28
rect 8019 -62 8053 -28
rect 8087 -62 8121 -28
<< mvnsubdiff >>
rect 8893 2899 8917 2933
rect 8951 2899 8991 2933
rect 9025 2899 9065 2933
rect 9099 2899 9139 2933
rect 9173 2899 9213 2933
rect 9247 2899 9287 2933
rect 9321 2899 9361 2933
rect 9395 2899 9435 2933
rect 9469 2899 9493 2933
rect -115 1362 -47 1396
rect -13 1362 22 1396
rect 56 1362 91 1396
rect 125 1362 160 1396
rect 194 1362 229 1396
rect 263 1362 298 1396
rect 332 1362 367 1396
rect 401 1362 436 1396
rect 470 1362 504 1396
rect 538 1362 572 1396
rect 606 1362 640 1396
rect 674 1362 708 1396
rect 742 1362 776 1396
rect 810 1362 858 1396
rect 892 1362 930 1396
rect 964 1362 1035 1396
rect -115 1327 -81 1362
rect -115 1258 -81 1293
rect -115 1189 -81 1224
rect -115 1120 -81 1155
rect -115 1051 -81 1086
rect 1001 1328 1035 1362
rect 1001 1239 1035 1294
rect 1001 1150 1035 1205
rect 1001 1062 1035 1116
rect 1001 1028 1069 1062
rect 1103 1028 1142 1062
rect 1176 1028 1215 1062
rect 1249 1028 1288 1062
rect 1322 1028 1361 1062
rect 1395 1028 1433 1062
rect 1467 1028 1505 1062
rect 1539 1028 1577 1062
rect 1611 1028 1649 1062
rect 1683 1028 1721 1062
rect 1755 1028 1793 1062
rect 1827 1028 1865 1062
rect 1899 1028 1937 1062
rect 1971 1028 2009 1062
rect 2043 1028 2081 1062
rect 2115 1028 2139 1062
rect -115 982 -81 1017
rect -115 913 -81 948
rect -115 844 -81 879
rect -115 775 -81 810
rect -115 706 -81 741
rect -115 637 -81 672
rect -115 567 -81 603
rect -115 497 -81 533
rect -115 427 -81 463
rect -115 357 -81 393
rect -115 287 -81 323
rect -115 217 -81 253
rect -115 147 -81 183
rect -115 77 -81 113
rect -115 7 -81 43
rect -115 -63 -81 -27
rect 2258 268 2292 292
rect 2258 196 2292 234
rect 2258 124 2292 162
rect 2258 51 2292 90
rect 2258 -22 2292 17
rect 2258 -80 2292 -56
rect -115 -121 -81 -97
<< psubdiffcont >>
rect 4262 850 4296 884
rect 4262 780 4296 814
rect 4262 710 4296 744
rect 4262 640 4296 674
rect 4262 570 4296 604
rect 4262 499 4296 533
rect 4262 428 4296 462
rect 4262 357 4296 391
rect 4262 286 4296 320
rect 4262 215 4296 249
rect 4262 144 4296 178
rect 4262 73 4296 107
rect 2657 23 2691 57
rect 2725 23 2759 57
rect 2793 23 2827 57
rect 2861 23 2895 57
rect 2929 23 2963 57
rect 2997 23 3031 57
rect 3065 23 3099 57
rect 3133 23 3167 57
rect 3201 23 3235 57
rect 3269 23 3303 57
rect 3337 23 3371 57
rect 3405 23 3439 57
rect 3473 23 3507 57
rect 3541 23 3575 57
rect 3609 23 3643 57
rect 3677 23 3711 57
rect 4262 2 4296 36
<< nsubdiffcont >>
rect 2357 1457 2391 1491
rect 2425 1457 2459 1491
rect 2493 1457 2527 1491
rect 2561 1457 2595 1491
rect 2629 1457 2663 1491
rect 2697 1457 2731 1491
rect 2765 1457 2799 1491
rect 2833 1457 2867 1491
rect 2901 1457 2935 1491
rect 2969 1457 3003 1491
rect 3037 1457 3071 1491
rect 3105 1457 3139 1491
rect 3173 1457 3207 1491
rect 3241 1457 3275 1491
rect 3309 1457 3343 1491
rect 3377 1457 3411 1491
rect 3445 1457 3479 1491
rect 3513 1457 3547 1491
rect 3581 1457 3615 1491
rect 3649 1457 3683 1491
<< mvpsubdiffcont >>
rect 6304 1452 6338 1486
rect 6372 1452 6406 1486
rect 6440 1452 6474 1486
rect 6508 1452 6542 1486
rect 6576 1452 6610 1486
rect 6644 1452 6678 1486
rect 6712 1452 6746 1486
rect 6780 1452 6814 1486
rect 6848 1452 6882 1486
rect 6916 1452 6950 1486
rect 6984 1452 7018 1486
rect 7052 1452 7086 1486
rect 7120 1452 7154 1486
rect 7188 1452 7222 1486
rect 7256 1452 7290 1486
rect 7324 1452 7358 1486
rect 7392 1452 7426 1486
rect 7460 1452 7494 1486
rect 7528 1452 7562 1486
rect 7596 1452 7630 1486
rect 7664 1452 7698 1486
rect 7732 1452 7766 1486
rect 7800 1452 7834 1486
rect 7868 1452 7902 1486
rect 7936 1452 7970 1486
rect 8004 1452 8038 1486
rect 8072 1452 8106 1486
rect 8140 1452 8174 1486
rect 8208 1452 8242 1486
rect 8276 1452 8310 1486
rect 8344 1452 8378 1486
rect 8412 1452 8446 1486
rect 8480 1452 8514 1486
rect 8548 1452 8582 1486
rect 8616 1452 8650 1486
rect 8684 1452 8718 1486
rect 8752 1452 8786 1486
rect 8820 1452 8854 1486
rect 8888 1452 8922 1486
rect 8956 1452 8990 1486
rect 9024 1452 9058 1486
rect 9092 1452 9126 1486
rect 9160 1452 9194 1486
rect 9228 1452 9262 1486
rect 9296 1452 9330 1486
rect 9364 1452 9398 1486
rect 9432 1452 9466 1486
rect 9500 1452 9534 1486
rect 9568 1452 9602 1486
rect 9636 1452 9670 1486
rect 9704 1452 9738 1486
rect 9772 1452 9806 1486
rect 9840 1452 9874 1486
rect 9908 1452 9942 1486
rect 9976 1452 10010 1486
rect 6236 1318 6270 1352
rect 6236 1250 6270 1284
rect 5159 1182 5193 1216
rect 5227 1182 5261 1216
rect 5295 1182 5329 1216
rect 5363 1182 5397 1216
rect 5431 1182 5465 1216
rect 5499 1182 5533 1216
rect 5567 1182 5601 1216
rect 5635 1182 5669 1216
rect 5703 1182 5737 1216
rect 5771 1182 5805 1216
rect 5839 1182 5873 1216
rect 5907 1182 5941 1216
rect 5975 1182 6009 1216
rect 6043 1182 6077 1216
rect 6165 1182 6199 1216
rect 10091 1384 10125 1418
rect 10091 1316 10125 1350
rect 10091 1248 10125 1282
rect 10091 1180 10125 1214
rect 10091 1112 10125 1146
rect 10091 1044 10125 1078
rect 10091 976 10125 1010
rect 10091 908 10125 942
rect 10091 840 10125 874
rect 10091 772 10125 806
rect 10091 704 10125 738
rect 10091 636 10125 670
rect 10091 568 10125 602
rect 10091 500 10125 534
rect 10091 432 10125 466
rect 10091 364 10125 398
rect 10091 296 10125 330
rect 10091 228 10125 262
rect 10091 160 10125 194
rect 10091 92 10125 126
rect 5071 -62 5105 -28
rect 5139 -62 5173 -28
rect 5207 -62 5241 -28
rect 5275 -62 5309 -28
rect 5343 -62 5377 -28
rect 5411 -62 5445 -28
rect 5479 -62 5513 -28
rect 5547 -62 5581 -28
rect 5615 -62 5649 -28
rect 5683 -62 5717 -28
rect 5751 -62 5785 -28
rect 5819 -62 5853 -28
rect 5887 -62 5921 -28
rect 5955 -62 5989 -28
rect 6023 -62 6057 -28
rect 6091 -62 6125 -28
rect 6159 -62 6193 -28
rect 6285 -62 6319 -28
rect 6353 -62 6387 -28
rect 6421 -62 6455 -28
rect 6489 -62 6523 -28
rect 6557 -62 6591 -28
rect 6625 -62 6659 -28
rect 6693 -62 6727 -28
rect 6761 -62 6795 -28
rect 6829 -62 6863 -28
rect 6897 -62 6931 -28
rect 6965 -62 6999 -28
rect 7033 -62 7067 -28
rect 7101 -62 7135 -28
rect 7169 -62 7203 -28
rect 7237 -62 7271 -28
rect 7305 -62 7339 -28
rect 7373 -62 7407 -28
rect 7441 -62 7475 -28
rect 7509 -62 7543 -28
rect 7577 -62 7611 -28
rect 7645 -62 7679 -28
rect 7713 -62 7747 -28
rect 7781 -62 7815 -28
rect 7849 -62 7883 -28
rect 7917 -62 7951 -28
rect 7985 -62 8019 -28
rect 8053 -62 8087 -28
<< mvnsubdiffcont >>
rect 8917 2899 8951 2933
rect 8991 2899 9025 2933
rect 9065 2899 9099 2933
rect 9139 2899 9173 2933
rect 9213 2899 9247 2933
rect 9287 2899 9321 2933
rect 9361 2899 9395 2933
rect 9435 2899 9469 2933
rect -47 1362 -13 1396
rect 22 1362 56 1396
rect 91 1362 125 1396
rect 160 1362 194 1396
rect 229 1362 263 1396
rect 298 1362 332 1396
rect 367 1362 401 1396
rect 436 1362 470 1396
rect 504 1362 538 1396
rect 572 1362 606 1396
rect 640 1362 674 1396
rect 708 1362 742 1396
rect 776 1362 810 1396
rect 858 1362 892 1396
rect 930 1362 964 1396
rect -115 1293 -81 1327
rect -115 1224 -81 1258
rect -115 1155 -81 1189
rect -115 1086 -81 1120
rect -115 1017 -81 1051
rect 1001 1294 1035 1328
rect 1001 1205 1035 1239
rect 1001 1116 1035 1150
rect 1069 1028 1103 1062
rect 1142 1028 1176 1062
rect 1215 1028 1249 1062
rect 1288 1028 1322 1062
rect 1361 1028 1395 1062
rect 1433 1028 1467 1062
rect 1505 1028 1539 1062
rect 1577 1028 1611 1062
rect 1649 1028 1683 1062
rect 1721 1028 1755 1062
rect 1793 1028 1827 1062
rect 1865 1028 1899 1062
rect 1937 1028 1971 1062
rect 2009 1028 2043 1062
rect 2081 1028 2115 1062
rect -115 948 -81 982
rect -115 879 -81 913
rect -115 810 -81 844
rect -115 741 -81 775
rect -115 672 -81 706
rect -115 603 -81 637
rect -115 533 -81 567
rect -115 463 -81 497
rect -115 393 -81 427
rect -115 323 -81 357
rect -115 253 -81 287
rect -115 183 -81 217
rect -115 113 -81 147
rect -115 43 -81 77
rect -115 -27 -81 7
rect -115 -97 -81 -63
rect 2258 234 2292 268
rect 2258 162 2292 196
rect 2258 90 2292 124
rect 2258 17 2292 51
rect 2258 -56 2292 -22
<< poly >>
rect 8795 2677 8861 2743
rect 8795 2643 8811 2677
rect 8845 2643 8861 2677
rect 8795 2609 8861 2643
rect 8795 2575 8811 2609
rect 8845 2575 8861 2609
rect 8795 2541 8861 2575
rect 8795 2507 8811 2541
rect 8845 2507 8861 2541
rect 8795 2487 8861 2507
rect 8790 2152 8856 2168
rect 8790 2118 8806 2152
rect 8840 2118 8856 2152
rect 8790 2018 8856 2118
rect 8790 1984 8806 2018
rect 8840 1984 8856 2018
rect 8790 1968 8856 1984
rect 4835 1572 5723 1588
rect 1075 1551 1141 1567
rect 1075 1517 1091 1551
rect 1125 1517 1141 1551
rect 1075 1474 1141 1517
rect 4264 1537 4520 1553
rect 4264 1503 4280 1537
rect 4314 1503 4375 1537
rect 4409 1503 4470 1537
rect 4504 1503 4520 1537
rect 4835 1538 4851 1572
rect 4885 1538 4920 1572
rect 4954 1538 4989 1572
rect 5023 1538 5058 1572
rect 5092 1538 5127 1572
rect 5161 1538 5196 1572
rect 5230 1538 5265 1572
rect 5299 1538 5333 1572
rect 5367 1538 5401 1572
rect 5435 1538 5469 1572
rect 5503 1538 5537 1572
rect 5571 1538 5605 1572
rect 5639 1538 5673 1572
rect 5707 1538 5723 1572
rect 4835 1522 5723 1538
rect 5779 1572 5959 1588
rect 5779 1538 5795 1572
rect 5829 1538 5909 1572
rect 5943 1538 5959 1572
rect 5779 1522 5959 1538
rect 1075 1440 1091 1474
rect 1125 1440 1141 1474
rect 4264 1487 4520 1503
rect 1075 1397 1141 1440
rect 1075 1363 1091 1397
rect 1125 1363 1141 1397
rect 1075 1319 1141 1363
rect 1075 1285 1091 1319
rect 1125 1285 1141 1319
rect 1075 1241 1141 1285
rect 1075 1207 1091 1241
rect 1125 1207 1141 1241
rect 1075 1191 1141 1207
rect 5188 1128 6112 1144
rect 5188 1094 5208 1128
rect 5242 1094 5276 1128
rect 5310 1094 5344 1128
rect 5378 1094 5412 1128
rect 5446 1094 5480 1128
rect 5514 1094 5548 1128
rect 5582 1094 5616 1128
rect 5650 1094 5684 1128
rect 5718 1094 5752 1128
rect 5786 1094 5820 1128
rect 5854 1094 5888 1128
rect 5922 1094 6112 1128
rect 5188 1078 6112 1094
rect 5969 1074 6112 1078
rect 3868 1014 3988 1030
rect 2366 731 2466 751
rect 2522 731 2622 751
rect 2366 715 2620 731
rect 2366 681 2382 715
rect 2416 681 2476 715
rect 2510 681 2570 715
rect 2604 681 2620 715
rect 2366 665 2620 681
rect 2802 630 2902 751
rect 2646 602 2902 630
rect 2646 568 2662 602
rect 2696 568 2757 602
rect 2791 568 2852 602
rect 2886 568 2902 602
rect 2646 518 2902 568
rect 2646 484 2662 518
rect 2696 484 2757 518
rect 2791 484 2852 518
rect 2886 484 2902 518
rect 2646 364 2902 484
rect 2958 642 3058 751
rect 3114 642 3214 751
rect 2958 602 3214 642
rect 2958 568 2974 602
rect 3008 568 3069 602
rect 3103 568 3164 602
rect 3198 568 3214 602
rect 2958 518 3214 568
rect 2958 484 2974 518
rect 3008 484 3069 518
rect 3103 484 3164 518
rect 3198 484 3214 518
rect 2958 458 3214 484
rect 2958 364 3058 458
rect 3114 364 3214 458
rect 3270 634 3370 751
rect 3426 634 3526 751
rect 3582 634 3682 751
rect 3270 602 3682 634
rect 3270 568 3286 602
rect 3320 568 3364 602
rect 3398 568 3442 602
rect 3476 568 3519 602
rect 3553 568 3596 602
rect 3630 568 3682 602
rect 3270 518 3682 568
rect 3270 484 3286 518
rect 3320 484 3364 518
rect 3398 484 3442 518
rect 3476 484 3519 518
rect 3553 484 3596 518
rect 3630 484 3682 518
rect 3270 433 3682 484
rect 3270 364 3370 433
rect 3426 364 3526 433
rect 3582 364 3682 433
rect 3868 725 3988 802
rect 3868 691 3913 725
rect 3947 691 3988 725
rect 3868 641 3988 691
rect 3868 607 3913 641
rect 3947 607 3988 641
rect 3868 557 3988 607
rect 3868 523 3913 557
rect 3947 523 3988 557
rect 3868 473 3988 523
rect 3868 439 3913 473
rect 3947 439 3988 473
rect 3868 389 3988 439
rect 3868 355 3913 389
rect 3947 355 3988 389
rect 3868 306 3988 355
rect 6400 728 8904 744
rect 6400 694 6416 728
rect 6450 694 6485 728
rect 6519 694 6554 728
rect 6588 694 6623 728
rect 6657 694 6692 728
rect 6726 694 6761 728
rect 6795 694 6830 728
rect 6864 694 6899 728
rect 6933 694 6968 728
rect 7002 694 7037 728
rect 7071 694 7106 728
rect 7140 694 7175 728
rect 7209 694 7244 728
rect 7278 694 7314 728
rect 7348 694 7384 728
rect 7418 694 7454 728
rect 7488 694 7524 728
rect 7558 694 7594 728
rect 7628 694 7664 728
rect 7698 694 7734 728
rect 7768 694 7804 728
rect 7838 694 7874 728
rect 7908 694 7944 728
rect 7978 694 8014 728
rect 8048 694 8084 728
rect 8118 694 8154 728
rect 8188 694 8224 728
rect 8258 694 8294 728
rect 8328 694 8364 728
rect 8398 694 8434 728
rect 8468 694 8504 728
rect 8538 694 8574 728
rect 8608 694 8644 728
rect 8678 694 8714 728
rect 8748 694 8784 728
rect 8818 694 8854 728
rect 8888 694 8904 728
rect 6400 678 8904 694
rect 8960 728 9960 744
rect 8960 694 8976 728
rect 9010 694 9047 728
rect 9081 694 9118 728
rect 9152 694 9190 728
rect 9224 694 9262 728
rect 9296 694 9334 728
rect 9368 694 9406 728
rect 9440 694 9478 728
rect 9512 694 9550 728
rect 9584 694 9622 728
rect 9656 694 9694 728
rect 9728 694 9766 728
rect 9800 694 9838 728
rect 9872 694 9910 728
rect 9944 694 9960 728
rect 8960 678 9960 694
rect 4434 363 4734 364
rect 4426 362 4865 363
rect 4426 347 4890 362
rect 4426 313 4532 347
rect 4566 313 4811 347
rect 4845 313 4890 347
rect 4426 307 4890 313
rect 4426 257 4626 307
rect 4730 297 4865 307
rect 4698 27 4898 43
rect 4698 -7 4746 27
rect 4780 -7 4816 27
rect 4850 -7 4898 27
rect 1124 -128 2128 -112
rect 4698 -117 4898 -7
rect 49 -152 857 -144
rect 68 -168 857 -152
rect 68 -202 88 -168
rect 122 -202 156 -168
rect 190 -202 224 -168
rect 258 -202 292 -168
rect 326 -202 360 -168
rect 394 -202 428 -168
rect 462 -202 496 -168
rect 530 -202 564 -168
rect 598 -202 632 -168
rect 666 -202 700 -168
rect 734 -202 768 -168
rect 802 -202 857 -168
rect 1124 -162 1190 -128
rect 1224 -162 1258 -128
rect 1292 -162 1326 -128
rect 1360 -162 1394 -128
rect 1428 -162 1462 -128
rect 1496 -162 1530 -128
rect 1564 -162 1598 -128
rect 1632 -162 1666 -128
rect 1700 -162 1734 -128
rect 1768 -162 1802 -128
rect 1836 -162 1870 -128
rect 1904 -162 1938 -128
rect 1972 -162 2006 -128
rect 2040 -162 2074 -128
rect 2108 -162 2128 -128
rect 1124 -178 2128 -162
rect 68 -218 857 -202
rect 1144 -475 1210 -459
rect 1144 -509 1160 -475
rect 1194 -509 1210 -475
rect 1144 -559 1210 -509
rect 1144 -593 1160 -559
rect 1194 -593 1210 -559
rect 675 -658 741 -642
rect 675 -692 691 -658
rect 725 -692 741 -658
rect 675 -792 741 -692
rect 675 -826 691 -792
rect 725 -826 741 -792
rect 675 -842 741 -826
rect 1144 -643 1210 -593
rect 1144 -677 1160 -643
rect 1194 -677 1210 -643
rect 1144 -726 1210 -677
rect 1144 -760 1160 -726
rect 1194 -760 1210 -726
rect 1144 -809 1210 -760
rect 1144 -843 1160 -809
rect 1194 -843 1210 -809
rect 1144 -859 1210 -843
<< polycont >>
rect 8811 2643 8845 2677
rect 8811 2575 8845 2609
rect 8811 2507 8845 2541
rect 8806 2118 8840 2152
rect 8806 1984 8840 2018
rect 1091 1517 1125 1551
rect 4280 1503 4314 1537
rect 4375 1503 4409 1537
rect 4470 1503 4504 1537
rect 4851 1538 4885 1572
rect 4920 1538 4954 1572
rect 4989 1538 5023 1572
rect 5058 1538 5092 1572
rect 5127 1538 5161 1572
rect 5196 1538 5230 1572
rect 5265 1538 5299 1572
rect 5333 1538 5367 1572
rect 5401 1538 5435 1572
rect 5469 1538 5503 1572
rect 5537 1538 5571 1572
rect 5605 1538 5639 1572
rect 5673 1538 5707 1572
rect 5795 1538 5829 1572
rect 5909 1538 5943 1572
rect 1091 1440 1125 1474
rect 1091 1363 1125 1397
rect 1091 1285 1125 1319
rect 1091 1207 1125 1241
rect 5208 1094 5242 1128
rect 5276 1094 5310 1128
rect 5344 1094 5378 1128
rect 5412 1094 5446 1128
rect 5480 1094 5514 1128
rect 5548 1094 5582 1128
rect 5616 1094 5650 1128
rect 5684 1094 5718 1128
rect 5752 1094 5786 1128
rect 5820 1094 5854 1128
rect 5888 1094 5922 1128
rect 2382 681 2416 715
rect 2476 681 2510 715
rect 2570 681 2604 715
rect 2662 568 2696 602
rect 2757 568 2791 602
rect 2852 568 2886 602
rect 2662 484 2696 518
rect 2757 484 2791 518
rect 2852 484 2886 518
rect 2974 568 3008 602
rect 3069 568 3103 602
rect 3164 568 3198 602
rect 2974 484 3008 518
rect 3069 484 3103 518
rect 3164 484 3198 518
rect 3286 568 3320 602
rect 3364 568 3398 602
rect 3442 568 3476 602
rect 3519 568 3553 602
rect 3596 568 3630 602
rect 3286 484 3320 518
rect 3364 484 3398 518
rect 3442 484 3476 518
rect 3519 484 3553 518
rect 3596 484 3630 518
rect 3913 691 3947 725
rect 3913 607 3947 641
rect 3913 523 3947 557
rect 3913 439 3947 473
rect 3913 355 3947 389
rect 6416 694 6450 728
rect 6485 694 6519 728
rect 6554 694 6588 728
rect 6623 694 6657 728
rect 6692 694 6726 728
rect 6761 694 6795 728
rect 6830 694 6864 728
rect 6899 694 6933 728
rect 6968 694 7002 728
rect 7037 694 7071 728
rect 7106 694 7140 728
rect 7175 694 7209 728
rect 7244 694 7278 728
rect 7314 694 7348 728
rect 7384 694 7418 728
rect 7454 694 7488 728
rect 7524 694 7558 728
rect 7594 694 7628 728
rect 7664 694 7698 728
rect 7734 694 7768 728
rect 7804 694 7838 728
rect 7874 694 7908 728
rect 7944 694 7978 728
rect 8014 694 8048 728
rect 8084 694 8118 728
rect 8154 694 8188 728
rect 8224 694 8258 728
rect 8294 694 8328 728
rect 8364 694 8398 728
rect 8434 694 8468 728
rect 8504 694 8538 728
rect 8574 694 8608 728
rect 8644 694 8678 728
rect 8714 694 8748 728
rect 8784 694 8818 728
rect 8854 694 8888 728
rect 8976 694 9010 728
rect 9047 694 9081 728
rect 9118 694 9152 728
rect 9190 694 9224 728
rect 9262 694 9296 728
rect 9334 694 9368 728
rect 9406 694 9440 728
rect 9478 694 9512 728
rect 9550 694 9584 728
rect 9622 694 9656 728
rect 9694 694 9728 728
rect 9766 694 9800 728
rect 9838 694 9872 728
rect 9910 694 9944 728
rect 4532 313 4566 347
rect 4811 313 4845 347
rect 4746 -7 4780 27
rect 4816 -7 4850 27
rect 88 -202 122 -168
rect 156 -202 190 -168
rect 224 -202 258 -168
rect 292 -202 326 -168
rect 360 -202 394 -168
rect 428 -202 462 -168
rect 496 -202 530 -168
rect 564 -202 598 -168
rect 632 -202 666 -168
rect 700 -202 734 -168
rect 768 -202 802 -168
rect 1190 -162 1224 -128
rect 1258 -162 1292 -128
rect 1326 -162 1360 -128
rect 1394 -162 1428 -128
rect 1462 -162 1496 -128
rect 1530 -162 1564 -128
rect 1598 -162 1632 -128
rect 1666 -162 1700 -128
rect 1734 -162 1768 -128
rect 1802 -162 1836 -128
rect 1870 -162 1904 -128
rect 1938 -162 1972 -128
rect 2006 -162 2040 -128
rect 2074 -162 2108 -128
rect 1160 -509 1194 -475
rect 1160 -593 1194 -559
rect 691 -692 725 -658
rect 691 -826 725 -792
rect 1160 -677 1194 -643
rect 1160 -760 1194 -726
rect 1160 -843 1194 -809
<< locali >>
rect 8893 2905 8917 2933
rect 8951 2905 8991 2933
rect 9025 2905 9065 2933
rect 9099 2905 9139 2933
rect 8951 2899 8974 2905
rect 9025 2899 9055 2905
rect 9099 2899 9136 2905
rect 9173 2899 9213 2933
rect 9247 2905 9287 2933
rect 9321 2905 9361 2933
rect 9395 2905 9435 2933
rect 9469 2905 9493 2933
rect 9251 2899 9287 2905
rect 9332 2899 9361 2905
rect 9413 2899 9435 2905
rect 8927 2871 8974 2899
rect 9008 2871 9055 2899
rect 9089 2871 9136 2899
rect 9170 2871 9217 2899
rect 9251 2871 9298 2899
rect 9332 2871 9379 2899
rect 9413 2871 9459 2899
rect 9132 2788 9260 2797
rect 9166 2754 9226 2788
rect 9132 2745 9260 2754
rect 8811 2677 8845 2743
rect 8811 2609 8845 2643
rect 8907 2632 9035 2641
rect 8941 2598 9001 2632
rect 8907 2589 9035 2598
rect 8811 2541 8845 2571
rect 8811 2487 8845 2499
rect 9132 2475 9260 2484
rect 9166 2441 9226 2475
rect 9132 2432 9260 2441
rect 8944 2179 8995 2213
rect 9029 2179 9079 2213
rect 9113 2179 9163 2213
rect 8806 2152 8840 2168
rect 8806 2074 8840 2118
rect 8839 2040 8840 2074
rect 8805 2018 8840 2040
rect 8805 2002 8806 2018
rect 8839 1968 8840 1984
rect 9186 1923 9252 1957
rect 9286 1923 9351 1957
rect 4264 1720 4520 1729
rect 4264 1686 4276 1720
rect 4310 1686 4375 1720
rect 4409 1686 4474 1720
rect 4508 1686 4520 1720
rect 1428 1578 1470 1612
rect 1504 1578 1546 1612
rect 1580 1578 1621 1612
rect 1091 1551 1125 1567
rect 1091 1474 1125 1517
rect 4264 1537 4520 1686
rect 4264 1503 4280 1537
rect 4314 1503 4375 1537
rect 4409 1503 4470 1537
rect 4504 1503 4520 1537
rect 4649 1674 4687 1708
rect 2333 1457 2345 1491
rect 2391 1457 2417 1491
rect 2459 1457 2489 1491
rect 2527 1457 2561 1491
rect 2595 1457 2629 1491
rect 2667 1457 2697 1491
rect 2739 1457 2765 1491
rect 2811 1457 2833 1491
rect 2883 1457 2901 1491
rect 2955 1457 2969 1491
rect 3027 1457 3037 1491
rect 3099 1457 3105 1491
rect 3171 1457 3173 1491
rect 3207 1457 3209 1491
rect 3275 1457 3281 1491
rect 3343 1457 3353 1491
rect 3411 1457 3425 1491
rect 3479 1457 3497 1491
rect 3547 1457 3569 1491
rect 3615 1457 3641 1491
rect 3683 1457 3738 1491
rect 1091 1397 1125 1440
rect -115 1362 -47 1396
rect -13 1362 22 1396
rect 56 1362 91 1396
rect 125 1362 160 1396
rect 194 1362 229 1396
rect 263 1362 298 1396
rect 332 1362 367 1396
rect 401 1362 436 1396
rect 470 1362 504 1396
rect 538 1362 572 1396
rect 606 1362 640 1396
rect 674 1362 708 1396
rect 742 1362 776 1396
rect 810 1362 858 1396
rect 892 1362 930 1396
rect 964 1362 1035 1396
rect -115 1327 -81 1362
rect 1001 1328 1035 1362
rect -115 1258 -81 1293
rect -115 1189 -81 1224
rect -115 1120 -81 1155
rect -115 1068 -81 1086
rect 517 1302 602 1305
rect 517 1268 543 1302
rect 577 1268 602 1302
rect 517 1197 602 1268
rect 517 1163 543 1197
rect 577 1163 602 1197
rect -115 982 -81 1017
rect -115 913 -81 945
rect -115 844 -81 856
rect -115 801 -81 810
rect 211 1034 220 1068
rect 254 1034 263 1068
rect 211 979 263 1034
rect 211 945 220 979
rect 254 945 263 979
rect 211 890 263 945
rect 211 856 220 890
rect 254 856 263 890
rect 211 801 263 856
rect 211 767 220 801
rect 254 767 263 801
rect -115 706 -81 741
rect -115 637 -81 672
rect -115 567 -81 603
rect -115 497 -81 533
rect -5 565 4 599
rect 38 565 47 599
rect -5 504 47 565
rect -5 470 4 504
rect 38 470 47 504
rect -115 427 -81 463
rect -115 357 -81 393
rect -115 287 -81 323
rect -115 217 -81 253
rect -115 147 -81 183
rect -115 77 -81 113
rect -115 7 -81 43
rect 427 154 436 188
rect 470 154 479 188
rect 427 102 479 154
rect 427 68 436 102
rect 470 68 479 102
rect 427 15 479 68
rect 427 -19 436 15
rect 470 -19 479 15
rect -115 -63 -81 -27
rect -115 -121 -81 -97
rect 517 -168 602 1163
rect 733 1302 818 1305
rect 733 1268 759 1302
rect 793 1268 818 1302
rect 733 1197 818 1268
rect 733 1163 759 1197
rect 793 1163 818 1197
rect 643 1034 652 1068
rect 686 1034 695 1068
rect 643 979 695 1034
rect 643 945 652 979
rect 686 945 695 979
rect 643 890 695 945
rect 643 856 652 890
rect 686 856 695 890
rect 643 801 695 856
rect 643 767 652 801
rect 686 767 695 801
rect 733 690 818 1163
rect 1001 1239 1035 1294
rect 1001 1150 1035 1205
rect 1091 1319 1125 1363
rect 1934 1362 1973 1396
rect 2007 1362 2046 1396
rect 2312 1365 2321 1399
rect 2355 1365 2364 1399
rect 1091 1241 1125 1263
rect 1091 1197 1125 1207
rect 2312 1318 2364 1365
rect 2312 1284 2321 1318
rect 2355 1284 2364 1318
rect 2312 1237 2364 1284
rect 2312 1203 2321 1237
rect 2355 1203 2364 1237
rect 1428 1146 1470 1180
rect 1504 1146 1546 1180
rect 1580 1146 1621 1180
rect 1001 1062 1035 1116
rect 1001 1028 1069 1062
rect 1103 1028 1142 1062
rect 1176 1028 1215 1062
rect 1249 1028 1288 1062
rect 1322 1028 1361 1062
rect 1395 1028 1433 1062
rect 1467 1028 1505 1062
rect 1539 1028 1577 1062
rect 1611 1028 1649 1062
rect 1683 1028 1721 1062
rect 1755 1028 1793 1062
rect 1827 1028 1865 1062
rect 1899 1028 1937 1062
rect 1971 1028 2009 1062
rect 2043 1028 2081 1062
rect 2115 1028 2139 1062
rect 1818 902 1827 936
rect 1861 902 1870 936
rect 1818 842 1870 902
rect 1818 808 1827 842
rect 1861 808 1870 842
rect 754 656 792 690
rect 733 -168 818 656
rect 1070 565 1079 599
rect 1113 565 1122 599
rect 1070 505 1122 565
rect 1070 471 1079 505
rect 1113 471 1122 505
rect 1382 565 1391 599
rect 1425 565 1434 599
rect 1382 505 1434 565
rect 1382 471 1391 505
rect 1425 471 1434 505
rect 1694 565 1703 599
rect 1737 565 1746 599
rect 1694 505 1746 565
rect 1694 471 1703 505
rect 1737 471 1746 505
rect 1226 337 1235 371
rect 1269 337 1278 371
rect 1226 277 1278 337
rect 1226 243 1235 277
rect 1269 243 1278 277
rect 1538 337 1547 371
rect 1581 337 1590 371
rect 1538 277 1590 337
rect 1538 243 1547 277
rect 1581 243 1590 277
rect 1818 188 1870 808
rect 2130 902 2139 936
rect 2173 902 2182 936
rect 2130 842 2182 902
rect 2130 808 2139 842
rect 2173 808 2182 842
rect 1974 702 1983 736
rect 2017 702 2026 736
rect 1974 642 2026 702
rect 1974 608 1983 642
rect 2017 608 2026 642
rect 859 154 868 188
rect 902 154 911 188
rect 859 102 911 154
rect 859 68 868 102
rect 902 68 911 102
rect 859 15 911 68
rect 859 -19 868 15
rect 902 -19 911 15
rect 1818 154 1827 188
rect 1861 154 1870 188
rect 1818 102 1870 154
rect 1818 68 1827 102
rect 1861 68 1870 102
rect 1818 15 1870 68
rect 1818 -19 1827 15
rect 1861 -19 1870 15
rect 2130 188 2182 808
rect 2468 810 2520 1387
rect 2624 1365 2633 1399
rect 2667 1365 2676 1399
rect 2624 1318 2676 1365
rect 2624 1284 2633 1318
rect 2667 1284 2676 1318
rect 2624 1237 2676 1284
rect 2624 1203 2633 1237
rect 2667 1203 2676 1237
rect 2748 895 2800 1387
rect 2904 1365 2913 1399
rect 2947 1365 2956 1399
rect 2904 1318 2956 1365
rect 2904 1284 2913 1318
rect 2947 1284 2956 1318
rect 2904 1237 2956 1284
rect 2904 1203 2913 1237
rect 2947 1203 2956 1237
rect 3216 1365 3225 1399
rect 3259 1365 3268 1399
rect 3216 1318 3268 1365
rect 3216 1284 3225 1318
rect 3259 1284 3268 1318
rect 3216 1237 3268 1284
rect 3216 1203 3225 1237
rect 3259 1203 3268 1237
rect 3528 1365 3537 1399
rect 3571 1365 3580 1399
rect 3528 1318 3580 1365
rect 3528 1284 3537 1318
rect 3571 1284 3580 1318
rect 3528 1237 3580 1284
rect 3528 1203 3537 1237
rect 3571 1203 3580 1237
rect 3823 908 3857 1256
rect 2748 861 2757 895
rect 2791 861 2800 895
rect 2468 749 2706 810
rect 2748 801 2800 861
rect 3069 836 3103 874
rect 3381 836 3415 874
rect 3693 836 3727 874
rect 3823 836 3857 874
rect 3999 1212 4033 1250
rect 4342 1249 4458 1441
rect 4342 1215 4349 1249
rect 4383 1215 4421 1249
rect 4455 1215 4458 1249
rect 4342 1214 4458 1215
rect 3999 824 4033 1178
rect 4615 1140 4723 1674
rect 4835 1538 4848 1572
rect 4885 1538 4920 1572
rect 4958 1538 4989 1572
rect 5034 1538 5058 1572
rect 5109 1538 5127 1572
rect 5184 1538 5196 1572
rect 5259 1538 5265 1572
rect 5299 1538 5300 1572
rect 5367 1538 5375 1572
rect 5435 1538 5450 1572
rect 5503 1538 5525 1572
rect 5571 1538 5600 1572
rect 5639 1538 5673 1572
rect 5709 1538 5723 1572
rect 5779 1538 5794 1572
rect 5829 1538 5905 1572
rect 5943 1538 5959 1572
rect 4790 1467 4918 1476
rect 4824 1433 4884 1467
rect 4790 1424 4918 1433
rect 5215 1467 5343 1476
rect 5249 1433 5309 1467
rect 5215 1424 5343 1433
rect 5578 1365 5684 1538
rect 5737 1467 5865 1476
rect 5771 1433 5831 1467
rect 5737 1424 5865 1433
rect 5970 1392 6076 1488
rect 4879 1340 5107 1349
rect 4879 1306 4979 1340
rect 5013 1306 5073 1340
rect 4879 1297 5107 1306
rect 5392 1340 5520 1349
rect 5426 1306 5486 1340
rect 5612 1331 5650 1365
rect 5978 1314 6076 1392
rect 5392 1297 5520 1306
rect 4615 1130 4701 1140
rect 4085 1027 4701 1130
rect 4879 1111 4931 1297
rect 6004 1280 6042 1314
rect 6236 1452 6304 1486
rect 6346 1452 6372 1486
rect 6419 1452 6440 1486
rect 6492 1452 6508 1486
rect 6565 1452 6576 1486
rect 6638 1452 6644 1486
rect 6711 1452 6712 1486
rect 6746 1452 6750 1486
rect 6814 1452 6823 1486
rect 6882 1452 6896 1486
rect 6950 1452 6969 1486
rect 7018 1452 7042 1486
rect 7086 1452 7115 1486
rect 7154 1452 7188 1486
rect 7222 1452 7256 1486
rect 7295 1452 7324 1486
rect 7368 1452 7392 1486
rect 7441 1452 7460 1486
rect 7514 1452 7528 1486
rect 7587 1452 7596 1486
rect 7660 1452 7664 1486
rect 7698 1452 7699 1486
rect 7766 1452 7772 1486
rect 7834 1452 7845 1486
rect 7902 1452 7918 1486
rect 7970 1452 7991 1486
rect 8038 1452 8064 1486
rect 8106 1452 8137 1486
rect 8174 1452 8208 1486
rect 8244 1452 8276 1486
rect 8317 1452 8344 1486
rect 8390 1452 8412 1486
rect 8463 1452 8480 1486
rect 8536 1452 8548 1486
rect 8609 1452 8616 1486
rect 8682 1452 8684 1486
rect 8718 1452 8721 1486
rect 8786 1452 8794 1486
rect 8854 1452 8867 1486
rect 8922 1452 8940 1486
rect 8990 1452 9013 1486
rect 9058 1452 9086 1486
rect 9126 1452 9159 1486
rect 9194 1452 9228 1486
rect 9266 1452 9296 1486
rect 9339 1452 9364 1486
rect 9412 1452 9432 1486
rect 9485 1452 9500 1486
rect 9558 1452 9568 1486
rect 9631 1452 9636 1486
rect 9738 1452 9743 1486
rect 9806 1452 9816 1486
rect 9874 1452 9889 1486
rect 9942 1452 9976 1486
rect 10016 1452 10125 1486
rect 6236 1414 6273 1452
rect 6236 1380 6239 1414
rect 10088 1418 10125 1452
rect 10088 1414 10091 1418
rect 10122 1380 10125 1384
rect 6236 1352 6273 1380
rect 6270 1339 6273 1352
rect 6236 1305 6239 1318
rect 6236 1284 6273 1305
rect 6270 1264 6273 1284
rect 5027 1216 5101 1231
rect 4745 1095 4931 1111
rect 4779 1061 4817 1095
rect 4851 1061 4931 1095
rect 5020 1197 5101 1216
rect 5135 1216 5175 1231
rect 5209 1216 5249 1231
rect 5283 1216 5323 1231
rect 5357 1216 5397 1231
rect 5135 1197 5159 1216
rect 5209 1197 5227 1216
rect 5283 1197 5295 1216
rect 5357 1197 5363 1216
rect 5020 1182 5159 1197
rect 5193 1182 5227 1197
rect 5261 1182 5295 1197
rect 5329 1182 5363 1197
rect 5431 1216 5472 1231
rect 5506 1216 5547 1231
rect 5581 1216 5622 1231
rect 5656 1216 5697 1231
rect 5731 1216 5772 1231
rect 5806 1216 5847 1231
rect 5881 1216 5922 1231
rect 6122 1216 6164 1231
rect 6236 1230 6239 1250
rect 6236 1216 6273 1230
rect 5397 1182 5431 1197
rect 5465 1197 5472 1216
rect 5533 1197 5547 1216
rect 5601 1197 5622 1216
rect 5669 1197 5697 1216
rect 5465 1182 5499 1197
rect 5533 1182 5567 1197
rect 5601 1182 5635 1197
rect 5669 1182 5703 1197
rect 5737 1182 5771 1216
rect 5806 1197 5839 1216
rect 5881 1197 5907 1216
rect 5956 1197 5975 1216
rect 5805 1182 5839 1197
rect 5873 1182 5907 1197
rect 5941 1182 5975 1197
rect 6009 1182 6043 1216
rect 6077 1197 6164 1216
rect 6077 1182 6165 1197
rect 6199 1189 6273 1216
rect 6355 1308 6389 1346
rect 6355 1236 6389 1274
rect 6867 1308 6901 1346
rect 6867 1236 6901 1274
rect 7379 1308 7413 1346
rect 7379 1236 7413 1274
rect 7891 1308 7925 1346
rect 7891 1236 7925 1274
rect 8403 1308 8437 1346
rect 8403 1236 8437 1274
rect 8915 1308 8949 1346
rect 8915 1236 8949 1274
rect 9267 1308 9301 1346
rect 9267 1236 9301 1274
rect 9619 1308 9653 1346
rect 9619 1236 9653 1274
rect 9971 1308 10005 1346
rect 9971 1236 10005 1274
rect 10088 1350 10125 1380
rect 10088 1342 10091 1350
rect 10122 1308 10125 1316
rect 10088 1282 10125 1308
rect 10088 1270 10091 1282
rect 10122 1236 10125 1248
rect 10088 1214 10125 1236
rect 6199 1182 6239 1189
rect 5020 1159 5061 1182
rect 5020 1125 5027 1159
rect 5020 1094 5061 1125
rect 5188 1094 5200 1128
rect 5242 1094 5272 1128
rect 5310 1094 5344 1128
rect 5378 1094 5412 1128
rect 5450 1094 5480 1128
rect 5522 1094 5548 1128
rect 5594 1094 5616 1128
rect 5666 1094 5684 1128
rect 5738 1094 5752 1128
rect 5810 1094 5820 1128
rect 5882 1094 5888 1128
rect 5954 1094 5969 1128
rect 6239 1114 6273 1155
rect 4745 1059 4931 1061
rect 5027 1079 5061 1094
rect 2748 767 2757 801
rect 2791 767 2800 801
rect 2231 681 2382 715
rect 2416 681 2476 715
rect 2510 681 2570 715
rect 2604 681 2620 715
rect 2231 636 2620 681
rect 2231 630 2309 636
rect 2231 596 2255 630
rect 2289 596 2309 630
rect 2654 602 2706 749
rect 2231 558 2309 596
rect 2231 524 2255 558
rect 2289 524 2309 558
rect 2231 506 2309 524
rect 2373 568 2662 602
rect 2696 568 2757 602
rect 2791 568 2852 602
rect 2886 568 2902 602
rect 2373 518 2902 568
rect 2373 484 2662 518
rect 2696 484 2757 518
rect 2791 484 2852 518
rect 2886 484 2902 518
rect 2958 590 2974 602
rect 2958 556 2964 590
rect 3008 568 3069 602
rect 3103 568 3164 602
rect 3198 568 3214 602
rect 2998 556 3214 568
rect 2958 518 3214 556
rect 2958 484 2964 518
rect 3008 484 3069 518
rect 3103 484 3164 518
rect 3198 484 3214 518
rect 3270 590 3286 602
rect 3270 556 3276 590
rect 3320 568 3364 602
rect 3398 568 3442 602
rect 3476 568 3519 602
rect 3553 568 3596 602
rect 3630 568 3646 602
rect 3310 556 3646 568
rect 3270 518 3646 556
rect 3270 484 3276 518
rect 3320 484 3364 518
rect 3398 484 3442 518
rect 3476 484 3519 518
rect 3553 484 3596 518
rect 3630 484 3646 518
rect 2373 297 2491 484
rect 2748 387 2757 421
rect 2791 387 2800 421
rect 2130 154 2139 188
rect 2173 154 2182 188
rect 2130 102 2182 154
rect 2130 68 2139 102
rect 2173 68 2182 102
rect 2130 15 2182 68
rect 2130 -19 2139 15
rect 2173 -19 2182 15
rect 2258 268 2292 292
rect 2258 196 2292 234
rect 2258 124 2292 162
rect 2258 51 2292 90
rect 2258 -22 2292 17
rect 2258 -80 2292 -56
rect 2373 281 2508 297
rect 2373 247 2385 281
rect 2419 247 2462 281
rect 2496 247 2508 281
rect 2373 231 2508 247
rect 2373 -33 2491 231
rect 2592 222 2644 330
rect 2748 327 2800 387
rect 2748 293 2757 327
rect 2791 293 2800 327
rect 2592 188 2601 222
rect 2635 188 2644 222
rect 2592 150 2644 188
rect 2592 116 2601 150
rect 2635 116 2644 150
rect 2904 222 2956 330
rect 3069 327 3103 365
rect 2904 188 2913 222
rect 2947 188 2956 222
rect 2904 150 2956 188
rect 2904 116 2913 150
rect 2947 116 2956 150
rect 3216 222 3268 330
rect 3381 310 3415 348
rect 3216 188 3225 222
rect 3259 188 3268 222
rect 3216 150 3268 188
rect 3216 116 3225 150
rect 3259 116 3268 150
rect 3528 222 3580 330
rect 3693 310 3727 348
rect 3823 283 3857 802
rect 3893 740 3975 743
rect 4085 740 4183 1027
rect 5027 999 5061 1045
rect 3893 725 4183 740
rect 3893 691 3913 725
rect 3947 691 4183 725
rect 3893 641 4183 691
rect 3893 607 3913 641
rect 3947 638 4183 641
rect 4262 884 4296 908
rect 4262 814 4296 850
rect 4262 744 4296 780
rect 4262 674 4296 710
rect 3947 607 3975 638
rect 3893 557 3975 607
rect 3893 523 3913 557
rect 3947 523 3975 557
rect 3893 473 3975 523
rect 3893 439 3913 473
rect 3947 439 3975 473
rect 3893 389 3975 439
rect 3893 355 3913 389
rect 3947 355 3975 389
rect 3893 336 3975 355
rect 4262 604 4296 640
rect 4262 533 4296 570
rect 4262 462 4296 499
rect 4262 412 4296 428
rect 4262 340 4296 357
rect 4262 285 4296 286
rect 3528 188 3537 222
rect 3571 188 3580 222
rect 3528 150 3580 188
rect 3528 116 3537 150
rect 3571 116 3580 150
rect 3992 249 4296 285
rect 3992 222 4262 249
rect 3992 188 3999 222
rect 4033 215 4262 222
rect 4033 188 4296 215
rect 3992 178 4296 188
rect 3992 150 4262 178
rect 3992 116 3999 150
rect 4033 144 4262 150
rect 4033 116 4296 144
rect 3992 107 4296 116
rect 3992 73 4262 107
rect 2593 23 2609 57
rect 2643 23 2657 57
rect 2715 23 2725 57
rect 2787 23 2793 57
rect 2859 23 2861 57
rect 2895 23 2897 57
rect 2963 23 2969 57
rect 3031 23 3041 57
rect 3099 23 3113 57
rect 3167 23 3185 57
rect 3235 23 3257 57
rect 3303 23 3329 57
rect 3371 23 3401 57
rect 3439 23 3473 57
rect 3507 23 3541 57
rect 3579 23 3609 57
rect 3651 23 3677 57
rect 3723 23 3735 57
rect 3992 36 4296 73
rect 4330 727 4432 951
rect 4901 917 4935 963
rect 6239 1039 6273 1080
rect 10088 1198 10091 1214
rect 10122 1164 10125 1180
rect 10088 1146 10125 1164
rect 10088 1126 10091 1146
rect 10122 1092 10125 1112
rect 10088 1078 10125 1092
rect 10088 1054 10091 1078
rect 10122 1020 10125 1044
rect 5027 920 5061 965
rect 5143 898 5177 948
rect 5455 898 5489 948
rect 6239 964 6273 1005
rect 6239 889 6273 930
rect 6239 814 6273 855
rect 6611 948 6645 986
rect 6611 876 6645 914
rect 7123 948 7157 986
rect 7123 876 7157 914
rect 7635 948 7669 986
rect 7635 876 7669 914
rect 8147 948 8181 986
rect 8147 876 8181 914
rect 8659 948 8693 986
rect 8659 876 8693 914
rect 9091 948 9125 986
rect 9091 876 9125 914
rect 9443 948 9477 986
rect 9443 876 9477 914
rect 9795 948 9829 986
rect 9795 876 9829 914
rect 10088 1010 10125 1020
rect 10088 982 10091 1010
rect 10122 948 10125 976
rect 10088 942 10125 948
rect 10088 910 10091 942
rect 10122 876 10125 908
rect 10088 874 10125 876
rect 10088 840 10091 874
rect 10088 838 10125 840
rect 10122 806 10125 838
rect 4330 693 4389 727
rect 4423 693 4432 727
rect 4330 647 4432 693
rect 4330 613 4389 647
rect 4423 613 4432 647
rect 4901 647 4935 693
rect 5967 691 6076 750
rect 6001 657 6039 691
rect 6073 657 6076 691
rect 4330 60 4432 613
rect 4630 526 4689 609
rect 4630 492 4645 526
rect 4679 492 4689 526
rect 4630 436 4689 492
rect 4630 402 4645 436
rect 4679 402 4689 436
rect 5299 508 5333 546
rect 5299 436 5333 474
rect 5611 508 5645 546
rect 5611 436 5645 474
rect 4477 313 4532 347
rect 4574 313 4586 347
rect 4630 334 4689 402
rect 3992 2 4262 36
rect 3992 -22 4296 2
rect 2407 -67 2445 -33
rect 2479 -67 2491 -33
rect 1124 -162 1146 -128
rect 1180 -162 1190 -128
rect 1252 -162 1258 -128
rect 1324 -162 1326 -128
rect 1360 -162 1362 -128
rect 1428 -162 1434 -128
rect 1496 -162 1506 -128
rect 1564 -162 1578 -128
rect 1632 -162 1650 -128
rect 1700 -162 1722 -128
rect 1768 -162 1794 -128
rect 1836 -162 1866 -128
rect 1904 -162 1938 -128
rect 1972 -162 2006 -128
rect 2044 -162 2074 -128
rect 2116 -162 2128 -128
rect 4631 -144 4689 334
rect 4730 313 4747 347
rect 4781 313 4811 347
rect 4853 313 4865 347
rect 5967 326 6076 657
rect 6375 728 8904 804
rect 6375 694 6414 728
rect 6450 694 6485 728
rect 6527 694 6554 728
rect 6606 694 6623 728
rect 6685 694 6692 728
rect 6726 694 6731 728
rect 6795 694 6811 728
rect 6864 694 6891 728
rect 6933 694 6968 728
rect 7005 694 7037 728
rect 7085 694 7106 728
rect 7165 694 7175 728
rect 7209 694 7244 728
rect 7278 694 7314 728
rect 7348 694 7384 728
rect 7418 694 7454 728
rect 7488 694 7514 728
rect 7558 694 7590 728
rect 7628 694 7664 728
rect 7700 694 7734 728
rect 7776 694 7804 728
rect 7852 694 7874 728
rect 7928 694 7944 728
rect 8005 694 8014 728
rect 8082 694 8084 728
rect 8118 694 8125 728
rect 8188 694 8202 728
rect 8258 694 8279 728
rect 8328 694 8356 728
rect 8398 694 8434 728
rect 8468 694 8504 728
rect 8538 694 8574 728
rect 8608 694 8644 728
rect 8678 694 8714 728
rect 8748 694 8784 728
rect 8818 694 8854 728
rect 8888 694 8904 728
rect 6375 618 8904 694
rect 8960 728 9972 804
rect 8960 694 8976 728
rect 9010 694 9047 728
rect 9081 694 9118 728
rect 9152 694 9190 728
rect 9224 694 9262 728
rect 9296 694 9334 728
rect 9368 694 9406 728
rect 9440 694 9478 728
rect 9512 694 9550 728
rect 9604 694 9622 728
rect 9656 694 9658 728
rect 9692 694 9694 728
rect 9728 694 9747 728
rect 9800 694 9836 728
rect 9872 694 9910 728
rect 9959 694 9972 728
rect 8960 618 9972 694
rect 10088 772 10091 804
rect 10088 766 10125 772
rect 10122 738 10125 766
rect 10088 704 10091 732
rect 10088 694 10125 704
rect 10122 670 10125 694
rect 10088 636 10091 660
rect 10088 622 10125 636
rect 10122 602 10125 622
rect 6123 508 6157 546
rect 6123 436 6157 474
rect 6611 508 6645 546
rect 6611 436 6645 474
rect 7123 508 7157 546
rect 7123 436 7157 474
rect 7635 508 7669 546
rect 7635 436 7669 474
rect 8147 508 8181 546
rect 8147 436 8181 474
rect 8659 508 8693 546
rect 8659 436 8693 474
rect 9091 508 9125 546
rect 9091 436 9125 474
rect 9443 508 9477 546
rect 9443 436 9477 474
rect 9795 508 9829 546
rect 9795 436 9829 474
rect 10088 568 10091 588
rect 10088 550 10125 568
rect 10122 534 10125 550
rect 10088 500 10091 516
rect 10088 478 10125 500
rect 10122 466 10125 478
rect 10088 432 10091 444
rect 10088 406 10125 432
rect 4730 27 4853 313
rect 5143 252 5177 290
rect 5143 180 5177 218
rect 4900 111 4909 145
rect 4943 111 4952 145
rect 4900 51 4952 111
rect 4730 -7 4746 27
rect 4780 -7 4816 27
rect 4850 -7 4866 27
rect 4900 17 4909 51
rect 4943 17 4952 51
rect 6001 292 6039 326
rect 6073 312 6076 326
rect 10122 398 10125 406
rect 10088 364 10091 372
rect 10088 334 10125 364
rect 10122 330 10125 334
rect 10088 296 10091 300
rect 5455 252 5489 290
rect 10088 262 10125 296
rect 5455 180 5489 218
rect 5867 148 5901 186
rect 5027 72 5061 139
rect 5867 76 5901 114
rect 6355 148 6389 186
rect 6355 76 6389 114
rect 6867 148 6901 186
rect 6867 76 6901 114
rect 7379 148 7413 186
rect 7379 76 7413 114
rect 7891 148 7925 186
rect 7891 76 7925 114
rect 8403 148 8437 186
rect 8403 76 8437 114
rect 8915 148 8949 186
rect 8915 76 8949 114
rect 9267 148 9301 186
rect 9267 76 9301 114
rect 9619 148 9653 186
rect 9619 76 9653 114
rect 9971 148 10005 186
rect 9971 76 10005 114
rect 10088 194 10125 228
rect 10088 190 10091 194
rect 10122 156 10125 160
rect 10088 126 10125 156
rect 10088 117 10091 126
rect 10122 83 10125 92
rect 10088 44 10125 83
rect 4903 -143 4943 17
rect 5027 -28 5061 38
rect 10122 10 10125 44
rect 10088 6 10125 10
rect 10088 -28 10122 6
rect 5027 -62 5071 -28
rect 5133 -62 5139 -28
rect 5206 -62 5207 -28
rect 5241 -62 5245 -28
rect 5309 -62 5318 -28
rect 5377 -62 5391 -28
rect 5445 -62 5464 -28
rect 5513 -62 5537 -28
rect 5581 -62 5610 -28
rect 5649 -62 5683 -28
rect 5717 -62 5751 -28
rect 5789 -62 5819 -28
rect 5861 -62 5887 -28
rect 5933 -62 5955 -28
rect 6005 -62 6023 -28
rect 6077 -62 6091 -28
rect 6149 -62 6159 -28
rect 6221 -62 6285 -28
rect 6345 -62 6353 -28
rect 6418 -62 6421 -28
rect 6455 -62 6457 -28
rect 6523 -62 6530 -28
rect 6591 -62 6603 -28
rect 6659 -62 6676 -28
rect 6727 -62 6749 -28
rect 6795 -62 6822 -28
rect 6863 -62 6895 -28
rect 6931 -62 6965 -28
rect 7002 -62 7033 -28
rect 7075 -62 7101 -28
rect 7148 -62 7169 -28
rect 7221 -62 7237 -28
rect 7294 -62 7305 -28
rect 7367 -62 7373 -28
rect 7440 -62 7441 -28
rect 7475 -62 7479 -28
rect 7543 -62 7552 -28
rect 7611 -62 7625 -28
rect 7679 -62 7698 -28
rect 7747 -62 7771 -28
rect 7815 -62 7844 -28
rect 7883 -62 7917 -28
rect 7951 -62 7985 -28
rect 8024 -62 8053 -28
rect 8097 -62 8136 -28
rect 8170 -62 8209 -28
rect 8243 -62 8282 -28
rect 8316 -62 8355 -28
rect 8389 -62 8428 -28
rect 8462 -62 8501 -28
rect 8535 -62 8574 -28
rect 8608 -62 8647 -28
rect 8681 -62 8720 -28
rect 8754 -62 8792 -28
rect 8826 -62 8864 -28
rect 8898 -62 8936 -28
rect 8970 -62 9008 -28
rect 9042 -62 9080 -28
rect 9114 -62 9152 -28
rect 9186 -62 9224 -28
rect 9258 -62 9296 -28
rect 9330 -62 9368 -28
rect 9402 -62 9440 -28
rect 9474 -62 9512 -28
rect 9546 -62 9584 -28
rect 9618 -62 9656 -28
rect 9690 -62 9728 -28
rect 9762 -62 9800 -28
rect 9834 -62 9872 -28
rect 9906 -62 9944 -28
rect 9978 -62 10016 -28
rect 10050 -62 10122 -28
rect 68 -202 80 -168
rect 122 -202 152 -168
rect 190 -202 224 -168
rect 258 -202 292 -168
rect 330 -202 360 -168
rect 402 -202 428 -168
rect 474 -202 496 -168
rect 546 -202 564 -168
rect 618 -202 632 -168
rect 690 -202 700 -168
rect 762 -202 768 -168
rect 834 -202 857 -168
rect 685 -255 1197 -241
rect 685 -289 703 -255
rect 737 -289 778 -255
rect 812 -289 853 -255
rect 887 -289 928 -255
rect 962 -289 1003 -255
rect 1037 -289 1077 -255
rect 1111 -289 1151 -255
rect 1185 -289 1197 -255
rect 685 -475 1197 -289
rect 685 -509 1160 -475
rect 1194 -509 1197 -475
rect 1242 -434 1420 -409
rect 1242 -468 1257 -434
rect 1291 -468 1329 -434
rect 1363 -468 1420 -434
rect 1242 -485 1420 -468
rect 685 -559 1197 -509
rect 685 -593 1160 -559
rect 1194 -593 1197 -559
rect -269 -631 -231 -597
rect 685 -643 1197 -593
rect 685 -658 1160 -643
rect 685 -692 691 -658
rect 725 -677 1160 -658
rect 1194 -677 1197 -643
rect 725 -692 1197 -677
rect 685 -726 1197 -692
rect 685 -760 1160 -726
rect 1194 -760 1197 -726
rect 685 -792 1197 -760
rect 685 -826 691 -792
rect 725 -809 1197 -792
rect 725 -826 1160 -809
rect 685 -843 1160 -826
rect 1194 -843 1197 -809
rect 685 -862 1197 -843
<< viali >>
rect 8893 2899 8917 2905
rect 8917 2899 8927 2905
rect 8974 2899 8991 2905
rect 8991 2899 9008 2905
rect 9055 2899 9065 2905
rect 9065 2899 9089 2905
rect 9136 2899 9139 2905
rect 9139 2899 9170 2905
rect 9217 2899 9247 2905
rect 9247 2899 9251 2905
rect 9298 2899 9321 2905
rect 9321 2899 9332 2905
rect 9379 2899 9395 2905
rect 9395 2899 9413 2905
rect 9459 2899 9469 2905
rect 9469 2899 9493 2905
rect 8893 2871 8927 2899
rect 8974 2871 9008 2899
rect 9055 2871 9089 2899
rect 9136 2871 9170 2899
rect 9217 2871 9251 2899
rect 9298 2871 9332 2899
rect 9379 2871 9413 2899
rect 9459 2871 9493 2899
rect 9132 2754 9166 2788
rect 9226 2754 9260 2788
rect 8811 2643 8845 2677
rect 8811 2575 8845 2605
rect 8907 2598 8941 2632
rect 9001 2598 9035 2632
rect 8811 2571 8845 2575
rect 8811 2507 8845 2533
rect 8811 2499 8845 2507
rect 9132 2441 9166 2475
rect 9226 2441 9260 2475
rect 8910 2179 8944 2213
rect 8995 2179 9029 2213
rect 9079 2179 9113 2213
rect 9163 2179 9197 2213
rect 8805 2040 8839 2074
rect 8805 1984 8806 2002
rect 8806 1984 8839 2002
rect 8805 1968 8839 1984
rect 9152 1923 9186 1957
rect 9252 1923 9286 1957
rect 9351 1923 9385 1957
rect 4276 1686 4310 1720
rect 4375 1686 4409 1720
rect 4474 1686 4508 1720
rect 1394 1578 1428 1612
rect 1470 1578 1504 1612
rect 1546 1578 1580 1612
rect 1621 1578 1655 1612
rect 4615 1674 4649 1708
rect 4687 1674 4721 1708
rect 2345 1457 2357 1491
rect 2357 1457 2379 1491
rect 2417 1457 2425 1491
rect 2425 1457 2451 1491
rect 2489 1457 2493 1491
rect 2493 1457 2523 1491
rect 2561 1457 2595 1491
rect 2633 1457 2663 1491
rect 2663 1457 2667 1491
rect 2705 1457 2731 1491
rect 2731 1457 2739 1491
rect 2777 1457 2799 1491
rect 2799 1457 2811 1491
rect 2849 1457 2867 1491
rect 2867 1457 2883 1491
rect 2921 1457 2935 1491
rect 2935 1457 2955 1491
rect 2993 1457 3003 1491
rect 3003 1457 3027 1491
rect 3065 1457 3071 1491
rect 3071 1457 3099 1491
rect 3137 1457 3139 1491
rect 3139 1457 3171 1491
rect 3209 1457 3241 1491
rect 3241 1457 3243 1491
rect 3281 1457 3309 1491
rect 3309 1457 3315 1491
rect 3353 1457 3377 1491
rect 3377 1457 3387 1491
rect 3425 1457 3445 1491
rect 3445 1457 3459 1491
rect 3497 1457 3513 1491
rect 3513 1457 3531 1491
rect 3569 1457 3581 1491
rect 3581 1457 3603 1491
rect 3641 1457 3649 1491
rect 3649 1457 3675 1491
rect 543 1268 577 1302
rect 543 1163 577 1197
rect -115 1051 -81 1068
rect -115 1034 -81 1051
rect -115 948 -81 979
rect -115 945 -81 948
rect -115 879 -81 890
rect -115 856 -81 879
rect -115 775 -81 801
rect -115 767 -81 775
rect 220 1034 254 1068
rect 220 945 254 979
rect 220 856 254 890
rect 220 767 254 801
rect 4 565 38 599
rect 4 470 38 504
rect 436 154 470 188
rect 436 68 470 102
rect 436 -19 470 15
rect 759 1268 793 1302
rect 759 1163 793 1197
rect 652 1034 686 1068
rect 652 945 686 979
rect 652 856 686 890
rect 652 767 686 801
rect 1900 1362 1934 1396
rect 1973 1362 2007 1396
rect 2046 1362 2080 1396
rect 2321 1365 2355 1399
rect 1091 1285 1125 1297
rect 1091 1263 1125 1285
rect 2321 1284 2355 1318
rect 2321 1203 2355 1237
rect 1091 1163 1125 1197
rect 1394 1146 1428 1180
rect 1470 1146 1504 1180
rect 1546 1146 1580 1180
rect 1621 1146 1655 1180
rect 1827 902 1861 936
rect 1827 808 1861 842
rect 720 656 754 690
rect 792 656 826 690
rect 1079 565 1113 599
rect 1079 471 1113 505
rect 1391 565 1425 599
rect 1391 471 1425 505
rect 1703 565 1737 599
rect 1703 471 1737 505
rect 1235 337 1269 371
rect 1235 243 1269 277
rect 1547 337 1581 371
rect 1547 243 1581 277
rect 2139 902 2173 936
rect 2139 808 2173 842
rect 1983 702 2017 736
rect 1983 608 2017 642
rect 868 154 902 188
rect 868 68 902 102
rect 868 -19 902 15
rect 1827 154 1861 188
rect 1827 68 1861 102
rect 1827 -19 1861 15
rect 2633 1365 2667 1399
rect 2633 1284 2667 1318
rect 2633 1203 2667 1237
rect 2913 1365 2947 1399
rect 2913 1284 2947 1318
rect 2913 1203 2947 1237
rect 3225 1365 3259 1399
rect 3225 1284 3259 1318
rect 3225 1203 3259 1237
rect 3537 1365 3571 1399
rect 3537 1284 3571 1318
rect 3537 1203 3571 1237
rect 2757 861 2791 895
rect 3069 874 3103 908
rect 3069 802 3103 836
rect 3381 874 3415 908
rect 3381 802 3415 836
rect 3693 874 3727 908
rect 3693 802 3727 836
rect 3823 874 3857 908
rect 3823 802 3857 836
rect 3999 1250 4033 1284
rect 4349 1215 4383 1249
rect 4421 1215 4455 1249
rect 3999 1178 4033 1212
rect 4848 1538 4851 1572
rect 4851 1538 4882 1572
rect 4924 1538 4954 1572
rect 4954 1538 4958 1572
rect 5000 1538 5023 1572
rect 5023 1538 5034 1572
rect 5075 1538 5092 1572
rect 5092 1538 5109 1572
rect 5150 1538 5161 1572
rect 5161 1538 5184 1572
rect 5225 1538 5230 1572
rect 5230 1538 5259 1572
rect 5300 1538 5333 1572
rect 5333 1538 5334 1572
rect 5375 1538 5401 1572
rect 5401 1538 5409 1572
rect 5450 1538 5469 1572
rect 5469 1538 5484 1572
rect 5525 1538 5537 1572
rect 5537 1538 5559 1572
rect 5600 1538 5605 1572
rect 5605 1538 5634 1572
rect 5675 1538 5707 1572
rect 5707 1538 5709 1572
rect 5794 1538 5795 1572
rect 5795 1538 5828 1572
rect 5905 1538 5909 1572
rect 5909 1538 5939 1572
rect 4790 1433 4824 1467
rect 4884 1433 4918 1467
rect 5215 1433 5249 1467
rect 5309 1433 5343 1467
rect 5737 1433 5771 1467
rect 5831 1433 5865 1467
rect 4979 1306 5013 1340
rect 5073 1306 5107 1340
rect 5392 1306 5426 1340
rect 5486 1306 5520 1340
rect 5578 1331 5612 1365
rect 5650 1331 5684 1365
rect 5970 1280 6004 1314
rect 6042 1280 6076 1314
rect 6312 1452 6338 1486
rect 6338 1452 6346 1486
rect 6385 1452 6406 1486
rect 6406 1452 6419 1486
rect 6458 1452 6474 1486
rect 6474 1452 6492 1486
rect 6531 1452 6542 1486
rect 6542 1452 6565 1486
rect 6604 1452 6610 1486
rect 6610 1452 6638 1486
rect 6677 1452 6678 1486
rect 6678 1452 6711 1486
rect 6750 1452 6780 1486
rect 6780 1452 6784 1486
rect 6823 1452 6848 1486
rect 6848 1452 6857 1486
rect 6896 1452 6916 1486
rect 6916 1452 6930 1486
rect 6969 1452 6984 1486
rect 6984 1452 7003 1486
rect 7042 1452 7052 1486
rect 7052 1452 7076 1486
rect 7115 1452 7120 1486
rect 7120 1452 7149 1486
rect 7188 1452 7222 1486
rect 7261 1452 7290 1486
rect 7290 1452 7295 1486
rect 7334 1452 7358 1486
rect 7358 1452 7368 1486
rect 7407 1452 7426 1486
rect 7426 1452 7441 1486
rect 7480 1452 7494 1486
rect 7494 1452 7514 1486
rect 7553 1452 7562 1486
rect 7562 1452 7587 1486
rect 7626 1452 7630 1486
rect 7630 1452 7660 1486
rect 7699 1452 7732 1486
rect 7732 1452 7733 1486
rect 7772 1452 7800 1486
rect 7800 1452 7806 1486
rect 7845 1452 7868 1486
rect 7868 1452 7879 1486
rect 7918 1452 7936 1486
rect 7936 1452 7952 1486
rect 7991 1452 8004 1486
rect 8004 1452 8025 1486
rect 8064 1452 8072 1486
rect 8072 1452 8098 1486
rect 8137 1452 8140 1486
rect 8140 1452 8171 1486
rect 8210 1452 8242 1486
rect 8242 1452 8244 1486
rect 8283 1452 8310 1486
rect 8310 1452 8317 1486
rect 8356 1452 8378 1486
rect 8378 1452 8390 1486
rect 8429 1452 8446 1486
rect 8446 1452 8463 1486
rect 8502 1452 8514 1486
rect 8514 1452 8536 1486
rect 8575 1452 8582 1486
rect 8582 1452 8609 1486
rect 8648 1452 8650 1486
rect 8650 1452 8682 1486
rect 8721 1452 8752 1486
rect 8752 1452 8755 1486
rect 8794 1452 8820 1486
rect 8820 1452 8828 1486
rect 8867 1452 8888 1486
rect 8888 1452 8901 1486
rect 8940 1452 8956 1486
rect 8956 1452 8974 1486
rect 9013 1452 9024 1486
rect 9024 1452 9047 1486
rect 9086 1452 9092 1486
rect 9092 1452 9120 1486
rect 9159 1452 9160 1486
rect 9160 1452 9193 1486
rect 9232 1452 9262 1486
rect 9262 1452 9266 1486
rect 9305 1452 9330 1486
rect 9330 1452 9339 1486
rect 9378 1452 9398 1486
rect 9398 1452 9412 1486
rect 9451 1452 9466 1486
rect 9466 1452 9485 1486
rect 9524 1452 9534 1486
rect 9534 1452 9558 1486
rect 9597 1452 9602 1486
rect 9602 1452 9631 1486
rect 9670 1452 9704 1486
rect 9743 1452 9772 1486
rect 9772 1452 9777 1486
rect 9816 1452 9840 1486
rect 9840 1452 9850 1486
rect 9889 1452 9908 1486
rect 9908 1452 9923 1486
rect 9982 1452 10010 1486
rect 10010 1452 10016 1486
rect 6239 1380 6273 1414
rect 10088 1384 10091 1414
rect 10091 1384 10122 1414
rect 10088 1380 10122 1384
rect 6239 1318 6270 1339
rect 6270 1318 6273 1339
rect 6239 1305 6273 1318
rect 6239 1250 6270 1264
rect 6270 1250 6273 1264
rect 4745 1061 4779 1095
rect 4817 1061 4851 1095
rect 5101 1197 5135 1231
rect 5175 1216 5209 1231
rect 5249 1216 5283 1231
rect 5323 1216 5357 1231
rect 5175 1197 5193 1216
rect 5193 1197 5209 1216
rect 5249 1197 5261 1216
rect 5261 1197 5283 1216
rect 5323 1197 5329 1216
rect 5329 1197 5357 1216
rect 5397 1197 5431 1231
rect 5472 1216 5506 1231
rect 5547 1216 5581 1231
rect 5622 1216 5656 1231
rect 5697 1216 5731 1231
rect 5772 1216 5806 1231
rect 5847 1216 5881 1231
rect 5922 1216 5956 1231
rect 6164 1216 6198 1231
rect 6239 1230 6273 1250
rect 5472 1197 5499 1216
rect 5499 1197 5506 1216
rect 5547 1197 5567 1216
rect 5567 1197 5581 1216
rect 5622 1197 5635 1216
rect 5635 1197 5656 1216
rect 5697 1197 5703 1216
rect 5703 1197 5731 1216
rect 5772 1197 5805 1216
rect 5805 1197 5806 1216
rect 5847 1197 5873 1216
rect 5873 1197 5881 1216
rect 5922 1197 5941 1216
rect 5941 1197 5956 1216
rect 6164 1197 6165 1216
rect 6165 1197 6198 1216
rect 6355 1346 6389 1380
rect 6355 1274 6389 1308
rect 6355 1202 6389 1236
rect 6867 1346 6901 1380
rect 6867 1274 6901 1308
rect 6867 1202 6901 1236
rect 7379 1346 7413 1380
rect 7379 1274 7413 1308
rect 7379 1202 7413 1236
rect 7891 1346 7925 1380
rect 7891 1274 7925 1308
rect 7891 1202 7925 1236
rect 8403 1346 8437 1380
rect 8403 1274 8437 1308
rect 8403 1202 8437 1236
rect 8915 1346 8949 1380
rect 8915 1274 8949 1308
rect 8915 1202 8949 1236
rect 9267 1346 9301 1380
rect 9267 1274 9301 1308
rect 9267 1202 9301 1236
rect 9619 1346 9653 1380
rect 9619 1274 9653 1308
rect 9619 1202 9653 1236
rect 9971 1346 10005 1380
rect 9971 1274 10005 1308
rect 9971 1202 10005 1236
rect 10088 1316 10091 1342
rect 10091 1316 10122 1342
rect 10088 1308 10122 1316
rect 10088 1248 10091 1270
rect 10091 1248 10122 1270
rect 10088 1236 10122 1248
rect 5027 1125 5061 1159
rect 6239 1155 6273 1189
rect 5200 1094 5208 1128
rect 5208 1094 5234 1128
rect 5272 1094 5276 1128
rect 5276 1094 5306 1128
rect 5344 1094 5378 1128
rect 5416 1094 5446 1128
rect 5446 1094 5450 1128
rect 5488 1094 5514 1128
rect 5514 1094 5522 1128
rect 5560 1094 5582 1128
rect 5582 1094 5594 1128
rect 5632 1094 5650 1128
rect 5650 1094 5666 1128
rect 5704 1094 5718 1128
rect 5718 1094 5738 1128
rect 5776 1094 5786 1128
rect 5786 1094 5810 1128
rect 5848 1094 5854 1128
rect 5854 1094 5882 1128
rect 5920 1094 5922 1128
rect 5922 1094 5954 1128
rect 5027 1045 5061 1079
rect 2757 767 2791 801
rect 2255 596 2289 630
rect 2255 524 2289 558
rect 2964 568 2974 590
rect 2974 568 2998 590
rect 2964 556 2998 568
rect 2964 484 2974 518
rect 2974 484 2998 518
rect 3276 568 3286 590
rect 3286 568 3310 590
rect 3276 556 3310 568
rect 3276 484 3286 518
rect 3286 484 3310 518
rect 2757 387 2791 421
rect 2139 154 2173 188
rect 2139 68 2173 102
rect 2139 -19 2173 15
rect 2385 247 2419 281
rect 2462 247 2496 281
rect 3069 365 3103 399
rect 2757 293 2791 327
rect 2601 188 2635 222
rect 2601 116 2635 150
rect 3381 348 3415 382
rect 3069 293 3103 327
rect 2913 188 2947 222
rect 2913 116 2947 150
rect 3693 348 3727 382
rect 3381 276 3415 310
rect 3225 188 3259 222
rect 3225 116 3259 150
rect 3693 276 3727 310
rect 4901 963 4935 997
rect 4262 391 4296 412
rect 4262 378 4296 391
rect 4262 320 4296 340
rect 4262 306 4296 320
rect 3537 188 3571 222
rect 3537 116 3571 150
rect 3999 188 4033 222
rect 3999 116 4033 150
rect 2609 23 2643 57
rect 2681 23 2691 57
rect 2691 23 2715 57
rect 2753 23 2759 57
rect 2759 23 2787 57
rect 2825 23 2827 57
rect 2827 23 2859 57
rect 2897 23 2929 57
rect 2929 23 2931 57
rect 2969 23 2997 57
rect 2997 23 3003 57
rect 3041 23 3065 57
rect 3065 23 3075 57
rect 3113 23 3133 57
rect 3133 23 3147 57
rect 3185 23 3201 57
rect 3201 23 3219 57
rect 3257 23 3269 57
rect 3269 23 3291 57
rect 3329 23 3337 57
rect 3337 23 3363 57
rect 3401 23 3405 57
rect 3405 23 3435 57
rect 3473 23 3507 57
rect 3545 23 3575 57
rect 3575 23 3579 57
rect 3617 23 3643 57
rect 3643 23 3651 57
rect 3689 23 3711 57
rect 3711 23 3723 57
rect 4901 883 4935 917
rect 5027 965 5061 999
rect 6239 1080 6273 1114
rect 6239 1005 6273 1039
rect 10088 1180 10091 1198
rect 10091 1180 10122 1198
rect 10088 1164 10122 1180
rect 10088 1112 10091 1126
rect 10091 1112 10122 1126
rect 10088 1092 10122 1112
rect 10088 1044 10091 1054
rect 10091 1044 10122 1054
rect 10088 1020 10122 1044
rect 5027 886 5061 920
rect 5143 948 5177 982
rect 5143 864 5177 898
rect 5455 948 5489 982
rect 5455 864 5489 898
rect 6239 930 6273 964
rect 6239 855 6273 889
rect 6611 986 6645 1020
rect 6611 914 6645 948
rect 6611 842 6645 876
rect 7123 986 7157 1020
rect 7123 914 7157 948
rect 7123 842 7157 876
rect 7635 986 7669 1020
rect 7635 914 7669 948
rect 7635 842 7669 876
rect 8147 986 8181 1020
rect 8147 914 8181 948
rect 8147 842 8181 876
rect 8659 986 8693 1020
rect 8659 914 8693 948
rect 8659 842 8693 876
rect 9091 986 9125 1020
rect 9091 914 9125 948
rect 9091 842 9125 876
rect 9443 986 9477 1020
rect 9443 914 9477 948
rect 9443 842 9477 876
rect 9795 986 9829 1020
rect 9795 914 9829 948
rect 9795 842 9829 876
rect 10088 976 10091 982
rect 10091 976 10122 982
rect 10088 948 10122 976
rect 10088 908 10091 910
rect 10091 908 10122 910
rect 10088 876 10122 908
rect 6239 780 6273 814
rect 10088 806 10122 838
rect 10088 804 10091 806
rect 10091 804 10122 806
rect 4389 693 4423 727
rect 4389 613 4423 647
rect 4901 693 4935 727
rect 4901 613 4935 647
rect 5967 657 6001 691
rect 6039 657 6073 691
rect 4645 492 4679 526
rect 4645 402 4679 436
rect 5299 546 5333 580
rect 5299 474 5333 508
rect 5299 402 5333 436
rect 5611 546 5645 580
rect 5611 474 5645 508
rect 5611 402 5645 436
rect 4540 313 4566 347
rect 4566 313 4574 347
rect 2373 -67 2407 -33
rect 2445 -67 2479 -33
rect 1146 -162 1180 -128
rect 1218 -162 1224 -128
rect 1224 -162 1252 -128
rect 1290 -162 1292 -128
rect 1292 -162 1324 -128
rect 1362 -162 1394 -128
rect 1394 -162 1396 -128
rect 1434 -162 1462 -128
rect 1462 -162 1468 -128
rect 1506 -162 1530 -128
rect 1530 -162 1540 -128
rect 1578 -162 1598 -128
rect 1598 -162 1612 -128
rect 1650 -162 1666 -128
rect 1666 -162 1684 -128
rect 1722 -162 1734 -128
rect 1734 -162 1756 -128
rect 1794 -162 1802 -128
rect 1802 -162 1828 -128
rect 1866 -162 1870 -128
rect 1870 -162 1900 -128
rect 1938 -162 1972 -128
rect 2010 -162 2040 -128
rect 2040 -162 2044 -128
rect 2082 -162 2108 -128
rect 2108 -162 2116 -128
rect 4747 313 4781 347
rect 4819 313 4845 347
rect 4845 313 4853 347
rect 6414 694 6416 728
rect 6416 694 6448 728
rect 6493 694 6519 728
rect 6519 694 6527 728
rect 6572 694 6588 728
rect 6588 694 6606 728
rect 6651 694 6657 728
rect 6657 694 6685 728
rect 6731 694 6761 728
rect 6761 694 6765 728
rect 6811 694 6830 728
rect 6830 694 6845 728
rect 6891 694 6899 728
rect 6899 694 6925 728
rect 6971 694 7002 728
rect 7002 694 7005 728
rect 7051 694 7071 728
rect 7071 694 7085 728
rect 7131 694 7140 728
rect 7140 694 7165 728
rect 7514 694 7524 728
rect 7524 694 7548 728
rect 7590 694 7594 728
rect 7594 694 7624 728
rect 7666 694 7698 728
rect 7698 694 7700 728
rect 7742 694 7768 728
rect 7768 694 7776 728
rect 7818 694 7838 728
rect 7838 694 7852 728
rect 7894 694 7908 728
rect 7908 694 7928 728
rect 7971 694 7978 728
rect 7978 694 8005 728
rect 8048 694 8082 728
rect 8125 694 8154 728
rect 8154 694 8159 728
rect 8202 694 8224 728
rect 8224 694 8236 728
rect 8279 694 8294 728
rect 8294 694 8313 728
rect 8356 694 8364 728
rect 8364 694 8390 728
rect 9570 694 9584 728
rect 9584 694 9604 728
rect 9658 694 9692 728
rect 9747 694 9766 728
rect 9766 694 9781 728
rect 9836 694 9838 728
rect 9838 694 9870 728
rect 9925 694 9944 728
rect 9944 694 9959 728
rect 10088 738 10122 766
rect 10088 732 10091 738
rect 10091 732 10122 738
rect 10088 670 10122 694
rect 10088 660 10091 670
rect 10091 660 10122 670
rect 10088 602 10122 622
rect 10088 588 10091 602
rect 10091 588 10122 602
rect 6123 546 6157 580
rect 6123 474 6157 508
rect 6123 402 6157 436
rect 6611 546 6645 580
rect 6611 474 6645 508
rect 6611 402 6645 436
rect 7123 546 7157 580
rect 7123 474 7157 508
rect 7123 402 7157 436
rect 7635 546 7669 580
rect 7635 474 7669 508
rect 7635 402 7669 436
rect 8147 546 8181 580
rect 8147 474 8181 508
rect 8147 402 8181 436
rect 8659 546 8693 580
rect 8659 474 8693 508
rect 8659 402 8693 436
rect 9091 546 9125 580
rect 9091 474 9125 508
rect 9091 402 9125 436
rect 9443 546 9477 580
rect 9443 474 9477 508
rect 9443 402 9477 436
rect 9795 546 9829 580
rect 9795 474 9829 508
rect 9795 402 9829 436
rect 10088 534 10122 550
rect 10088 516 10091 534
rect 10091 516 10122 534
rect 10088 466 10122 478
rect 10088 444 10091 466
rect 10091 444 10122 466
rect 5143 290 5177 324
rect 5143 218 5177 252
rect 4909 111 4943 145
rect 4909 17 4943 51
rect 5027 139 5061 173
rect 5143 146 5177 180
rect 5455 290 5489 324
rect 5967 292 6001 326
rect 6039 292 6073 326
rect 10088 398 10122 406
rect 10088 372 10091 398
rect 10091 372 10122 398
rect 10088 330 10122 334
rect 10088 300 10091 330
rect 10091 300 10122 330
rect 5455 218 5489 252
rect 10088 228 10091 262
rect 10091 228 10122 262
rect 5455 146 5489 180
rect 5867 186 5901 220
rect 5027 38 5061 72
rect 5867 114 5901 148
rect 5867 42 5901 76
rect 6355 186 6389 220
rect 6355 114 6389 148
rect 6355 42 6389 76
rect 6867 186 6901 220
rect 6867 114 6901 148
rect 6867 42 6901 76
rect 7379 186 7413 220
rect 7379 114 7413 148
rect 7379 42 7413 76
rect 7891 186 7925 220
rect 7891 114 7925 148
rect 7891 42 7925 76
rect 8403 186 8437 220
rect 8403 114 8437 148
rect 8403 42 8437 76
rect 8915 186 8949 220
rect 8915 114 8949 148
rect 8915 42 8949 76
rect 9267 186 9301 220
rect 9267 114 9301 148
rect 9267 42 9301 76
rect 9619 186 9653 220
rect 9619 114 9653 148
rect 9619 42 9653 76
rect 9971 186 10005 220
rect 9971 114 10005 148
rect 9971 42 10005 76
rect 10088 160 10091 190
rect 10091 160 10122 190
rect 10088 156 10122 160
rect 10088 92 10091 117
rect 10091 92 10122 117
rect 10088 83 10122 92
rect 10088 10 10122 44
rect 5099 -62 5105 -28
rect 5105 -62 5133 -28
rect 5172 -62 5173 -28
rect 5173 -62 5206 -28
rect 5245 -62 5275 -28
rect 5275 -62 5279 -28
rect 5318 -62 5343 -28
rect 5343 -62 5352 -28
rect 5391 -62 5411 -28
rect 5411 -62 5425 -28
rect 5464 -62 5479 -28
rect 5479 -62 5498 -28
rect 5537 -62 5547 -28
rect 5547 -62 5571 -28
rect 5610 -62 5615 -28
rect 5615 -62 5644 -28
rect 5683 -62 5717 -28
rect 5755 -62 5785 -28
rect 5785 -62 5789 -28
rect 5827 -62 5853 -28
rect 5853 -62 5861 -28
rect 5899 -62 5921 -28
rect 5921 -62 5933 -28
rect 5971 -62 5989 -28
rect 5989 -62 6005 -28
rect 6043 -62 6057 -28
rect 6057 -62 6077 -28
rect 6115 -62 6125 -28
rect 6125 -62 6149 -28
rect 6187 -62 6193 -28
rect 6193 -62 6221 -28
rect 6311 -62 6319 -28
rect 6319 -62 6345 -28
rect 6384 -62 6387 -28
rect 6387 -62 6418 -28
rect 6457 -62 6489 -28
rect 6489 -62 6491 -28
rect 6530 -62 6557 -28
rect 6557 -62 6564 -28
rect 6603 -62 6625 -28
rect 6625 -62 6637 -28
rect 6676 -62 6693 -28
rect 6693 -62 6710 -28
rect 6749 -62 6761 -28
rect 6761 -62 6783 -28
rect 6822 -62 6829 -28
rect 6829 -62 6856 -28
rect 6895 -62 6897 -28
rect 6897 -62 6929 -28
rect 6968 -62 6999 -28
rect 6999 -62 7002 -28
rect 7041 -62 7067 -28
rect 7067 -62 7075 -28
rect 7114 -62 7135 -28
rect 7135 -62 7148 -28
rect 7187 -62 7203 -28
rect 7203 -62 7221 -28
rect 7260 -62 7271 -28
rect 7271 -62 7294 -28
rect 7333 -62 7339 -28
rect 7339 -62 7367 -28
rect 7406 -62 7407 -28
rect 7407 -62 7440 -28
rect 7479 -62 7509 -28
rect 7509 -62 7513 -28
rect 7552 -62 7577 -28
rect 7577 -62 7586 -28
rect 7625 -62 7645 -28
rect 7645 -62 7659 -28
rect 7698 -62 7713 -28
rect 7713 -62 7732 -28
rect 7771 -62 7781 -28
rect 7781 -62 7805 -28
rect 7844 -62 7849 -28
rect 7849 -62 7878 -28
rect 7917 -62 7951 -28
rect 7990 -62 8019 -28
rect 8019 -62 8024 -28
rect 8063 -62 8087 -28
rect 8087 -62 8097 -28
rect 8136 -62 8170 -28
rect 8209 -62 8243 -28
rect 8282 -62 8316 -28
rect 8355 -62 8389 -28
rect 8428 -62 8462 -28
rect 8501 -62 8535 -28
rect 8574 -62 8608 -28
rect 8647 -62 8681 -28
rect 8720 -62 8754 -28
rect 8792 -62 8826 -28
rect 8864 -62 8898 -28
rect 8936 -62 8970 -28
rect 9008 -62 9042 -28
rect 9080 -62 9114 -28
rect 9152 -62 9186 -28
rect 9224 -62 9258 -28
rect 9296 -62 9330 -28
rect 9368 -62 9402 -28
rect 9440 -62 9474 -28
rect 9512 -62 9546 -28
rect 9584 -62 9618 -28
rect 9656 -62 9690 -28
rect 9728 -62 9762 -28
rect 9800 -62 9834 -28
rect 9872 -62 9906 -28
rect 9944 -62 9978 -28
rect 10016 -62 10050 -28
rect 80 -202 88 -168
rect 88 -202 114 -168
rect 152 -202 156 -168
rect 156 -202 186 -168
rect 224 -202 258 -168
rect 296 -202 326 -168
rect 326 -202 330 -168
rect 368 -202 394 -168
rect 394 -202 402 -168
rect 440 -202 462 -168
rect 462 -202 474 -168
rect 512 -202 530 -168
rect 530 -202 546 -168
rect 584 -202 598 -168
rect 598 -202 618 -168
rect 656 -202 666 -168
rect 666 -202 690 -168
rect 728 -202 734 -168
rect 734 -202 762 -168
rect 800 -202 802 -168
rect 802 -202 834 -168
rect 703 -289 737 -255
rect 778 -289 812 -255
rect 853 -289 887 -255
rect 928 -289 962 -255
rect 1003 -289 1037 -255
rect 1077 -289 1111 -255
rect 1151 -289 1185 -255
rect 1257 -468 1291 -434
rect 1329 -468 1363 -434
rect -303 -631 -269 -597
rect -231 -631 -197 -597
<< metal1 >>
tri 6950 3543 6988 3581 se
rect 6988 3575 7040 3581
tri 6067 3469 6141 3543 se
rect 6141 3523 6988 3543
rect 6141 3511 7040 3523
rect 6141 3491 6988 3511
tri 6141 3469 6163 3491 nw
tri 6950 3469 6972 3491 ne
rect 6972 3469 6988 3491
tri 6032 3434 6067 3469 se
rect 5372 3428 5424 3434
tri 5997 3399 6032 3434 se
rect 6032 3399 6067 3434
rect 5372 3364 5424 3376
tri 5424 3358 5465 3399 sw
tri 5993 3395 5997 3399 se
rect 5997 3395 6067 3399
tri 6067 3395 6141 3469 nw
tri 6972 3453 6988 3469 ne
rect 6988 3453 7040 3459
tri 5956 3358 5993 3395 se
rect 5993 3358 6030 3395
tri 6030 3358 6067 3395 nw
rect 5424 3312 5978 3358
rect 5372 3306 5978 3312
tri 5978 3306 6030 3358 nw
rect 7520 2859 7526 2911
rect 7578 2859 7642 2911
rect 7694 2905 9505 2911
rect 7694 2871 8893 2905
rect 8927 2871 8974 2905
rect 9008 2871 9055 2905
rect 9089 2871 9136 2905
rect 9170 2871 9217 2905
rect 9251 2871 9298 2905
rect 9332 2871 9379 2905
rect 9413 2871 9459 2905
rect 9493 2871 9505 2905
rect 7694 2865 9505 2871
rect 7694 2859 7700 2865
tri 7700 2859 7706 2865 nw
rect 9120 2797 9312 2803
rect 9120 2788 9260 2797
rect 9120 2754 9132 2788
rect 9166 2754 9226 2788
rect 9120 2745 9260 2754
rect 8799 2677 8857 2743
rect 8799 2643 8811 2677
rect 8845 2643 8857 2677
rect 9120 2719 9312 2745
rect 9120 2667 9260 2719
rect 8799 2605 8857 2643
rect 8799 2571 8811 2605
rect 8845 2571 8857 2605
tri 8771 2533 8799 2561 se
rect 8799 2533 8857 2571
rect 8895 2632 9047 2647
rect 8895 2598 8907 2632
rect 8941 2598 9001 2632
rect 9035 2598 9047 2632
rect 8895 2583 9047 2598
tri 8895 2539 8939 2583 ne
tri 8740 2502 8771 2533 se
rect 8771 2502 8811 2533
rect 8668 2499 8811 2502
rect 8845 2499 8857 2533
rect 8668 2450 8857 2499
rect 8668 2441 8769 2450
tri 8769 2441 8778 2450 nw
rect 7151 2369 8497 2375
rect 7203 2323 8497 2369
rect 8549 2323 8561 2375
rect 8613 2323 8619 2375
rect 7151 2305 7203 2317
rect 7151 2247 7203 2253
tri 7203 2247 7279 2323 nw
tri 8637 2002 8668 2033 se
rect 8668 2011 8720 2441
tri 8720 2392 8769 2441 nw
tri 8899 2392 8939 2432 se
rect 8939 2406 9003 2583
tri 9003 2539 9047 2583 nw
rect 9120 2641 9312 2667
rect 9120 2589 9260 2641
rect 9120 2563 9312 2589
rect 9120 2511 9260 2563
rect 9120 2484 9312 2511
rect 9120 2475 9260 2484
rect 9120 2441 9132 2475
rect 9166 2441 9226 2475
rect 9120 2432 9260 2441
rect 9120 2426 9312 2432
rect 8939 2392 8972 2406
tri 8882 2375 8899 2392 se
rect 8899 2375 8972 2392
tri 8972 2375 9003 2406 nw
rect 8762 2323 8768 2375
rect 8820 2323 8832 2375
rect 8884 2323 8920 2375
tri 8920 2323 8972 2375 nw
rect 8763 2167 8769 2219
rect 8821 2167 8833 2219
rect 8885 2213 9209 2219
rect 8885 2179 8910 2213
rect 8944 2179 8995 2213
rect 9029 2179 9079 2213
rect 9113 2179 9163 2213
rect 9197 2179 9209 2213
rect 8885 2173 9209 2179
rect 8885 2167 8891 2173
tri 8891 2167 8897 2173 nw
rect 8668 2002 8711 2011
tri 8711 2002 8720 2011 nw
rect 8799 2074 8845 2086
rect 8799 2040 8805 2074
rect 8839 2040 8845 2074
rect 8799 2002 8845 2040
tri 8603 1968 8637 2002 se
rect 8637 1968 8677 2002
tri 8677 1968 8711 2002 nw
rect 8799 1968 8805 2002
rect 8839 1968 8845 2002
tri 8594 1959 8603 1968 se
rect 8603 1959 8668 1968
tri 8668 1959 8677 1968 nw
tri 8592 1957 8594 1959 se
rect 8594 1957 8666 1959
tri 8666 1957 8668 1959 nw
tri 8798 1957 8799 1958 se
rect 8799 1957 8845 1968
tri 8588 1953 8592 1957 se
rect 8592 1953 8632 1957
tri 7114 1923 7144 1953 se
rect 7144 1923 8632 1953
tri 8632 1923 8666 1957 nw
tri 8764 1923 8798 1957 se
rect 8798 1938 8845 1957
rect 8798 1923 8830 1938
tri 8830 1923 8845 1938 nw
rect 9137 2040 9585 2046
rect 9137 1988 9456 2040
rect 9508 1988 9532 2040
rect 9584 1988 9585 2040
rect 9137 1972 9585 1988
rect 9137 1957 9456 1972
rect 9137 1923 9152 1957
rect 9186 1923 9252 1957
rect 9286 1923 9351 1957
rect 9385 1923 9456 1957
tri 7070 1879 7114 1923 se
rect 7114 1901 8610 1923
tri 8610 1901 8632 1923 nw
tri 8742 1901 8764 1923 se
rect 8764 1901 8799 1923
rect 7114 1879 7144 1901
tri 7144 1879 7166 1901 nw
tri 8733 1892 8742 1901 se
rect 8742 1892 8799 1901
tri 8799 1892 8830 1923 nw
rect 9137 1920 9456 1923
rect 9508 1920 9532 1972
rect 9584 1920 9585 1972
rect 9137 1914 9585 1920
tri 8720 1879 8733 1892 se
rect 8733 1879 8763 1892
tri 6996 1805 7070 1879 se
tri 7070 1805 7144 1879 nw
tri 8697 1856 8720 1879 se
rect 8720 1856 8763 1879
tri 8763 1856 8799 1892 nw
tri 7151 1805 7202 1856 se
rect 7202 1810 8717 1856
tri 8717 1810 8763 1856 nw
tri 6985 1794 6996 1805 se
rect 6996 1794 7007 1805
tri 4506 1738 4562 1794 se
rect 4562 1742 7007 1794
tri 7007 1742 7070 1805 nw
tri 7136 1790 7151 1805 se
rect 7151 1790 7202 1805
tri 7202 1790 7222 1810 nw
tri 7088 1742 7136 1790 se
rect 4562 1738 4571 1742
rect 2129 1732 2181 1738
tri 4497 1729 4506 1738 se
rect 4506 1729 4571 1738
tri 4571 1729 4584 1742 nw
tri 7075 1729 7088 1742 se
rect 7088 1729 7136 1742
tri 2181 1686 2185 1690 sw
rect 2181 1680 2185 1686
rect 2129 1674 2185 1680
tri 2185 1674 2197 1686 sw
rect 4164 1677 4170 1729
rect 4222 1677 4234 1729
rect 4286 1720 4550 1729
rect 4310 1686 4375 1720
rect 4409 1686 4474 1720
rect 4508 1708 4550 1720
tri 4550 1708 4571 1729 nw
tri 7070 1724 7075 1729 se
rect 7075 1724 7136 1729
tri 7136 1724 7202 1790 nw
tri 7060 1714 7070 1724 se
rect 7070 1714 7080 1724
rect 4603 1708 7080 1714
rect 4508 1686 4520 1708
rect 4286 1677 4520 1686
tri 4520 1678 4550 1708 nw
rect 4603 1674 4615 1708
rect 4649 1674 4687 1708
rect 4721 1674 7080 1708
rect 2129 1668 2197 1674
rect 1382 1612 1667 1618
rect 1382 1578 1394 1612
rect 1428 1578 1470 1612
rect 1504 1578 1546 1612
rect 1580 1578 1621 1612
rect 1655 1578 1667 1612
rect 2181 1638 2197 1668
tri 2197 1638 2233 1674 sw
rect 4603 1668 7080 1674
tri 7080 1668 7136 1724 nw
tri 7409 1638 7425 1654 se
rect 7425 1648 7477 1654
rect 2181 1616 7425 1638
rect 2129 1610 7425 1616
tri 7393 1578 7425 1610 ne
tri 7477 1638 7493 1654 sw
tri 9800 1638 9811 1649 se
rect 9811 1643 9863 1649
rect 7477 1610 9811 1638
rect 7425 1584 7477 1596
rect 512 1302 1131 1314
rect 512 1268 543 1302
rect 577 1268 759 1302
rect 793 1297 1131 1302
rect 793 1268 1091 1297
rect 512 1263 1091 1268
rect 1125 1263 1131 1297
rect 512 1197 1131 1263
rect 512 1163 543 1197
rect 577 1163 759 1197
rect 793 1163 1091 1197
rect 1125 1163 1131 1197
rect 512 1151 1131 1163
rect 1382 1180 1667 1578
rect 4836 1572 5721 1578
rect 4836 1538 4848 1572
rect 4882 1538 4924 1572
rect 4958 1538 5000 1572
rect 5034 1538 5075 1572
rect 5109 1538 5150 1572
rect 5184 1538 5225 1572
rect 5259 1538 5300 1572
rect 5334 1538 5375 1572
rect 5409 1538 5450 1572
rect 5484 1538 5525 1572
rect 5559 1538 5600 1572
rect 5634 1538 5675 1572
rect 5709 1538 5721 1572
rect 4836 1532 5721 1538
rect 5782 1572 5951 1578
rect 5782 1538 5794 1572
rect 5828 1538 5905 1572
rect 5939 1538 5951 1572
rect 5782 1532 5951 1538
tri 6049 1532 6095 1578 se
rect 6095 1532 7074 1578
tri 5770 1506 5782 1518 se
rect 5782 1506 5889 1532
rect 2253 1500 4610 1506
rect 2253 1491 4433 1500
rect 2253 1457 2345 1491
rect 2379 1457 2417 1491
rect 2451 1457 2489 1491
rect 2523 1457 2561 1491
rect 2595 1457 2633 1491
rect 2667 1457 2705 1491
rect 2739 1457 2777 1491
rect 2811 1457 2849 1491
rect 2883 1457 2921 1491
rect 2955 1457 2993 1491
rect 3027 1457 3065 1491
rect 3099 1457 3137 1491
rect 3171 1457 3209 1491
rect 3243 1457 3281 1491
rect 3315 1457 3353 1491
rect 3387 1457 3425 1491
rect 3459 1457 3497 1491
rect 3531 1457 3569 1491
rect 3603 1457 3641 1491
rect 3675 1457 4433 1491
rect 2253 1448 4433 1457
rect 4485 1448 4557 1500
rect 4609 1448 4610 1500
tri 5750 1486 5770 1506 se
rect 5770 1486 5889 1506
tri 5889 1488 5933 1532 nw
tri 6029 1512 6049 1532 se
rect 6049 1512 6095 1532
tri 6095 1512 6115 1532 nw
tri 7062 1526 7068 1532 ne
rect 7068 1526 7074 1532
rect 7126 1526 7158 1578
rect 7210 1526 7242 1578
rect 7294 1526 7326 1578
rect 7378 1526 7384 1578
tri 7477 1578 7509 1610 nw
tri 9764 1578 9796 1610 ne
rect 9796 1591 9811 1610
rect 9796 1579 9863 1591
rect 9796 1578 9811 1579
tri 9796 1563 9811 1578 ne
rect 7425 1526 7477 1532
rect 9811 1521 9863 1527
tri 6005 1488 6029 1512 se
rect 6029 1488 6069 1512
tri 6003 1486 6005 1488 se
rect 6005 1486 6069 1488
tri 6069 1486 6095 1512 nw
rect 6233 1486 10128 1492
tri 5746 1482 5750 1486 se
rect 5750 1482 5889 1486
rect 2253 1424 4610 1448
rect 1382 1146 1394 1180
rect 1428 1146 1470 1180
rect 1504 1146 1546 1180
rect 1580 1146 1621 1180
rect 1655 1146 1667 1180
rect 1382 1140 1667 1146
rect 1888 1396 2092 1402
rect 1888 1362 1900 1396
rect 1934 1362 1973 1396
rect 2007 1362 2046 1396
rect 2080 1362 2092 1396
rect -121 1074 1568 1080
rect -121 1068 1376 1074
rect -121 1034 -115 1068
rect -81 1034 220 1068
rect 254 1034 652 1068
rect 686 1034 1376 1068
rect -121 1022 1376 1034
rect 1428 1022 1446 1074
rect 1498 1022 1516 1074
rect 1888 1039 2092 1362
rect 2253 1399 4433 1424
rect 2253 1365 2321 1399
rect 2355 1365 2633 1399
rect 2667 1365 2913 1399
rect 2947 1365 3225 1399
rect 3259 1365 3537 1399
rect 3571 1372 4433 1399
rect 4485 1372 4557 1424
rect 4609 1372 4610 1424
rect 4778 1467 5889 1482
rect 4778 1433 4790 1467
rect 4824 1433 4884 1467
rect 4918 1433 5215 1467
rect 5249 1433 5309 1467
rect 5343 1433 5737 1467
rect 5771 1433 5831 1467
rect 5865 1433 5889 1467
tri 5969 1452 6003 1486 se
rect 6003 1452 6035 1486
tri 6035 1452 6069 1486 nw
rect 6233 1452 6312 1486
rect 6346 1452 6385 1486
rect 6419 1452 6458 1486
rect 6492 1452 6531 1486
rect 6565 1452 6604 1486
rect 6638 1452 6677 1486
rect 6711 1452 6750 1486
rect 6784 1452 6823 1486
rect 6857 1452 6896 1486
rect 6930 1452 6969 1486
rect 7003 1452 7042 1486
rect 7076 1452 7115 1486
rect 7149 1452 7188 1486
rect 7222 1452 7261 1486
rect 7295 1452 7334 1486
rect 7368 1452 7407 1486
rect 7441 1452 7480 1486
rect 7514 1452 7553 1486
rect 7587 1452 7626 1486
rect 7660 1452 7699 1486
rect 7733 1452 7772 1486
rect 7806 1452 7845 1486
rect 7879 1452 7918 1486
rect 7952 1452 7991 1486
rect 8025 1452 8064 1486
rect 8098 1452 8137 1486
rect 8171 1452 8210 1486
rect 8244 1452 8283 1486
rect 8317 1452 8356 1486
rect 8390 1452 8429 1486
rect 8463 1452 8502 1486
rect 8536 1452 8575 1486
rect 8609 1452 8648 1486
rect 8682 1452 8721 1486
rect 8755 1452 8794 1486
rect 8828 1452 8867 1486
rect 8901 1452 8940 1486
rect 8974 1452 9013 1486
rect 9047 1452 9086 1486
rect 9120 1452 9159 1486
rect 9193 1452 9232 1486
rect 9266 1452 9305 1486
rect 9339 1452 9378 1486
rect 9412 1452 9451 1486
rect 9485 1452 9524 1486
rect 9558 1452 9597 1486
rect 9631 1452 9670 1486
rect 9704 1452 9743 1486
rect 9777 1452 9816 1486
rect 9850 1452 9889 1486
rect 9923 1452 9982 1486
rect 10016 1452 10128 1486
tri 5963 1446 5969 1452 se
rect 5969 1446 6029 1452
tri 6029 1446 6035 1452 nw
rect 6233 1446 10128 1452
rect 4778 1418 5889 1433
tri 5935 1418 5963 1446 se
rect 5963 1418 5997 1446
tri 5931 1414 5935 1418 se
rect 5935 1414 5997 1418
tri 5997 1414 6029 1446 nw
rect 6233 1414 6298 1446
tri 6298 1414 6330 1446 nw
tri 10034 1414 10066 1446 ne
rect 10066 1414 10128 1446
tri 5897 1380 5931 1414 se
rect 5931 1380 5963 1414
tri 5963 1380 5997 1414 nw
rect 6233 1380 6239 1414
rect 6273 1380 6279 1414
tri 6279 1395 6298 1414 nw
tri 10066 1398 10082 1414 ne
rect 3571 1365 4610 1372
tri 5888 1371 5897 1380 se
rect 5897 1371 5929 1380
rect 2253 1348 4610 1365
rect 5566 1365 5929 1371
rect 2253 1318 4433 1348
rect 2253 1284 2321 1318
rect 2355 1284 2633 1318
rect 2667 1284 2913 1318
rect 2947 1284 3225 1318
rect 3259 1284 3537 1318
rect 3571 1296 4433 1318
rect 4485 1296 4557 1348
rect 4609 1296 4610 1348
rect 3571 1289 4610 1296
rect 4967 1349 5532 1355
rect 4967 1340 5361 1349
rect 5413 1340 5425 1349
rect 5477 1340 5532 1349
rect 4967 1306 4979 1340
rect 5013 1306 5073 1340
rect 5107 1306 5361 1340
rect 5477 1306 5486 1340
rect 5520 1306 5532 1340
rect 5566 1331 5578 1365
rect 5612 1331 5650 1365
rect 5684 1346 5929 1365
tri 5929 1346 5963 1380 nw
rect 5684 1342 5925 1346
tri 5925 1342 5929 1346 nw
rect 5684 1339 5922 1342
tri 5922 1339 5925 1342 nw
rect 6233 1339 6279 1380
rect 5684 1331 5908 1339
rect 5566 1325 5908 1331
tri 5908 1325 5922 1339 nw
tri 6228 1325 6233 1330 se
rect 6233 1325 6239 1339
tri 6223 1320 6228 1325 se
rect 6228 1320 6239 1325
rect 4967 1297 5361 1306
rect 5413 1297 5425 1306
rect 5477 1297 5532 1306
rect 4967 1291 5532 1297
rect 5958 1314 6088 1320
rect 3571 1284 4203 1289
rect 2253 1250 3999 1284
rect 4033 1280 4203 1284
tri 4203 1280 4212 1289 nw
rect 5958 1280 5970 1314
rect 6004 1280 6042 1314
rect 6076 1280 6088 1314
tri 6208 1305 6223 1320 se
rect 6223 1305 6239 1320
rect 6273 1305 6279 1339
rect 4033 1274 4197 1280
tri 4197 1274 4203 1280 nw
rect 5958 1274 6088 1280
tri 6177 1274 6208 1305 se
rect 6208 1274 6279 1305
rect 4033 1270 4193 1274
tri 4193 1270 4197 1274 nw
tri 5972 1270 5976 1274 ne
rect 5976 1270 6084 1274
tri 6084 1270 6088 1274 nw
tri 6173 1270 6177 1274 se
rect 6177 1270 6279 1274
rect 4033 1264 4187 1270
tri 4187 1264 4193 1270 nw
tri 5976 1264 5982 1270 ne
rect 5982 1264 6078 1270
tri 6078 1264 6084 1270 nw
tri 6167 1264 6173 1270 se
rect 6173 1264 6279 1270
rect 4033 1250 4172 1264
rect 2253 1249 4172 1250
tri 4172 1249 4187 1264 nw
tri 5982 1255 5991 1264 ne
rect 5991 1255 6045 1264
rect 4337 1249 4843 1255
rect 2253 1237 4138 1249
rect 2253 1203 2321 1237
rect 2355 1203 2633 1237
rect 2667 1203 2913 1237
rect 2947 1203 3225 1237
rect 3259 1203 3537 1237
rect 3571 1215 4138 1237
tri 4138 1215 4172 1249 nw
rect 4337 1215 4349 1249
rect 4383 1215 4421 1249
rect 4455 1231 4843 1249
tri 4843 1231 4867 1255 sw
tri 5991 1249 5997 1255 ne
rect 5021 1231 5968 1237
rect 4455 1223 4867 1231
tri 4867 1223 4875 1231 sw
rect 4455 1215 4875 1223
rect 3571 1212 4120 1215
rect 3571 1203 3999 1212
rect 2253 1182 3999 1203
tri 3569 1178 3573 1182 ne
rect 3573 1178 3999 1182
rect 4033 1197 4120 1212
tri 4120 1197 4138 1215 nw
rect 4337 1209 4875 1215
tri 4823 1197 4835 1209 ne
rect 4835 1197 4875 1209
tri 4875 1197 4901 1223 sw
rect 5021 1197 5101 1231
rect 5135 1197 5175 1231
rect 5209 1197 5249 1231
rect 5283 1197 5323 1231
rect 5357 1197 5397 1231
rect 5431 1197 5472 1231
rect 5506 1197 5547 1231
rect 5581 1197 5622 1231
rect 5656 1197 5697 1231
rect 5731 1197 5772 1231
rect 5806 1197 5847 1231
rect 5881 1197 5922 1231
rect 5956 1197 5968 1231
rect 4033 1189 4112 1197
tri 4112 1189 4120 1197 nw
tri 4835 1189 4843 1197 ne
rect 4843 1189 4901 1197
tri 4901 1189 4909 1197 sw
rect 5021 1191 5968 1197
rect 5997 1231 6045 1255
tri 6045 1231 6078 1264 nw
tri 6140 1237 6167 1264 se
rect 6167 1237 6239 1264
rect 6110 1231 6239 1237
rect 5021 1189 5125 1191
tri 5125 1189 5127 1191 nw
rect 4033 1178 4088 1189
tri 3573 1165 3586 1178 ne
rect 3586 1165 4088 1178
tri 4088 1165 4112 1189 nw
tri 4843 1165 4867 1189 ne
rect 4867 1165 4909 1189
tri 4867 1159 4873 1165 ne
rect 4873 1159 4909 1165
tri 4909 1159 4939 1189 sw
rect 5021 1159 5091 1189
tri 4873 1157 4875 1159 ne
rect 4875 1157 4939 1159
tri 4939 1157 4941 1159 sw
tri 4875 1137 4895 1157 ne
tri 2392 1095 2406 1109 se
rect 2406 1095 4863 1109
tri 2358 1061 2392 1095 se
rect 2392 1061 4745 1095
rect 4779 1061 4817 1095
rect 4851 1061 4863 1095
tri 2342 1045 2358 1061 se
rect 2358 1045 4863 1061
tri 2341 1044 2342 1045 se
rect 2342 1044 2426 1045
tri 2092 1039 2097 1044 sw
tri 2336 1039 2341 1044 se
rect 2341 1039 2426 1044
tri 2426 1039 2432 1045 nw
rect -121 1009 1568 1022
rect -121 979 1376 1009
rect -121 945 -115 979
rect -81 945 220 979
rect 254 945 652 979
rect 686 957 1376 979
rect 1428 957 1446 1009
rect 1498 957 1516 1009
tri 1869 1005 1888 1024 se
rect 1888 1005 2097 1039
tri 2097 1005 2131 1039 sw
tri 2316 1019 2336 1039 se
rect 2336 1019 2406 1039
tri 2406 1019 2426 1039 nw
tri 2302 1005 2316 1019 se
rect 2316 1005 2392 1019
tri 2392 1005 2406 1019 nw
tri 1863 999 1869 1005 se
rect 1869 999 2131 1005
tri 2131 999 2137 1005 sw
tri 2296 999 2302 1005 se
rect 2302 999 2386 1005
tri 2386 999 2392 1005 nw
tri 2481 999 2484 1002 se
rect 2484 999 4706 1002
tri 4706 999 4709 1002 sw
tri 1861 997 1863 999 se
rect 1863 997 2137 999
tri 2137 997 2139 999 sw
tri 2294 997 2296 999 se
rect 2296 997 2384 999
tri 2384 997 2386 999 nw
tri 2479 997 2481 999 se
rect 2481 997 4709 999
tri 4709 997 4711 999 sw
rect 4895 997 4941 1157
tri 1827 963 1861 997 se
rect 1861 963 2139 997
tri 2139 963 2173 997 sw
tri 2286 989 2294 997 se
rect 2294 989 2350 997
rect 686 945 1568 957
rect -121 944 1568 945
rect -121 892 1376 944
rect 1428 892 1446 944
rect 1498 892 1516 944
rect -121 890 1568 892
rect -121 856 -115 890
rect -81 856 220 890
rect 254 856 652 890
rect 686 879 1568 890
rect 686 856 1376 879
rect -121 827 1376 856
rect 1428 827 1446 879
rect 1498 827 1516 879
rect -121 814 1568 827
rect -121 801 1376 814
rect -121 767 -115 801
rect -81 767 220 801
rect 254 767 652 801
rect 686 767 1376 801
rect -121 762 1376 767
rect 1428 762 1446 814
rect 1498 762 1516 814
tri 1812 948 1827 963 se
rect 1827 948 2173 963
tri 2173 948 2188 963 sw
rect 1812 936 2188 948
rect 1812 902 1827 936
rect 1861 902 2139 936
rect 2173 902 2188 936
rect 1812 842 2188 902
rect 1812 808 1827 842
rect 1861 808 2139 842
rect 2173 808 2188 842
rect 1812 796 2188 808
tri 2284 802 2286 804 se
rect 2286 802 2350 989
tri 2350 963 2384 997 nw
tri 2445 963 2479 997 se
rect 2479 969 4711 997
tri 4711 969 4739 997 sw
rect 2479 963 4739 969
tri 4739 963 4745 969 sw
rect 4895 963 4901 997
rect 4935 963 4941 997
tri 2430 948 2445 963 se
rect 2445 950 4745 963
rect 2445 948 2504 950
tri 2504 948 2506 950 nw
tri 4684 948 4686 950 ne
rect 4686 948 4745 950
tri 4745 948 4760 963 sw
tri 2283 801 2284 802 se
rect 2284 801 2350 802
tri 2278 796 2283 801 se
rect 2283 796 2350 801
tri 2249 767 2278 796 se
rect 2278 778 2350 796
rect 2278 767 2339 778
tri 2339 767 2350 778 nw
tri 2414 932 2430 948 se
rect 2430 932 2488 948
tri 2488 932 2504 948 nw
tri 4686 932 4702 948 ne
rect 4702 932 4760 948
rect 2414 930 2486 932
tri 2486 930 2488 932 nw
tri 4702 930 4704 932 ne
rect 4704 930 4760 932
tri 4760 930 4778 948 sw
rect 2414 920 2476 930
tri 2476 920 2486 930 nw
tri 4704 922 4712 930 ne
rect 4712 922 4778 930
tri 4208 920 4210 922 se
rect 4210 920 4262 922
tri 4712 920 4714 922 ne
rect 4714 920 4778 922
tri 4778 920 4788 930 sw
rect 2414 917 2473 920
tri 2473 917 2476 920 nw
tri 2248 766 2249 767 se
rect 2249 766 2338 767
tri 2338 766 2339 767 nw
rect -121 755 1568 762
tri 2237 755 2248 766 se
rect 2248 755 2320 766
tri 2230 748 2237 755 se
rect 2237 748 2320 755
tri 2320 748 2338 766 nw
rect 1968 736 2304 748
rect 1968 702 1983 736
rect 2017 732 2304 736
tri 2304 732 2320 748 nw
rect 2017 728 2300 732
tri 2300 728 2304 732 nw
rect 2017 727 2299 728
tri 2299 727 2300 728 nw
rect 2017 702 2265 727
rect 708 693 1810 696
tri 1810 693 1813 696 sw
rect 1968 693 2265 702
tri 2265 693 2299 727 nw
rect 708 691 1813 693
tri 1813 691 1815 693 sw
rect 1968 691 2263 693
tri 2263 691 2265 693 nw
rect 708 690 1815 691
rect 708 656 720 690
rect 754 656 792 690
rect 826 657 1815 690
tri 1815 657 1849 691 sw
rect 1968 684 2256 691
tri 2256 684 2263 691 nw
rect 1968 657 2075 684
tri 2075 657 2102 684 nw
rect 826 656 1849 657
rect 708 650 1849 656
tri 1782 647 1785 650 ne
rect 1785 647 1849 650
tri 1849 647 1859 657 sw
rect 1968 647 2065 657
tri 2065 647 2075 657 nw
tri 1785 642 1790 647 ne
rect 1790 642 1859 647
tri 1859 642 1864 647 sw
rect 1968 642 2048 647
tri 1790 611 1821 642 ne
rect 1821 611 1864 642
rect -242 605 1752 611
tri 1821 608 1824 611 ne
rect 1824 608 1864 611
tri 1864 608 1898 642 sw
rect 1968 608 1983 642
rect 2017 630 2048 642
tri 2048 630 2065 647 nw
rect 2129 636 2295 642
rect 2017 608 2032 630
tri 2032 614 2048 630 nw
rect -242 553 -237 605
rect -185 599 1752 605
rect -185 565 4 599
rect 38 565 1079 599
rect 1113 565 1391 599
rect 1425 565 1703 599
rect 1737 565 1752 599
tri 1824 596 1836 608 ne
rect 1836 596 1898 608
tri 1898 596 1910 608 sw
rect 1968 596 2032 608
tri 1836 590 1842 596 ne
rect 1842 590 1910 596
tri 1910 590 1916 596 sw
tri 1842 583 1849 590 ne
rect 1849 583 1916 590
tri 1916 583 1923 590 sw
rect 2181 630 2295 636
rect 2181 596 2255 630
rect 2289 596 2295 630
rect 2181 584 2295 596
rect -185 553 1752 565
tri 1849 558 1874 583 ne
rect 1874 558 1923 583
tri 1923 558 1948 583 sw
rect 2129 570 2295 584
rect -242 516 1752 553
tri 1874 524 1908 558 ne
rect 1908 524 1948 558
tri 1948 524 1982 558 sw
tri 1908 518 1914 524 ne
rect 1914 518 1982 524
tri 1982 518 1988 524 sw
rect 2181 558 2295 570
rect 2181 524 2255 558
rect 2289 524 2295 558
rect 2181 518 2295 524
rect -242 464 -237 516
rect -185 505 1752 516
tri 1914 509 1923 518 ne
rect 1923 509 1988 518
tri 1988 509 1997 518 sw
rect 2129 512 2295 518
rect -185 504 1079 505
rect -185 470 4 504
rect 38 471 1079 504
rect 1113 471 1391 505
rect 1425 471 1703 505
rect 1737 471 1752 505
tri 1923 484 1948 509 ne
rect 1948 484 1997 509
tri 1997 484 2022 509 sw
tri 2398 484 2414 500 se
rect 2414 484 2466 917
tri 2466 910 2473 917 nw
rect 3063 908 3109 920
tri 1948 474 1958 484 ne
rect 1958 474 2022 484
tri 2022 474 2032 484 sw
tri 2388 474 2398 484 se
rect 2398 478 2466 484
rect 2398 474 2462 478
tri 2462 474 2466 478 nw
rect 2742 895 2806 907
rect 2742 861 2757 895
rect 2791 861 2806 895
rect 2742 801 2806 861
rect 2742 767 2757 801
rect 2791 767 2806 801
rect 2742 657 2806 767
rect 3063 874 3069 908
rect 3103 874 3109 908
rect 3063 836 3109 874
rect 3063 802 3069 836
rect 3103 802 3109 836
rect 3063 693 3109 802
rect 3375 908 3421 920
rect 3375 874 3381 908
rect 3415 874 3421 908
rect 3375 838 3421 874
rect 3687 908 3733 920
rect 3687 874 3693 908
rect 3727 874 3733 908
tri 3421 838 3423 840 sw
rect 3375 836 3423 838
tri 3423 836 3425 838 sw
rect 3687 836 3733 874
rect 3375 802 3381 836
rect 3415 802 3425 836
tri 3425 802 3459 836 sw
tri 3674 802 3687 815 se
rect 3687 802 3693 836
rect 3727 802 3733 836
rect 3375 790 3459 802
tri 3459 790 3471 802 sw
tri 3662 790 3674 802 se
rect 3674 790 3733 802
rect 3817 917 3863 920
tri 3863 917 3866 920 sw
tri 4205 917 4208 920 se
rect 4208 917 4262 920
tri 4714 917 4717 920 ne
rect 4717 917 4788 920
tri 4788 917 4791 920 sw
rect 4895 917 4941 963
rect 3817 908 3866 917
rect 3817 874 3823 908
rect 3857 883 3866 908
tri 3866 883 3900 917 sw
tri 4171 883 4205 917 se
rect 4205 916 4262 917
rect 4205 883 4210 916
rect 3857 878 3900 883
tri 3900 878 3905 883 sw
tri 4166 878 4171 883 se
rect 4171 878 4210 883
rect 3857 874 4210 878
rect 3817 864 4210 874
tri 4717 895 4739 917 ne
rect 4739 895 4791 917
tri 4791 895 4813 917 sw
tri 4739 883 4751 895 ne
rect 4751 883 4813 895
tri 4813 883 4825 895 sw
rect 4895 883 4901 917
rect 4935 883 4941 917
tri 4751 864 4770 883 ne
rect 4770 864 4825 883
tri 4825 864 4844 883 sw
rect 4895 871 4941 883
rect 5021 1125 5027 1159
rect 5061 1155 5091 1159
tri 5091 1155 5125 1189 nw
rect 5061 1125 5067 1155
tri 5067 1131 5091 1155 nw
rect 5021 1079 5067 1125
rect 5188 1128 5969 1140
rect 5188 1094 5200 1128
rect 5234 1094 5272 1128
rect 5306 1094 5344 1128
rect 5378 1094 5416 1128
rect 5450 1094 5488 1128
rect 5522 1094 5560 1128
rect 5594 1094 5632 1128
rect 5666 1094 5704 1128
rect 5738 1094 5776 1128
rect 5810 1094 5848 1128
rect 5882 1094 5920 1128
rect 5954 1094 5969 1128
rect 5188 1082 5969 1094
tri 5682 1080 5684 1082 ne
rect 5684 1080 5916 1082
tri 5916 1080 5918 1082 nw
rect 5021 1045 5027 1079
rect 5061 1045 5067 1079
tri 5684 1054 5710 1080 ne
rect 5710 1054 5890 1080
tri 5890 1054 5916 1080 nw
rect 5021 999 5067 1045
tri 5710 1039 5725 1054 ne
rect 5725 1039 5875 1054
tri 5875 1039 5890 1054 nw
tri 5725 1029 5735 1039 ne
rect 5021 965 5027 999
rect 5061 965 5067 999
rect 5021 920 5067 965
rect 5021 886 5027 920
rect 5061 886 5067 920
rect 5021 874 5067 886
rect 5137 982 5495 994
rect 5137 948 5143 982
rect 5177 948 5455 982
rect 5489 948 5495 982
rect 5137 898 5495 948
rect 5137 864 5143 898
rect 5177 864 5455 898
rect 5489 864 5495 898
rect 5735 930 5843 1039
tri 5843 1007 5875 1039 nw
rect 5735 914 5827 930
tri 5827 914 5843 930 nw
rect 5735 910 5823 914
tri 5823 910 5827 914 nw
rect 5735 896 5809 910
tri 5809 896 5823 910 nw
tri 5728 889 5735 896 se
rect 5735 889 5802 896
tri 5802 889 5809 896 nw
rect 3817 852 4262 864
tri 4770 855 4779 864 ne
rect 4779 855 4844 864
tri 4844 855 4853 864 sw
rect 3817 836 4210 852
rect 3817 802 3823 836
rect 3857 832 4210 836
rect 3857 814 3887 832
tri 3887 814 3905 832 nw
tri 4172 814 4190 832 ne
rect 4190 814 4210 832
rect 3857 802 3863 814
rect 3375 780 3471 790
tri 3471 780 3481 790 sw
tri 3652 780 3662 790 se
rect 3662 780 3733 790
tri 3733 780 3749 796 sw
rect 3817 790 3863 802
tri 3863 790 3887 814 nw
tri 4190 794 4210 814 ne
tri 4779 842 4792 855 ne
rect 4792 842 4853 855
tri 4853 842 4866 855 sw
rect 5137 852 5495 864
tri 5694 855 5728 889 se
rect 5728 855 5768 889
tri 5768 855 5802 889 nw
tri 5691 852 5694 855 se
rect 5694 852 5755 855
tri 5681 842 5691 852 se
rect 5691 842 5755 852
tri 5755 842 5768 855 nw
tri 4792 838 4796 842 ne
rect 4796 838 4866 842
tri 4866 838 4870 842 sw
tri 5677 838 5681 842 se
rect 5681 838 5751 842
tri 5751 838 5755 842 nw
tri 4796 821 4813 838 ne
rect 4813 821 4870 838
tri 4870 821 4887 838 sw
tri 5661 822 5677 838 se
rect 5677 822 5735 838
tri 5735 822 5751 838 nw
tri 5660 821 5661 822 se
rect 5661 821 5727 822
tri 4813 814 4820 821 ne
rect 4820 814 5727 821
tri 5727 814 5735 822 nw
rect 4210 794 4262 800
tri 4820 794 4840 814 ne
rect 4840 794 5693 814
tri 4840 790 4844 794 ne
rect 4844 790 5693 794
tri 4844 780 4854 790 ne
rect 4854 780 5693 790
tri 5693 780 5727 814 nw
rect 3375 779 3481 780
tri 3481 779 3482 780 sw
tri 3651 779 3652 780 se
rect 3652 779 3749 780
rect 3375 766 3749 779
tri 3749 766 3763 780 sw
tri 4854 769 4865 780 ne
rect 4865 769 5682 780
tri 5682 769 5693 780 nw
rect 3375 760 3763 766
tri 3763 760 3769 766 sw
rect 3375 733 3733 760
tri 3635 732 3636 733 ne
rect 3636 732 3733 733
tri 3636 728 3640 732 ne
rect 3640 728 3733 732
tri 3640 727 3641 728 ne
rect 3641 727 3733 728
rect 4383 727 4941 739
tri 5990 732 5997 739 se
rect 5997 732 6043 1231
tri 6043 1229 6045 1231 nw
rect 6110 1197 6164 1231
rect 6198 1230 6239 1231
rect 6273 1230 6279 1264
rect 6198 1197 6279 1230
rect 6110 1191 6279 1197
tri 6139 1189 6141 1191 ne
rect 6141 1189 6279 1191
rect 6349 1380 10011 1392
rect 6349 1346 6355 1380
rect 6389 1346 6867 1380
rect 6901 1346 7379 1380
rect 7413 1346 7891 1380
rect 7925 1346 8403 1380
rect 8437 1346 8915 1380
rect 8949 1346 9267 1380
rect 9301 1346 9619 1380
rect 9653 1346 9971 1380
rect 10005 1346 10011 1380
rect 6349 1308 10011 1346
rect 6349 1274 6355 1308
rect 6389 1274 6867 1308
rect 6901 1274 7379 1308
rect 7413 1274 7891 1308
rect 7925 1274 8403 1308
rect 8437 1274 8915 1308
rect 8949 1274 9267 1308
rect 9301 1274 9619 1308
rect 9653 1274 9971 1308
rect 10005 1274 10011 1308
rect 6349 1236 10011 1274
rect 6349 1202 6355 1236
rect 6389 1202 6867 1236
rect 6901 1202 7379 1236
rect 7413 1202 7891 1236
rect 7925 1202 8403 1236
rect 8437 1202 8915 1236
rect 8949 1202 9267 1236
rect 9301 1202 9619 1236
rect 9653 1202 9971 1236
rect 10005 1202 10011 1236
rect 6349 1190 10011 1202
rect 10082 1380 10088 1414
rect 10122 1380 10128 1414
rect 10082 1342 10128 1380
rect 10082 1308 10088 1342
rect 10122 1308 10128 1342
rect 10082 1270 10128 1308
rect 10082 1236 10088 1270
rect 10122 1236 10128 1270
rect 10082 1198 10128 1236
tri 6141 1155 6175 1189 ne
rect 6175 1155 6239 1189
rect 6273 1155 6279 1189
tri 8587 1164 8613 1190 ne
rect 8613 1164 9162 1190
tri 9162 1164 9188 1190 nw
rect 10082 1164 10088 1198
rect 10122 1164 10128 1198
tri 6175 1126 6204 1155 ne
rect 6204 1126 6279 1155
tri 8613 1126 8651 1164 ne
rect 8651 1126 9124 1164
tri 9124 1126 9162 1164 nw
tri 10061 1126 10082 1147 se
rect 10082 1126 10128 1164
tri 6204 1114 6216 1126 ne
rect 6216 1114 6279 1126
tri 6216 1097 6233 1114 ne
rect 6233 1080 6239 1114
rect 6273 1080 6279 1114
tri 8651 1092 8685 1126 ne
rect 8685 1092 9090 1126
tri 9090 1092 9124 1126 nw
tri 10027 1092 10061 1126 se
rect 10061 1092 10088 1126
rect 10122 1092 10128 1126
rect 6233 1039 6279 1080
tri 8685 1054 8723 1092 ne
rect 8723 1054 9052 1092
tri 9052 1054 9090 1092 nw
tri 9989 1054 10027 1092 se
rect 10027 1054 10128 1092
tri 8723 1043 8734 1054 ne
rect 6233 1005 6239 1039
rect 6273 1005 6279 1039
rect 6233 964 6279 1005
rect 6233 930 6239 964
rect 6273 930 6279 964
rect 6233 889 6279 930
rect 6233 855 6239 889
rect 6273 855 6279 889
rect 6233 814 6279 855
rect 6460 1020 7780 1032
rect 6460 986 6611 1020
rect 6645 986 7123 1020
rect 7157 986 7635 1020
rect 7669 986 7780 1020
rect 6460 948 7780 986
rect 6460 914 6611 948
rect 6645 914 7123 948
rect 7157 914 7635 948
rect 7669 914 7780 948
rect 6460 876 7780 914
rect 6460 842 6611 876
rect 6645 842 7123 876
rect 7157 842 7635 876
rect 7669 842 7780 876
rect 6460 830 7780 842
rect 8117 1020 8699 1032
rect 8117 986 8147 1020
rect 8181 986 8659 1020
rect 8693 986 8699 1020
rect 8117 948 8699 986
rect 8117 914 8147 948
rect 8181 914 8659 948
rect 8693 914 8699 948
rect 8117 876 8699 914
rect 8117 842 8147 876
rect 8181 842 8659 876
rect 8693 842 8699 876
rect 8117 830 8699 842
rect 6233 780 6239 814
rect 6273 780 6279 814
tri 7192 804 7218 830 ne
rect 7218 804 7465 830
tri 7465 804 7491 830 nw
tri 8433 804 8459 830 ne
rect 8459 804 8699 830
rect 6233 768 6279 780
tri 7218 778 7244 804 ne
tri 6043 732 6050 739 sw
tri 5986 728 5990 732 se
rect 5990 728 6050 732
tri 6050 728 6054 732 sw
rect 6402 728 7177 734
tri 3641 696 3672 727 ne
rect 3672 696 3751 727
tri 3109 693 3112 696 sw
tri 3672 693 3675 696 ne
rect 3675 693 3751 696
tri 3751 693 3785 727 nw
rect 4383 693 4389 727
rect 4423 693 4901 727
rect 4935 693 4941 727
rect 3063 691 3112 693
tri 3112 691 3114 693 sw
tri 3675 691 3677 693 ne
rect 3677 691 3749 693
tri 3749 691 3751 693 nw
tri 2806 657 2833 684 sw
rect 3063 657 3114 691
tri 3114 657 3148 691 sw
tri 3677 681 3687 691 ne
rect 2742 647 2833 657
tri 2833 647 2843 657 sw
rect 3063 647 3148 657
tri 3148 647 3158 657 sw
rect 2742 614 2843 647
tri 2843 614 2876 647 sw
rect 2742 590 3020 614
rect 2742 556 2964 590
rect 2998 556 3020 590
rect 2742 518 3020 556
rect 2742 484 2964 518
rect 2998 484 3020 518
rect 38 470 1752 471
rect -185 464 1752 470
rect -242 458 1752 464
tri 1958 458 1974 474 ne
rect 1974 458 2032 474
tri 1974 444 1988 458 ne
rect 1988 444 2032 458
tri 2032 444 2062 474 sw
tri 2358 444 2388 474 se
rect 2388 444 2432 474
tri 2432 444 2462 474 nw
rect 2742 472 3020 484
rect 3063 613 3158 647
tri 3158 613 3192 647 sw
rect 3063 602 3192 613
tri 3192 602 3203 613 sw
rect 3063 590 3316 602
rect 3063 556 3276 590
rect 3310 556 3316 590
rect 3063 518 3316 556
rect 3063 484 3276 518
rect 3310 484 3316 518
tri 3682 492 3687 497 se
rect 3687 492 3733 691
tri 3733 675 3749 691 nw
rect 4383 647 4941 693
tri 5955 697 5986 728 se
rect 5986 697 6054 728
tri 6054 697 6085 728 sw
rect 5955 691 6085 697
rect 5955 657 5967 691
rect 6001 657 6039 691
rect 6073 657 6085 691
rect 6402 694 6414 728
rect 6448 694 6493 728
rect 6527 694 6572 728
rect 6606 694 6651 728
rect 6685 694 6731 728
rect 6765 694 6811 728
rect 6845 694 6891 728
rect 6925 694 6971 728
rect 7005 694 7051 728
rect 7085 694 7131 728
rect 7165 694 7177 728
rect 6402 688 7177 694
rect 5955 651 6085 657
rect 4383 613 4389 647
rect 4423 613 4901 647
rect 4935 613 4941 647
tri 7223 622 7244 643 se
rect 7244 622 7439 804
tri 7439 778 7465 804 nw
tri 8459 778 8485 804 ne
rect 8485 778 8699 804
tri 8485 766 8497 778 ne
rect 8497 766 8699 778
tri 8497 755 8508 766 ne
tri 8333 734 8336 737 se
rect 8336 734 8342 737
rect 7502 728 8342 734
rect 7502 694 7514 728
rect 7548 694 7590 728
rect 7624 694 7666 728
rect 7700 694 7742 728
rect 7776 694 7818 728
rect 7852 694 7894 728
rect 7928 694 7971 728
rect 8005 694 8048 728
rect 8082 694 8125 728
rect 8159 694 8202 728
rect 8236 694 8279 728
rect 8313 694 8342 728
rect 7502 688 8342 694
tri 8333 685 8336 688 ne
rect 8336 685 8342 688
rect 8394 685 8406 737
rect 8458 685 8464 737
tri 8499 660 8508 669 se
rect 8508 660 8699 766
tri 8482 643 8499 660 se
rect 8499 643 8699 660
tri 7439 622 7460 643 sw
tri 8461 622 8482 643 se
rect 8482 622 8699 643
rect 4383 601 4941 613
tri 7202 601 7223 622 se
rect 7223 601 7460 622
tri 7193 592 7202 601 se
rect 7202 592 7460 601
tri 7460 592 7490 622 sw
tri 8431 592 8461 622 se
rect 8461 592 8699 622
tri 5077 588 5081 592 se
rect 5081 588 7810 592
tri 5069 580 5077 588 se
rect 5077 580 7810 588
tri 5035 546 5069 580 se
rect 5069 546 5299 580
rect 5333 546 5611 580
rect 5645 546 6123 580
rect 6157 546 6611 580
rect 6645 546 7123 580
rect 7157 546 7635 580
rect 7669 546 7810 580
tri 5028 539 5035 546 se
rect 5035 539 7810 546
rect 3063 472 3316 484
tri 3664 474 3682 492 se
rect 3682 474 3733 492
tri 3662 472 3664 474 se
rect 3664 472 3733 474
rect 2742 444 2848 472
tri 2848 444 2876 472 nw
rect 3063 444 3177 472
tri 3177 444 3205 472 nw
tri 3634 444 3662 472 se
rect 3662 444 3733 472
tri 1988 436 1996 444 ne
rect 1996 436 2062 444
tri 2062 436 2070 444 sw
tri 2350 436 2358 444 se
rect 2358 436 2424 444
tri 2424 436 2432 444 nw
rect 2742 436 2840 444
tri 2840 436 2848 444 nw
rect 3063 436 3169 444
tri 3169 436 3177 444 nw
tri 3626 436 3634 444 se
rect 3634 436 3733 444
tri 1996 435 1997 436 ne
rect 1997 435 2070 436
tri 2070 435 2071 436 sw
tri 2349 435 2350 436 se
rect 2350 435 2423 436
tri 2423 435 2424 436 nw
tri 1997 421 2011 435 ne
rect 2011 421 2409 435
tri 2409 421 2423 435 nw
rect 2742 421 2816 436
tri 2011 387 2045 421 ne
rect 2045 387 2375 421
tri 2375 387 2409 421 nw
rect 2742 387 2757 421
rect 2791 412 2816 421
tri 2816 412 2840 436 nw
rect 3063 412 3145 436
tri 3145 412 3169 436 nw
tri 3602 412 3626 436 se
rect 3626 412 3733 436
rect 4636 526 7810 539
rect 4636 492 4645 526
rect 4679 508 7810 526
rect 4679 492 5299 508
rect 4636 474 5299 492
rect 5333 474 5611 508
rect 5645 474 6123 508
rect 6157 474 6611 508
rect 6645 474 7123 508
rect 7157 474 7635 508
rect 7669 474 7810 508
rect 4636 436 7810 474
tri 4136 412 4148 424 se
rect 4148 412 4302 424
rect 2791 387 2806 412
tri 2806 402 2816 412 nw
tri 2045 383 2049 387 ne
rect 2049 383 2371 387
tri 2371 383 2375 387 nw
rect 1220 371 1636 383
rect 1220 337 1235 371
rect 1269 337 1547 371
rect 1581 365 1636 371
tri 1636 365 1654 383 sw
rect 1581 348 1654 365
tri 1654 348 1671 365 sw
rect 1581 347 1671 348
tri 1671 347 1672 348 sw
rect 1581 340 1672 347
tri 1672 340 1679 347 sw
rect 1581 337 1679 340
rect 1220 327 1679 337
tri 1679 327 1692 340 sw
rect 2742 327 2806 387
rect 1220 297 1692 327
tri 1692 297 1722 327 sw
rect 1220 281 2508 297
rect 2742 293 2757 327
rect 2791 293 2806 327
rect 2742 281 2806 293
rect 3063 399 3115 412
rect 3063 365 3069 399
rect 3103 382 3115 399
tri 3115 382 3145 412 nw
tri 3584 394 3602 412 se
rect 3602 394 3733 412
rect 3375 382 3733 394
rect 3103 365 3109 382
tri 3109 376 3115 382 nw
rect 3063 327 3109 365
rect 3063 293 3069 327
rect 3103 293 3109 327
rect 3063 281 3109 293
rect 3375 348 3381 382
rect 3415 348 3693 382
rect 3727 348 3733 382
tri 4102 378 4136 412 se
rect 4136 378 4262 412
rect 4296 378 4302 412
rect 4636 402 4645 436
rect 4679 402 5299 436
rect 5333 402 5611 436
rect 5645 402 6123 436
rect 6157 402 6611 436
rect 6645 402 7123 436
rect 7157 402 7635 436
rect 7669 402 7810 436
rect 4636 390 7810 402
rect 7811 391 7812 591
rect 8112 391 8113 591
rect 8114 580 8699 592
rect 8114 546 8147 580
rect 8181 546 8659 580
rect 8693 546 8699 580
rect 8114 508 8699 546
rect 8114 474 8147 508
rect 8181 474 8659 508
rect 8693 474 8699 508
rect 8114 436 8699 474
rect 8114 402 8147 436
rect 8181 402 8659 436
rect 8693 402 8699 436
rect 8114 390 8699 402
tri 4096 372 4102 378 se
rect 4102 372 4302 378
tri 8724 372 8734 382 se
rect 8734 372 9035 1054
tri 9035 1037 9052 1054 nw
tri 9972 1037 9989 1054 se
rect 9989 1037 10088 1054
tri 9967 1032 9972 1037 se
rect 9972 1032 10088 1037
rect 9085 1020 10088 1032
rect 10122 1020 10128 1054
rect 9085 986 9091 1020
rect 9125 986 9443 1020
rect 9477 986 9795 1020
rect 9829 986 10128 1020
rect 9085 982 10128 986
rect 9085 948 10088 982
rect 10122 948 10128 982
rect 9085 914 9091 948
rect 9125 914 9443 948
rect 9477 914 9795 948
rect 9829 914 10128 948
rect 9085 910 10128 914
rect 9085 876 10088 910
rect 10122 876 10128 910
rect 9085 842 9091 876
rect 9125 842 9443 876
rect 9477 842 9795 876
rect 9829 842 10128 876
rect 9085 838 10128 842
rect 9085 830 10088 838
tri 9085 804 9111 830 ne
rect 9111 804 9280 830
tri 9280 804 9306 830 nw
tri 9992 804 10018 830 ne
rect 10018 804 10088 830
rect 10122 804 10128 838
tri 9111 766 9149 804 ne
rect 9149 766 9242 804
tri 9242 766 9280 804 nw
tri 10018 773 10049 804 ne
rect 10049 773 10128 804
tri 9804 766 9811 773 se
rect 9811 767 9863 773
tri 9149 761 9154 766 ne
tri 9153 660 9154 661 se
rect 9154 660 9237 766
tri 9237 761 9242 766 nw
tri 9799 761 9804 766 se
rect 9804 761 9811 766
tri 9772 734 9799 761 se
rect 9799 734 9811 761
rect 9558 728 9811 734
tri 9863 766 9870 773 sw
tri 10049 766 10056 773 ne
rect 10056 766 10128 773
rect 9863 734 9870 766
tri 9870 734 9902 766 sw
tri 10056 740 10082 766 ne
rect 9863 728 9971 734
rect 9558 694 9570 728
rect 9604 694 9658 728
rect 9692 694 9747 728
rect 9781 715 9811 728
rect 9781 703 9836 715
rect 9781 694 9811 703
rect 9870 694 9925 728
rect 9959 694 9971 728
rect 9558 688 9811 694
tri 9772 678 9782 688 ne
rect 9782 678 9811 688
tri 9237 660 9255 678 sw
tri 9782 660 9800 678 ne
rect 9800 660 9811 678
tri 9115 622 9153 660 se
rect 9153 622 9255 660
tri 9255 622 9293 660 sw
tri 9800 649 9811 660 ne
rect 9863 688 9971 694
rect 10082 732 10088 766
rect 10122 732 10128 766
rect 10082 694 10128 732
rect 9863 660 9874 688
tri 9874 660 9902 688 nw
tri 10060 660 10082 682 se
rect 10082 660 10088 694
rect 10122 660 10128 694
rect 9811 645 9863 651
tri 9863 649 9874 660 nw
tri 10049 649 10060 660 se
rect 10060 649 10128 660
tri 10045 645 10049 649 se
rect 10049 645 10128 649
tri 10022 622 10045 645 se
rect 10045 622 10128 645
tri 9085 592 9115 622 se
rect 9115 592 9293 622
tri 9293 592 9323 622 sw
tri 9992 592 10022 622 se
rect 10022 592 10088 622
rect 9085 588 10088 592
rect 10122 588 10128 622
rect 9085 580 10128 588
rect 9085 546 9091 580
rect 9125 546 9443 580
rect 9477 546 9795 580
rect 9829 550 10128 580
rect 9829 546 10088 550
rect 9085 516 10088 546
rect 10122 516 10128 550
rect 9085 508 10128 516
rect 9085 474 9091 508
rect 9125 474 9443 508
rect 9477 474 9795 508
rect 9829 478 10128 508
rect 9829 474 10088 478
rect 9085 444 10088 474
rect 10122 444 10128 478
rect 9085 436 10128 444
rect 9085 402 9091 436
rect 9125 402 9443 436
rect 9477 402 9795 436
rect 9829 406 10128 436
rect 9829 402 10088 406
rect 9085 390 10088 402
tri 9950 382 9958 390 ne
rect 9958 382 10088 390
tri 9035 372 9045 382 sw
tri 9958 372 9968 382 ne
rect 9968 372 10088 382
rect 10122 372 10128 406
rect 3375 310 3733 348
tri 4071 347 4096 372 se
rect 4096 347 4302 372
tri 8711 359 8724 372 se
rect 8724 359 9045 372
tri 4427 347 4439 359 se
rect 4439 347 5066 359
tri 4064 340 4071 347 se
rect 4071 340 4302 347
rect 1220 277 2385 281
rect 1220 243 1235 277
rect 1269 243 1547 277
rect 1581 247 2385 277
rect 2419 247 2462 281
rect 2496 247 2508 281
rect 3375 276 3381 310
rect 3415 276 3693 310
rect 3727 276 3733 310
tri 4030 306 4064 340 se
rect 4064 306 4262 340
rect 4296 306 4302 340
tri 4393 313 4427 347 se
rect 4427 313 4540 347
rect 4574 313 4747 347
rect 4781 313 4819 347
rect 4853 336 5066 347
tri 5066 336 5089 359 sw
tri 8688 336 8711 359 se
rect 8711 336 9045 359
rect 4853 326 8446 336
rect 4853 324 5967 326
rect 4853 313 5143 324
tri 4014 290 4030 306 se
rect 4030 294 4302 306
tri 4374 294 4393 313 se
rect 4393 301 5143 313
rect 4393 294 4452 301
rect 4030 290 4188 294
tri 4188 290 4192 294 nw
tri 4370 290 4374 294 se
rect 4374 290 4452 294
tri 4452 290 4463 301 nw
tri 4967 290 4978 301 ne
rect 4978 290 5143 301
rect 5177 290 5455 324
rect 5489 292 5967 324
rect 6001 292 6039 326
rect 6073 292 8446 326
rect 5489 290 8446 292
rect 3375 264 3733 276
tri 3988 264 4014 290 se
rect 4014 264 4160 290
tri 3986 262 3988 264 se
rect 3988 262 4160 264
tri 4160 262 4188 290 nw
tri 4357 277 4370 290 se
rect 4370 277 4439 290
tri 4439 277 4452 290 nw
tri 4978 278 4990 290 ne
rect 4990 284 8446 290
rect 8498 284 8510 336
rect 8562 284 8572 336
tri 8686 334 8688 336 se
rect 8688 334 9045 336
tri 9045 334 9083 372 sw
tri 9968 334 10006 372 ne
rect 10006 334 10128 372
tri 8652 300 8686 334 se
rect 8686 300 9083 334
tri 9083 300 9117 334 sw
tri 10006 300 10040 334 ne
rect 10040 300 10088 334
rect 10122 300 10128 334
rect 4990 278 8572 284
tri 8630 278 8652 300 se
rect 8652 278 9117 300
tri 5093 277 5094 278 ne
rect 5094 277 5523 278
tri 4342 262 4357 277 se
rect 4357 262 4424 277
tri 4424 262 4439 277 nw
tri 5094 262 5109 277 ne
rect 5109 262 5523 277
tri 5523 262 5539 278 nw
tri 8614 262 8630 278 se
rect 8630 262 9117 278
tri 9117 262 9155 300 sw
tri 10040 262 10078 300 ne
rect 10078 262 10128 300
tri 3976 252 3986 262 se
rect 3986 252 4150 262
tri 4150 252 4160 262 nw
tri 4332 252 4342 262 se
rect 4342 252 4414 262
tri 4414 252 4424 262 nw
tri 5109 252 5119 262 ne
rect 5119 252 5495 262
tri 3974 250 3976 252 se
rect 3976 250 4148 252
tri 4148 250 4150 252 nw
tri 4330 250 4332 252 se
rect 4332 250 4380 252
rect 1581 243 2508 247
rect 1220 231 2508 243
tri 3958 234 3974 250 se
rect 3974 234 4116 250
tri 2317 222 2326 231 ne
rect 2326 222 2499 231
tri 2499 222 2508 231 nw
rect 2550 222 4116 234
tri 2326 200 2348 222 ne
rect 2348 200 2465 222
rect 421 194 2188 200
rect 421 188 1027 194
rect 421 154 436 188
rect 470 154 868 188
rect 902 154 1027 188
rect 421 142 1027 154
rect 1079 188 2188 194
tri 2348 188 2360 200 ne
rect 2360 188 2465 200
tri 2465 188 2499 222 nw
rect 2550 188 2601 222
rect 2635 188 2913 222
rect 2947 188 3225 222
rect 3259 188 3537 222
rect 3571 188 3999 222
rect 4033 218 4116 222
tri 4116 218 4148 250 nw
tri 4298 218 4330 250 se
rect 4330 218 4380 250
tri 4380 218 4414 252 nw
tri 5119 234 5137 252 ne
rect 5137 218 5143 252
rect 5177 218 5455 252
rect 5489 218 5495 252
tri 5495 234 5523 262 nw
tri 8586 234 8614 262 se
rect 8614 234 9155 262
tri 8584 232 8586 234 se
rect 8586 232 9155 234
tri 9155 232 9185 262 sw
tri 10078 258 10082 262 ne
rect 4033 188 4087 218
tri 4087 189 4116 218 nw
tri 4275 195 4298 218 se
rect 4298 195 4357 218
tri 4357 195 4380 218 nw
tri 4269 189 4275 195 se
rect 4275 189 4348 195
rect 1079 154 1827 188
rect 1861 154 2139 188
rect 2173 154 2188 188
tri 2360 186 2362 188 ne
rect 2362 186 2463 188
tri 2463 186 2465 188 nw
tri 2362 180 2368 186 ne
rect 2368 180 2457 186
tri 2457 180 2463 186 nw
tri 2368 173 2375 180 ne
rect 2375 173 2450 180
tri 2450 173 2457 180 nw
tri 2375 170 2378 173 ne
rect 1079 142 2188 154
rect 421 117 2188 142
rect 421 102 1027 117
rect 421 68 436 102
rect 470 68 868 102
rect 902 68 1027 102
rect 421 65 1027 68
rect 1079 102 2188 117
rect 1079 68 1827 102
rect 1861 68 2139 102
rect 2173 68 2188 102
rect 1079 65 2188 68
rect 421 39 2188 65
rect 421 15 1027 39
rect 421 -19 436 15
rect 470 -19 868 15
rect 902 -13 1027 15
rect 1079 15 2188 39
tri 2370 23 2378 31 se
rect 2378 23 2447 173
tri 2447 170 2450 173 nw
rect 2550 150 4087 188
tri 4266 186 4269 189 se
rect 4269 186 4348 189
tri 4348 186 4357 195 nw
tri 4260 180 4266 186 se
rect 4266 180 4342 186
tri 4342 180 4348 186 nw
tri 4253 173 4260 180 se
rect 4260 173 4335 180
tri 4335 173 4342 180 nw
rect 5021 173 5067 185
rect 2550 116 2601 150
rect 2635 116 2913 150
rect 2947 116 3225 150
rect 3259 116 3537 150
rect 3571 116 3999 150
rect 4033 116 4087 150
tri 4225 145 4253 173 se
rect 4253 145 4307 173
tri 4307 145 4335 173 nw
rect 2550 57 4087 116
tri 2447 23 2455 31 sw
rect 2550 23 2609 57
rect 2643 23 2681 57
rect 2715 23 2753 57
rect 2787 23 2825 57
rect 2859 23 2897 57
rect 2931 23 2969 57
rect 3003 23 3041 57
rect 3075 23 3113 57
rect 3147 23 3185 57
rect 3219 23 3257 57
rect 3291 23 3329 57
rect 3363 23 3401 57
rect 3435 23 3473 57
rect 3507 23 3545 57
rect 3579 23 3617 57
rect 3651 23 3689 57
rect 3723 23 4087 57
tri 2364 17 2370 23 se
rect 2370 17 2455 23
tri 2455 17 2461 23 sw
rect 1079 -13 1827 15
rect 902 -19 1827 -13
rect 1861 -19 2139 15
rect 2173 -19 2188 15
tri 2357 10 2364 17 se
rect 2364 10 2461 17
tri 2461 10 2468 17 sw
rect 2550 11 4087 23
tri 4207 127 4225 145 se
rect 4225 127 4289 145
tri 4289 127 4307 145 nw
rect 4207 111 4273 127
tri 4273 111 4289 127 nw
tri 4202 17 4207 22 se
rect 4207 17 4265 111
tri 4265 103 4273 111 nw
rect 4438 105 4444 157
rect 4496 105 4551 157
rect 4603 145 4958 157
rect 4603 111 4909 145
rect 4943 111 4958 145
rect 4603 105 4958 111
tri 4196 11 4202 17 se
rect 4202 11 4265 17
tri 4195 10 4196 11 se
rect 4196 10 4265 11
rect 421 -31 2188 -19
tri 2320 -27 2357 10 se
rect 2357 -27 2468 10
tri 2468 -27 2505 10 sw
tri 4158 -27 4195 10 se
rect 4195 -23 4265 10
rect 4438 59 4958 105
rect 4438 7 4444 59
rect 4496 7 4551 59
rect 4603 51 4958 59
rect 4603 17 4909 51
rect 4943 17 4958 51
rect 4603 7 4958 17
rect 4438 5 4958 7
rect 5021 139 5027 173
rect 5061 139 5067 173
rect 5021 72 5067 139
rect 5137 180 5495 218
rect 5137 146 5143 180
rect 5177 146 5455 180
rect 5489 146 5495 180
rect 5137 134 5495 146
rect 5861 220 10011 232
rect 5861 186 5867 220
rect 5901 186 6355 220
rect 6389 186 6867 220
rect 6901 186 7379 220
rect 7413 186 7891 220
rect 7925 186 8403 220
rect 8437 186 8915 220
rect 8949 186 9267 220
rect 9301 186 9619 220
rect 9653 186 9971 220
rect 10005 186 10011 220
rect 5861 148 10011 186
rect 5021 38 5027 72
rect 5061 42 5067 72
rect 5861 114 5867 148
rect 5901 114 6355 148
rect 6389 114 6867 148
rect 6901 114 7379 148
rect 7413 114 7891 148
rect 7925 114 8403 148
rect 8437 114 8915 148
rect 8949 114 9267 148
rect 9301 114 9619 148
rect 9653 114 9971 148
rect 10005 114 10011 148
rect 5861 76 10011 114
tri 5067 42 5070 45 sw
rect 5861 42 5867 76
rect 5901 42 6355 76
rect 6389 42 6867 76
rect 6901 42 7379 76
rect 7413 42 7891 76
rect 7925 42 8403 76
rect 8437 42 8915 76
rect 8949 42 9267 76
rect 9301 42 9619 76
rect 9653 42 9971 76
rect 10005 42 10011 76
rect 5061 38 5070 42
rect 5021 10 5070 38
tri 5070 10 5102 42 sw
rect 5861 30 10011 42
rect 10082 228 10088 262
rect 10122 228 10128 262
rect 10082 190 10128 228
rect 10082 156 10088 190
rect 10122 156 10128 190
rect 10082 117 10128 156
rect 10082 83 10088 117
rect 10122 83 10128 117
rect 10082 44 10128 83
rect 10082 10 10088 44
rect 10122 10 10128 44
rect 4195 -27 4260 -23
tri 2319 -28 2320 -27 se
rect 2320 -28 4260 -27
tri 4260 -28 4265 -23 nw
rect 5021 -22 5102 10
tri 5102 -22 5134 10 sw
rect 10082 -22 10128 10
rect 5021 -28 10128 -22
tri 2317 -30 2319 -28 se
rect 2319 -30 4226 -28
tri 2316 -31 2317 -30 se
rect 2317 -31 4226 -30
tri 2314 -33 2316 -31 se
rect 2316 -33 4226 -31
tri 2280 -67 2314 -33 se
rect 2314 -67 2373 -33
rect 2407 -67 2445 -33
rect 2479 -62 4226 -33
tri 4226 -62 4260 -28 nw
rect 5021 -62 5099 -28
rect 5133 -62 5172 -28
rect 5206 -62 5245 -28
rect 5279 -62 5318 -28
rect 5352 -62 5391 -28
rect 5425 -62 5464 -28
rect 5498 -62 5537 -28
rect 5571 -62 5610 -28
rect 5644 -62 5683 -28
rect 5717 -62 5755 -28
rect 5789 -62 5827 -28
rect 5861 -62 5899 -28
rect 5933 -62 5971 -28
rect 6005 -62 6043 -28
rect 6077 -62 6115 -28
rect 6149 -62 6187 -28
rect 6221 -62 6311 -28
rect 6345 -62 6384 -28
rect 6418 -62 6457 -28
rect 6491 -62 6530 -28
rect 6564 -62 6603 -28
rect 6637 -62 6676 -28
rect 6710 -62 6749 -28
rect 6783 -62 6822 -28
rect 6856 -62 6895 -28
rect 6929 -62 6968 -28
rect 7002 -62 7041 -28
rect 7075 -62 7114 -28
rect 7148 -62 7187 -28
rect 7221 -62 7260 -28
rect 7294 -62 7333 -28
rect 7367 -62 7406 -28
rect 7440 -62 7479 -28
rect 7513 -62 7552 -28
rect 7586 -62 7625 -28
rect 7659 -62 7698 -28
rect 7732 -62 7771 -28
rect 7805 -62 7844 -28
rect 7878 -62 7917 -28
rect 7951 -62 7990 -28
rect 8024 -62 8063 -28
rect 8097 -62 8136 -28
rect 8170 -62 8209 -28
rect 8243 -62 8282 -28
rect 8316 -62 8355 -28
rect 8389 -62 8428 -28
rect 8462 -62 8501 -28
rect 8535 -62 8574 -28
rect 8608 -62 8647 -28
rect 8681 -62 8720 -28
rect 8754 -62 8792 -28
rect 8826 -62 8864 -28
rect 8898 -62 8936 -28
rect 8970 -62 9008 -28
rect 9042 -62 9080 -28
rect 9114 -62 9152 -28
rect 9186 -62 9224 -28
rect 9258 -62 9296 -28
rect 9330 -62 9368 -28
rect 9402 -62 9440 -28
rect 9474 -62 9512 -28
rect 9546 -62 9584 -28
rect 9618 -62 9656 -28
rect 9690 -62 9728 -28
rect 9762 -62 9800 -28
rect 9834 -62 9872 -28
rect 9906 -62 9944 -28
rect 9978 -62 10016 -28
rect 10050 -62 10128 -28
rect 2479 -67 4215 -62
tri 2254 -93 2280 -67 se
rect 2280 -73 4215 -67
tri 4215 -73 4226 -62 nw
rect 5021 -68 10128 -62
rect 2280 -93 2320 -73
tri 2320 -93 2340 -73 nw
tri 2231 -116 2254 -93 se
tri 914 -128 926 -116 se
rect 926 -128 2128 -116
tri 886 -156 914 -128 se
rect 914 -156 1146 -128
rect 68 -162 1146 -156
rect 1180 -162 1218 -128
rect 1252 -162 1290 -128
rect 1324 -162 1362 -128
rect 1396 -162 1434 -128
rect 1468 -162 1506 -128
rect 1540 -162 1578 -128
rect 1612 -162 1650 -128
rect 1684 -162 1722 -128
rect 1756 -162 1794 -128
rect 1828 -162 1866 -128
rect 1900 -162 1938 -128
rect 1972 -162 2010 -128
rect 2044 -162 2082 -128
rect 2116 -162 2128 -128
tri 2188 -159 2231 -116 se
rect 2231 -159 2254 -116
tri 2254 -159 2320 -93 nw
rect 68 -168 2128 -162
rect 68 -202 80 -168
rect 114 -202 152 -168
rect 186 -202 224 -168
rect 258 -202 296 -168
rect 330 -202 368 -168
rect 402 -202 440 -168
rect 474 -202 512 -168
rect 546 -202 584 -168
rect 618 -202 656 -168
rect 690 -202 728 -168
rect 762 -202 800 -168
rect 834 -174 2128 -168
tri 2173 -174 2188 -159 se
rect 2188 -174 2209 -159
rect 834 -202 922 -174
rect 68 -214 922 -202
tri 922 -214 962 -174 nw
tri 2143 -204 2173 -174 se
rect 2173 -204 2209 -174
tri 2209 -204 2254 -159 nw
tri 1245 -214 1255 -204 se
rect 1255 -214 2177 -204
tri 1212 -247 1245 -214 se
rect 1245 -236 2177 -214
tri 2177 -236 2209 -204 nw
rect 1245 -247 1276 -236
tri 1276 -247 1287 -236 nw
rect 691 -255 1226 -247
rect 691 -289 703 -255
rect 737 -289 778 -255
rect 812 -289 853 -255
rect 887 -289 928 -255
rect 962 -289 1003 -255
rect 1037 -289 1077 -255
rect 1111 -289 1151 -255
rect 1185 -289 1226 -255
rect 691 -297 1226 -289
tri 1226 -297 1276 -247 nw
tri 9246 -297 9260 -283 se
rect 9260 -289 9312 -283
tri 9232 -311 9246 -297 se
rect 9246 -311 9260 -297
rect 8440 -363 8446 -311
rect 8498 -363 8510 -311
rect 8562 -341 9260 -311
rect 8562 -353 9312 -341
rect 8562 -363 9260 -353
tri 9212 -411 9260 -363 ne
rect 9260 -411 9312 -405
rect 949 -480 955 -428
rect 1007 -480 1021 -428
rect 1073 -434 1375 -428
rect 1073 -468 1257 -434
rect 1291 -468 1329 -434
rect 1363 -468 1375 -434
rect 1073 -474 1375 -468
rect 1073 -480 1079 -474
tri 1079 -480 1085 -474 nw
rect -237 -513 -185 -507
tri -315 -591 -237 -513 se
rect -237 -579 -185 -565
rect -315 -597 -237 -591
tri 1960 -582 1970 -572 se
rect 1970 -578 2022 -572
rect -315 -631 -303 -597
rect -269 -631 -237 -597
rect -315 -637 -185 -631
tri 2022 -582 2032 -572 sw
rect 1970 -642 2022 -630
rect 1970 -700 2022 -694
rect 9 -864 647 -847
tri 647 -864 664 -847 sw
tri -51 -952 9 -892 ne
rect 9 -952 1411 -864
rect 1144 -1054 1171 -952
tri 1171 -1054 1273 -952 nw
tri -258 -1390 9 -1123 se
rect 7425 -1240 7705 -1234
rect 7477 -1292 7705 -1240
rect 7425 -1304 7705 -1292
rect 7477 -1314 7705 -1304
tri 7705 -1314 7785 -1234 sw
tri 8398 -1314 8410 -1302 se
rect 7477 -1356 8423 -1314
rect 7425 -1362 8423 -1356
<< rmetal1 >>
rect 7810 591 7812 592
rect 7810 391 7811 591
rect 7810 390 7812 391
rect 8112 591 8114 592
rect 8113 391 8114 591
rect 8112 390 8114 391
<< via1 >>
rect 6988 3523 7040 3575
rect 5372 3376 5424 3428
rect 5372 3312 5424 3364
rect 6988 3459 7040 3511
rect 7526 2859 7578 2911
rect 7642 2859 7694 2911
rect 9260 2745 9312 2797
rect 9260 2667 9312 2719
rect 7151 2317 7203 2369
rect 8497 2323 8549 2375
rect 8561 2323 8613 2375
rect 7151 2253 7203 2305
rect 9260 2589 9312 2641
rect 9260 2511 9312 2563
rect 9260 2432 9312 2484
rect 8768 2323 8820 2375
rect 8832 2323 8884 2375
rect 8769 2167 8821 2219
rect 8833 2167 8885 2219
rect 9456 1988 9508 2040
rect 9532 1988 9584 2040
rect 9456 1920 9508 1972
rect 9532 1920 9584 1972
rect 2129 1680 2181 1732
rect 4170 1677 4222 1729
rect 4234 1720 4286 1729
rect 4234 1686 4276 1720
rect 4276 1686 4286 1720
rect 4234 1677 4286 1686
rect 2129 1616 2181 1668
rect 7425 1596 7477 1648
rect 4433 1448 4485 1500
rect 4557 1448 4609 1500
rect 7074 1526 7126 1578
rect 7158 1526 7210 1578
rect 7242 1526 7294 1578
rect 7326 1526 7378 1578
rect 7425 1532 7477 1584
rect 9811 1591 9863 1643
rect 9811 1527 9863 1579
rect 1376 1022 1428 1074
rect 1446 1022 1498 1074
rect 1516 1022 1568 1074
rect 4433 1372 4485 1424
rect 4557 1372 4609 1424
rect 4433 1296 4485 1348
rect 4557 1296 4609 1348
rect 5361 1340 5413 1349
rect 5425 1340 5477 1349
rect 5361 1306 5392 1340
rect 5392 1306 5413 1340
rect 5425 1306 5426 1340
rect 5426 1306 5477 1340
rect 5361 1297 5413 1306
rect 5425 1297 5477 1306
rect 1376 957 1428 1009
rect 1446 957 1498 1009
rect 1516 957 1568 1009
rect 1376 892 1428 944
rect 1446 892 1498 944
rect 1516 892 1568 944
rect 1376 827 1428 879
rect 1446 827 1498 879
rect 1516 827 1568 879
rect 1376 762 1428 814
rect 1446 762 1498 814
rect 1516 762 1568 814
rect -237 553 -185 605
rect 2129 584 2181 636
rect 2129 518 2181 570
rect -237 464 -185 516
rect 4210 864 4262 916
rect 4210 800 4262 852
rect 8342 728 8394 737
rect 8342 694 8356 728
rect 8356 694 8390 728
rect 8390 694 8394 728
rect 8342 685 8394 694
rect 8406 685 8458 737
rect 9811 728 9863 767
rect 9811 715 9836 728
rect 9836 715 9863 728
rect 9811 694 9836 703
rect 9836 694 9863 703
rect 9811 651 9863 694
rect 8446 284 8498 336
rect 8510 284 8562 336
rect 1027 142 1079 194
rect 1027 65 1079 117
rect 1027 -13 1079 39
rect 4444 105 4496 157
rect 4551 105 4603 157
rect 4444 7 4496 59
rect 4551 7 4603 59
rect 8446 -363 8498 -311
rect 8510 -363 8562 -311
rect 9260 -341 9312 -289
rect 9260 -405 9312 -353
rect 955 -480 1007 -428
rect 1021 -480 1073 -428
rect -237 -565 -185 -513
rect -237 -597 -185 -579
rect -237 -631 -231 -597
rect -231 -631 -197 -597
rect -197 -631 -185 -597
rect 1970 -630 2022 -578
rect 1970 -694 2022 -642
rect 7425 -1292 7477 -1240
rect 7425 -1356 7477 -1304
<< metal2 >>
rect 6988 3575 7040 3581
rect 6988 3511 7040 3523
rect 6988 3453 7040 3459
tri 6988 3452 6989 3453 ne
rect 5372 3428 5424 3434
rect 5372 3364 5424 3376
rect 5372 2970 5424 3312
tri 5372 2918 5424 2970 ne
tri 5424 2933 5483 2992 sw
rect 5424 2918 5483 2933
tri 5424 2911 5431 2918 ne
rect 2129 1732 2181 1738
rect 2129 1668 2181 1680
rect 4164 1677 4170 1729
rect 4222 1677 4234 1729
rect 4286 1677 4292 1729
tri 4164 1648 4193 1677 ne
rect 4193 1648 4263 1677
tri 4263 1648 4292 1677 nw
tri 4193 1631 4210 1648 ne
rect 1376 1074 1568 1080
rect 1428 1022 1446 1074
rect 1498 1022 1516 1074
rect 1376 1009 1568 1022
rect 1428 957 1446 1009
rect 1498 957 1516 1009
rect 1376 944 1568 957
rect 1428 892 1446 944
rect 1498 892 1516 944
rect 1376 879 1568 892
rect 1428 827 1446 879
rect 1498 827 1516 879
rect 1376 814 1568 827
rect 1428 762 1446 814
rect 1498 762 1516 814
rect 1376 756 1568 762
rect 2129 636 2181 1616
rect 4210 916 4262 1648
tri 4262 1647 4263 1648 nw
rect 4210 852 4262 864
rect 4210 794 4262 800
rect 4433 1500 4609 1506
rect 4485 1448 4557 1500
rect 4433 1424 4609 1448
rect 4485 1372 4557 1424
rect 4433 1348 4609 1372
rect 4485 1296 4557 1348
rect -237 605 -185 611
rect -237 516 -185 553
rect -237 -513 -185 464
rect 2129 570 2181 584
rect 1027 194 1079 200
rect 1027 117 1079 142
rect 1027 39 1079 65
tri 1014 -363 1027 -350 se
rect 1027 -363 1079 -13
tri 2055 -109 2129 -35 se
rect 2129 -57 2181 518
rect 4433 157 4609 1296
tri 5355 1355 5431 1431 se
rect 5431 1355 5483 2918
rect 6989 2566 7040 3453
rect 7520 2859 7526 2911
rect 7578 2859 7642 2911
rect 7694 2859 7700 2911
rect 9260 2797 9312 2803
rect 9260 2719 9312 2745
rect 9260 2641 9312 2667
tri 7040 2566 7041 2567 sw
rect 6989 2563 7041 2566
tri 7041 2563 7044 2566 sw
rect 9260 2563 9312 2589
rect 6989 2537 7044 2563
tri 6989 2511 7015 2537 ne
rect 7015 2511 7044 2537
tri 7044 2511 7096 2563 sw
tri 7015 2485 7041 2511 ne
rect 7041 2485 7096 2511
tri 7096 2485 7122 2511 sw
tri 7041 2484 7042 2485 ne
rect 7042 2484 7122 2485
tri 7122 2484 7123 2485 sw
rect 9260 2484 9312 2511
tri 7042 2432 7094 2484 ne
rect 7094 2432 7123 2484
tri 7123 2432 7175 2484 sw
tri 7094 2404 7122 2432 ne
rect 7122 2404 7175 2432
tri 7175 2404 7203 2432 sw
tri 7122 2375 7151 2404 ne
rect 7151 2369 7203 2404
rect 8491 2323 8497 2375
rect 8549 2323 8561 2375
rect 8613 2323 8768 2375
rect 8820 2323 8832 2375
rect 8884 2323 8890 2375
rect 7151 2305 7203 2317
rect 7151 2247 7203 2253
rect 8763 2167 8769 2219
rect 8821 2167 8833 2219
rect 8885 2167 8891 2219
tri 8763 2110 8820 2167 ne
rect 7425 1648 7477 1654
rect 7425 1584 7477 1596
rect 7068 1526 7074 1578
rect 7126 1526 7158 1578
rect 7210 1526 7242 1578
rect 7294 1526 7326 1578
rect 7378 1526 7384 1578
rect 5355 1349 5483 1355
rect 5355 1297 5361 1349
rect 5413 1297 5425 1349
rect 5477 1297 5483 1349
rect 5355 1291 5483 1297
rect 4433 105 4444 157
rect 4496 105 4551 157
rect 4603 105 4609 157
rect 4433 59 4609 105
rect 4433 7 4444 59
rect 4496 7 4551 59
rect 4603 7 4609 59
rect 4433 6 4609 7
tri 2129 -109 2181 -57 nw
tri 1981 -183 2055 -109 se
tri 2055 -183 2129 -109 nw
tri 972 -405 1014 -363 se
rect 1014 -405 1079 -363
tri 949 -428 972 -405 se
rect 972 -428 1079 -405
rect 949 -480 955 -428
rect 1007 -480 1021 -428
rect 1073 -480 1079 -428
tri 1970 -194 1981 -183 se
rect 1981 -194 2022 -183
rect -237 -579 -185 -565
rect -237 -637 -185 -631
rect 1970 -578 2022 -194
tri 2022 -216 2055 -183 nw
rect 1970 -642 2022 -630
rect 1970 -700 2022 -694
rect 7425 -1240 7477 1532
tri 8746 788 8820 862 se
rect 8820 840 8872 2167
tri 8872 2148 8891 2167 nw
tri 8820 788 8872 840 nw
tri 8725 767 8746 788 se
rect 8746 767 8799 788
tri 8799 767 8820 788 nw
tri 8695 737 8725 767 se
rect 8725 737 8769 767
tri 8769 737 8799 767 nw
rect 8336 685 8342 737
rect 8394 685 8406 737
rect 8458 715 8747 737
tri 8747 715 8769 737 nw
rect 8458 703 8735 715
tri 8735 703 8747 715 nw
rect 8458 685 8717 703
tri 8717 685 8735 703 nw
rect 8440 284 8446 336
rect 8498 284 8510 336
rect 8562 284 8568 336
tri 8440 246 8478 284 ne
tri 8462 -289 8478 -273 se
rect 8478 -289 8530 284
tri 8530 246 8568 284 nw
tri 8530 -289 8546 -273 sw
rect 9260 -289 9312 2432
rect 9456 2040 9584 2046
rect 9508 1988 9532 2040
rect 9456 1972 9584 1988
rect 9508 1920 9532 1972
rect 9456 1914 9584 1920
rect 9811 1643 9863 1649
rect 9811 1579 9863 1591
rect 9811 767 9863 1527
rect 9811 703 9863 715
rect 9811 645 9863 651
tri 8440 -311 8462 -289 se
rect 8462 -311 8546 -289
tri 8546 -311 8568 -289 sw
rect 8440 -363 8446 -311
rect 8498 -363 8510 -311
rect 8562 -363 8568 -311
rect 9260 -353 9312 -341
rect 9260 -411 9312 -405
rect 7425 -1304 7477 -1292
rect 7425 -1362 7477 -1356
use nfet_CDNS_524688791851224  nfet_CDNS_524688791851224_0
timestamp 1704896540
transform -1 0 4626 0 1 75
box -98 -32 282 182
use nfet_CDNS_524688791851225  nfet_CDNS_524688791851225_0
timestamp 1704896540
transform -1 0 4898 0 1 -138
box -82 -32 282 116
use nfet_CDNS_524688791851226  nfet_CDNS_524688791851226_0
timestamp 1704896540
transform -1 0 4898 0 1 75
box -82 -32 282 232
use nfet_CDNS_524688791851227  nfet_CDNS_524688791851227_0
timestamp 1704896540
transform -1 0 4890 0 1 394
box -82 -32 538 632
use nfet_CDNS_524688791851228  nfet_CDNS_524688791851228_0
timestamp 1704896540
transform 1 0 5779 0 1 1290
box -82 -32 262 232
use nfet_CDNS_524688791851229  nfet_CDNS_524688791851229_0
timestamp 1704896540
transform 1 0 4835 0 1 1290
box -82 -32 970 232
use nfet_CDNS_524688791851230  nfet_CDNS_524688791851230_0
timestamp 1704896540
transform 0 -1 9488 1 0 1968
box -82 -32 282 632
use nfet_CDNS_524688791851231  nfet_CDNS_524688791851231_0
timestamp 1704896540
transform 1 0 3270 0 1 132
box -82 -32 494 232
use nfet_CDNS_524688791851232  nfet_CDNS_524688791851232_0
timestamp 1704896540
transform 1 0 2958 0 1 132
box -82 -32 338 232
use nfet_CDNS_524688791851233  nfet_CDNS_524688791851233_0
timestamp 1704896540
transform 1 0 2646 0 1 132
box -82 -32 338 232
use nfet_CDNS_524688791851234  nfet_CDNS_524688791851234_0
timestamp 1704896540
transform -1 0 5600 0 1 46
box -82 -32 494 1032
use nfet_CDNS_524688791851235  nfet_CDNS_524688791851235_0
timestamp 1704896540
transform -1 0 6112 0 1 46
box -82 -32 538 1032
use nfet_CDNS_524688791851236  nfet_CDNS_524688791851236_0
timestamp 1704896540
transform 1 0 8960 0 -1 1376
box -82 -32 1082 632
use nfet_CDNS_524688791851236  nfet_CDNS_524688791851236_1
timestamp 1704896540
transform 1 0 8960 0 1 46
box -82 -32 1082 632
use nfet_CDNS_524688791851237  nfet_CDNS_524688791851237_0
timestamp 1704896540
transform 1 0 6400 0 -1 1376
box -82 -32 2586 632
use nfet_CDNS_524688791851237  nfet_CDNS_524688791851237_1
timestamp 1704896540
transform 1 0 6400 0 1 46
box -82 -32 2586 632
use pfet_CDNS_524688791851212  pfet_CDNS_524688791851212_0
timestamp 1704896540
transform 0 1 -357 1 0 -842
box -119 -66 322 1066
use pfet_CDNS_524688791851213  pfet_CDNS_524688791851213_0
timestamp 1704896540
transform 0 -1 1392 -1 0 -459
box -122 -66 519 216
use pfet_CDNS_524688791851214  pfet_CDNS_524688791851214_0
timestamp 1704896540
transform 1 0 4263 0 1 1305
box -119 -66 375 216
use pfet_CDNS_524688791851215  pfet_CDNS_524688791851215_0
timestamp 1704896540
transform 0 -1 2173 1 0 1191
box -122 -66 498 1066
use pfet_CDNS_524688791851216  pfet_CDNS_524688791851216_0
timestamp 1704896540
transform 1 0 3270 0 -1 1383
box -122 -66 534 666
use pfet_CDNS_524688791851217  pfet_CDNS_524688791851217_0
timestamp 1704896540
transform 1 0 2802 0 -1 1383
box -122 -66 222 666
use pfet_CDNS_524688791851218  pfet_CDNS_524688791851218_0
timestamp 1704896540
transform 1 0 2366 0 -1 1383
box -122 -66 378 666
use pfet_CDNS_524688791851218  pfet_CDNS_524688791851218_1
timestamp 1704896540
transform 1 0 2958 0 -1 1383
box -122 -66 378 666
use pfet_CDNS_524688791851219  pfet_CDNS_524688791851219_0
timestamp 1704896540
transform 0 1 8893 1 0 2487
box -122 -66 378 666
use pfet_CDNS_524688791851220  pfet_CDNS_524688791851220_0
timestamp 1704896540
transform 1 0 1872 0 -1 920
box -122 -66 378 1066
use pfet_CDNS_524688791851221  pfet_CDNS_524688791851221_0
timestamp 1704896540
transform 1 0 1124 0 -1 920
box -122 -66 690 1066
use pfet_CDNS_524688791851222  pfet_CDNS_524688791851222_0
timestamp 1704896540
transform 1 0 49 0 1 -112
box -122 -66 282 1466
use pfet_CDNS_524688791851223  pfet_CDNS_524688791851223_0
timestamp 1704896540
transform 1 0 265 0 1 -112
box -122 -66 714 1466
use sky130_fd_io__hvsbt_inv_x1_sio  sky130_fd_io__hvsbt_inv_x1_sio_0
timestamp 1704896540
transform -1 0 4107 0 1 306
box 0 -192 358 1016
use sky130_fd_io__tk_em1o_CDNS_524688791851211  sky130_fd_io__tk_em1o_CDNS_524688791851211_0
timestamp 1704896540
transform 1 0 7758 0 1 390
box 0 0 1 1
<< labels >>
flabel comment s 5942 1116 5942 1116 0 FreeSans 400 180 0 0 in_h
flabel comment s 9819 707 9819 707 0 FreeSans 440 180 0 0 en_h
flabel comment s 8472 725 8472 725 0 FreeSans 400 180 0 0 in_vt
flabel metal1 s 9224 1942 9224 1942 0 FreeSans 200 0 0 0 vgnd
flabel metal1 s 4991 1326 4991 1326 0 FreeSans 200 0 0 0 a
flabel metal1 s 9195 2534 9195 2534 0 FreeSans 200 0 0 0 b
flabel metal1 s 8967 2614 8967 2614 0 FreeSans 200 0 0 0 a
flabel metal1 s 8831 2622 8831 2622 0 FreeSans 200 90 0 0 vtrip_sel_h
flabel metal1 s 1454 1300 1454 1300 3 FreeSans 520 0 0 0 vcc_io
flabel metal1 s 956 -904 956 -904 0 FreeSans 44 0 0 0 vgnd
flabel metal1 s 5292 1544 5336 1572 3 FreeSans 520 0 0 0 vpwr
port 3 nsew
flabel metal1 s 3235 571 3287 588 3 FreeSans 520 0 0 0 out_h_n
port 4 nsew
flabel metal1 s 85 861 205 981 3 FreeSans 520 0 0 0 vcc_io
port 2 nsew
flabel metal1 s 4715 118 4715 118 0 FreeSans 440 0 0 0 vcc_io
flabel metal1 s 9643 441 9836 553 3 FreeSans 520 0 0 0 vgnd
port 1 nsew
flabel metal1 s 9655 497 9655 497 3 FreeSans 520 0 0 0 vgnd
flabel metal1 s 9643 867 9836 979 3 FreeSans 520 0 0 0 vgnd
port 1 nsew
flabel metal1 s 1383 317 1383 317 0 FreeSans 200 0 0 0 b
flabel metal1 s 9636 692 9691 724 3 FreeSans 520 0 0 0 en_h
port 8 nsew
flabel metal1 s 8256 693 8326 727 3 FreeSans 520 0 0 0 in_vt
port 5 nsew
flabel metal1 s 3939 122 3939 122 0 FreeSans 200 0 0 0 vgnd
flabel metal1 s 5803 1111 5803 1111 3 FreeSans 520 0 0 0 in_h
flabel metal1 s 3693 474 3731 581 3 FreeSans 520 0 0 0 out_h
port 7 nsew
flabel metal1 s 2817 1338 2817 1338 3 FreeSans 520 0 0 0 vcc_io
flabel metal1 s 2652 73 2772 193 3 FreeSans 520 0 0 0 vgnd
port 1 nsew
flabel locali s 3909 664 3955 701 3 FreeSans 520 0 0 0 vtrip_sel_h_n
port 9 nsew
flabel locali s 9396 2924 9396 2924 0 FreeSans 200 0 0 0 vcc_io
flabel locali s 3835 801 3835 801 3 FreeSans 520 90 0 0 vtrip_sel_h
<< properties >>
string GDS_END 85750782
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85638434
string path 245.925 16.125 245.925 19.325 
<< end >>
