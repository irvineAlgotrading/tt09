magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< pwell >>
rect -76 -26 204 1426
<< nmos >>
rect 0 0 36 1400
rect 92 0 128 1400
<< ndiff >>
rect -50 0 0 1400
rect 128 0 178 1400
<< poly >>
rect 0 1400 36 1432
rect 0 -32 36 0
rect 92 1400 128 1432
rect 92 -32 128 0
<< locali >>
rect -45 -4 -11 1354
rect 47 -4 81 1354
rect 139 -4 173 1354
use DFL1sd2_CDNS_55959141808679  DFL1sd2_CDNS_55959141808679_0
timestamp 1704896540
transform -1 0 0 0 1 0
box -26 -26 82 1426
use DFL1sd2_CDNS_55959141808679  DFL1sd2_CDNS_55959141808679_1
timestamp 1704896540
transform 1 0 36 0 1 0
box -26 -26 82 1426
use DFL1sd2_CDNS_55959141808679  DFL1sd2_CDNS_55959141808679_2
timestamp 1704896540
transform 1 0 128 0 1 0
box -26 -26 82 1426
<< labels >>
flabel comment s 156 675 156 675 0 FreeSans 300 0 0 0 S
flabel comment s 64 675 64 675 0 FreeSans 300 0 0 0 D
flabel comment s -28 675 -28 675 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 2733002
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 2731678
<< end >>
