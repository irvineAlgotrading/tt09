magic
tech sky130B
timestamp 1704896540
<< pwell >>
rect -13 -13 72 960
<< ndiff >>
rect 0 941 59 947
rect 0 6 4 941
rect 55 6 59 941
rect 0 0 59 6
<< ndiffc >>
rect 4 6 55 941
<< locali >>
rect 4 941 55 949
rect 4 -2 55 6
<< properties >>
string GDS_END 34406062
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 34402282
<< end >>
