magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< pwell >>
rect -68 -26 1803 92
<< ndiff >>
rect -42 50 0 66
rect -42 16 -34 50
rect -42 0 0 16
rect 1735 50 1777 66
rect 1769 16 1777 50
rect 1735 0 1777 16
<< ndiffc >>
rect -34 16 0 50
rect 1735 16 1769 50
<< ndiffres >>
rect 0 0 1735 66
<< locali >>
rect -34 50 0 66
rect -34 0 0 16
rect 1735 50 1769 66
rect 1735 0 1769 16
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_0
timestamp 1704896540
transform -1 0 8 0 1 4
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_1
timestamp 1704896540
transform 1 0 1727 0 1 4
box 0 0 1 1
<< properties >>
string GDS_END 79940140
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 79939638
<< end >>
