magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -38 261 498 582
<< pwell >>
rect 1 21 459 203
rect 29 -17 63 21
<< locali >>
rect 167 409 267 493
rect 17 133 65 398
rect 99 367 267 409
rect 99 165 133 367
rect 167 283 247 333
rect 305 323 345 481
rect 281 289 345 323
rect 167 199 201 283
rect 281 249 317 289
rect 244 215 317 249
rect 351 215 443 255
rect 99 129 169 165
<< obsli1 >>
rect 0 527 460 561
rect 27 435 69 527
rect 379 291 443 527
rect 237 165 443 173
rect 203 139 443 165
rect 203 95 269 139
rect 17 59 269 95
rect 307 17 341 105
rect 375 56 443 139
rect 0 -17 460 17
<< metal1 >>
rect 0 496 460 592
rect 0 -48 460 48
<< labels >>
rlabel locali s 351 215 443 255 6 A1
port 1 nsew signal input
rlabel locali s 244 215 317 249 6 A2
port 2 nsew signal input
rlabel locali s 281 249 317 289 6 A2
port 2 nsew signal input
rlabel locali s 281 289 345 323 6 A2
port 2 nsew signal input
rlabel locali s 305 323 345 481 6 A2
port 2 nsew signal input
rlabel locali s 17 133 65 398 6 B1
port 3 nsew signal input
rlabel locali s 167 199 201 283 6 B2
port 4 nsew signal input
rlabel locali s 167 283 247 333 6 B2
port 4 nsew signal input
rlabel metal1 s 0 -48 460 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1 21 459 203 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 498 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 460 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 99 129 169 165 6 Y
port 9 nsew signal output
rlabel locali s 99 165 133 367 6 Y
port 9 nsew signal output
rlabel locali s 99 367 267 409 6 Y
port 9 nsew signal output
rlabel locali s 167 409 267 493 6 Y
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 460 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1375324
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1370488
<< end >>
