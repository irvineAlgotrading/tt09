magic
tech sky130A
timestamp 1704896540
<< properties >>
string GDS_END 92017378
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 92016610
<< end >>
