magic
tech sky130B
timestamp 1704896540
<< viali >>
rect 0 0 161 53
<< metal1 >>
rect -6 53 167 56
rect -6 0 0 53
rect 161 0 167 53
rect -6 -3 167 0
<< properties >>
string GDS_END 95638648
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 95637876
<< end >>
