magic
tech sky130A
magscale 1 2
timestamp 1704896540
use sky130_fd_pr__hvdfm1sd2__example_5595914180849  sky130_fd_pr__hvdfm1sd2__example_5595914180849_0
timestamp 1704896540
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd__example_5595914180848  sky130_fd_pr__hvdfm1sd__example_5595914180848_0
timestamp 1704896540
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd__example_5595914180848  sky130_fd_pr__hvdfm1sd__example_5595914180848_1
timestamp 1704896540
transform 1 0 256 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 74523238
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 74521668
<< end >>
