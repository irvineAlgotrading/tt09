magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< obsli1 >>
rect 214 200 14555 39939
<< obsm1 >>
rect 222 194 14724 39945
<< metal2 >>
rect 187 38112 13440 39015
rect 2824 37931 3019 38112
rect 187 37917 3019 37931
rect 187 37011 2824 37917
rect 187 37005 3054 37011
rect 2824 36781 3054 37005
rect 187 36771 3064 36781
rect 187 36758 3162 36771
rect 3064 36673 3162 36758
rect 3162 36571 3264 36673
rect 3264 36445 3390 36571
rect 3390 36296 3539 36445
rect 187 34556 11592 36296
rect 3211 34231 3536 34556
rect 2824 34214 3211 34231
rect 187 33844 3211 34214
rect 12222 34225 14858 37065
rect 187 31696 2824 33844
rect 12222 32491 14858 32497
rect 11505 31774 14858 32491
rect 187 29956 11341 31696
rect 3212 29631 3537 29956
rect 12222 29631 14858 31774
rect 2824 29449 3212 29631
rect 3361 29622 14858 29631
rect 187 29243 3212 29449
rect 3361 29342 3650 29622
rect 187 13550 2824 29243
rect 12222 27891 14858 27897
rect 11502 27171 14858 27891
rect 12222 25025 14858 27171
rect 12222 23291 14858 23297
rect 11495 22564 14858 23291
rect 12222 20425 14858 22564
rect 12222 18691 14858 18697
rect 11513 17982 14858 18691
rect 12222 15825 14858 17982
rect 4964 15123 14858 15133
rect 4724 15121 14858 15123
rect 4724 14883 4964 15121
rect 3682 14831 14858 14883
rect 4730 14611 4964 14831
rect 4730 14597 14858 14611
rect 3230 13296 3533 13599
rect 187 11556 11342 13296
rect 3212 11231 3537 11556
rect 12222 11231 14858 14097
rect 2824 10857 3212 11231
rect 3492 11219 14858 11231
rect 187 10843 3212 10857
rect 3492 10953 3770 11219
rect 187 8476 2824 9105
rect 187 8070 10840 8476
rect 3629 7735 3978 8070
rect 187 7721 3978 7735
rect 3205 7297 3629 7721
rect 10515 7756 10829 8070
rect 10829 7670 10934 7756
rect 10829 7651 11383 7670
rect 3041 7147 3205 7297
rect 187 7133 3205 7147
rect 10934 7223 11383 7651
rect 187 5863 3041 7133
rect 12222 6191 14858 9497
rect 187 5854 3764 5863
rect 3041 5140 3764 5854
rect 187 2480 7379 5140
rect 4879 2212 5640 2480
rect 11163 5132 14858 6191
rect 187 1719 5640 2212
rect 187 1513 4879 1719
rect 187 411 4879 985
rect 99 0 4879 411
rect 5179 0 5579 197
rect 10078 0 14858 5132
<< obsm2 >>
rect 99 38056 131 38112
rect 99 37987 2768 38056
rect 99 36949 131 37987
rect 13496 38056 14858 38112
rect 3075 37861 14858 38056
rect 2880 37121 14858 37861
rect 2880 37067 12166 37121
rect 99 36837 2768 36949
rect 99 36702 131 36837
rect 3110 36837 12166 37067
rect 3120 36827 12166 36837
rect 99 36617 3008 36702
rect 3218 36729 12166 36827
rect 99 36515 3106 36617
rect 3320 36627 12166 36729
rect 99 36389 3208 36515
rect 3446 36501 12166 36627
rect 99 36352 3334 36389
rect 99 34500 131 36352
rect 3595 36352 12166 36501
rect 99 34287 3155 34500
rect 99 34270 2768 34287
rect 99 29900 131 34270
rect 11648 34500 12166 36352
rect 3592 34175 12166 34500
rect 3267 34169 12166 34175
rect 3267 33788 14858 34169
rect 2880 32553 14858 33788
rect 2880 32547 12166 32553
rect 2880 31752 11449 32547
rect 11397 31718 11449 31752
rect 99 29687 3156 29900
rect 99 29505 2768 29687
rect 11397 29900 12166 31718
rect 3593 29687 12166 29900
rect 99 13494 131 29505
rect 3268 29286 3305 29575
rect 3706 29286 14858 29566
rect 3268 29187 14858 29286
rect 2880 27953 14858 29187
rect 2880 27947 12166 27953
rect 2880 27115 11446 27947
rect 2880 24969 12166 27115
rect 2880 23353 14858 24969
rect 2880 23347 12166 23353
rect 2880 22508 11439 23347
rect 2880 20369 12166 22508
rect 2880 18753 14858 20369
rect 2880 18747 12166 18753
rect 2880 17926 11457 18747
rect 2880 15769 12166 17926
rect 2880 15189 14858 15769
rect 2880 15179 4908 15189
rect 2880 14939 4668 15179
rect 2880 14775 3626 14939
rect 5020 14939 14858 15065
rect 2880 14541 4674 14775
rect 5020 14667 14858 14775
rect 2880 14153 14858 14541
rect 2880 13655 12166 14153
rect 2880 13494 3174 13655
rect 99 13352 3174 13494
rect 99 11500 131 13352
rect 3589 13352 12166 13655
rect 99 11287 3156 11500
rect 99 10913 2768 11287
rect 11398 11500 12166 13352
rect 3593 11287 12166 11500
rect 99 10787 131 10913
rect 3268 10897 3436 11175
rect 3826 10897 14858 11163
rect 3268 10787 14858 10897
rect 99 9553 14858 10787
rect 99 9161 12166 9553
rect 99 8014 131 9161
rect 2880 8532 12166 9161
rect 99 7791 3573 8014
rect 99 7665 131 7791
rect 99 7353 3149 7665
rect 99 7203 2985 7353
rect 4034 7700 10459 8014
rect 10896 8014 12166 8532
rect 10885 7812 12166 8014
rect 4034 7665 10773 7700
rect 3685 7595 10773 7665
rect 10990 7726 12166 7812
rect 99 5798 131 7203
rect 3685 7241 10878 7595
rect 3261 7167 10878 7241
rect 11439 7167 12166 7726
rect 3261 7077 12166 7167
rect 3097 6247 12166 7077
rect 3097 5919 11107 6247
rect 99 5196 2985 5798
rect 99 2424 131 5196
rect 3820 5196 11107 5919
rect 7435 5188 11107 5196
rect 99 2268 4823 2424
rect 99 1457 131 2268
rect 7435 2424 10022 5188
rect 5696 1663 10022 2424
rect 4935 1457 10022 1663
rect 99 1041 10022 1457
rect 99 467 131 1041
tri 155 467 187 499 se
tri 99 411 155 467 se
rect 155 411 187 467
rect 4935 253 10022 1041
rect 4935 197 5123 253
rect 5635 197 10022 253
<< metal3 >>
rect 5179 0 7379 2485
rect 7578 0 9778 2476
<< obsm3 >>
rect 2525 2565 12298 39015
rect 2525 2476 5099 2565
rect 7459 2556 12298 2565
rect 7459 2476 7498 2556
rect 9858 2476 12298 2556
<< labels >>
rlabel metal3 s 5179 0 7379 2485 6 src_bdy_hvc
port 1 nsew ground bidirectional
rlabel metal2 s 99 0 4879 411 6 src_bdy_hvc
port 1 nsew ground bidirectional
rlabel metal2 s 187 411 4879 985 6 src_bdy_hvc
port 1 nsew ground bidirectional
rlabel metal2 s 4879 1719 5640 2480 6 src_bdy_hvc
port 1 nsew ground bidirectional
rlabel metal2 s 187 1513 4879 2212 6 src_bdy_hvc
port 1 nsew ground bidirectional
rlabel metal2 s 187 2480 7379 5140 6 src_bdy_hvc
port 1 nsew ground bidirectional
rlabel metal2 s 187 5854 3041 5863 6 src_bdy_hvc
port 1 nsew ground bidirectional
rlabel metal2 s 3041 5140 3764 5863 6 src_bdy_hvc
port 1 nsew ground bidirectional
rlabel metal2 s 187 5863 3041 7133 6 src_bdy_hvc
port 1 nsew ground bidirectional
rlabel metal2 s 187 7133 3041 7147 6 src_bdy_hvc
port 1 nsew ground bidirectional
rlabel metal2 s 3041 7133 3205 7297 6 src_bdy_hvc
port 1 nsew ground bidirectional
rlabel metal2 s 3205 7297 3629 7721 6 src_bdy_hvc
port 1 nsew ground bidirectional
rlabel metal2 s 187 7721 3629 7735 6 src_bdy_hvc
port 1 nsew ground bidirectional
rlabel metal2 s 3629 7721 3978 8070 6 src_bdy_hvc
port 1 nsew ground bidirectional
rlabel metal2 s 10934 7223 11383 7651 6 src_bdy_hvc
port 1 nsew ground bidirectional
rlabel metal2 s 10515 7756 10829 8070 6 src_bdy_hvc
port 1 nsew ground bidirectional
rlabel metal2 s 10829 7651 10934 7756 6 src_bdy_hvc
port 1 nsew ground bidirectional
rlabel metal2 s 10934 7651 11383 7670 6 src_bdy_hvc
port 1 nsew ground bidirectional
rlabel metal2 s 187 8070 10840 8476 6 src_bdy_hvc
port 1 nsew ground bidirectional
rlabel metal2 s 187 8476 2824 9105 6 src_bdy_hvc
port 1 nsew ground bidirectional
rlabel metal2 s 3212 11231 3537 11556 6 src_bdy_hvc
port 1 nsew ground bidirectional
rlabel metal2 s 2824 10843 3212 11231 6 src_bdy_hvc
port 1 nsew ground bidirectional
rlabel metal2 s 187 10843 2824 10857 6 src_bdy_hvc
port 1 nsew ground bidirectional
rlabel metal2 s 187 11556 11342 13296 6 src_bdy_hvc
port 1 nsew ground bidirectional
rlabel metal2 s 187 13550 2824 29449 6 src_bdy_hvc
port 1 nsew ground bidirectional
rlabel metal2 s 3230 13296 3533 13599 6 src_bdy_hvc
port 1 nsew ground bidirectional
rlabel metal2 s 3212 29631 3537 29956 6 src_bdy_hvc
port 1 nsew ground bidirectional
rlabel metal2 s 2824 29243 3212 29631 6 src_bdy_hvc
port 1 nsew ground bidirectional
rlabel metal2 s 187 29956 11341 31696 6 src_bdy_hvc
port 1 nsew ground bidirectional
rlabel metal2 s 187 31696 2824 33466 6 src_bdy_hvc
port 1 nsew ground bidirectional
rlabel metal2 s 3211 34231 3536 34556 6 src_bdy_hvc
port 1 nsew ground bidirectional
rlabel metal2 s 2824 33844 3211 34231 6 src_bdy_hvc
port 1 nsew ground bidirectional
rlabel metal2 s 187 33466 2824 34214 6 src_bdy_hvc
port 1 nsew ground bidirectional
rlabel metal2 s 187 34556 11592 36296 6 src_bdy_hvc
port 1 nsew ground bidirectional
rlabel metal2 s 187 36758 3064 36771 6 src_bdy_hvc
port 1 nsew ground bidirectional
rlabel metal2 s 3064 36673 3162 36771 6 src_bdy_hvc
port 1 nsew ground bidirectional
rlabel metal2 s 3162 36571 3264 36673 6 src_bdy_hvc
port 1 nsew ground bidirectional
rlabel metal2 s 3264 36445 3390 36571 6 src_bdy_hvc
port 1 nsew ground bidirectional
rlabel metal2 s 3390 36296 3539 36445 6 src_bdy_hvc
port 1 nsew ground bidirectional
rlabel metal2 s 187 36771 3064 36781 6 src_bdy_hvc
port 1 nsew ground bidirectional
rlabel metal2 s 187 37005 2824 37011 6 src_bdy_hvc
port 1 nsew ground bidirectional
rlabel metal2 s 2824 36781 3054 37011 6 src_bdy_hvc
port 1 nsew ground bidirectional
rlabel metal2 s 187 37011 2824 37917 6 src_bdy_hvc
port 1 nsew ground bidirectional
rlabel metal2 s 2824 37917 3019 38112 6 src_bdy_hvc
port 1 nsew ground bidirectional
rlabel metal2 s 187 37917 2824 37931 6 src_bdy_hvc
port 1 nsew ground bidirectional
rlabel metal2 s 187 38112 13440 39015 6 src_bdy_hvc
port 1 nsew ground bidirectional
rlabel metal3 s 7578 0 9778 2476 6 drn_hvc
port 2 nsew power bidirectional
rlabel metal2 s 10078 0 14858 5132 6 drn_hvc
port 2 nsew power bidirectional
rlabel metal2 s 11163 5132 12222 6191 6 drn_hvc
port 2 nsew power bidirectional
rlabel metal2 s 12222 5132 14858 9497 6 drn_hvc
port 2 nsew power bidirectional
rlabel metal2 s 3770 11219 14858 11231 6 drn_hvc
port 2 nsew power bidirectional
rlabel metal2 s 3492 10953 3770 11231 6 drn_hvc
port 2 nsew power bidirectional
rlabel metal2 s 12222 11231 14858 14097 6 drn_hvc
port 2 nsew power bidirectional
rlabel metal2 s 4730 14597 4964 14831 6 drn_hvc
port 2 nsew power bidirectional
rlabel metal2 s 4964 14597 14858 14611 6 drn_hvc
port 2 nsew power bidirectional
rlabel metal2 s 3682 14831 14858 14883 6 drn_hvc
port 2 nsew power bidirectional
rlabel metal2 s 4964 15121 14858 15133 6 drn_hvc
port 2 nsew power bidirectional
rlabel metal2 s 4724 14883 4964 15123 6 drn_hvc
port 2 nsew power bidirectional
rlabel metal2 s 12222 15825 14858 17792 6 drn_hvc
port 2 nsew power bidirectional
rlabel metal2 s 11513 17982 12222 18691 6 drn_hvc
port 2 nsew power bidirectional
rlabel metal2 s 12222 17792 14858 18697 6 drn_hvc
port 2 nsew power bidirectional
rlabel metal2 s 12222 20425 14858 22392 6 drn_hvc
port 2 nsew power bidirectional
rlabel metal2 s 11495 22564 12222 23291 6 drn_hvc
port 2 nsew power bidirectional
rlabel metal2 s 12222 22392 14858 23297 6 drn_hvc
port 2 nsew power bidirectional
rlabel metal2 s 12222 25025 14858 26992 6 drn_hvc
port 2 nsew power bidirectional
rlabel metal2 s 11502 27171 12222 27891 6 drn_hvc
port 2 nsew power bidirectional
rlabel metal2 s 12222 26992 14858 27897 6 drn_hvc
port 2 nsew power bidirectional
rlabel metal2 s 3650 29622 14858 29631 6 drn_hvc
port 2 nsew power bidirectional
rlabel metal2 s 3361 29342 3650 29631 6 drn_hvc
port 2 nsew power bidirectional
rlabel metal2 s 12222 29631 14858 31606 6 drn_hvc
port 2 nsew power bidirectional
rlabel metal2 s 11505 31774 12222 32491 6 drn_hvc
port 2 nsew power bidirectional
rlabel metal2 s 12222 31606 14858 32497 6 drn_hvc
port 2 nsew power bidirectional
rlabel metal2 s 12222 34225 14858 37065 6 drn_hvc
port 2 nsew power bidirectional
rlabel metal2 s 5179 0 5579 197 6 ogc_hvc
port 3 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 15000 40000
string LEFclass BLOCK
string LEFsymmetry R90
string LEFview TRUE
string GDS_END 38322748
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 34527630
<< end >>
