magic
tech sky130B
timestamp 1704896540
<< metal1 >>
rect 0 0 3 58
rect 189 0 192 58
<< via1 >>
rect 3 0 189 58
<< metal2 >>
rect 0 0 3 58
rect 189 0 192 58
<< properties >>
string GDS_END 85516634
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85515734
<< end >>
