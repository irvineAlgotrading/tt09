magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -36 -36 92 236
<< pdiff >>
rect 0 182 56 200
rect 0 148 11 182
rect 45 148 56 182
rect 0 114 56 148
rect 0 80 11 114
rect 45 80 56 114
rect 0 46 56 80
rect 0 12 11 46
rect 45 12 56 46
rect 0 0 56 12
<< pdiffc >>
rect 11 148 45 182
rect 11 80 45 114
rect 11 12 45 46
<< locali >>
rect 11 182 45 198
rect 11 114 45 140
rect 11 46 45 68
<< viali >>
rect 11 148 45 174
rect 11 140 45 148
rect 11 80 45 102
rect 11 68 45 80
rect 11 12 45 30
rect 11 -4 45 12
<< metal1 >>
rect 5 174 51 186
rect 5 140 11 174
rect 45 140 51 174
rect 5 102 51 140
rect 5 68 11 102
rect 45 68 51 102
rect 5 30 51 68
rect 5 -4 11 30
rect 45 -4 51 30
rect 5 -16 51 -4
<< properties >>
string GDS_END 6086264
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 6085556
<< end >>
