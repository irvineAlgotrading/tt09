magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< metal2 >>
rect 0 9025 536 9034
rect 0 0 536 9
<< via2 >>
rect 0 9 536 9025
<< metal3 >>
rect -5 9025 541 9030
rect -5 9 0 9025
rect 536 9 541 9025
rect -5 4 541 9
<< properties >>
string GDS_END 93578804
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 93528048
<< end >>
