magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< metal2 >>
rect 0 145 296 154
rect 0 0 296 9
<< via2 >>
rect 0 9 296 145
<< metal3 >>
rect -5 145 301 150
rect -5 9 0 145
rect 296 9 301 145
rect -5 4 301 9
<< properties >>
string GDS_END 87512382
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 87511738
<< end >>
