magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -266 -66 562 666
<< mvpmos >>
rect 0 0 120 600
rect 176 0 296 600
<< mvpdiff >>
rect -50 0 0 600
rect 296 0 346 600
<< poly >>
rect 0 600 120 632
rect 0 -32 120 0
rect 176 600 296 632
rect 176 -32 296 0
<< locali >>
rect -113 -4 -11 550
rect 131 -4 165 538
rect 307 -4 409 550
use DFL1sd2_CDNS_5246887918535  DFL1sd2_CDNS_5246887918535_0
timestamp 1704896540
transform 1 0 120 0 1 0
box -36 -36 92 636
use hvDFTPL1s_CDNS_52468879185914  hvDFTPL1s_CDNS_52468879185914_0
timestamp 1704896540
transform -1 0 0 0 1 0
box -36 -36 236 636
use hvDFTPL1s_CDNS_52468879185914  hvDFTPL1s_CDNS_52468879185914_1
timestamp 1704896540
transform 1 0 296 0 1 0
box -36 -36 236 636
<< labels >>
flabel comment s -62 273 -62 273 0 FreeSans 300 0 0 0 S
flabel comment s 148 267 148 267 0 FreeSans 300 0 0 0 D
flabel comment s 358 273 358 273 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 80520826
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 80519308
<< end >>
