magic
tech sky130B
timestamp 1704896540
<< metal1 >>
rect 0 0 3 410
rect 61 0 64 410
<< via1 >>
rect 3 0 61 410
<< metal2 >>
rect 0 0 3 410
rect 61 0 64 410
<< properties >>
string GDS_END 79840504
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 79838708
<< end >>
