magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -36 538 404 1177
<< pwell >>
rect 232 25 334 159
<< psubdiff >>
rect 258 109 308 133
rect 258 75 266 109
rect 300 75 308 109
rect 258 51 308 75
<< nsubdiff >>
rect 258 1045 308 1069
rect 258 1011 266 1045
rect 300 1011 308 1045
rect 258 987 308 1011
<< psubdiffcont >>
rect 266 75 300 109
<< nsubdiffcont >>
rect 266 1011 300 1045
<< poly >>
rect 114 555 144 819
rect 48 539 144 555
rect 48 505 64 539
rect 98 505 144 539
rect 48 489 144 505
rect 114 149 144 489
<< polycont >>
rect 64 505 98 539
<< locali >>
rect 0 1103 368 1137
rect 62 924 96 1103
rect 266 1045 300 1103
rect 266 995 300 1011
rect 64 539 98 555
rect 64 489 98 505
rect 162 539 196 990
rect 162 505 213 539
rect 162 54 196 505
rect 266 109 300 125
rect 62 17 96 54
rect 266 17 300 75
rect 0 -17 368 17
use contact_12  contact_12_0
timestamp 1704896540
transform 1 0 48 0 1 489
box 0 0 1 1
use contact_23  contact_23_0
timestamp 1704896540
transform 1 0 258 0 1 987
box 0 0 1 1
use contact_24  contact_24_0
timestamp 1704896540
transform 1 0 258 0 1 51
box 0 0 1 1
use nmos_m1_w0_360_sli_dli_da_p  nmos_m1_w0_360_sli_dli_da_p_0
timestamp 1704896540
transform 1 0 54 0 1 51
box -26 -26 176 98
use pmos_m1_w1_120_sli_dli_da_p  pmos_m1_w1_120_sli_dli_da_p_0
timestamp 1704896540
transform 1 0 54 0 1 845
box -59 -54 209 278
<< labels >>
rlabel locali s 196 522 196 522 4 Z
port 2 nsew
rlabel locali s 81 522 81 522 4 A
port 1 nsew
rlabel locali s 184 1120 184 1120 4 vdd
port 3 nsew
rlabel locali s 184 0 184 0 4 gnd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 368 1120
string GDS_END 3595660
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 3593942
<< end >>
