magic
tech sky130A
timestamp 1704896540
<< metal1 >>
rect 0 0 3 314
rect 61 0 64 314
<< via1 >>
rect 3 0 61 314
<< metal2 >>
rect 0 0 3 314
rect 61 0 64 314
<< properties >>
string GDS_END 85848684
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85847272
<< end >>
