magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< pwell >>
rect -26 -26 226 226
<< ndiff >>
rect 0 182 60 200
rect 0 148 11 182
rect 45 148 60 182
rect 0 114 60 148
rect 0 80 11 114
rect 45 80 60 114
rect 0 46 60 80
rect 0 12 11 46
rect 45 12 60 46
rect 0 0 60 12
<< ndiffc >>
rect 11 148 45 182
rect 11 80 45 114
rect 11 12 45 46
<< psubdiff >>
rect 60 126 200 200
rect 60 92 79 126
rect 113 92 200 126
rect 60 58 200 92
rect 60 24 79 58
rect 113 24 200 58
rect 60 0 200 24
<< psubdiffcont >>
rect 79 92 113 126
rect 79 24 113 58
<< locali >>
rect 11 182 113 198
rect 45 148 113 182
rect 11 126 113 148
rect 11 114 79 126
rect 45 92 79 114
rect 45 80 113 92
rect 11 58 113 80
rect 11 46 79 58
rect 45 24 79 46
rect 45 12 113 24
rect 11 -4 113 12
<< properties >>
string GDS_END 80534290
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 80533582
<< end >>
