magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect 286 1012 904 2076
rect 286 1004 900 1012
<< pwell >>
rect 801 -66 887 586
<< nsubdiff >>
rect 834 2016 868 2040
rect 834 1946 868 1982
rect 834 1876 868 1912
rect 834 1806 868 1842
rect 834 1736 868 1772
rect 834 1666 868 1702
rect 834 1596 868 1632
rect 834 1526 868 1562
rect 834 1456 868 1492
rect 834 1386 868 1422
rect 834 1316 868 1352
rect 834 1246 868 1282
rect 834 1176 868 1212
rect 834 1106 868 1142
rect 834 1048 868 1072
<< mvpsubdiff >>
rect 827 536 861 560
rect 827 462 861 502
rect 827 388 861 428
rect 827 314 861 354
rect 827 240 861 280
rect 827 166 861 206
rect 827 92 861 132
rect 827 18 861 58
rect 827 -40 861 -16
<< nsubdiffcont >>
rect 834 1982 868 2016
rect 834 1912 868 1946
rect 834 1842 868 1876
rect 834 1772 868 1806
rect 834 1702 868 1736
rect 834 1632 868 1666
rect 834 1562 868 1596
rect 834 1492 868 1526
rect 834 1422 868 1456
rect 834 1352 868 1386
rect 834 1282 868 1316
rect 834 1212 868 1246
rect 834 1142 868 1176
rect 834 1072 868 1106
<< mvpsubdiffcont >>
rect 827 502 861 536
rect 827 428 861 462
rect 827 354 861 388
rect 827 280 861 314
rect 827 206 861 240
rect 827 132 861 166
rect 827 58 861 92
rect 827 -16 861 18
<< poly >>
rect 369 2122 503 2138
rect 369 2088 385 2122
rect 419 2088 453 2122
rect 487 2088 503 2122
rect 369 2072 503 2088
rect 375 2066 411 2072
rect 467 2066 503 2072
rect 375 1008 411 1014
rect 467 1008 503 1014
rect 664 1008 700 1014
rect 370 992 504 1008
rect 370 958 386 992
rect 420 958 454 992
rect 488 958 504 992
rect 370 942 504 958
rect 572 992 706 1008
rect 572 958 588 992
rect 622 958 656 992
rect 690 958 706 992
rect 572 942 706 958
rect 572 936 608 942
<< polycont >>
rect 385 2088 419 2122
rect 453 2088 487 2122
rect 386 958 420 992
rect 454 958 488 992
rect 588 958 622 992
rect 656 958 690 992
<< locali >>
rect 369 2088 385 2122
rect 419 2088 453 2122
rect 487 2088 503 2122
rect 326 1926 340 2044
rect 422 1982 456 2020
rect 715 1982 749 2020
rect 834 2016 868 2040
rect 272 1892 340 1926
rect 326 1415 340 1892
rect 255 1381 340 1415
rect 326 1094 340 1381
rect 834 1946 868 1982
rect 834 1876 868 1912
rect 834 1806 868 1842
rect 834 1736 868 1772
rect 834 1666 868 1702
rect 834 1596 868 1632
rect 834 1526 868 1562
rect 834 1456 868 1492
rect 834 1386 868 1422
rect 834 1316 868 1352
rect 834 1246 868 1282
rect 834 1176 868 1212
rect 834 1106 868 1142
rect 422 1060 456 1094
rect 711 1060 745 1094
rect 422 1026 745 1060
rect 834 1048 868 1072
rect 370 958 386 992
rect 420 958 454 992
rect 488 958 504 992
rect 572 958 588 992
rect 622 958 656 992
rect 690 958 706 992
rect 619 833 653 871
rect 527 750 561 788
rect 619 761 653 799
rect 711 750 745 788
rect 412 602 446 636
rect 827 536 861 560
rect 359 430 393 468
rect 359 358 393 396
rect 827 462 861 502
rect 827 388 861 428
rect 827 314 861 354
rect 827 240 861 280
rect 183 128 217 166
rect 183 56 217 94
rect 535 128 569 166
rect 535 56 569 94
rect 827 166 861 206
rect 827 92 861 132
rect 359 -12 393 22
rect 711 -12 745 22
rect 359 -46 745 -12
rect 827 18 861 58
rect 827 -40 861 -16
<< viali >>
rect 422 2020 456 2054
rect 422 1948 456 1982
rect 715 2020 749 2054
rect 715 1948 749 1982
rect 619 871 653 905
rect 527 788 561 822
rect 527 716 561 750
rect 619 799 653 833
rect 619 727 653 761
rect 711 788 745 822
rect 711 716 745 750
rect 359 468 393 502
rect 359 396 393 430
rect 359 324 393 358
rect 183 166 217 200
rect 183 94 217 128
rect 183 22 217 56
rect 535 166 569 200
rect 535 94 569 128
rect 535 22 569 56
<< metal1 >>
rect 509 2174 601 2202
rect 310 1536 370 2174
tri 535 2149 560 2174 ne
tri 548 2060 560 2072 se
rect 560 2060 601 2174
rect 407 2059 471 2060
rect 407 2007 413 2059
rect 465 2007 471 2059
tri 542 2054 548 2060 se
rect 548 2054 601 2060
tri 531 2043 542 2054 se
rect 542 2043 601 2054
rect 407 1995 471 2007
rect 407 1943 413 1995
rect 465 1943 471 1995
rect 407 1942 471 1943
rect 310 1500 334 1536
tri 334 1500 370 1536 nw
rect 546 1121 601 2043
rect 703 2059 767 2060
rect 703 2007 709 2059
rect 761 2007 767 2059
rect 703 1995 767 2007
rect 703 1943 709 1995
rect 761 1943 767 1995
rect 703 1942 767 1943
rect 635 1129 669 1164
tri 613 1031 629 1047 se
rect 629 1031 675 1101
rect 613 1027 675 1031
rect 613 905 659 1027
tri 659 1011 675 1027 nw
rect 613 871 619 905
rect 653 871 659 905
rect 521 822 567 834
rect 521 788 527 822
rect 561 788 567 822
rect 521 750 567 788
rect 521 716 527 750
rect 561 716 567 750
rect 521 687 567 716
rect 613 833 659 871
rect 613 799 619 833
rect 653 799 659 833
rect 613 761 659 799
rect 613 727 619 761
rect 653 727 659 761
rect 613 715 659 727
rect 705 822 751 834
rect 705 788 711 822
rect 745 788 751 822
rect 705 750 751 788
rect 705 716 711 750
rect 745 716 751 750
tri 567 687 592 712 sw
tri 680 687 705 712 se
rect 705 687 751 716
rect 521 641 751 687
tri 680 616 705 641 ne
rect 705 552 751 641
rect 816 562 868 568
tri 680 514 705 539 se
rect 353 502 705 514
rect 353 468 359 502
rect 393 468 705 502
rect 353 430 705 468
rect 353 396 359 430
rect 393 396 705 430
rect 353 358 705 396
rect 353 324 359 358
rect 393 324 705 358
rect 353 312 705 324
tri 680 287 705 312 ne
rect 816 498 868 510
rect 177 200 575 212
rect 177 166 183 200
rect 217 166 535 200
rect 569 166 575 200
rect 177 128 575 166
rect 177 94 183 128
rect 217 94 535 128
rect 569 94 575 128
rect 177 56 575 94
rect 177 22 183 56
rect 217 22 535 56
rect 569 22 575 56
rect 177 10 575 22
rect 816 -7 868 446
<< via1 >>
rect 413 2054 465 2059
rect 413 2020 422 2054
rect 422 2020 456 2054
rect 456 2020 465 2054
rect 413 2007 465 2020
rect 413 1982 465 1995
rect 413 1948 422 1982
rect 422 1948 456 1982
rect 456 1948 465 1982
rect 413 1943 465 1948
rect 709 2054 761 2059
rect 709 2020 715 2054
rect 715 2020 749 2054
rect 749 2020 761 2054
rect 709 2007 761 2020
rect 709 1982 761 1995
rect 709 1948 715 1982
rect 715 1948 749 1982
rect 749 1948 761 1982
rect 709 1943 761 1948
rect 816 510 868 562
rect 816 446 868 498
<< metal2 >>
rect 407 2007 413 2059
rect 465 2007 709 2059
rect 761 2007 767 2059
rect 407 1995 767 2007
rect 407 1943 413 1995
rect 465 1943 709 1995
rect 761 1943 767 1995
rect -27 562 868 568
rect -27 510 816 562
rect -27 498 868 510
rect -27 446 816 498
rect -27 440 868 446
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_0
timestamp 1704896540
transform 1 0 715 0 -1 2054
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_1
timestamp 1704896540
transform 1 0 422 0 -1 2054
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1704896540
transform 0 -1 745 -1 0 822
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1704896540
transform 0 -1 561 -1 0 822
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1704896540
transform 0 -1 653 -1 0 905
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_1
timestamp 1704896540
transform 0 1 183 1 0 22
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_2
timestamp 1704896540
transform 0 1 535 1 0 22
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_3
timestamp 1704896540
transform 0 1 359 1 0 324
box 0 0 1 1
use L1M1_CDNS_52468879185195  L1M1_CDNS_52468879185195_0
timestamp 1704896540
transform 0 1 711 -1 0 557
box -12 -6 550 40
use L1M1_CDNS_52468879185195  L1M1_CDNS_52468879185195_1
timestamp 1704896540
transform 0 1 827 1 0 5
box -12 -6 550 40
use L1M1_CDNS_52468879185381  L1M1_CDNS_52468879185381_0
timestamp 1704896540
transform 0 -1 547 -1 0 2031
box -12 -6 910 40
use L1M1_CDNS_52468879185381  L1M1_CDNS_52468879185381_1
timestamp 1704896540
transform 0 -1 364 -1 0 2031
box -12 -6 910 40
use L1M1_CDNS_52468879185381  L1M1_CDNS_52468879185381_2
timestamp 1704896540
transform 0 -1 669 1 0 1094
box -12 -6 910 40
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1704896540
transform 0 -1 868 1 0 440
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_0
timestamp 1704896540
transform -1 0 767 0 1 1943
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_1
timestamp 1704896540
transform -1 0 471 0 1 1943
box 0 0 1 1
use nfet_CDNS_524688791851204  nfet_CDNS_524688791851204_0
timestamp 1704896540
transform -1 0 700 0 -1 560
box -79 -26 551 626
use nfet_CDNS_524688791851205  nfet_CDNS_524688791851205_0
timestamp 1704896540
transform 1 0 572 0 1 720
box -79 -26 207 226
use pfet_CDNS_524688791851196  pfet_CDNS_524688791851196_0
timestamp 1704896540
transform -1 0 503 0 -1 2040
box -89 -36 217 1036
use pfet_CDNS_524688791851206  pfet_CDNS_524688791851206_0
timestamp 1704896540
transform -1 0 700 0 -1 2040
box -89 -36 125 1036
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_0
timestamp 1704896540
transform 0 -1 706 1 0 942
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_1
timestamp 1704896540
transform 0 -1 504 1 0 942
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_2
timestamp 1704896540
transform 0 -1 503 1 0 2072
box 0 0 1 1
use PYL1_CDNS_524688791851203  PYL1_CDNS_524688791851203_0
timestamp 1704896540
transform 0 -1 701 -1 0 652
box 0 0 66 474
<< labels >>
flabel metal1 s 430 79 494 119 0 FreeSans 200 180 0 0 vgnd
port 2 nsew
flabel metal1 s 635 1129 669 1164 0 FreeSans 600 0 0 0 out
port 1 nsew
flabel locali s 622 958 656 992 0 FreeSans 600 0 0 0 in
port 4 nsew
flabel locali s 420 959 454 992 0 FreeSans 600 0 0 0 ie_n
port 5 nsew
flabel locali s 412 602 446 636 0 FreeSans 600 180 0 0 ie
port 6 nsew
<< properties >>
string GDS_END 85774804
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85768466
string path 21.275 51.650 21.275 25.550 
<< end >>
