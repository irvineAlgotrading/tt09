magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -38 261 1786 582
<< pwell >>
rect 1 201 1433 203
rect 1 23 1744 201
rect 1 21 289 23
rect 747 21 937 23
rect 1348 21 1744 23
rect 30 -17 64 21
<< scnmos >>
rect 87 47 117 177
rect 171 47 201 177
rect 278 93 308 177
rect 501 49 531 177
rect 589 49 619 177
rect 831 47 861 177
rect 1017 49 1047 177
rect 1168 49 1198 133
rect 1327 49 1357 177
rect 1447 47 1477 167
rect 1547 47 1577 175
rect 1631 47 1661 175
<< scpmoshvt >>
rect 91 297 121 497
rect 175 297 205 497
rect 278 297 308 425
rect 488 325 518 493
rect 585 297 615 465
rect 797 297 827 497
rect 1017 297 1047 465
rect 1168 297 1198 425
rect 1343 329 1373 457
rect 1446 329 1476 497
rect 1547 297 1577 497
rect 1631 297 1661 497
<< ndiff >>
rect 27 129 87 177
rect 27 95 35 129
rect 69 95 87 129
rect 27 47 87 95
rect 117 129 171 177
rect 117 95 127 129
rect 161 95 171 129
rect 117 47 171 95
rect 201 93 278 177
rect 308 169 393 177
rect 308 135 347 169
rect 381 135 393 169
rect 308 93 393 135
rect 447 165 501 177
rect 447 131 457 165
rect 491 131 501 165
rect 201 89 263 93
rect 201 55 211 89
rect 245 55 263 89
rect 201 47 263 55
rect 447 49 501 131
rect 531 91 589 177
rect 531 57 543 91
rect 577 57 589 91
rect 531 49 589 57
rect 619 91 689 177
rect 619 57 643 91
rect 677 57 689 91
rect 619 49 689 57
rect 773 157 831 177
rect 773 123 787 157
rect 821 123 831 157
rect 773 89 831 123
rect 773 55 787 89
rect 821 55 831 89
rect 773 47 831 55
rect 861 165 913 177
rect 861 131 871 165
rect 905 131 913 165
rect 861 124 913 131
rect 861 47 911 124
rect 967 104 1017 177
rect 965 97 1017 104
rect 965 63 973 97
rect 1007 63 1017 97
rect 965 49 1017 63
rect 1047 133 1147 177
rect 1223 169 1327 177
rect 1223 135 1269 169
rect 1303 135 1327 169
rect 1223 133 1327 135
rect 1047 126 1168 133
rect 1047 92 1057 126
rect 1091 92 1168 126
rect 1047 49 1168 92
rect 1198 49 1327 133
rect 1357 167 1407 177
rect 1497 167 1547 175
rect 1357 93 1447 167
rect 1357 59 1369 93
rect 1403 59 1447 93
rect 1357 49 1447 59
rect 1374 47 1447 49
rect 1477 142 1547 167
rect 1477 108 1503 142
rect 1537 108 1547 142
rect 1477 47 1547 108
rect 1577 97 1631 175
rect 1577 63 1587 97
rect 1621 63 1631 97
rect 1577 47 1631 63
rect 1661 101 1718 175
rect 1661 67 1671 101
rect 1705 67 1718 101
rect 1661 47 1718 67
<< pdiff >>
rect 27 485 91 497
rect 27 451 35 485
rect 69 451 91 485
rect 27 417 91 451
rect 27 383 35 417
rect 69 383 91 417
rect 27 349 91 383
rect 27 315 35 349
rect 69 315 91 349
rect 27 297 91 315
rect 121 477 175 497
rect 121 443 131 477
rect 165 443 175 477
rect 121 409 175 443
rect 121 375 131 409
rect 165 375 175 409
rect 121 341 175 375
rect 121 307 131 341
rect 165 307 175 341
rect 121 297 175 307
rect 205 477 263 497
rect 205 443 216 477
rect 250 443 263 477
rect 205 425 263 443
rect 205 297 278 425
rect 308 341 364 425
rect 308 307 318 341
rect 352 307 364 341
rect 423 413 488 493
rect 423 379 444 413
rect 478 379 488 413
rect 423 325 488 379
rect 518 481 570 493
rect 518 447 528 481
rect 562 465 570 481
rect 745 481 797 497
rect 562 447 585 465
rect 518 325 585 447
rect 308 297 364 307
rect 535 297 585 325
rect 615 423 691 465
rect 745 447 753 481
rect 787 447 797 481
rect 745 435 797 447
rect 615 339 692 423
rect 615 305 646 339
rect 680 305 692 339
rect 615 297 692 305
rect 746 297 797 435
rect 827 343 879 497
rect 827 309 837 343
rect 871 309 879 343
rect 827 297 879 309
rect 933 405 1017 465
rect 933 371 941 405
rect 975 371 1017 405
rect 933 297 1017 371
rect 1047 425 1146 465
rect 1388 489 1446 497
rect 1388 457 1400 489
rect 1258 425 1343 457
rect 1047 409 1168 425
rect 1047 375 1097 409
rect 1131 375 1168 409
rect 1047 341 1168 375
rect 1047 307 1097 341
rect 1131 307 1168 341
rect 1047 297 1168 307
rect 1198 421 1343 425
rect 1198 387 1299 421
rect 1333 387 1343 421
rect 1198 329 1343 387
rect 1373 455 1400 457
rect 1434 455 1446 489
rect 1373 329 1446 455
rect 1476 341 1547 497
rect 1476 329 1503 341
rect 1198 297 1293 329
rect 1491 307 1503 329
rect 1537 307 1547 341
rect 1491 297 1547 307
rect 1577 489 1631 497
rect 1577 455 1587 489
rect 1621 455 1631 489
rect 1577 297 1631 455
rect 1661 477 1718 497
rect 1661 443 1672 477
rect 1706 443 1718 477
rect 1661 409 1718 443
rect 1661 375 1672 409
rect 1706 375 1718 409
rect 1661 297 1718 375
<< ndiffc >>
rect 35 95 69 129
rect 127 95 161 129
rect 347 135 381 169
rect 457 131 491 165
rect 211 55 245 89
rect 543 57 577 91
rect 643 57 677 91
rect 787 123 821 157
rect 787 55 821 89
rect 871 131 905 165
rect 973 63 1007 97
rect 1269 135 1303 169
rect 1057 92 1091 126
rect 1369 59 1403 93
rect 1503 108 1537 142
rect 1587 63 1621 97
rect 1671 67 1705 101
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 131 443 165 477
rect 131 375 165 409
rect 131 307 165 341
rect 216 443 250 477
rect 318 307 352 341
rect 444 379 478 413
rect 528 447 562 481
rect 753 447 787 481
rect 646 305 680 339
rect 837 309 871 343
rect 941 371 975 405
rect 1097 375 1131 409
rect 1097 307 1131 341
rect 1299 387 1333 421
rect 1400 455 1434 489
rect 1503 307 1537 341
rect 1587 455 1621 489
rect 1672 443 1706 477
rect 1672 375 1706 409
<< poly >>
rect 91 497 121 523
rect 175 497 205 523
rect 488 493 518 519
rect 278 425 308 483
rect 585 465 615 504
rect 797 497 827 523
rect 91 265 121 297
rect 175 265 205 297
rect 278 265 308 297
rect 488 271 518 325
rect 1017 493 1373 523
rect 1446 497 1476 523
rect 1547 497 1577 523
rect 1631 497 1661 523
rect 1017 465 1047 493
rect 1343 457 1373 493
rect 1168 425 1198 451
rect 488 265 531 271
rect 585 265 615 297
rect 87 249 236 265
rect 87 215 192 249
rect 226 215 236 249
rect 87 199 236 215
rect 278 249 531 265
rect 278 215 458 249
rect 492 215 531 249
rect 278 199 531 215
rect 573 249 627 265
rect 573 215 583 249
rect 617 215 627 249
rect 797 247 827 297
rect 1017 247 1047 297
rect 1168 265 1198 297
rect 1343 265 1373 329
rect 797 217 1047 247
rect 573 199 627 215
rect 87 177 117 199
rect 171 177 201 199
rect 278 177 308 199
rect 501 177 531 199
rect 589 177 619 199
rect 831 177 861 217
rect 1017 177 1047 217
rect 1089 249 1198 265
rect 1089 215 1099 249
rect 1133 215 1198 249
rect 1089 199 1198 215
rect 278 67 308 93
rect 87 21 117 47
rect 171 21 201 47
rect 501 21 531 49
rect 589 21 619 49
rect 1168 133 1198 199
rect 1327 249 1381 265
rect 1446 256 1476 329
rect 1547 265 1577 297
rect 1631 265 1661 297
rect 1446 255 1477 256
rect 1327 215 1337 249
rect 1371 215 1381 249
rect 1327 199 1381 215
rect 1423 239 1477 255
rect 1423 205 1433 239
rect 1467 205 1477 239
rect 1327 177 1357 199
rect 1423 189 1477 205
rect 1519 249 1577 265
rect 1519 215 1529 249
rect 1563 215 1577 249
rect 1519 199 1577 215
rect 1619 249 1673 265
rect 1619 215 1629 249
rect 1663 215 1673 249
rect 1619 199 1673 215
rect 1447 167 1477 189
rect 1547 175 1577 199
rect 1631 175 1661 199
rect 831 21 861 47
rect 1017 21 1047 49
rect 1168 23 1198 49
rect 1327 21 1357 49
rect 1447 21 1477 47
rect 1547 21 1577 47
rect 1631 21 1661 47
<< polycont >>
rect 192 215 226 249
rect 458 215 492 249
rect 583 215 617 249
rect 1099 215 1133 249
rect 1337 215 1371 249
rect 1433 205 1467 239
rect 1529 215 1563 249
rect 1629 215 1663 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 17 485 75 527
rect 17 451 35 485
rect 69 451 75 485
rect 17 417 75 451
rect 17 383 35 417
rect 69 383 75 417
rect 17 349 75 383
rect 17 315 35 349
rect 69 315 75 349
rect 17 298 75 315
rect 109 477 165 493
rect 109 443 131 477
rect 199 477 266 527
rect 737 481 803 527
rect 1571 489 1638 527
rect 199 443 216 477
rect 250 443 266 477
rect 302 447 528 481
rect 562 447 596 481
rect 737 447 753 481
rect 787 447 803 481
rect 870 455 1400 489
rect 1434 455 1489 489
rect 1571 455 1587 489
rect 1621 455 1638 489
rect 1672 477 1731 493
rect 109 409 165 443
rect 302 409 336 447
rect 870 413 904 455
rect 109 375 131 409
rect 109 341 165 375
rect 109 307 131 341
rect 109 288 165 307
rect 199 375 336 409
rect 404 379 444 413
rect 478 379 904 413
rect 941 405 975 421
rect 109 185 158 288
rect 199 265 233 375
rect 279 307 318 341
rect 352 307 596 341
rect 192 249 233 265
rect 226 215 233 249
rect 192 199 233 215
rect 17 129 75 147
rect 17 95 35 129
rect 69 95 75 129
rect 17 17 75 95
rect 109 129 161 185
rect 198 173 233 199
rect 198 139 313 173
rect 109 95 127 129
rect 109 70 161 95
rect 195 89 245 105
rect 195 55 211 89
rect 195 17 245 55
rect 279 85 313 139
rect 347 169 381 307
rect 562 265 596 307
rect 630 305 646 339
rect 680 323 707 339
rect 651 289 673 305
rect 651 275 707 289
rect 415 249 528 265
rect 415 215 458 249
rect 492 215 528 249
rect 562 249 617 265
rect 562 215 583 249
rect 562 199 617 215
rect 347 119 381 135
rect 441 165 517 181
rect 441 131 457 165
rect 491 159 517 165
rect 651 159 685 275
rect 741 241 775 379
rect 821 309 837 343
rect 871 309 905 343
rect 821 289 905 309
rect 491 131 685 159
rect 441 125 685 131
rect 719 207 775 241
rect 719 91 753 207
rect 857 187 905 289
rect 506 85 543 91
rect 279 57 543 85
rect 577 57 593 91
rect 627 57 643 91
rect 677 57 753 91
rect 787 157 821 173
rect 787 89 821 123
rect 279 51 593 57
rect 891 165 905 187
rect 857 131 871 153
rect 857 83 905 131
rect 941 119 975 371
rect 1009 178 1043 455
rect 1706 443 1731 477
rect 1672 421 1731 443
rect 1079 375 1097 409
rect 1131 375 1162 409
rect 1079 341 1162 375
rect 1079 307 1097 341
rect 1131 323 1162 341
rect 1269 387 1299 421
rect 1333 409 1731 421
rect 1333 387 1672 409
rect 1131 307 1133 323
rect 1079 289 1133 307
rect 1167 289 1235 323
rect 1082 249 1167 254
rect 1082 215 1099 249
rect 1133 215 1167 249
rect 1082 199 1167 215
rect 1125 187 1167 199
rect 1009 165 1051 178
rect 1009 144 1091 165
rect 1017 131 1091 144
rect 1057 126 1091 131
rect 1125 153 1133 187
rect 1125 126 1167 153
rect 941 85 949 119
rect 787 17 821 55
rect 941 63 973 85
rect 1007 63 1023 97
rect 1057 64 1091 92
rect 1201 85 1235 289
rect 1269 169 1303 387
rect 1634 375 1672 387
rect 1706 375 1731 409
rect 1337 289 1453 323
rect 1487 307 1503 341
rect 1537 307 1651 341
rect 1487 299 1651 307
rect 1337 249 1371 289
rect 1617 265 1651 299
rect 1337 199 1371 215
rect 1405 239 1467 255
rect 1405 205 1433 239
rect 1501 249 1583 265
rect 1501 215 1529 249
rect 1563 215 1583 249
rect 1617 249 1663 265
rect 1617 215 1629 249
rect 1405 189 1467 205
rect 1617 199 1663 215
rect 1405 187 1446 189
rect 1405 153 1409 187
rect 1443 153 1446 187
rect 1617 181 1651 199
rect 1405 146 1446 153
rect 1503 150 1651 181
rect 1495 147 1651 150
rect 1269 119 1303 135
rect 1495 142 1553 147
rect 1495 119 1503 142
rect 1337 85 1369 93
rect 941 53 1023 63
rect 1201 59 1369 85
rect 1403 59 1430 93
rect 1495 85 1501 119
rect 1537 108 1553 142
rect 1697 117 1731 375
rect 1535 85 1553 108
rect 1495 59 1553 85
rect 1587 97 1621 113
rect 1201 51 1430 59
rect 1587 17 1621 63
rect 1671 101 1731 117
rect 1705 67 1731 101
rect 1671 51 1731 67
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 673 305 680 323
rect 680 305 707 323
rect 673 289 707 305
rect 857 165 891 187
rect 857 153 871 165
rect 871 153 891 165
rect 1133 289 1167 323
rect 1133 153 1167 187
rect 949 97 983 119
rect 949 85 973 97
rect 973 85 983 97
rect 1409 153 1443 187
rect 1501 108 1503 119
rect 1503 108 1535 119
rect 1501 85 1535 108
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
<< metal1 >>
rect 0 561 1748 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1748 561
rect 0 496 1748 527
rect 661 323 719 329
rect 661 289 673 323
rect 707 320 719 323
rect 1121 323 1179 329
rect 1121 320 1133 323
rect 707 292 1133 320
rect 707 289 719 292
rect 661 283 719 289
rect 1121 289 1133 292
rect 1167 289 1179 323
rect 1121 283 1179 289
rect 845 187 903 193
rect 845 153 857 187
rect 891 184 903 187
rect 1121 187 1179 193
rect 1121 184 1133 187
rect 891 156 1133 184
rect 891 153 903 156
rect 845 147 903 153
rect 1121 153 1133 156
rect 1167 184 1179 187
rect 1397 187 1455 193
rect 1397 184 1409 187
rect 1167 156 1409 184
rect 1167 153 1179 156
rect 1121 147 1179 153
rect 1397 153 1409 156
rect 1443 153 1455 187
rect 1397 147 1455 153
rect 937 119 995 125
rect 937 85 949 119
rect 983 116 995 119
rect 1489 119 1547 125
rect 1489 116 1501 119
rect 983 88 1501 116
rect 983 85 995 88
rect 937 79 995 85
rect 1489 85 1501 88
rect 1535 85 1547 119
rect 1489 79 1547 85
rect 0 17 1748 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1748 17
rect 0 -48 1748 -17
<< labels >>
flabel locali s 121 357 155 391 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 1409 289 1443 323 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 489 221 523 255 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 1501 221 1535 255 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 hkscl5hdv1_xnor3_1
flabel comment s 0 544 0 544 3 FreeSans 200 0 0 0 HHNEC
rlabel metal1 s 0 -48 1748 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1748 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1748 544
string GDS_END 592498
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 580320
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 8.740 0.000 
<< end >>
