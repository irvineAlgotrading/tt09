magic
tech sky130A
timestamp 1704896540
<< metal1 >>
rect 0 0 3 26
rect 29 0 35 26
rect 61 0 67 26
rect 93 0 99 26
rect 125 0 131 26
rect 157 0 163 26
rect 189 0 195 26
rect 221 0 227 26
rect 253 0 259 26
rect 285 0 291 26
rect 317 0 323 26
rect 349 0 355 26
rect 381 0 387 26
rect 413 0 419 26
rect 445 0 451 26
rect 477 0 483 26
rect 509 0 515 26
rect 541 0 547 26
rect 573 0 579 26
rect 605 0 611 26
rect 637 0 643 26
rect 669 0 675 26
rect 701 0 707 26
rect 733 0 739 26
rect 765 0 771 26
rect 797 0 803 26
rect 829 0 835 26
rect 861 0 867 26
rect 893 0 899 26
rect 925 0 931 26
rect 957 0 963 26
rect 989 0 995 26
rect 1021 0 1027 26
rect 1053 0 1059 26
rect 1085 0 1091 26
rect 1117 0 1123 26
rect 1149 0 1155 26
rect 1181 0 1187 26
rect 1213 0 1219 26
rect 1245 0 1251 26
rect 1277 0 1283 26
rect 1309 0 1315 26
rect 1341 0 1347 26
rect 1373 0 1379 26
rect 1405 0 1411 26
rect 1437 0 1443 26
rect 1469 0 1475 26
rect 1501 0 1507 26
rect 1533 0 1539 26
rect 1565 0 1571 26
rect 1597 0 1603 26
rect 1629 0 1635 26
rect 1661 0 1667 26
rect 1693 0 1699 26
rect 1725 0 1731 26
rect 1757 0 1763 26
rect 1789 0 1795 26
rect 1821 0 1827 26
rect 1853 0 1859 26
rect 1885 0 1891 26
rect 1917 0 1923 26
rect 1949 0 1955 26
rect 1981 0 1987 26
rect 2013 0 2019 26
rect 2045 0 2051 26
rect 2077 0 2083 26
rect 2109 0 2115 26
rect 2141 0 2147 26
rect 2173 0 2179 26
rect 2205 0 2211 26
rect 2237 0 2243 26
rect 2269 0 2275 26
rect 2301 0 2307 26
rect 2333 0 2339 26
rect 2365 0 2371 26
rect 2397 0 2403 26
rect 2429 0 2435 26
rect 2461 0 2467 26
rect 2493 0 2499 26
rect 2525 0 2531 26
rect 2557 0 2563 26
rect 2589 0 2595 26
rect 2621 0 2627 26
rect 2653 0 2659 26
rect 2685 0 2691 26
rect 2717 0 2723 26
rect 2749 0 2755 26
rect 2781 0 2787 26
rect 2813 0 2819 26
rect 2845 0 2851 26
rect 2877 0 2883 26
rect 2909 0 2915 26
rect 2941 0 2947 26
rect 2973 0 2979 26
rect 3005 0 3011 26
rect 3037 0 3043 26
rect 3069 0 3075 26
rect 3101 0 3107 26
rect 3133 0 3139 26
rect 3165 0 3171 26
rect 3197 0 3203 26
rect 3229 0 3235 26
rect 3261 0 3267 26
rect 3293 0 3299 26
rect 3325 0 3331 26
rect 3357 0 3363 26
rect 3389 0 3395 26
rect 3421 0 3427 26
rect 3453 0 3459 26
rect 3485 0 3491 26
rect 3517 0 3523 26
rect 3549 0 3555 26
rect 3581 0 3587 26
rect 3613 0 3619 26
rect 3645 0 3651 26
rect 3677 0 3683 26
rect 3709 0 3715 26
rect 3741 0 3747 26
rect 3773 0 3779 26
rect 3805 0 3811 26
rect 3837 0 3843 26
rect 3869 0 3875 26
rect 3901 0 3907 26
rect 3933 0 3939 26
rect 3965 0 3971 26
rect 3997 0 4003 26
rect 4029 0 4035 26
rect 4061 0 4067 26
rect 4093 0 4099 26
rect 4125 0 4131 26
rect 4157 0 4163 26
rect 4189 0 4195 26
rect 4221 0 4227 26
rect 4253 0 4259 26
rect 4285 0 4291 26
rect 4317 0 4323 26
rect 4349 0 4355 26
rect 4381 0 4387 26
rect 4413 0 4419 26
rect 4445 0 4451 26
rect 4477 0 4483 26
rect 4509 0 4515 26
rect 4541 0 4547 26
rect 4573 0 4579 26
rect 4605 0 4611 26
rect 4637 0 4643 26
rect 4669 0 4675 26
rect 4701 0 4707 26
rect 4733 0 4739 26
rect 4765 0 4771 26
rect 4797 0 4803 26
rect 4829 0 4835 26
rect 4861 0 4867 26
rect 4893 0 4899 26
rect 4925 0 4931 26
rect 4957 0 4963 26
rect 4989 0 4995 26
rect 5021 0 5027 26
rect 5053 0 5059 26
rect 5085 0 5091 26
rect 5117 0 5123 26
rect 5149 0 5155 26
rect 5181 0 5187 26
rect 5213 0 5219 26
rect 5245 0 5251 26
rect 5277 0 5283 26
rect 5309 0 5315 26
rect 5341 0 5347 26
rect 5373 0 5379 26
rect 5405 0 5411 26
rect 5437 0 5443 26
rect 5469 0 5475 26
rect 5501 0 5507 26
rect 5533 0 5539 26
rect 5565 0 5571 26
rect 5597 0 5603 26
rect 5629 0 5635 26
rect 5661 0 5667 26
rect 5693 0 5699 26
rect 5725 0 5731 26
rect 5757 0 5763 26
rect 5789 0 5795 26
rect 5821 0 5827 26
rect 5853 0 5859 26
rect 5885 0 5891 26
rect 5917 0 5923 26
rect 5949 0 5955 26
rect 5981 0 5987 26
rect 6013 0 6019 26
rect 6045 0 6051 26
rect 6077 0 6083 26
rect 6109 0 6115 26
rect 6141 0 6147 26
rect 6173 0 6179 26
rect 6205 0 6211 26
rect 6237 0 6243 26
rect 6269 0 6275 26
rect 6301 0 6307 26
rect 6333 0 6339 26
rect 6365 0 6371 26
rect 6397 0 6403 26
rect 6429 0 6435 26
rect 6461 0 6467 26
rect 6493 0 6499 26
rect 6525 0 6531 26
rect 6557 0 6563 26
rect 6589 0 6595 26
rect 6621 0 6627 26
rect 6653 0 6659 26
rect 6685 0 6691 26
rect 6717 0 6723 26
rect 6749 0 6755 26
rect 6781 0 6787 26
rect 6813 0 6819 26
rect 6845 0 6851 26
rect 6877 0 6883 26
rect 6909 0 6915 26
rect 6941 0 6947 26
rect 6973 0 6979 26
rect 7005 0 7011 26
rect 7037 0 7043 26
rect 7069 0 7075 26
rect 7101 0 7107 26
rect 7133 0 7139 26
rect 7165 0 7171 26
rect 7197 0 7203 26
rect 7229 0 7235 26
rect 7261 0 7267 26
rect 7293 0 7299 26
rect 7325 0 7331 26
rect 7357 0 7363 26
rect 7389 0 7395 26
rect 7421 0 7427 26
rect 7453 0 7459 26
rect 7485 0 7491 26
rect 7517 0 7523 26
rect 7549 0 7555 26
rect 7581 0 7587 26
rect 7613 0 7619 26
rect 7645 0 7651 26
rect 7677 0 7683 26
rect 7709 0 7715 26
rect 7741 0 7747 26
rect 7773 0 7779 26
rect 7805 0 7811 26
rect 7837 0 7843 26
rect 7869 0 7875 26
rect 7901 0 7907 26
rect 7933 0 7939 26
rect 7965 0 7971 26
rect 7997 0 8003 26
rect 8029 0 8035 26
rect 8061 0 8067 26
rect 8093 0 8099 26
rect 8125 0 8131 26
rect 8157 0 8163 26
rect 8189 0 8195 26
rect 8221 0 8227 26
rect 8253 0 8259 26
rect 8285 0 8291 26
rect 8317 0 8323 26
rect 8349 0 8355 26
rect 8381 0 8387 26
rect 8413 0 8419 26
rect 8445 0 8451 26
rect 8477 0 8483 26
rect 8509 0 8515 26
rect 8541 0 8547 26
rect 8573 0 8579 26
rect 8605 0 8611 26
rect 8637 0 8643 26
rect 8669 0 8675 26
rect 8701 0 8707 26
rect 8733 0 8739 26
rect 8765 0 8771 26
rect 8797 0 8803 26
rect 8829 0 8835 26
rect 8861 0 8867 26
rect 8893 0 8899 26
rect 8925 0 8931 26
rect 8957 0 8963 26
rect 8989 0 8995 26
rect 9021 0 9027 26
rect 9053 0 9059 26
rect 9085 0 9091 26
rect 9117 0 9123 26
rect 9149 0 9155 26
rect 9181 0 9187 26
rect 9213 0 9219 26
rect 9245 0 9251 26
rect 9277 0 9283 26
rect 9309 0 9315 26
rect 9341 0 9347 26
rect 9373 0 9379 26
rect 9405 0 9411 26
rect 9437 0 9443 26
rect 9469 0 9475 26
rect 9501 0 9507 26
rect 9533 0 9539 26
rect 9565 0 9571 26
rect 9597 0 9603 26
rect 9629 0 9635 26
rect 9661 0 9667 26
rect 9693 0 9699 26
rect 9725 0 9731 26
rect 9757 0 9763 26
rect 9789 0 9795 26
rect 9821 0 9827 26
rect 9853 0 9859 26
rect 9885 0 9891 26
rect 9917 0 9923 26
rect 9949 0 9955 26
rect 9981 0 9987 26
rect 10013 0 10019 26
rect 10045 0 10051 26
rect 10077 0 10083 26
rect 10109 0 10115 26
rect 10141 0 10147 26
rect 10173 0 10179 26
rect 10205 0 10211 26
rect 10237 0 10243 26
rect 10269 0 10275 26
rect 10301 0 10304 26
<< via1 >>
rect 3 0 29 26
rect 35 0 61 26
rect 67 0 93 26
rect 99 0 125 26
rect 131 0 157 26
rect 163 0 189 26
rect 195 0 221 26
rect 227 0 253 26
rect 259 0 285 26
rect 291 0 317 26
rect 323 0 349 26
rect 355 0 381 26
rect 387 0 413 26
rect 419 0 445 26
rect 451 0 477 26
rect 483 0 509 26
rect 515 0 541 26
rect 547 0 573 26
rect 579 0 605 26
rect 611 0 637 26
rect 643 0 669 26
rect 675 0 701 26
rect 707 0 733 26
rect 739 0 765 26
rect 771 0 797 26
rect 803 0 829 26
rect 835 0 861 26
rect 867 0 893 26
rect 899 0 925 26
rect 931 0 957 26
rect 963 0 989 26
rect 995 0 1021 26
rect 1027 0 1053 26
rect 1059 0 1085 26
rect 1091 0 1117 26
rect 1123 0 1149 26
rect 1155 0 1181 26
rect 1187 0 1213 26
rect 1219 0 1245 26
rect 1251 0 1277 26
rect 1283 0 1309 26
rect 1315 0 1341 26
rect 1347 0 1373 26
rect 1379 0 1405 26
rect 1411 0 1437 26
rect 1443 0 1469 26
rect 1475 0 1501 26
rect 1507 0 1533 26
rect 1539 0 1565 26
rect 1571 0 1597 26
rect 1603 0 1629 26
rect 1635 0 1661 26
rect 1667 0 1693 26
rect 1699 0 1725 26
rect 1731 0 1757 26
rect 1763 0 1789 26
rect 1795 0 1821 26
rect 1827 0 1853 26
rect 1859 0 1885 26
rect 1891 0 1917 26
rect 1923 0 1949 26
rect 1955 0 1981 26
rect 1987 0 2013 26
rect 2019 0 2045 26
rect 2051 0 2077 26
rect 2083 0 2109 26
rect 2115 0 2141 26
rect 2147 0 2173 26
rect 2179 0 2205 26
rect 2211 0 2237 26
rect 2243 0 2269 26
rect 2275 0 2301 26
rect 2307 0 2333 26
rect 2339 0 2365 26
rect 2371 0 2397 26
rect 2403 0 2429 26
rect 2435 0 2461 26
rect 2467 0 2493 26
rect 2499 0 2525 26
rect 2531 0 2557 26
rect 2563 0 2589 26
rect 2595 0 2621 26
rect 2627 0 2653 26
rect 2659 0 2685 26
rect 2691 0 2717 26
rect 2723 0 2749 26
rect 2755 0 2781 26
rect 2787 0 2813 26
rect 2819 0 2845 26
rect 2851 0 2877 26
rect 2883 0 2909 26
rect 2915 0 2941 26
rect 2947 0 2973 26
rect 2979 0 3005 26
rect 3011 0 3037 26
rect 3043 0 3069 26
rect 3075 0 3101 26
rect 3107 0 3133 26
rect 3139 0 3165 26
rect 3171 0 3197 26
rect 3203 0 3229 26
rect 3235 0 3261 26
rect 3267 0 3293 26
rect 3299 0 3325 26
rect 3331 0 3357 26
rect 3363 0 3389 26
rect 3395 0 3421 26
rect 3427 0 3453 26
rect 3459 0 3485 26
rect 3491 0 3517 26
rect 3523 0 3549 26
rect 3555 0 3581 26
rect 3587 0 3613 26
rect 3619 0 3645 26
rect 3651 0 3677 26
rect 3683 0 3709 26
rect 3715 0 3741 26
rect 3747 0 3773 26
rect 3779 0 3805 26
rect 3811 0 3837 26
rect 3843 0 3869 26
rect 3875 0 3901 26
rect 3907 0 3933 26
rect 3939 0 3965 26
rect 3971 0 3997 26
rect 4003 0 4029 26
rect 4035 0 4061 26
rect 4067 0 4093 26
rect 4099 0 4125 26
rect 4131 0 4157 26
rect 4163 0 4189 26
rect 4195 0 4221 26
rect 4227 0 4253 26
rect 4259 0 4285 26
rect 4291 0 4317 26
rect 4323 0 4349 26
rect 4355 0 4381 26
rect 4387 0 4413 26
rect 4419 0 4445 26
rect 4451 0 4477 26
rect 4483 0 4509 26
rect 4515 0 4541 26
rect 4547 0 4573 26
rect 4579 0 4605 26
rect 4611 0 4637 26
rect 4643 0 4669 26
rect 4675 0 4701 26
rect 4707 0 4733 26
rect 4739 0 4765 26
rect 4771 0 4797 26
rect 4803 0 4829 26
rect 4835 0 4861 26
rect 4867 0 4893 26
rect 4899 0 4925 26
rect 4931 0 4957 26
rect 4963 0 4989 26
rect 4995 0 5021 26
rect 5027 0 5053 26
rect 5059 0 5085 26
rect 5091 0 5117 26
rect 5123 0 5149 26
rect 5155 0 5181 26
rect 5187 0 5213 26
rect 5219 0 5245 26
rect 5251 0 5277 26
rect 5283 0 5309 26
rect 5315 0 5341 26
rect 5347 0 5373 26
rect 5379 0 5405 26
rect 5411 0 5437 26
rect 5443 0 5469 26
rect 5475 0 5501 26
rect 5507 0 5533 26
rect 5539 0 5565 26
rect 5571 0 5597 26
rect 5603 0 5629 26
rect 5635 0 5661 26
rect 5667 0 5693 26
rect 5699 0 5725 26
rect 5731 0 5757 26
rect 5763 0 5789 26
rect 5795 0 5821 26
rect 5827 0 5853 26
rect 5859 0 5885 26
rect 5891 0 5917 26
rect 5923 0 5949 26
rect 5955 0 5981 26
rect 5987 0 6013 26
rect 6019 0 6045 26
rect 6051 0 6077 26
rect 6083 0 6109 26
rect 6115 0 6141 26
rect 6147 0 6173 26
rect 6179 0 6205 26
rect 6211 0 6237 26
rect 6243 0 6269 26
rect 6275 0 6301 26
rect 6307 0 6333 26
rect 6339 0 6365 26
rect 6371 0 6397 26
rect 6403 0 6429 26
rect 6435 0 6461 26
rect 6467 0 6493 26
rect 6499 0 6525 26
rect 6531 0 6557 26
rect 6563 0 6589 26
rect 6595 0 6621 26
rect 6627 0 6653 26
rect 6659 0 6685 26
rect 6691 0 6717 26
rect 6723 0 6749 26
rect 6755 0 6781 26
rect 6787 0 6813 26
rect 6819 0 6845 26
rect 6851 0 6877 26
rect 6883 0 6909 26
rect 6915 0 6941 26
rect 6947 0 6973 26
rect 6979 0 7005 26
rect 7011 0 7037 26
rect 7043 0 7069 26
rect 7075 0 7101 26
rect 7107 0 7133 26
rect 7139 0 7165 26
rect 7171 0 7197 26
rect 7203 0 7229 26
rect 7235 0 7261 26
rect 7267 0 7293 26
rect 7299 0 7325 26
rect 7331 0 7357 26
rect 7363 0 7389 26
rect 7395 0 7421 26
rect 7427 0 7453 26
rect 7459 0 7485 26
rect 7491 0 7517 26
rect 7523 0 7549 26
rect 7555 0 7581 26
rect 7587 0 7613 26
rect 7619 0 7645 26
rect 7651 0 7677 26
rect 7683 0 7709 26
rect 7715 0 7741 26
rect 7747 0 7773 26
rect 7779 0 7805 26
rect 7811 0 7837 26
rect 7843 0 7869 26
rect 7875 0 7901 26
rect 7907 0 7933 26
rect 7939 0 7965 26
rect 7971 0 7997 26
rect 8003 0 8029 26
rect 8035 0 8061 26
rect 8067 0 8093 26
rect 8099 0 8125 26
rect 8131 0 8157 26
rect 8163 0 8189 26
rect 8195 0 8221 26
rect 8227 0 8253 26
rect 8259 0 8285 26
rect 8291 0 8317 26
rect 8323 0 8349 26
rect 8355 0 8381 26
rect 8387 0 8413 26
rect 8419 0 8445 26
rect 8451 0 8477 26
rect 8483 0 8509 26
rect 8515 0 8541 26
rect 8547 0 8573 26
rect 8579 0 8605 26
rect 8611 0 8637 26
rect 8643 0 8669 26
rect 8675 0 8701 26
rect 8707 0 8733 26
rect 8739 0 8765 26
rect 8771 0 8797 26
rect 8803 0 8829 26
rect 8835 0 8861 26
rect 8867 0 8893 26
rect 8899 0 8925 26
rect 8931 0 8957 26
rect 8963 0 8989 26
rect 8995 0 9021 26
rect 9027 0 9053 26
rect 9059 0 9085 26
rect 9091 0 9117 26
rect 9123 0 9149 26
rect 9155 0 9181 26
rect 9187 0 9213 26
rect 9219 0 9245 26
rect 9251 0 9277 26
rect 9283 0 9309 26
rect 9315 0 9341 26
rect 9347 0 9373 26
rect 9379 0 9405 26
rect 9411 0 9437 26
rect 9443 0 9469 26
rect 9475 0 9501 26
rect 9507 0 9533 26
rect 9539 0 9565 26
rect 9571 0 9597 26
rect 9603 0 9629 26
rect 9635 0 9661 26
rect 9667 0 9693 26
rect 9699 0 9725 26
rect 9731 0 9757 26
rect 9763 0 9789 26
rect 9795 0 9821 26
rect 9827 0 9853 26
rect 9859 0 9885 26
rect 9891 0 9917 26
rect 9923 0 9949 26
rect 9955 0 9981 26
rect 9987 0 10013 26
rect 10019 0 10045 26
rect 10051 0 10077 26
rect 10083 0 10109 26
rect 10115 0 10141 26
rect 10147 0 10173 26
rect 10179 0 10205 26
rect 10211 0 10237 26
rect 10243 0 10269 26
rect 10275 0 10301 26
<< metal2 >>
rect 0 0 3 26
rect 29 0 35 26
rect 61 0 67 26
rect 93 0 99 26
rect 125 0 131 26
rect 157 0 163 26
rect 189 0 195 26
rect 221 0 227 26
rect 253 0 259 26
rect 285 0 291 26
rect 317 0 323 26
rect 349 0 355 26
rect 381 0 387 26
rect 413 0 419 26
rect 445 0 451 26
rect 477 0 483 26
rect 509 0 515 26
rect 541 0 547 26
rect 573 0 579 26
rect 605 0 611 26
rect 637 0 643 26
rect 669 0 675 26
rect 701 0 707 26
rect 733 0 739 26
rect 765 0 771 26
rect 797 0 803 26
rect 829 0 835 26
rect 861 0 867 26
rect 893 0 899 26
rect 925 0 931 26
rect 957 0 963 26
rect 989 0 995 26
rect 1021 0 1027 26
rect 1053 0 1059 26
rect 1085 0 1091 26
rect 1117 0 1123 26
rect 1149 0 1155 26
rect 1181 0 1187 26
rect 1213 0 1219 26
rect 1245 0 1251 26
rect 1277 0 1283 26
rect 1309 0 1315 26
rect 1341 0 1347 26
rect 1373 0 1379 26
rect 1405 0 1411 26
rect 1437 0 1443 26
rect 1469 0 1475 26
rect 1501 0 1507 26
rect 1533 0 1539 26
rect 1565 0 1571 26
rect 1597 0 1603 26
rect 1629 0 1635 26
rect 1661 0 1667 26
rect 1693 0 1699 26
rect 1725 0 1731 26
rect 1757 0 1763 26
rect 1789 0 1795 26
rect 1821 0 1827 26
rect 1853 0 1859 26
rect 1885 0 1891 26
rect 1917 0 1923 26
rect 1949 0 1955 26
rect 1981 0 1987 26
rect 2013 0 2019 26
rect 2045 0 2051 26
rect 2077 0 2083 26
rect 2109 0 2115 26
rect 2141 0 2147 26
rect 2173 0 2179 26
rect 2205 0 2211 26
rect 2237 0 2243 26
rect 2269 0 2275 26
rect 2301 0 2307 26
rect 2333 0 2339 26
rect 2365 0 2371 26
rect 2397 0 2403 26
rect 2429 0 2435 26
rect 2461 0 2467 26
rect 2493 0 2499 26
rect 2525 0 2531 26
rect 2557 0 2563 26
rect 2589 0 2595 26
rect 2621 0 2627 26
rect 2653 0 2659 26
rect 2685 0 2691 26
rect 2717 0 2723 26
rect 2749 0 2755 26
rect 2781 0 2787 26
rect 2813 0 2819 26
rect 2845 0 2851 26
rect 2877 0 2883 26
rect 2909 0 2915 26
rect 2941 0 2947 26
rect 2973 0 2979 26
rect 3005 0 3011 26
rect 3037 0 3043 26
rect 3069 0 3075 26
rect 3101 0 3107 26
rect 3133 0 3139 26
rect 3165 0 3171 26
rect 3197 0 3203 26
rect 3229 0 3235 26
rect 3261 0 3267 26
rect 3293 0 3299 26
rect 3325 0 3331 26
rect 3357 0 3363 26
rect 3389 0 3395 26
rect 3421 0 3427 26
rect 3453 0 3459 26
rect 3485 0 3491 26
rect 3517 0 3523 26
rect 3549 0 3555 26
rect 3581 0 3587 26
rect 3613 0 3619 26
rect 3645 0 3651 26
rect 3677 0 3683 26
rect 3709 0 3715 26
rect 3741 0 3747 26
rect 3773 0 3779 26
rect 3805 0 3811 26
rect 3837 0 3843 26
rect 3869 0 3875 26
rect 3901 0 3907 26
rect 3933 0 3939 26
rect 3965 0 3971 26
rect 3997 0 4003 26
rect 4029 0 4035 26
rect 4061 0 4067 26
rect 4093 0 4099 26
rect 4125 0 4131 26
rect 4157 0 4163 26
rect 4189 0 4195 26
rect 4221 0 4227 26
rect 4253 0 4259 26
rect 4285 0 4291 26
rect 4317 0 4323 26
rect 4349 0 4355 26
rect 4381 0 4387 26
rect 4413 0 4419 26
rect 4445 0 4451 26
rect 4477 0 4483 26
rect 4509 0 4515 26
rect 4541 0 4547 26
rect 4573 0 4579 26
rect 4605 0 4611 26
rect 4637 0 4643 26
rect 4669 0 4675 26
rect 4701 0 4707 26
rect 4733 0 4739 26
rect 4765 0 4771 26
rect 4797 0 4803 26
rect 4829 0 4835 26
rect 4861 0 4867 26
rect 4893 0 4899 26
rect 4925 0 4931 26
rect 4957 0 4963 26
rect 4989 0 4995 26
rect 5021 0 5027 26
rect 5053 0 5059 26
rect 5085 0 5091 26
rect 5117 0 5123 26
rect 5149 0 5155 26
rect 5181 0 5187 26
rect 5213 0 5219 26
rect 5245 0 5251 26
rect 5277 0 5283 26
rect 5309 0 5315 26
rect 5341 0 5347 26
rect 5373 0 5379 26
rect 5405 0 5411 26
rect 5437 0 5443 26
rect 5469 0 5475 26
rect 5501 0 5507 26
rect 5533 0 5539 26
rect 5565 0 5571 26
rect 5597 0 5603 26
rect 5629 0 5635 26
rect 5661 0 5667 26
rect 5693 0 5699 26
rect 5725 0 5731 26
rect 5757 0 5763 26
rect 5789 0 5795 26
rect 5821 0 5827 26
rect 5853 0 5859 26
rect 5885 0 5891 26
rect 5917 0 5923 26
rect 5949 0 5955 26
rect 5981 0 5987 26
rect 6013 0 6019 26
rect 6045 0 6051 26
rect 6077 0 6083 26
rect 6109 0 6115 26
rect 6141 0 6147 26
rect 6173 0 6179 26
rect 6205 0 6211 26
rect 6237 0 6243 26
rect 6269 0 6275 26
rect 6301 0 6307 26
rect 6333 0 6339 26
rect 6365 0 6371 26
rect 6397 0 6403 26
rect 6429 0 6435 26
rect 6461 0 6467 26
rect 6493 0 6499 26
rect 6525 0 6531 26
rect 6557 0 6563 26
rect 6589 0 6595 26
rect 6621 0 6627 26
rect 6653 0 6659 26
rect 6685 0 6691 26
rect 6717 0 6723 26
rect 6749 0 6755 26
rect 6781 0 6787 26
rect 6813 0 6819 26
rect 6845 0 6851 26
rect 6877 0 6883 26
rect 6909 0 6915 26
rect 6941 0 6947 26
rect 6973 0 6979 26
rect 7005 0 7011 26
rect 7037 0 7043 26
rect 7069 0 7075 26
rect 7101 0 7107 26
rect 7133 0 7139 26
rect 7165 0 7171 26
rect 7197 0 7203 26
rect 7229 0 7235 26
rect 7261 0 7267 26
rect 7293 0 7299 26
rect 7325 0 7331 26
rect 7357 0 7363 26
rect 7389 0 7395 26
rect 7421 0 7427 26
rect 7453 0 7459 26
rect 7485 0 7491 26
rect 7517 0 7523 26
rect 7549 0 7555 26
rect 7581 0 7587 26
rect 7613 0 7619 26
rect 7645 0 7651 26
rect 7677 0 7683 26
rect 7709 0 7715 26
rect 7741 0 7747 26
rect 7773 0 7779 26
rect 7805 0 7811 26
rect 7837 0 7843 26
rect 7869 0 7875 26
rect 7901 0 7907 26
rect 7933 0 7939 26
rect 7965 0 7971 26
rect 7997 0 8003 26
rect 8029 0 8035 26
rect 8061 0 8067 26
rect 8093 0 8099 26
rect 8125 0 8131 26
rect 8157 0 8163 26
rect 8189 0 8195 26
rect 8221 0 8227 26
rect 8253 0 8259 26
rect 8285 0 8291 26
rect 8317 0 8323 26
rect 8349 0 8355 26
rect 8381 0 8387 26
rect 8413 0 8419 26
rect 8445 0 8451 26
rect 8477 0 8483 26
rect 8509 0 8515 26
rect 8541 0 8547 26
rect 8573 0 8579 26
rect 8605 0 8611 26
rect 8637 0 8643 26
rect 8669 0 8675 26
rect 8701 0 8707 26
rect 8733 0 8739 26
rect 8765 0 8771 26
rect 8797 0 8803 26
rect 8829 0 8835 26
rect 8861 0 8867 26
rect 8893 0 8899 26
rect 8925 0 8931 26
rect 8957 0 8963 26
rect 8989 0 8995 26
rect 9021 0 9027 26
rect 9053 0 9059 26
rect 9085 0 9091 26
rect 9117 0 9123 26
rect 9149 0 9155 26
rect 9181 0 9187 26
rect 9213 0 9219 26
rect 9245 0 9251 26
rect 9277 0 9283 26
rect 9309 0 9315 26
rect 9341 0 9347 26
rect 9373 0 9379 26
rect 9405 0 9411 26
rect 9437 0 9443 26
rect 9469 0 9475 26
rect 9501 0 9507 26
rect 9533 0 9539 26
rect 9565 0 9571 26
rect 9597 0 9603 26
rect 9629 0 9635 26
rect 9661 0 9667 26
rect 9693 0 9699 26
rect 9725 0 9731 26
rect 9757 0 9763 26
rect 9789 0 9795 26
rect 9821 0 9827 26
rect 9853 0 9859 26
rect 9885 0 9891 26
rect 9917 0 9923 26
rect 9949 0 9955 26
rect 9981 0 9987 26
rect 10013 0 10019 26
rect 10045 0 10051 26
rect 10077 0 10083 26
rect 10109 0 10115 26
rect 10141 0 10147 26
rect 10173 0 10179 26
rect 10205 0 10211 26
rect 10237 0 10243 26
rect 10269 0 10275 26
rect 10301 0 10304 26
<< properties >>
string GDS_END 78509354
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 78488614
<< end >>
