magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< dnwell >>
rect 1279 8376 8627 11090
rect 1279 7302 4481 8376
rect 1279 439 4110 7302
<< nwell >>
rect 1199 10980 8707 11170
rect -59 10810 8707 10980
rect -59 379 111 10810
rect 1199 7389 1559 10810
rect 8347 8296 8707 10810
rect 1199 7219 4195 7389
rect 1199 2171 1559 7219
rect 4025 2171 4195 7219
rect 1199 2001 4195 2171
rect 1199 1771 1559 2001
rect 4025 1771 4195 2001
rect 1199 379 4195 1771
rect -59 359 4195 379
rect -59 209 1369 359
<< pwell >>
rect 171 10496 1139 10726
rect 171 8729 259 10496
rect 1051 8729 1139 10496
rect 171 8481 1139 8729
rect 171 6714 259 8481
rect 1051 6714 1139 8481
rect 171 6466 1139 6714
rect 171 4699 259 6466
rect 1051 4699 1139 6466
rect 171 4451 1139 4699
rect 171 2684 259 4451
rect 1051 2684 1139 4451
rect 171 2436 1139 2684
rect 171 669 259 2436
rect 1051 669 1139 2436
rect 171 439 1139 669
rect 1663 10662 8287 10750
rect 1663 8804 1751 10662
rect 8199 8804 8287 10662
rect 1619 8716 8287 8804
rect 1619 7537 1707 8716
rect 1619 7449 4165 7537
rect 1619 7049 3965 7137
rect 1619 2319 1707 7049
rect 3877 2319 3965 7049
rect 1619 2231 3965 2319
<< mvndiff >>
rect 307 10582 373 10590
rect 307 10548 323 10582
rect 357 10548 373 10582
rect 307 10522 373 10548
rect 433 10582 499 10590
rect 433 10548 449 10582
rect 483 10548 499 10582
rect 433 10522 499 10548
rect 559 10582 625 10590
rect 559 10548 575 10582
rect 609 10548 625 10582
rect 559 10522 625 10548
rect 685 10582 751 10590
rect 685 10548 701 10582
rect 735 10548 751 10582
rect 685 10522 751 10548
rect 811 10582 877 10590
rect 811 10548 827 10582
rect 861 10548 877 10582
rect 811 10522 877 10548
rect 937 10582 1003 10590
rect 937 10548 953 10582
rect 987 10548 1003 10582
rect 937 10522 1003 10548
rect 307 8677 373 8703
rect 307 8643 323 8677
rect 357 8643 373 8677
rect 307 8635 373 8643
rect 433 8677 499 8703
rect 433 8643 449 8677
rect 483 8643 499 8677
rect 433 8635 499 8643
rect 559 8677 625 8703
rect 559 8643 575 8677
rect 609 8643 625 8677
rect 559 8635 625 8643
rect 685 8677 751 8703
rect 685 8643 701 8677
rect 735 8643 751 8677
rect 685 8635 751 8643
rect 811 8677 877 8703
rect 811 8643 827 8677
rect 861 8643 877 8677
rect 811 8635 877 8643
rect 937 8677 1003 8703
rect 937 8643 953 8677
rect 987 8643 1003 8677
rect 937 8635 1003 8643
rect 307 8567 373 8575
rect 307 8533 323 8567
rect 357 8533 373 8567
rect 307 8507 373 8533
rect 433 8567 499 8575
rect 433 8533 449 8567
rect 483 8533 499 8567
rect 433 8507 499 8533
rect 559 8567 625 8575
rect 559 8533 575 8567
rect 609 8533 625 8567
rect 559 8507 625 8533
rect 685 8567 751 8575
rect 685 8533 701 8567
rect 735 8533 751 8567
rect 685 8507 751 8533
rect 811 8567 877 8575
rect 811 8533 827 8567
rect 861 8533 877 8567
rect 811 8507 877 8533
rect 937 8567 1003 8575
rect 937 8533 953 8567
rect 987 8533 1003 8567
rect 937 8507 1003 8533
rect 307 6662 373 6688
rect 307 6628 323 6662
rect 357 6628 373 6662
rect 307 6620 373 6628
rect 433 6662 499 6688
rect 433 6628 449 6662
rect 483 6628 499 6662
rect 433 6620 499 6628
rect 559 6662 625 6688
rect 559 6628 575 6662
rect 609 6628 625 6662
rect 559 6620 625 6628
rect 685 6662 751 6688
rect 685 6628 701 6662
rect 735 6628 751 6662
rect 685 6620 751 6628
rect 811 6662 877 6688
rect 811 6628 827 6662
rect 861 6628 877 6662
rect 811 6620 877 6628
rect 937 6662 1003 6688
rect 937 6628 953 6662
rect 987 6628 1003 6662
rect 937 6620 1003 6628
rect 307 6552 373 6560
rect 307 6518 323 6552
rect 357 6518 373 6552
rect 307 6492 373 6518
rect 433 6552 499 6560
rect 433 6518 449 6552
rect 483 6518 499 6552
rect 433 6492 499 6518
rect 559 6552 625 6560
rect 559 6518 575 6552
rect 609 6518 625 6552
rect 559 6492 625 6518
rect 685 6552 751 6560
rect 685 6518 701 6552
rect 735 6518 751 6552
rect 685 6492 751 6518
rect 811 6552 877 6560
rect 811 6518 827 6552
rect 861 6518 877 6552
rect 811 6492 877 6518
rect 937 6552 1003 6560
rect 937 6518 953 6552
rect 987 6518 1003 6552
rect 937 6492 1003 6518
rect 307 4647 373 4673
rect 307 4613 323 4647
rect 357 4613 373 4647
rect 307 4605 373 4613
rect 433 4647 499 4673
rect 433 4613 449 4647
rect 483 4613 499 4647
rect 433 4605 499 4613
rect 559 4647 625 4673
rect 559 4613 575 4647
rect 609 4613 625 4647
rect 559 4605 625 4613
rect 685 4647 751 4673
rect 685 4613 701 4647
rect 735 4613 751 4647
rect 685 4605 751 4613
rect 811 4647 877 4673
rect 811 4613 827 4647
rect 861 4613 877 4647
rect 811 4605 877 4613
rect 937 4647 1003 4673
rect 937 4613 953 4647
rect 987 4613 1003 4647
rect 937 4605 1003 4613
rect 307 4537 373 4545
rect 307 4503 323 4537
rect 357 4503 373 4537
rect 307 4477 373 4503
rect 433 4537 499 4545
rect 433 4503 449 4537
rect 483 4503 499 4537
rect 433 4477 499 4503
rect 559 4537 625 4545
rect 559 4503 575 4537
rect 609 4503 625 4537
rect 559 4477 625 4503
rect 685 4537 751 4545
rect 685 4503 701 4537
rect 735 4503 751 4537
rect 685 4477 751 4503
rect 811 4537 877 4545
rect 811 4503 827 4537
rect 861 4503 877 4537
rect 811 4477 877 4503
rect 937 4537 1003 4545
rect 937 4503 953 4537
rect 987 4503 1003 4537
rect 937 4477 1003 4503
rect 307 2632 373 2658
rect 307 2598 323 2632
rect 357 2598 373 2632
rect 307 2590 373 2598
rect 433 2632 499 2658
rect 433 2598 449 2632
rect 483 2598 499 2632
rect 433 2590 499 2598
rect 559 2632 625 2658
rect 559 2598 575 2632
rect 609 2598 625 2632
rect 559 2590 625 2598
rect 685 2632 751 2658
rect 685 2598 701 2632
rect 735 2598 751 2632
rect 685 2590 751 2598
rect 811 2632 877 2658
rect 811 2598 827 2632
rect 861 2598 877 2632
rect 811 2590 877 2598
rect 937 2632 1003 2658
rect 937 2598 953 2632
rect 987 2598 1003 2632
rect 937 2590 1003 2598
rect 307 2522 373 2530
rect 307 2488 323 2522
rect 357 2488 373 2522
rect 307 2462 373 2488
rect 433 2522 499 2530
rect 433 2488 449 2522
rect 483 2488 499 2522
rect 433 2462 499 2488
rect 559 2522 625 2530
rect 559 2488 575 2522
rect 609 2488 625 2522
rect 559 2462 625 2488
rect 685 2522 751 2530
rect 685 2488 701 2522
rect 735 2488 751 2522
rect 685 2462 751 2488
rect 811 2522 877 2530
rect 811 2488 827 2522
rect 861 2488 877 2522
rect 811 2462 877 2488
rect 937 2522 1003 2530
rect 937 2488 953 2522
rect 987 2488 1003 2522
rect 937 2462 1003 2488
rect 307 617 373 643
rect 307 583 323 617
rect 357 583 373 617
rect 307 575 373 583
rect 433 617 499 643
rect 433 583 449 617
rect 483 583 499 617
rect 433 575 499 583
rect 559 617 625 643
rect 559 583 575 617
rect 609 583 625 617
rect 559 575 625 583
rect 685 617 751 643
rect 685 583 701 617
rect 735 583 751 617
rect 685 575 751 583
rect 811 617 877 643
rect 811 583 827 617
rect 861 583 877 617
rect 811 575 877 583
rect 937 617 1003 643
rect 937 583 953 617
rect 987 583 1003 617
rect 937 575 1003 583
<< mvndiffc >>
rect 323 10548 357 10582
rect 449 10548 483 10582
rect 575 10548 609 10582
rect 701 10548 735 10582
rect 827 10548 861 10582
rect 953 10548 987 10582
rect 323 8643 357 8677
rect 449 8643 483 8677
rect 575 8643 609 8677
rect 701 8643 735 8677
rect 827 8643 861 8677
rect 953 8643 987 8677
rect 323 8533 357 8567
rect 449 8533 483 8567
rect 575 8533 609 8567
rect 701 8533 735 8567
rect 827 8533 861 8567
rect 953 8533 987 8567
rect 323 6628 357 6662
rect 449 6628 483 6662
rect 575 6628 609 6662
rect 701 6628 735 6662
rect 827 6628 861 6662
rect 953 6628 987 6662
rect 323 6518 357 6552
rect 449 6518 483 6552
rect 575 6518 609 6552
rect 701 6518 735 6552
rect 827 6518 861 6552
rect 953 6518 987 6552
rect 323 4613 357 4647
rect 449 4613 483 4647
rect 575 4613 609 4647
rect 701 4613 735 4647
rect 827 4613 861 4647
rect 953 4613 987 4647
rect 323 4503 357 4537
rect 449 4503 483 4537
rect 575 4503 609 4537
rect 701 4503 735 4537
rect 827 4503 861 4537
rect 953 4503 987 4537
rect 323 2598 357 2632
rect 449 2598 483 2632
rect 575 2598 609 2632
rect 701 2598 735 2632
rect 827 2598 861 2632
rect 953 2598 987 2632
rect 323 2488 357 2522
rect 449 2488 483 2522
rect 575 2488 609 2522
rect 701 2488 735 2522
rect 827 2488 861 2522
rect 953 2488 987 2522
rect 323 583 357 617
rect 449 583 483 617
rect 575 583 609 617
rect 701 583 735 617
rect 827 583 861 617
rect 953 583 987 617
<< mvpsubdiff >>
rect 197 10699 1113 10700
rect 197 10666 297 10699
rect 197 10632 198 10666
rect 232 10665 297 10666
rect 331 10665 365 10699
rect 399 10665 433 10699
rect 467 10665 501 10699
rect 535 10665 569 10699
rect 603 10665 637 10699
rect 671 10665 705 10699
rect 739 10665 773 10699
rect 807 10665 841 10699
rect 875 10665 909 10699
rect 943 10665 977 10699
rect 1011 10665 1045 10699
rect 1079 10665 1113 10699
rect 232 10664 1113 10665
rect 232 10632 233 10664
rect 197 10598 233 10632
rect 197 10564 198 10598
rect 232 10564 233 10598
rect 1077 10597 1113 10664
rect 197 10530 233 10564
rect 197 10496 198 10530
rect 232 10496 233 10530
rect 1077 10563 1078 10597
rect 1112 10563 1113 10597
rect 1077 10529 1113 10563
rect 197 10462 233 10496
rect 197 10428 198 10462
rect 232 10428 233 10462
rect 197 10394 233 10428
rect 197 10360 198 10394
rect 232 10360 233 10394
rect 197 10326 233 10360
rect 197 10292 198 10326
rect 232 10292 233 10326
rect 197 10258 233 10292
rect 197 10224 198 10258
rect 232 10224 233 10258
rect 197 10190 233 10224
rect 197 10156 198 10190
rect 232 10156 233 10190
rect 197 10122 233 10156
rect 197 10088 198 10122
rect 232 10088 233 10122
rect 197 10054 233 10088
rect 197 10020 198 10054
rect 232 10020 233 10054
rect 197 9986 233 10020
rect 197 9952 198 9986
rect 232 9952 233 9986
rect 197 9918 233 9952
rect 197 9884 198 9918
rect 232 9884 233 9918
rect 197 9850 233 9884
rect 197 9816 198 9850
rect 232 9816 233 9850
rect 197 9782 233 9816
rect 197 9748 198 9782
rect 232 9748 233 9782
rect 197 9714 233 9748
rect 197 9680 198 9714
rect 232 9680 233 9714
rect 197 9646 233 9680
rect 197 9612 198 9646
rect 232 9612 233 9646
rect 197 9578 233 9612
rect 197 9544 198 9578
rect 232 9544 233 9578
rect 197 9510 233 9544
rect 197 9476 198 9510
rect 232 9476 233 9510
rect 197 9442 233 9476
rect 197 9408 198 9442
rect 232 9408 233 9442
rect 197 9374 233 9408
rect 197 9340 198 9374
rect 232 9340 233 9374
rect 197 9306 233 9340
rect 197 9272 198 9306
rect 232 9272 233 9306
rect 197 9238 233 9272
rect 197 9204 198 9238
rect 232 9204 233 9238
rect 197 9170 233 9204
rect 197 9136 198 9170
rect 232 9136 233 9170
rect 197 9102 233 9136
rect 197 9068 198 9102
rect 232 9068 233 9102
rect 197 9034 233 9068
rect 197 9000 198 9034
rect 232 9000 233 9034
rect 197 8966 233 9000
rect 197 8932 198 8966
rect 232 8932 233 8966
rect 197 8898 233 8932
rect 197 8864 198 8898
rect 232 8864 233 8898
rect 197 8830 233 8864
rect 197 8796 198 8830
rect 232 8796 233 8830
rect 197 8762 233 8796
rect 197 8728 198 8762
rect 232 8728 233 8762
rect 197 8694 233 8728
rect 1077 10495 1078 10529
rect 1112 10495 1113 10529
rect 1077 10461 1113 10495
rect 1077 10427 1078 10461
rect 1112 10427 1113 10461
rect 1077 10393 1113 10427
rect 1077 10359 1078 10393
rect 1112 10359 1113 10393
rect 1077 10325 1113 10359
rect 1077 10291 1078 10325
rect 1112 10291 1113 10325
rect 1077 10257 1113 10291
rect 1077 10223 1078 10257
rect 1112 10223 1113 10257
rect 1077 10189 1113 10223
rect 1077 10155 1078 10189
rect 1112 10155 1113 10189
rect 1077 10121 1113 10155
rect 1077 10087 1078 10121
rect 1112 10087 1113 10121
rect 1077 10053 1113 10087
rect 1077 10019 1078 10053
rect 1112 10019 1113 10053
rect 1077 9985 1113 10019
rect 1077 9951 1078 9985
rect 1112 9951 1113 9985
rect 1077 9917 1113 9951
rect 1077 9883 1078 9917
rect 1112 9883 1113 9917
rect 1077 9849 1113 9883
rect 1077 9815 1078 9849
rect 1112 9815 1113 9849
rect 1077 9781 1113 9815
rect 1077 9747 1078 9781
rect 1112 9747 1113 9781
rect 1077 9713 1113 9747
rect 1077 9679 1078 9713
rect 1112 9679 1113 9713
rect 1077 9645 1113 9679
rect 1077 9611 1078 9645
rect 1112 9611 1113 9645
rect 1077 9577 1113 9611
rect 1077 9543 1078 9577
rect 1112 9543 1113 9577
rect 1077 9509 1113 9543
rect 1077 9475 1078 9509
rect 1112 9475 1113 9509
rect 1077 9441 1113 9475
rect 1077 9407 1078 9441
rect 1112 9407 1113 9441
rect 1077 9373 1113 9407
rect 1077 9339 1078 9373
rect 1112 9339 1113 9373
rect 1077 9305 1113 9339
rect 1077 9271 1078 9305
rect 1112 9271 1113 9305
rect 1077 9237 1113 9271
rect 1077 9203 1078 9237
rect 1112 9203 1113 9237
rect 1077 9169 1113 9203
rect 1077 9135 1078 9169
rect 1112 9135 1113 9169
rect 1077 9101 1113 9135
rect 1077 9067 1078 9101
rect 1112 9067 1113 9101
rect 1077 9033 1113 9067
rect 1077 8999 1078 9033
rect 1112 8999 1113 9033
rect 1077 8965 1113 8999
rect 1077 8931 1078 8965
rect 1112 8931 1113 8965
rect 1077 8897 1113 8931
rect 1077 8863 1078 8897
rect 1112 8863 1113 8897
rect 1077 8829 1113 8863
rect 1077 8795 1078 8829
rect 1112 8795 1113 8829
rect 1077 8761 1113 8795
rect 1077 8727 1078 8761
rect 1112 8727 1113 8761
rect 197 8660 198 8694
rect 232 8660 233 8694
rect 197 8626 233 8660
rect 1077 8693 1113 8727
rect 1077 8659 1078 8693
rect 1112 8659 1113 8693
rect 197 8592 198 8626
rect 232 8592 233 8626
rect 197 8558 233 8592
rect 1077 8625 1113 8659
rect 1077 8591 1078 8625
rect 1112 8591 1113 8625
rect 197 8524 198 8558
rect 232 8524 233 8558
rect 197 8490 233 8524
rect 1077 8557 1113 8591
rect 1077 8523 1078 8557
rect 1112 8523 1113 8557
rect 197 8456 198 8490
rect 232 8456 233 8490
rect 197 8422 233 8456
rect 197 8388 198 8422
rect 232 8388 233 8422
rect 197 8354 233 8388
rect 197 8320 198 8354
rect 232 8320 233 8354
rect 197 8286 233 8320
rect 197 8252 198 8286
rect 232 8252 233 8286
rect 197 8218 233 8252
rect 197 8184 198 8218
rect 232 8184 233 8218
rect 197 8150 233 8184
rect 197 8116 198 8150
rect 232 8116 233 8150
rect 197 8082 233 8116
rect 197 8048 198 8082
rect 232 8048 233 8082
rect 197 8014 233 8048
rect 197 7980 198 8014
rect 232 7980 233 8014
rect 197 7946 233 7980
rect 197 7912 198 7946
rect 232 7912 233 7946
rect 197 7878 233 7912
rect 197 7844 198 7878
rect 232 7844 233 7878
rect 197 7810 233 7844
rect 197 7776 198 7810
rect 232 7776 233 7810
rect 197 7742 233 7776
rect 197 7708 198 7742
rect 232 7708 233 7742
rect 197 7674 233 7708
rect 197 7640 198 7674
rect 232 7640 233 7674
rect 197 7606 233 7640
rect 197 7572 198 7606
rect 232 7572 233 7606
rect 197 7538 233 7572
rect 197 7504 198 7538
rect 232 7504 233 7538
rect 197 7470 233 7504
rect 197 7436 198 7470
rect 232 7436 233 7470
rect 197 7402 233 7436
rect 197 7368 198 7402
rect 232 7368 233 7402
rect 197 7334 233 7368
rect 197 7300 198 7334
rect 232 7300 233 7334
rect 197 7266 233 7300
rect 197 7232 198 7266
rect 232 7232 233 7266
rect 197 7198 233 7232
rect 197 7164 198 7198
rect 232 7164 233 7198
rect 197 7130 233 7164
rect 197 7096 198 7130
rect 232 7096 233 7130
rect 197 7062 233 7096
rect 197 7028 198 7062
rect 232 7028 233 7062
rect 197 6994 233 7028
rect 197 6960 198 6994
rect 232 6960 233 6994
rect 197 6926 233 6960
rect 197 6892 198 6926
rect 232 6892 233 6926
rect 197 6858 233 6892
rect 197 6824 198 6858
rect 232 6824 233 6858
rect 197 6790 233 6824
rect 197 6756 198 6790
rect 232 6756 233 6790
rect 197 6722 233 6756
rect 197 6688 198 6722
rect 232 6688 233 6722
rect 1077 8489 1113 8523
rect 1077 8455 1078 8489
rect 1112 8455 1113 8489
rect 1077 8421 1113 8455
rect 1077 8387 1078 8421
rect 1112 8387 1113 8421
rect 1077 8353 1113 8387
rect 1077 8319 1078 8353
rect 1112 8319 1113 8353
rect 1077 8285 1113 8319
rect 1077 8251 1078 8285
rect 1112 8251 1113 8285
rect 1077 8217 1113 8251
rect 1077 8183 1078 8217
rect 1112 8183 1113 8217
rect 1077 8149 1113 8183
rect 1077 8115 1078 8149
rect 1112 8115 1113 8149
rect 1077 8081 1113 8115
rect 1077 8047 1078 8081
rect 1112 8047 1113 8081
rect 1077 8013 1113 8047
rect 1077 7979 1078 8013
rect 1112 7979 1113 8013
rect 1077 7945 1113 7979
rect 1077 7911 1078 7945
rect 1112 7911 1113 7945
rect 1077 7877 1113 7911
rect 1077 7843 1078 7877
rect 1112 7843 1113 7877
rect 1077 7809 1113 7843
rect 1077 7775 1078 7809
rect 1112 7775 1113 7809
rect 1077 7741 1113 7775
rect 1077 7707 1078 7741
rect 1112 7707 1113 7741
rect 1077 7673 1113 7707
rect 1077 7639 1078 7673
rect 1112 7639 1113 7673
rect 1077 7605 1113 7639
rect 1077 7571 1078 7605
rect 1112 7571 1113 7605
rect 1077 7537 1113 7571
rect 1077 7503 1078 7537
rect 1112 7503 1113 7537
rect 1077 7469 1113 7503
rect 1077 7435 1078 7469
rect 1112 7435 1113 7469
rect 1077 7401 1113 7435
rect 1077 7367 1078 7401
rect 1112 7367 1113 7401
rect 1077 7333 1113 7367
rect 1077 7299 1078 7333
rect 1112 7299 1113 7333
rect 1077 7265 1113 7299
rect 1077 7231 1078 7265
rect 1112 7231 1113 7265
rect 1077 7197 1113 7231
rect 1077 7163 1078 7197
rect 1112 7163 1113 7197
rect 1077 7129 1113 7163
rect 1077 7095 1078 7129
rect 1112 7095 1113 7129
rect 1077 7061 1113 7095
rect 1077 7027 1078 7061
rect 1112 7027 1113 7061
rect 1077 6993 1113 7027
rect 1077 6959 1078 6993
rect 1112 6959 1113 6993
rect 1077 6925 1113 6959
rect 1077 6891 1078 6925
rect 1112 6891 1113 6925
rect 1077 6857 1113 6891
rect 1077 6823 1078 6857
rect 1112 6823 1113 6857
rect 1077 6789 1113 6823
rect 1077 6755 1078 6789
rect 1112 6755 1113 6789
rect 1077 6721 1113 6755
rect 197 6654 233 6688
rect 197 6620 198 6654
rect 232 6620 233 6654
rect 1077 6687 1078 6721
rect 1112 6687 1113 6721
rect 1077 6653 1113 6687
rect 197 6586 233 6620
rect 197 6552 198 6586
rect 232 6552 233 6586
rect 1077 6619 1078 6653
rect 1112 6619 1113 6653
rect 1077 6585 1113 6619
rect 197 6518 233 6552
rect 197 6484 198 6518
rect 232 6484 233 6518
rect 1077 6551 1078 6585
rect 1112 6551 1113 6585
rect 1077 6517 1113 6551
rect 197 6450 233 6484
rect 197 6416 198 6450
rect 232 6416 233 6450
rect 197 6382 233 6416
rect 197 6348 198 6382
rect 232 6348 233 6382
rect 197 6314 233 6348
rect 197 6280 198 6314
rect 232 6280 233 6314
rect 197 6246 233 6280
rect 197 6212 198 6246
rect 232 6212 233 6246
rect 197 6178 233 6212
rect 197 6144 198 6178
rect 232 6144 233 6178
rect 197 6110 233 6144
rect 197 6076 198 6110
rect 232 6076 233 6110
rect 197 6042 233 6076
rect 197 6008 198 6042
rect 232 6008 233 6042
rect 197 5974 233 6008
rect 197 5940 198 5974
rect 232 5940 233 5974
rect 197 5906 233 5940
rect 197 5872 198 5906
rect 232 5872 233 5906
rect 197 5838 233 5872
rect 197 5804 198 5838
rect 232 5804 233 5838
rect 197 5770 233 5804
rect 197 5736 198 5770
rect 232 5736 233 5770
rect 197 5702 233 5736
rect 197 5668 198 5702
rect 232 5668 233 5702
rect 197 5634 233 5668
rect 197 5600 198 5634
rect 232 5600 233 5634
rect 197 5566 233 5600
rect 197 5532 198 5566
rect 232 5532 233 5566
rect 197 5498 233 5532
rect 197 5464 198 5498
rect 232 5464 233 5498
rect 197 5430 233 5464
rect 197 5396 198 5430
rect 232 5396 233 5430
rect 197 5362 233 5396
rect 197 5328 198 5362
rect 232 5328 233 5362
rect 197 5294 233 5328
rect 197 5260 198 5294
rect 232 5260 233 5294
rect 197 5226 233 5260
rect 197 5192 198 5226
rect 232 5192 233 5226
rect 197 5158 233 5192
rect 197 5124 198 5158
rect 232 5124 233 5158
rect 197 5090 233 5124
rect 197 5056 198 5090
rect 232 5056 233 5090
rect 197 5022 233 5056
rect 197 4988 198 5022
rect 232 4988 233 5022
rect 197 4954 233 4988
rect 197 4920 198 4954
rect 232 4920 233 4954
rect 197 4886 233 4920
rect 197 4852 198 4886
rect 232 4852 233 4886
rect 197 4818 233 4852
rect 197 4784 198 4818
rect 232 4784 233 4818
rect 197 4750 233 4784
rect 197 4716 198 4750
rect 232 4716 233 4750
rect 197 4682 233 4716
rect 197 4648 198 4682
rect 232 4648 233 4682
rect 1077 6483 1078 6517
rect 1112 6483 1113 6517
rect 1077 6449 1113 6483
rect 1077 6415 1078 6449
rect 1112 6415 1113 6449
rect 1077 6381 1113 6415
rect 1077 6347 1078 6381
rect 1112 6347 1113 6381
rect 1077 6313 1113 6347
rect 1077 6279 1078 6313
rect 1112 6279 1113 6313
rect 1077 6245 1113 6279
rect 1077 6211 1078 6245
rect 1112 6211 1113 6245
rect 1077 6177 1113 6211
rect 1077 6143 1078 6177
rect 1112 6143 1113 6177
rect 1077 6109 1113 6143
rect 1077 6075 1078 6109
rect 1112 6075 1113 6109
rect 1077 6041 1113 6075
rect 1077 6007 1078 6041
rect 1112 6007 1113 6041
rect 1077 5973 1113 6007
rect 1077 5939 1078 5973
rect 1112 5939 1113 5973
rect 1077 5905 1113 5939
rect 1077 5871 1078 5905
rect 1112 5871 1113 5905
rect 1077 5837 1113 5871
rect 1077 5803 1078 5837
rect 1112 5803 1113 5837
rect 1077 5769 1113 5803
rect 1077 5735 1078 5769
rect 1112 5735 1113 5769
rect 1077 5701 1113 5735
rect 1077 5667 1078 5701
rect 1112 5667 1113 5701
rect 1077 5633 1113 5667
rect 1077 5599 1078 5633
rect 1112 5599 1113 5633
rect 1077 5565 1113 5599
rect 1077 5531 1078 5565
rect 1112 5531 1113 5565
rect 1077 5497 1113 5531
rect 1077 5463 1078 5497
rect 1112 5463 1113 5497
rect 1077 5429 1113 5463
rect 1077 5395 1078 5429
rect 1112 5395 1113 5429
rect 1077 5361 1113 5395
rect 1077 5327 1078 5361
rect 1112 5327 1113 5361
rect 1077 5293 1113 5327
rect 1077 5259 1078 5293
rect 1112 5259 1113 5293
rect 1077 5225 1113 5259
rect 1077 5191 1078 5225
rect 1112 5191 1113 5225
rect 1077 5157 1113 5191
rect 1077 5123 1078 5157
rect 1112 5123 1113 5157
rect 1077 5089 1113 5123
rect 1077 5055 1078 5089
rect 1112 5055 1113 5089
rect 1077 5021 1113 5055
rect 1077 4987 1078 5021
rect 1112 4987 1113 5021
rect 1077 4953 1113 4987
rect 1077 4919 1078 4953
rect 1112 4919 1113 4953
rect 1077 4885 1113 4919
rect 1077 4851 1078 4885
rect 1112 4851 1113 4885
rect 1077 4817 1113 4851
rect 1077 4783 1078 4817
rect 1112 4783 1113 4817
rect 1077 4749 1113 4783
rect 1077 4715 1078 4749
rect 1112 4715 1113 4749
rect 1077 4681 1113 4715
rect 197 4614 233 4648
rect 197 4580 198 4614
rect 232 4580 233 4614
rect 1077 4647 1078 4681
rect 1112 4647 1113 4681
rect 1077 4613 1113 4647
rect 197 4546 233 4580
rect 197 4512 198 4546
rect 232 4512 233 4546
rect 1077 4579 1078 4613
rect 1112 4579 1113 4613
rect 1077 4545 1113 4579
rect 197 4478 233 4512
rect 197 4444 198 4478
rect 232 4444 233 4478
rect 1077 4511 1078 4545
rect 1112 4511 1113 4545
rect 1077 4477 1113 4511
rect 197 4410 233 4444
rect 197 4376 198 4410
rect 232 4376 233 4410
rect 197 4342 233 4376
rect 197 4308 198 4342
rect 232 4308 233 4342
rect 197 4274 233 4308
rect 197 4240 198 4274
rect 232 4240 233 4274
rect 197 4206 233 4240
rect 197 4172 198 4206
rect 232 4172 233 4206
rect 197 4138 233 4172
rect 197 4104 198 4138
rect 232 4104 233 4138
rect 197 4070 233 4104
rect 197 4036 198 4070
rect 232 4036 233 4070
rect 197 4002 233 4036
rect 197 3968 198 4002
rect 232 3968 233 4002
rect 197 3934 233 3968
rect 197 3900 198 3934
rect 232 3900 233 3934
rect 197 3866 233 3900
rect 197 3832 198 3866
rect 232 3832 233 3866
rect 197 3798 233 3832
rect 197 3764 198 3798
rect 232 3764 233 3798
rect 197 3730 233 3764
rect 197 3696 198 3730
rect 232 3696 233 3730
rect 197 3662 233 3696
rect 197 3628 198 3662
rect 232 3628 233 3662
rect 197 3594 233 3628
rect 197 3560 198 3594
rect 232 3560 233 3594
rect 197 3526 233 3560
rect 197 3492 198 3526
rect 232 3492 233 3526
rect 197 3458 233 3492
rect 197 3424 198 3458
rect 232 3424 233 3458
rect 197 3390 233 3424
rect 197 3356 198 3390
rect 232 3356 233 3390
rect 197 3322 233 3356
rect 197 3288 198 3322
rect 232 3288 233 3322
rect 197 3254 233 3288
rect 197 3220 198 3254
rect 232 3220 233 3254
rect 197 3186 233 3220
rect 197 3152 198 3186
rect 232 3152 233 3186
rect 197 3118 233 3152
rect 197 3084 198 3118
rect 232 3084 233 3118
rect 197 3050 233 3084
rect 197 3016 198 3050
rect 232 3016 233 3050
rect 197 2982 233 3016
rect 197 2948 198 2982
rect 232 2948 233 2982
rect 197 2914 233 2948
rect 197 2880 198 2914
rect 232 2880 233 2914
rect 197 2846 233 2880
rect 197 2812 198 2846
rect 232 2812 233 2846
rect 197 2778 233 2812
rect 197 2744 198 2778
rect 232 2744 233 2778
rect 197 2710 233 2744
rect 197 2676 198 2710
rect 232 2676 233 2710
rect 197 2642 233 2676
rect 1077 4443 1078 4477
rect 1112 4443 1113 4477
rect 1077 4409 1113 4443
rect 1077 4375 1078 4409
rect 1112 4375 1113 4409
rect 1077 4341 1113 4375
rect 1077 4307 1078 4341
rect 1112 4307 1113 4341
rect 1077 4273 1113 4307
rect 1077 4239 1078 4273
rect 1112 4239 1113 4273
rect 1077 4205 1113 4239
rect 1077 4171 1078 4205
rect 1112 4171 1113 4205
rect 1077 4137 1113 4171
rect 1077 4103 1078 4137
rect 1112 4103 1113 4137
rect 1077 4069 1113 4103
rect 1077 4035 1078 4069
rect 1112 4035 1113 4069
rect 1077 4001 1113 4035
rect 1077 3967 1078 4001
rect 1112 3967 1113 4001
rect 1077 3933 1113 3967
rect 1077 3899 1078 3933
rect 1112 3899 1113 3933
rect 1077 3865 1113 3899
rect 1077 3831 1078 3865
rect 1112 3831 1113 3865
rect 1077 3797 1113 3831
rect 1077 3763 1078 3797
rect 1112 3763 1113 3797
rect 1077 3729 1113 3763
rect 1077 3695 1078 3729
rect 1112 3695 1113 3729
rect 1077 3661 1113 3695
rect 1077 3627 1078 3661
rect 1112 3627 1113 3661
rect 1077 3593 1113 3627
rect 1077 3559 1078 3593
rect 1112 3559 1113 3593
rect 1077 3525 1113 3559
rect 1077 3491 1078 3525
rect 1112 3491 1113 3525
rect 1077 3457 1113 3491
rect 1077 3423 1078 3457
rect 1112 3423 1113 3457
rect 1077 3389 1113 3423
rect 1077 3355 1078 3389
rect 1112 3355 1113 3389
rect 1077 3321 1113 3355
rect 1077 3287 1078 3321
rect 1112 3287 1113 3321
rect 1077 3253 1113 3287
rect 1077 3219 1078 3253
rect 1112 3219 1113 3253
rect 1077 3185 1113 3219
rect 1077 3151 1078 3185
rect 1112 3151 1113 3185
rect 1077 3117 1113 3151
rect 1077 3083 1078 3117
rect 1112 3083 1113 3117
rect 1077 3049 1113 3083
rect 1077 3015 1078 3049
rect 1112 3015 1113 3049
rect 1077 2981 1113 3015
rect 1077 2947 1078 2981
rect 1112 2947 1113 2981
rect 1077 2913 1113 2947
rect 1077 2879 1078 2913
rect 1112 2879 1113 2913
rect 1077 2845 1113 2879
rect 1077 2811 1078 2845
rect 1112 2811 1113 2845
rect 1077 2777 1113 2811
rect 1077 2743 1078 2777
rect 1112 2743 1113 2777
rect 1077 2709 1113 2743
rect 1077 2675 1078 2709
rect 1112 2675 1113 2709
rect 197 2608 198 2642
rect 232 2608 233 2642
rect 197 2574 233 2608
rect 1077 2641 1113 2675
rect 1077 2607 1078 2641
rect 1112 2607 1113 2641
rect 197 2540 198 2574
rect 232 2540 233 2574
rect 197 2506 233 2540
rect 1077 2573 1113 2607
rect 1077 2539 1078 2573
rect 1112 2539 1113 2573
rect 197 2472 198 2506
rect 232 2472 233 2506
rect 197 2438 233 2472
rect 1077 2505 1113 2539
rect 1077 2471 1078 2505
rect 1112 2471 1113 2505
rect 197 2404 198 2438
rect 232 2404 233 2438
rect 197 2370 233 2404
rect 197 2336 198 2370
rect 232 2336 233 2370
rect 197 2302 233 2336
rect 197 2268 198 2302
rect 232 2268 233 2302
rect 197 2234 233 2268
rect 197 2200 198 2234
rect 232 2200 233 2234
rect 197 2166 233 2200
rect 197 2132 198 2166
rect 232 2132 233 2166
rect 197 2098 233 2132
rect 197 2064 198 2098
rect 232 2064 233 2098
rect 197 2030 233 2064
rect 197 1996 198 2030
rect 232 1996 233 2030
rect 197 1962 233 1996
rect 197 1928 198 1962
rect 232 1928 233 1962
rect 197 1894 233 1928
rect 197 1860 198 1894
rect 232 1860 233 1894
rect 197 1826 233 1860
rect 197 1792 198 1826
rect 232 1792 233 1826
rect 197 1758 233 1792
rect 197 1724 198 1758
rect 232 1724 233 1758
rect 197 1690 233 1724
rect 197 1656 198 1690
rect 232 1656 233 1690
rect 197 1622 233 1656
rect 197 1588 198 1622
rect 232 1588 233 1622
rect 197 1554 233 1588
rect 197 1520 198 1554
rect 232 1520 233 1554
rect 197 1486 233 1520
rect 197 1452 198 1486
rect 232 1452 233 1486
rect 197 1418 233 1452
rect 197 1384 198 1418
rect 232 1384 233 1418
rect 197 1350 233 1384
rect 197 1316 198 1350
rect 232 1316 233 1350
rect 197 1282 233 1316
rect 197 1248 198 1282
rect 232 1248 233 1282
rect 197 1214 233 1248
rect 197 1180 198 1214
rect 232 1180 233 1214
rect 197 1146 233 1180
rect 197 1112 198 1146
rect 232 1112 233 1146
rect 197 1078 233 1112
rect 197 1044 198 1078
rect 232 1044 233 1078
rect 197 1010 233 1044
rect 197 976 198 1010
rect 232 976 233 1010
rect 197 942 233 976
rect 197 908 198 942
rect 232 908 233 942
rect 197 874 233 908
rect 197 840 198 874
rect 232 840 233 874
rect 197 806 233 840
rect 197 772 198 806
rect 232 772 233 806
rect 197 738 233 772
rect 197 704 198 738
rect 232 704 233 738
rect 197 670 233 704
rect 197 636 198 670
rect 232 636 233 670
rect 1077 2437 1113 2471
rect 1077 2403 1078 2437
rect 1112 2403 1113 2437
rect 1077 2369 1113 2403
rect 1077 2335 1078 2369
rect 1112 2335 1113 2369
rect 1077 2301 1113 2335
rect 1077 2267 1078 2301
rect 1112 2267 1113 2301
rect 1077 2233 1113 2267
rect 1077 2199 1078 2233
rect 1112 2199 1113 2233
rect 1077 2165 1113 2199
rect 1077 2131 1078 2165
rect 1112 2131 1113 2165
rect 1077 2097 1113 2131
rect 1077 2063 1078 2097
rect 1112 2063 1113 2097
rect 1077 2029 1113 2063
rect 1077 1995 1078 2029
rect 1112 1995 1113 2029
rect 1077 1961 1113 1995
rect 1077 1927 1078 1961
rect 1112 1927 1113 1961
rect 1077 1893 1113 1927
rect 1077 1859 1078 1893
rect 1112 1859 1113 1893
rect 1077 1825 1113 1859
rect 1077 1791 1078 1825
rect 1112 1791 1113 1825
rect 1077 1757 1113 1791
rect 1077 1723 1078 1757
rect 1112 1723 1113 1757
rect 1077 1689 1113 1723
rect 1077 1655 1078 1689
rect 1112 1655 1113 1689
rect 1077 1621 1113 1655
rect 1077 1587 1078 1621
rect 1112 1587 1113 1621
rect 1077 1553 1113 1587
rect 1077 1519 1078 1553
rect 1112 1519 1113 1553
rect 1077 1485 1113 1519
rect 1077 1451 1078 1485
rect 1112 1451 1113 1485
rect 1077 1417 1113 1451
rect 1077 1383 1078 1417
rect 1112 1383 1113 1417
rect 1077 1349 1113 1383
rect 1077 1315 1078 1349
rect 1112 1315 1113 1349
rect 1077 1281 1113 1315
rect 1077 1247 1078 1281
rect 1112 1247 1113 1281
rect 1077 1213 1113 1247
rect 1077 1179 1078 1213
rect 1112 1179 1113 1213
rect 1077 1145 1113 1179
rect 1077 1111 1078 1145
rect 1112 1111 1113 1145
rect 1077 1077 1113 1111
rect 1077 1043 1078 1077
rect 1112 1043 1113 1077
rect 1077 1009 1113 1043
rect 1077 975 1078 1009
rect 1112 975 1113 1009
rect 1077 941 1113 975
rect 1077 907 1078 941
rect 1112 907 1113 941
rect 1077 873 1113 907
rect 1077 839 1078 873
rect 1112 839 1113 873
rect 1077 805 1113 839
rect 1077 771 1078 805
rect 1112 771 1113 805
rect 1077 737 1113 771
rect 1077 703 1078 737
rect 1112 703 1113 737
rect 1077 669 1113 703
rect 197 602 233 636
rect 197 568 198 602
rect 232 568 233 602
rect 1077 635 1078 669
rect 1112 635 1113 669
rect 1077 601 1113 635
rect 197 501 233 568
rect 1077 567 1078 601
rect 1112 567 1113 601
rect 1077 533 1113 567
rect 1077 501 1078 533
rect 197 500 1078 501
rect 197 466 231 500
rect 265 466 299 500
rect 333 466 367 500
rect 401 466 435 500
rect 469 466 503 500
rect 537 466 571 500
rect 605 466 639 500
rect 673 466 707 500
rect 741 466 775 500
rect 809 466 843 500
rect 877 466 911 500
rect 945 466 979 500
rect 1013 499 1078 500
rect 1112 499 1113 533
rect 1013 466 1113 499
rect 197 465 1113 466
rect 1689 10723 8261 10724
rect 1689 10690 1801 10723
rect 1689 10656 1690 10690
rect 1724 10689 1801 10690
rect 1835 10689 1869 10723
rect 1903 10689 1937 10723
rect 1971 10689 2005 10723
rect 2039 10689 2073 10723
rect 2107 10689 2141 10723
rect 2175 10689 2209 10723
rect 2243 10689 2277 10723
rect 2311 10689 2345 10723
rect 2379 10689 2413 10723
rect 2447 10689 2481 10723
rect 2515 10689 2549 10723
rect 2583 10689 2617 10723
rect 2651 10689 2685 10723
rect 2719 10689 2753 10723
rect 2787 10689 2821 10723
rect 2855 10689 2889 10723
rect 2923 10689 2957 10723
rect 2991 10689 3025 10723
rect 3059 10689 3093 10723
rect 3127 10689 3161 10723
rect 3195 10689 3229 10723
rect 3263 10689 3297 10723
rect 3331 10689 3365 10723
rect 3399 10689 3433 10723
rect 3467 10689 3501 10723
rect 3535 10689 3569 10723
rect 3603 10689 3637 10723
rect 3671 10689 3705 10723
rect 3739 10689 3773 10723
rect 3807 10689 3841 10723
rect 3875 10689 3909 10723
rect 3943 10689 3977 10723
rect 4011 10689 4045 10723
rect 4079 10689 4113 10723
rect 4147 10689 4181 10723
rect 4215 10689 4249 10723
rect 4283 10689 4317 10723
rect 4351 10689 4385 10723
rect 4419 10689 4453 10723
rect 4487 10689 4521 10723
rect 4555 10689 4589 10723
rect 4623 10689 4657 10723
rect 4691 10689 4725 10723
rect 4759 10689 4793 10723
rect 4827 10689 4861 10723
rect 4895 10689 4929 10723
rect 4963 10689 4997 10723
rect 5031 10689 5065 10723
rect 5099 10689 5133 10723
rect 5167 10689 5201 10723
rect 5235 10689 5269 10723
rect 5303 10689 5337 10723
rect 5371 10689 5405 10723
rect 5439 10689 5473 10723
rect 5507 10689 5541 10723
rect 5575 10689 5609 10723
rect 5643 10689 5677 10723
rect 5711 10689 5745 10723
rect 5779 10689 5813 10723
rect 5847 10689 5881 10723
rect 5915 10689 5949 10723
rect 5983 10689 6017 10723
rect 6051 10689 6085 10723
rect 6119 10689 6153 10723
rect 6187 10689 6221 10723
rect 6255 10689 6289 10723
rect 6323 10689 6357 10723
rect 6391 10689 6425 10723
rect 6459 10689 6493 10723
rect 6527 10689 6561 10723
rect 6595 10689 6629 10723
rect 6663 10689 6697 10723
rect 6731 10689 6765 10723
rect 6799 10689 6833 10723
rect 6867 10689 6901 10723
rect 6935 10689 6969 10723
rect 7003 10689 7037 10723
rect 7071 10689 7105 10723
rect 7139 10689 7173 10723
rect 7207 10689 7241 10723
rect 7275 10689 7309 10723
rect 7343 10689 7377 10723
rect 7411 10689 7445 10723
rect 7479 10689 7513 10723
rect 7547 10689 7581 10723
rect 7615 10689 7649 10723
rect 7683 10689 7717 10723
rect 7751 10689 7785 10723
rect 7819 10689 7853 10723
rect 7887 10689 7921 10723
rect 7955 10689 7989 10723
rect 8023 10689 8057 10723
rect 8091 10689 8125 10723
rect 8159 10689 8193 10723
rect 8227 10689 8261 10723
rect 1724 10688 8261 10689
rect 1724 10656 1725 10688
rect 1689 10622 1725 10656
rect 1689 10588 1690 10622
rect 1724 10588 1725 10622
rect 1689 10554 1725 10588
rect 8225 10646 8261 10688
rect 8225 10612 8226 10646
rect 8260 10612 8261 10646
rect 8225 10578 8261 10612
rect 1689 10520 1690 10554
rect 1724 10520 1725 10554
rect 1689 10486 1725 10520
rect 1689 10452 1690 10486
rect 1724 10452 1725 10486
rect 1689 10418 1725 10452
rect 1689 10384 1690 10418
rect 1724 10384 1725 10418
rect 1689 10350 1725 10384
rect 1689 10316 1690 10350
rect 1724 10316 1725 10350
rect 1689 10282 1725 10316
rect 1689 10248 1690 10282
rect 1724 10248 1725 10282
rect 1689 10214 1725 10248
rect 1689 10180 1690 10214
rect 1724 10180 1725 10214
rect 1689 10146 1725 10180
rect 1689 10112 1690 10146
rect 1724 10112 1725 10146
rect 1689 10078 1725 10112
rect 1689 10044 1690 10078
rect 1724 10044 1725 10078
rect 1689 10010 1725 10044
rect 1689 9976 1690 10010
rect 1724 9976 1725 10010
rect 1689 9942 1725 9976
rect 1689 9908 1690 9942
rect 1724 9908 1725 9942
rect 1689 9874 1725 9908
rect 1689 9840 1690 9874
rect 1724 9840 1725 9874
rect 1689 9806 1725 9840
rect 1689 9772 1690 9806
rect 1724 9772 1725 9806
rect 1689 9738 1725 9772
rect 8225 10544 8226 10578
rect 8260 10544 8261 10578
rect 8225 10510 8261 10544
rect 8225 10476 8226 10510
rect 8260 10476 8261 10510
rect 8225 10442 8261 10476
rect 8225 10408 8226 10442
rect 8260 10408 8261 10442
rect 8225 10374 8261 10408
rect 8225 10340 8226 10374
rect 8260 10340 8261 10374
rect 8225 10306 8261 10340
rect 8225 10272 8226 10306
rect 8260 10272 8261 10306
rect 8225 10238 8261 10272
rect 8225 10204 8226 10238
rect 8260 10204 8261 10238
rect 8225 10170 8261 10204
rect 8225 10136 8226 10170
rect 8260 10136 8261 10170
rect 8225 10102 8261 10136
rect 8225 10068 8226 10102
rect 8260 10068 8261 10102
rect 8225 10034 8261 10068
rect 8225 10000 8226 10034
rect 8260 10000 8261 10034
rect 8225 9966 8261 10000
rect 8225 9932 8226 9966
rect 8260 9932 8261 9966
rect 8225 9898 8261 9932
rect 8225 9864 8226 9898
rect 8260 9864 8261 9898
rect 8225 9830 8261 9864
rect 8225 9796 8226 9830
rect 8260 9796 8261 9830
rect 8225 9762 8261 9796
rect 1689 9704 1690 9738
rect 1724 9704 1725 9738
rect 8225 9728 8226 9762
rect 8260 9728 8261 9762
rect 1689 9670 1725 9704
rect 1689 9636 1690 9670
rect 1724 9636 1725 9670
rect 1689 9602 1725 9636
rect 1689 9568 1690 9602
rect 1724 9568 1725 9602
rect 1689 9534 1725 9568
rect 1689 9500 1690 9534
rect 1724 9500 1725 9534
rect 1689 9466 1725 9500
rect 1689 9432 1690 9466
rect 1724 9432 1725 9466
rect 1689 9398 1725 9432
rect 1689 9364 1690 9398
rect 1724 9364 1725 9398
rect 1689 9330 1725 9364
rect 1689 9296 1690 9330
rect 1724 9296 1725 9330
rect 1689 9262 1725 9296
rect 1689 9228 1690 9262
rect 1724 9228 1725 9262
rect 1689 9194 1725 9228
rect 1689 9160 1690 9194
rect 1724 9160 1725 9194
rect 1689 9126 1725 9160
rect 1689 9092 1690 9126
rect 1724 9092 1725 9126
rect 1689 9058 1725 9092
rect 1689 9024 1690 9058
rect 1724 9024 1725 9058
rect 1689 8990 1725 9024
rect 1689 8956 1690 8990
rect 1724 8956 1725 8990
rect 1689 8922 1725 8956
rect 1689 8888 1690 8922
rect 1724 8888 1725 8922
rect 8225 9694 8261 9728
rect 8225 9660 8226 9694
rect 8260 9660 8261 9694
rect 8225 9626 8261 9660
rect 8225 9592 8226 9626
rect 8260 9592 8261 9626
rect 8225 9558 8261 9592
rect 8225 9524 8226 9558
rect 8260 9524 8261 9558
rect 8225 9490 8261 9524
rect 8225 9456 8226 9490
rect 8260 9456 8261 9490
rect 8225 9422 8261 9456
rect 8225 9388 8226 9422
rect 8260 9388 8261 9422
rect 8225 9354 8261 9388
rect 8225 9320 8226 9354
rect 8260 9320 8261 9354
rect 8225 9286 8261 9320
rect 8225 9252 8226 9286
rect 8260 9252 8261 9286
rect 8225 9218 8261 9252
rect 8225 9184 8226 9218
rect 8260 9184 8261 9218
rect 8225 9150 8261 9184
rect 8225 9116 8226 9150
rect 8260 9116 8261 9150
rect 8225 9082 8261 9116
rect 8225 9048 8226 9082
rect 8260 9048 8261 9082
rect 8225 9014 8261 9048
rect 8225 8980 8226 9014
rect 8260 8980 8261 9014
rect 8225 8946 8261 8980
rect 8225 8912 8226 8946
rect 8260 8912 8261 8946
rect 1689 8778 1725 8888
rect 8225 8878 8261 8912
rect 8225 8844 8226 8878
rect 8260 8844 8261 8878
rect 8225 8810 8261 8844
rect 8225 8778 8226 8810
rect 1645 8777 8226 8778
rect 1645 8744 1723 8777
rect 1645 8710 1646 8744
rect 1680 8743 1723 8744
rect 1757 8743 1791 8777
rect 1825 8743 1859 8777
rect 1893 8743 1927 8777
rect 1961 8743 1995 8777
rect 2029 8743 2063 8777
rect 2097 8743 2131 8777
rect 2165 8743 2199 8777
rect 2233 8743 2267 8777
rect 2301 8743 2335 8777
rect 2369 8743 2403 8777
rect 2437 8743 2471 8777
rect 2505 8743 2539 8777
rect 2573 8743 2607 8777
rect 2641 8743 2675 8777
rect 2709 8743 2743 8777
rect 2777 8743 2811 8777
rect 2845 8743 2879 8777
rect 2913 8743 2947 8777
rect 2981 8743 3015 8777
rect 3049 8743 3083 8777
rect 3117 8743 3151 8777
rect 3185 8743 3219 8777
rect 3253 8743 3287 8777
rect 3321 8743 3355 8777
rect 3389 8743 3423 8777
rect 3457 8743 3491 8777
rect 3525 8743 3559 8777
rect 3593 8743 3627 8777
rect 3661 8743 3695 8777
rect 3729 8743 3763 8777
rect 3797 8743 3831 8777
rect 3865 8743 3899 8777
rect 3933 8743 3967 8777
rect 4001 8743 4035 8777
rect 4069 8743 4103 8777
rect 4137 8743 4171 8777
rect 4205 8743 4239 8777
rect 4273 8743 4307 8777
rect 4341 8743 4375 8777
rect 4409 8743 4443 8777
rect 4477 8743 4511 8777
rect 4545 8743 4579 8777
rect 4613 8743 4647 8777
rect 4681 8743 4715 8777
rect 4749 8743 4783 8777
rect 4817 8743 4851 8777
rect 4885 8743 4919 8777
rect 4953 8743 4987 8777
rect 5021 8743 5055 8777
rect 5089 8743 5123 8777
rect 5157 8743 5191 8777
rect 5225 8743 5259 8777
rect 5293 8743 5327 8777
rect 5361 8743 5395 8777
rect 5429 8743 5463 8777
rect 5497 8743 5531 8777
rect 5565 8743 5599 8777
rect 5633 8743 5667 8777
rect 5701 8743 5735 8777
rect 5769 8743 5803 8777
rect 5837 8743 5871 8777
rect 5905 8743 5939 8777
rect 5973 8743 6007 8777
rect 6041 8743 6075 8777
rect 6109 8743 6143 8777
rect 6177 8743 6211 8777
rect 6245 8743 6279 8777
rect 6313 8743 6347 8777
rect 6381 8743 6415 8777
rect 6449 8743 6483 8777
rect 6517 8743 6551 8777
rect 6585 8743 6619 8777
rect 6653 8743 6687 8777
rect 6721 8743 6755 8777
rect 6789 8743 6823 8777
rect 6857 8743 6891 8777
rect 6925 8743 6959 8777
rect 6993 8743 7027 8777
rect 7061 8743 7095 8777
rect 7129 8743 7163 8777
rect 7197 8743 7231 8777
rect 7265 8743 7299 8777
rect 7333 8743 7367 8777
rect 7401 8743 7435 8777
rect 7469 8743 7503 8777
rect 7537 8743 7571 8777
rect 7605 8743 7639 8777
rect 7673 8743 7707 8777
rect 7741 8743 7775 8777
rect 7809 8743 7843 8777
rect 7877 8743 7911 8777
rect 7945 8743 7979 8777
rect 8013 8743 8047 8777
rect 8081 8743 8115 8777
rect 8149 8776 8226 8777
rect 8260 8776 8261 8810
rect 8149 8743 8261 8776
rect 1680 8742 8261 8743
rect 1680 8710 1681 8742
rect 1645 8676 1681 8710
rect 1645 8642 1646 8676
rect 1680 8642 1681 8676
rect 1645 8608 1681 8642
rect 1645 8574 1646 8608
rect 1680 8574 1681 8608
rect 1645 8540 1681 8574
rect 1645 8506 1646 8540
rect 1680 8506 1681 8540
rect 1645 8472 1681 8506
rect 1645 8438 1646 8472
rect 1680 8438 1681 8472
rect 1645 8404 1681 8438
rect 1645 8370 1646 8404
rect 1680 8370 1681 8404
rect 1645 8336 1681 8370
rect 1645 8302 1646 8336
rect 1680 8302 1681 8336
rect 1645 8268 1681 8302
rect 1645 8234 1646 8268
rect 1680 8234 1681 8268
rect 1645 8200 1681 8234
rect 1645 8166 1646 8200
rect 1680 8166 1681 8200
rect 1645 8132 1681 8166
rect 1645 8098 1646 8132
rect 1680 8098 1681 8132
rect 1645 8064 1681 8098
rect 1645 8030 1646 8064
rect 1680 8030 1681 8064
rect 1645 7996 1681 8030
rect 1645 7962 1646 7996
rect 1680 7962 1681 7996
rect 1645 7928 1681 7962
rect 1645 7894 1646 7928
rect 1680 7894 1681 7928
rect 1645 7860 1681 7894
rect 1645 7826 1646 7860
rect 1680 7826 1681 7860
rect 1645 7792 1681 7826
rect 1645 7758 1646 7792
rect 1680 7758 1681 7792
rect 1645 7724 1681 7758
rect 1645 7690 1646 7724
rect 1680 7690 1681 7724
rect 1645 7656 1681 7690
rect 1645 7622 1646 7656
rect 1680 7622 1681 7656
rect 1645 7588 1681 7622
rect 1645 7554 1646 7588
rect 1680 7554 1681 7588
rect 1645 7511 1681 7554
rect 1645 7510 4139 7511
rect 1645 7476 1679 7510
rect 1713 7476 1747 7510
rect 1781 7476 1815 7510
rect 1849 7476 1883 7510
rect 1917 7476 1951 7510
rect 1985 7476 2019 7510
rect 2053 7476 2087 7510
rect 2121 7476 2155 7510
rect 2189 7476 2223 7510
rect 2257 7476 2291 7510
rect 2325 7476 2359 7510
rect 2393 7476 2427 7510
rect 2461 7476 2495 7510
rect 2529 7476 2563 7510
rect 2597 7476 2631 7510
rect 2665 7476 2699 7510
rect 2733 7476 2767 7510
rect 2801 7476 2835 7510
rect 2869 7476 2903 7510
rect 2937 7476 2971 7510
rect 3005 7476 3039 7510
rect 3073 7476 3107 7510
rect 3141 7476 3175 7510
rect 3209 7476 3243 7510
rect 3277 7476 3311 7510
rect 3345 7476 3379 7510
rect 3413 7476 3447 7510
rect 3481 7476 3515 7510
rect 3549 7476 3583 7510
rect 3617 7476 3651 7510
rect 3685 7476 3719 7510
rect 3753 7476 3787 7510
rect 3821 7476 3855 7510
rect 3889 7476 3923 7510
rect 3957 7476 3991 7510
rect 4025 7476 4059 7510
rect 4093 7476 4139 7510
rect 1645 7475 4139 7476
rect 1645 7110 3939 7111
rect 1645 7077 1763 7110
rect 1645 7043 1646 7077
rect 1680 7076 1763 7077
rect 1797 7076 1831 7110
rect 1865 7076 1899 7110
rect 1933 7076 1967 7110
rect 2001 7076 2035 7110
rect 2069 7076 2103 7110
rect 2137 7076 2171 7110
rect 2205 7076 2239 7110
rect 2273 7076 2307 7110
rect 2341 7076 2375 7110
rect 2409 7076 2443 7110
rect 2477 7076 2511 7110
rect 2545 7076 2579 7110
rect 2613 7076 2647 7110
rect 2681 7076 2715 7110
rect 2749 7076 2783 7110
rect 2817 7076 2851 7110
rect 2885 7076 2919 7110
rect 2953 7076 2987 7110
rect 3021 7076 3055 7110
rect 3089 7076 3123 7110
rect 3157 7076 3191 7110
rect 3225 7076 3259 7110
rect 3293 7076 3327 7110
rect 3361 7076 3395 7110
rect 3429 7076 3463 7110
rect 3497 7076 3531 7110
rect 3565 7076 3599 7110
rect 3633 7076 3667 7110
rect 3701 7076 3735 7110
rect 3769 7076 3803 7110
rect 3837 7076 3871 7110
rect 3905 7076 3939 7110
rect 1680 7075 3939 7076
rect 1680 7043 1681 7075
rect 1645 7009 1681 7043
rect 1645 6975 1646 7009
rect 1680 6975 1681 7009
rect 1645 6941 1681 6975
rect 3903 7035 3939 7075
rect 3903 7001 3904 7035
rect 3938 7001 3939 7035
rect 1645 6907 1646 6941
rect 1680 6907 1681 6941
rect 1645 6873 1681 6907
rect 1645 6839 1646 6873
rect 1680 6839 1681 6873
rect 1645 6805 1681 6839
rect 1645 6771 1646 6805
rect 1680 6771 1681 6805
rect 1645 6737 1681 6771
rect 1645 6703 1646 6737
rect 1680 6703 1681 6737
rect 1645 6669 1681 6703
rect 1645 6635 1646 6669
rect 1680 6635 1681 6669
rect 1645 6601 1681 6635
rect 1645 6567 1646 6601
rect 1680 6567 1681 6601
rect 1645 6533 1681 6567
rect 1645 6499 1646 6533
rect 1680 6499 1681 6533
rect 1645 6465 1681 6499
rect 1645 6431 1646 6465
rect 1680 6431 1681 6465
rect 1645 6397 1681 6431
rect 1645 6363 1646 6397
rect 1680 6363 1681 6397
rect 1645 6329 1681 6363
rect 1645 6295 1646 6329
rect 1680 6295 1681 6329
rect 1645 6261 1681 6295
rect 1645 6227 1646 6261
rect 1680 6227 1681 6261
rect 1645 6193 1681 6227
rect 1645 6159 1646 6193
rect 1680 6159 1681 6193
rect 1645 6125 1681 6159
rect 1645 6091 1646 6125
rect 1680 6091 1681 6125
rect 1645 6057 1681 6091
rect 1645 6023 1646 6057
rect 1680 6023 1681 6057
rect 1645 5989 1681 6023
rect 1645 5955 1646 5989
rect 1680 5955 1681 5989
rect 1645 5921 1681 5955
rect 1645 5887 1646 5921
rect 1680 5887 1681 5921
rect 3903 6967 3939 7001
rect 3903 6933 3904 6967
rect 3938 6933 3939 6967
rect 3903 6899 3939 6933
rect 3903 6865 3904 6899
rect 3938 6865 3939 6899
rect 3903 6831 3939 6865
rect 3903 6797 3904 6831
rect 3938 6797 3939 6831
rect 3903 6763 3939 6797
rect 3903 6729 3904 6763
rect 3938 6729 3939 6763
rect 3903 6695 3939 6729
rect 3903 6661 3904 6695
rect 3938 6661 3939 6695
rect 3903 6627 3939 6661
rect 3903 6593 3904 6627
rect 3938 6593 3939 6627
rect 3903 6559 3939 6593
rect 3903 6525 3904 6559
rect 3938 6525 3939 6559
rect 3903 6491 3939 6525
rect 3903 6457 3904 6491
rect 3938 6457 3939 6491
rect 3903 6423 3939 6457
rect 3903 6389 3904 6423
rect 3938 6389 3939 6423
rect 3903 6355 3939 6389
rect 3903 6321 3904 6355
rect 3938 6321 3939 6355
rect 3903 6287 3939 6321
rect 3903 6253 3904 6287
rect 3938 6253 3939 6287
rect 3903 6219 3939 6253
rect 3903 6185 3904 6219
rect 3938 6185 3939 6219
rect 3903 6151 3939 6185
rect 3903 6117 3904 6151
rect 3938 6117 3939 6151
rect 3903 6083 3939 6117
rect 3903 6049 3904 6083
rect 3938 6049 3939 6083
rect 3903 6015 3939 6049
rect 3903 5981 3904 6015
rect 3938 5981 3939 6015
rect 3903 5947 3939 5981
rect 3903 5913 3904 5947
rect 3938 5913 3939 5947
rect 1645 5853 1681 5887
rect 1645 5819 1646 5853
rect 1680 5819 1681 5853
rect 3903 5879 3939 5913
rect 1645 5785 1681 5819
rect 1645 5751 1646 5785
rect 1680 5751 1681 5785
rect 3903 5845 3904 5879
rect 3938 5845 3939 5879
rect 3903 5811 3939 5845
rect 3903 5777 3904 5811
rect 3938 5777 3939 5811
rect 1645 5717 1681 5751
rect 1645 5683 1646 5717
rect 1680 5683 1681 5717
rect 1645 5649 1681 5683
rect 1645 5615 1646 5649
rect 1680 5615 1681 5649
rect 1645 5581 1681 5615
rect 1645 5547 1646 5581
rect 1680 5547 1681 5581
rect 1645 5513 1681 5547
rect 1645 5479 1646 5513
rect 1680 5479 1681 5513
rect 1645 5445 1681 5479
rect 1645 5411 1646 5445
rect 1680 5411 1681 5445
rect 1645 5377 1681 5411
rect 1645 5343 1646 5377
rect 1680 5343 1681 5377
rect 1645 5309 1681 5343
rect 1645 5275 1646 5309
rect 1680 5275 1681 5309
rect 1645 5241 1681 5275
rect 1645 5207 1646 5241
rect 1680 5207 1681 5241
rect 1645 5173 1681 5207
rect 1645 5139 1646 5173
rect 1680 5139 1681 5173
rect 1645 5105 1681 5139
rect 1645 5071 1646 5105
rect 1680 5071 1681 5105
rect 1645 5037 1681 5071
rect 1645 5003 1646 5037
rect 1680 5003 1681 5037
rect 1645 4969 1681 5003
rect 1645 4935 1646 4969
rect 1680 4935 1681 4969
rect 1645 4901 1681 4935
rect 1645 4867 1646 4901
rect 1680 4867 1681 4901
rect 1645 4833 1681 4867
rect 1645 4799 1646 4833
rect 1680 4799 1681 4833
rect 1645 4765 1681 4799
rect 1645 4731 1646 4765
rect 1680 4731 1681 4765
rect 1645 4697 1681 4731
rect 3903 5743 3939 5777
rect 3903 5709 3904 5743
rect 3938 5709 3939 5743
rect 3903 5675 3939 5709
rect 3903 5641 3904 5675
rect 3938 5641 3939 5675
rect 3903 5607 3939 5641
rect 3903 5573 3904 5607
rect 3938 5573 3939 5607
rect 3903 5539 3939 5573
rect 3903 5505 3904 5539
rect 3938 5505 3939 5539
rect 3903 5471 3939 5505
rect 3903 5437 3904 5471
rect 3938 5437 3939 5471
rect 3903 5403 3939 5437
rect 3903 5369 3904 5403
rect 3938 5369 3939 5403
rect 3903 5335 3939 5369
rect 3903 5301 3904 5335
rect 3938 5301 3939 5335
rect 3903 5267 3939 5301
rect 3903 5233 3904 5267
rect 3938 5233 3939 5267
rect 3903 5199 3939 5233
rect 3903 5165 3904 5199
rect 3938 5165 3939 5199
rect 3903 5131 3939 5165
rect 3903 5097 3904 5131
rect 3938 5097 3939 5131
rect 3903 5063 3939 5097
rect 3903 5029 3904 5063
rect 3938 5029 3939 5063
rect 3903 4995 3939 5029
rect 3903 4961 3904 4995
rect 3938 4961 3939 4995
rect 3903 4927 3939 4961
rect 3903 4893 3904 4927
rect 3938 4893 3939 4927
rect 3903 4859 3939 4893
rect 3903 4825 3904 4859
rect 3938 4825 3939 4859
rect 3903 4791 3939 4825
rect 3903 4757 3904 4791
rect 3938 4757 3939 4791
rect 3903 4723 3939 4757
rect 1645 4663 1646 4697
rect 1680 4663 1681 4697
rect 1645 4629 1681 4663
rect 3903 4689 3904 4723
rect 3938 4689 3939 4723
rect 1645 4595 1646 4629
rect 1680 4595 1681 4629
rect 1645 4561 1681 4595
rect 3903 4655 3939 4689
rect 3903 4621 3904 4655
rect 3938 4621 3939 4655
rect 3903 4587 3939 4621
rect 1645 4527 1646 4561
rect 1680 4527 1681 4561
rect 1645 4493 1681 4527
rect 1645 4459 1646 4493
rect 1680 4459 1681 4493
rect 1645 4425 1681 4459
rect 1645 4391 1646 4425
rect 1680 4391 1681 4425
rect 1645 4357 1681 4391
rect 1645 4323 1646 4357
rect 1680 4323 1681 4357
rect 1645 4289 1681 4323
rect 1645 4255 1646 4289
rect 1680 4255 1681 4289
rect 1645 4221 1681 4255
rect 1645 4187 1646 4221
rect 1680 4187 1681 4221
rect 1645 4153 1681 4187
rect 1645 4119 1646 4153
rect 1680 4119 1681 4153
rect 1645 4085 1681 4119
rect 1645 4051 1646 4085
rect 1680 4051 1681 4085
rect 1645 4017 1681 4051
rect 1645 3983 1646 4017
rect 1680 3983 1681 4017
rect 1645 3949 1681 3983
rect 1645 3915 1646 3949
rect 1680 3915 1681 3949
rect 1645 3881 1681 3915
rect 1645 3847 1646 3881
rect 1680 3847 1681 3881
rect 1645 3813 1681 3847
rect 1645 3779 1646 3813
rect 1680 3779 1681 3813
rect 1645 3745 1681 3779
rect 1645 3711 1646 3745
rect 1680 3711 1681 3745
rect 1645 3677 1681 3711
rect 1645 3643 1646 3677
rect 1680 3643 1681 3677
rect 1645 3609 1681 3643
rect 1645 3575 1646 3609
rect 1680 3575 1681 3609
rect 1645 3541 1681 3575
rect 1645 3507 1646 3541
rect 1680 3507 1681 3541
rect 3903 4553 3904 4587
rect 3938 4553 3939 4587
rect 3903 4519 3939 4553
rect 3903 4485 3904 4519
rect 3938 4485 3939 4519
rect 3903 4451 3939 4485
rect 3903 4417 3904 4451
rect 3938 4417 3939 4451
rect 3903 4383 3939 4417
rect 3903 4349 3904 4383
rect 3938 4349 3939 4383
rect 3903 4315 3939 4349
rect 3903 4281 3904 4315
rect 3938 4281 3939 4315
rect 3903 4247 3939 4281
rect 3903 4213 3904 4247
rect 3938 4213 3939 4247
rect 3903 4179 3939 4213
rect 3903 4145 3904 4179
rect 3938 4145 3939 4179
rect 3903 4111 3939 4145
rect 3903 4077 3904 4111
rect 3938 4077 3939 4111
rect 3903 4043 3939 4077
rect 3903 4009 3904 4043
rect 3938 4009 3939 4043
rect 3903 3975 3939 4009
rect 3903 3941 3904 3975
rect 3938 3941 3939 3975
rect 3903 3907 3939 3941
rect 3903 3873 3904 3907
rect 3938 3873 3939 3907
rect 3903 3839 3939 3873
rect 3903 3805 3904 3839
rect 3938 3805 3939 3839
rect 3903 3771 3939 3805
rect 3903 3737 3904 3771
rect 3938 3737 3939 3771
rect 3903 3703 3939 3737
rect 3903 3669 3904 3703
rect 3938 3669 3939 3703
rect 3903 3635 3939 3669
rect 3903 3601 3904 3635
rect 3938 3601 3939 3635
rect 3903 3567 3939 3601
rect 3903 3533 3904 3567
rect 3938 3533 3939 3567
rect 1645 3473 1681 3507
rect 1645 3439 1646 3473
rect 1680 3439 1681 3473
rect 1645 3405 1681 3439
rect 1645 3371 1646 3405
rect 1680 3371 1681 3405
rect 1645 3337 1681 3371
rect 1645 3303 1646 3337
rect 1680 3303 1681 3337
rect 1645 3269 1681 3303
rect 1645 3235 1646 3269
rect 1680 3235 1681 3269
rect 1645 3201 1681 3235
rect 1645 3167 1646 3201
rect 1680 3167 1681 3201
rect 1645 3133 1681 3167
rect 1645 3099 1646 3133
rect 1680 3099 1681 3133
rect 1645 3065 1681 3099
rect 1645 3031 1646 3065
rect 1680 3031 1681 3065
rect 1645 2997 1681 3031
rect 1645 2963 1646 2997
rect 1680 2963 1681 2997
rect 1645 2929 1681 2963
rect 1645 2895 1646 2929
rect 1680 2895 1681 2929
rect 1645 2861 1681 2895
rect 1645 2827 1646 2861
rect 1680 2827 1681 2861
rect 1645 2793 1681 2827
rect 1645 2759 1646 2793
rect 1680 2759 1681 2793
rect 1645 2725 1681 2759
rect 1645 2691 1646 2725
rect 1680 2691 1681 2725
rect 1645 2657 1681 2691
rect 1645 2623 1646 2657
rect 1680 2623 1681 2657
rect 1645 2589 1681 2623
rect 1645 2555 1646 2589
rect 1680 2555 1681 2589
rect 1645 2521 1681 2555
rect 1645 2487 1646 2521
rect 1680 2487 1681 2521
rect 1645 2453 1681 2487
rect 1645 2419 1646 2453
rect 1680 2419 1681 2453
rect 1645 2293 1681 2419
rect 3903 3277 3939 3533
rect 3903 3243 3904 3277
rect 3938 3243 3939 3277
rect 3903 3209 3939 3243
rect 3903 3175 3904 3209
rect 3938 3175 3939 3209
rect 3903 3141 3939 3175
rect 3903 3107 3904 3141
rect 3938 3107 3939 3141
rect 3903 3073 3939 3107
rect 3903 3039 3904 3073
rect 3938 3039 3939 3073
rect 3903 3005 3939 3039
rect 3903 2971 3904 3005
rect 3938 2971 3939 3005
rect 3903 2937 3939 2971
rect 3903 2903 3904 2937
rect 3938 2903 3939 2937
rect 3903 2869 3939 2903
rect 3903 2835 3904 2869
rect 3938 2835 3939 2869
rect 3903 2801 3939 2835
rect 3903 2767 3904 2801
rect 3938 2767 3939 2801
rect 3903 2733 3939 2767
rect 3903 2699 3904 2733
rect 3938 2699 3939 2733
rect 3903 2665 3939 2699
rect 3903 2631 3904 2665
rect 3938 2631 3939 2665
rect 3903 2597 3939 2631
rect 3903 2563 3904 2597
rect 3938 2563 3939 2597
rect 3903 2529 3939 2563
rect 3903 2495 3904 2529
rect 3938 2495 3939 2529
rect 3903 2461 3939 2495
rect 3903 2427 3904 2461
rect 3938 2427 3939 2461
rect 3903 2393 3939 2427
rect 3903 2359 3904 2393
rect 3938 2359 3939 2393
rect 3903 2325 3939 2359
rect 3903 2293 3904 2325
rect 1645 2292 3904 2293
rect 1645 2258 1679 2292
rect 1713 2258 1747 2292
rect 1781 2258 1815 2292
rect 1849 2258 1883 2292
rect 1917 2258 1951 2292
rect 1985 2258 2019 2292
rect 2053 2258 2087 2292
rect 2121 2258 2155 2292
rect 2189 2258 2223 2292
rect 2257 2258 2291 2292
rect 2325 2258 2359 2292
rect 2393 2258 2427 2292
rect 2461 2258 2495 2292
rect 2529 2258 2563 2292
rect 2597 2258 2631 2292
rect 2665 2258 2699 2292
rect 2733 2258 2767 2292
rect 2801 2258 2835 2292
rect 2869 2258 2903 2292
rect 2937 2258 2971 2292
rect 3005 2258 3039 2292
rect 3073 2258 3107 2292
rect 3141 2258 3175 2292
rect 3209 2258 3243 2292
rect 3277 2258 3311 2292
rect 3345 2258 3379 2292
rect 3413 2258 3447 2292
rect 3481 2258 3515 2292
rect 3549 2258 3583 2292
rect 3617 2258 3651 2292
rect 3685 2258 3719 2292
rect 3753 2258 3787 2292
rect 3821 2291 3904 2292
rect 3938 2291 3939 2325
rect 3821 2258 3939 2291
rect 1645 2257 3939 2258
<< mvnsubdiff >>
rect 8 10912 8450 10913
rect 8 10878 42 10912
rect 76 10878 110 10912
rect 144 10878 178 10912
rect 212 10878 246 10912
rect 280 10878 314 10912
rect 348 10878 382 10912
rect 416 10878 450 10912
rect 484 10878 518 10912
rect 552 10878 586 10912
rect 620 10878 654 10912
rect 688 10878 722 10912
rect 756 10878 790 10912
rect 824 10878 858 10912
rect 892 10878 926 10912
rect 960 10878 994 10912
rect 1028 10878 1062 10912
rect 1096 10878 1130 10912
rect 1164 10878 1198 10912
rect 1232 10878 1266 10912
rect 1300 10878 1334 10912
rect 1368 10879 1582 10912
rect 1368 10878 1457 10879
rect 8 10877 1457 10878
rect 8 10789 44 10877
rect 8 10755 9 10789
rect 43 10755 44 10789
rect 8 10721 44 10755
rect 8 10687 9 10721
rect 43 10687 44 10721
rect 1456 10845 1457 10877
rect 1491 10878 1582 10879
rect 1616 10878 1650 10912
rect 1684 10878 1718 10912
rect 1752 10878 1786 10912
rect 1820 10878 1854 10912
rect 1888 10878 1922 10912
rect 1956 10878 1990 10912
rect 2024 10878 2058 10912
rect 2092 10878 2126 10912
rect 2160 10878 2194 10912
rect 2228 10878 2262 10912
rect 2296 10878 2330 10912
rect 2364 10878 2398 10912
rect 2432 10878 2466 10912
rect 2500 10878 2534 10912
rect 2568 10878 2602 10912
rect 2636 10878 2670 10912
rect 2704 10878 2738 10912
rect 2772 10878 2806 10912
rect 2840 10878 2874 10912
rect 2908 10878 2942 10912
rect 2976 10878 3010 10912
rect 3044 10878 3078 10912
rect 3112 10878 3146 10912
rect 3180 10878 3214 10912
rect 3248 10878 3282 10912
rect 3316 10878 3350 10912
rect 3384 10878 3418 10912
rect 3452 10878 3486 10912
rect 3520 10878 3554 10912
rect 3588 10878 3622 10912
rect 3656 10878 3690 10912
rect 3724 10878 3758 10912
rect 3792 10878 3826 10912
rect 3860 10878 3894 10912
rect 3928 10878 3962 10912
rect 3996 10878 4030 10912
rect 4064 10878 4098 10912
rect 4132 10878 4166 10912
rect 4200 10878 4234 10912
rect 4268 10878 4302 10912
rect 4336 10878 4370 10912
rect 4404 10878 4438 10912
rect 4472 10878 4506 10912
rect 4540 10878 4574 10912
rect 4608 10878 4642 10912
rect 4676 10878 4710 10912
rect 4744 10878 4778 10912
rect 4812 10878 4846 10912
rect 4880 10878 4914 10912
rect 4948 10878 4982 10912
rect 5016 10878 5050 10912
rect 5084 10878 5118 10912
rect 5152 10878 5186 10912
rect 5220 10878 5254 10912
rect 5288 10878 5322 10912
rect 5356 10878 5390 10912
rect 5424 10878 5458 10912
rect 5492 10878 5526 10912
rect 5560 10878 5594 10912
rect 5628 10878 5662 10912
rect 5696 10878 5730 10912
rect 5764 10878 5798 10912
rect 5832 10878 5866 10912
rect 5900 10878 5934 10912
rect 5968 10878 6002 10912
rect 6036 10878 6070 10912
rect 6104 10878 6138 10912
rect 6172 10878 6206 10912
rect 6240 10878 6274 10912
rect 6308 10878 6342 10912
rect 6376 10878 6410 10912
rect 6444 10878 6478 10912
rect 6512 10878 6546 10912
rect 6580 10878 6614 10912
rect 6648 10878 6682 10912
rect 6716 10878 6750 10912
rect 6784 10878 6818 10912
rect 6852 10878 6886 10912
rect 6920 10878 6954 10912
rect 6988 10878 7022 10912
rect 7056 10878 7090 10912
rect 7124 10878 7158 10912
rect 7192 10878 7226 10912
rect 7260 10878 7294 10912
rect 7328 10878 7362 10912
rect 7396 10878 7430 10912
rect 7464 10878 7498 10912
rect 7532 10878 7566 10912
rect 7600 10878 7634 10912
rect 7668 10878 7702 10912
rect 7736 10878 7770 10912
rect 7804 10878 7838 10912
rect 7872 10878 7906 10912
rect 7940 10878 7974 10912
rect 8008 10878 8042 10912
rect 8076 10878 8110 10912
rect 8144 10878 8178 10912
rect 8212 10878 8246 10912
rect 8280 10878 8314 10912
rect 8348 10878 8382 10912
rect 8416 10878 8450 10912
rect 1491 10877 8450 10878
rect 1491 10845 1492 10877
rect 1456 10811 1492 10845
rect 1456 10777 1457 10811
rect 1491 10777 1492 10811
rect 1456 10743 1492 10777
rect 1456 10709 1457 10743
rect 1491 10709 1492 10743
rect 8414 10819 8450 10877
rect 8414 10785 8415 10819
rect 8449 10785 8450 10819
rect 8414 10751 8450 10785
rect 8 10653 44 10687
rect 8 10619 9 10653
rect 43 10619 44 10653
rect 8 10585 44 10619
rect 8 10551 9 10585
rect 43 10551 44 10585
rect 8 10517 44 10551
rect 8 10483 9 10517
rect 43 10483 44 10517
rect 8 10449 44 10483
rect 8 10415 9 10449
rect 43 10415 44 10449
rect 8 10381 44 10415
rect 8 10347 9 10381
rect 43 10347 44 10381
rect 8 10313 44 10347
rect 8 10279 9 10313
rect 43 10279 44 10313
rect 8 10245 44 10279
rect 8 10211 9 10245
rect 43 10211 44 10245
rect 8 10177 44 10211
rect 8 10143 9 10177
rect 43 10143 44 10177
rect 8 10109 44 10143
rect 8 10075 9 10109
rect 43 10075 44 10109
rect 8 10041 44 10075
rect 8 10007 9 10041
rect 43 10007 44 10041
rect 8 9973 44 10007
rect 8 9939 9 9973
rect 43 9939 44 9973
rect 8 9905 44 9939
rect 8 9871 9 9905
rect 43 9871 44 9905
rect 8 9837 44 9871
rect 8 9803 9 9837
rect 43 9803 44 9837
rect 8 9769 44 9803
rect 8 9735 9 9769
rect 43 9735 44 9769
rect 8 9701 44 9735
rect 8 9667 9 9701
rect 43 9667 44 9701
rect 8 9633 44 9667
rect 8 9599 9 9633
rect 43 9599 44 9633
rect 8 9565 44 9599
rect 8 9531 9 9565
rect 43 9531 44 9565
rect 8 9497 44 9531
rect 8 9463 9 9497
rect 43 9463 44 9497
rect 8 9429 44 9463
rect 8 9395 9 9429
rect 43 9395 44 9429
rect 8 9361 44 9395
rect 8 9327 9 9361
rect 43 9327 44 9361
rect 8 9293 44 9327
rect 8 9259 9 9293
rect 43 9259 44 9293
rect 8 9225 44 9259
rect 8 9191 9 9225
rect 43 9191 44 9225
rect 8 9157 44 9191
rect 8 9123 9 9157
rect 43 9123 44 9157
rect 8 9089 44 9123
rect 8 9055 9 9089
rect 43 9055 44 9089
rect 8 9021 44 9055
rect 8 8987 9 9021
rect 43 8987 44 9021
rect 8 8953 44 8987
rect 8 8919 9 8953
rect 43 8919 44 8953
rect 8 8885 44 8919
rect 8 8851 9 8885
rect 43 8851 44 8885
rect 8 8817 44 8851
rect 8 8783 9 8817
rect 43 8783 44 8817
rect 8 8749 44 8783
rect 8 8715 9 8749
rect 43 8715 44 8749
rect 8 8681 44 8715
rect 8 8647 9 8681
rect 43 8647 44 8681
rect 8 8613 44 8647
rect 8 8579 9 8613
rect 43 8579 44 8613
rect 8 8545 44 8579
rect 8 8511 9 8545
rect 43 8511 44 8545
rect 8 8477 44 8511
rect 8 8443 9 8477
rect 43 8443 44 8477
rect 8 8409 44 8443
rect 8 8375 9 8409
rect 43 8375 44 8409
rect 8 8341 44 8375
rect 8 8307 9 8341
rect 43 8307 44 8341
rect 8 8273 44 8307
rect 8 8239 9 8273
rect 43 8239 44 8273
rect 8 8205 44 8239
rect 8 8171 9 8205
rect 43 8171 44 8205
rect 8 8137 44 8171
rect 8 8103 9 8137
rect 43 8103 44 8137
rect 8 8069 44 8103
rect 8 8035 9 8069
rect 43 8035 44 8069
rect 8 8001 44 8035
rect 8 7967 9 8001
rect 43 7967 44 8001
rect 8 7933 44 7967
rect 8 7899 9 7933
rect 43 7899 44 7933
rect 8 7865 44 7899
rect 8 7831 9 7865
rect 43 7831 44 7865
rect 8 7797 44 7831
rect 8 7763 9 7797
rect 43 7763 44 7797
rect 8 7729 44 7763
rect 8 7695 9 7729
rect 43 7695 44 7729
rect 8 7661 44 7695
rect 8 7627 9 7661
rect 43 7627 44 7661
rect 8 7593 44 7627
rect 8 7559 9 7593
rect 43 7559 44 7593
rect 8 7525 44 7559
rect 8 7491 9 7525
rect 43 7491 44 7525
rect 8 7457 44 7491
rect 8 7423 9 7457
rect 43 7423 44 7457
rect 8 7389 44 7423
rect 8 7355 9 7389
rect 43 7355 44 7389
rect 8 7321 44 7355
rect 8 7287 9 7321
rect 43 7287 44 7321
rect 8 7253 44 7287
rect 8 7219 9 7253
rect 43 7219 44 7253
rect 8 7185 44 7219
rect 8 7151 9 7185
rect 43 7151 44 7185
rect 8 7117 44 7151
rect 8 7083 9 7117
rect 43 7083 44 7117
rect 8 7049 44 7083
rect 8 7015 9 7049
rect 43 7015 44 7049
rect 8 6981 44 7015
rect 8 6947 9 6981
rect 43 6947 44 6981
rect 8 6913 44 6947
rect 8 6879 9 6913
rect 43 6879 44 6913
rect 8 6845 44 6879
rect 8 6811 9 6845
rect 43 6811 44 6845
rect 8 6777 44 6811
rect 8 6743 9 6777
rect 43 6743 44 6777
rect 8 6709 44 6743
rect 8 6675 9 6709
rect 43 6675 44 6709
rect 8 6641 44 6675
rect 8 6607 9 6641
rect 43 6607 44 6641
rect 8 6573 44 6607
rect 8 6539 9 6573
rect 43 6539 44 6573
rect 8 6505 44 6539
rect 8 6471 9 6505
rect 43 6471 44 6505
rect 8 6437 44 6471
rect 8 6403 9 6437
rect 43 6403 44 6437
rect 8 6369 44 6403
rect 8 6335 9 6369
rect 43 6335 44 6369
rect 8 6301 44 6335
rect 8 6267 9 6301
rect 43 6267 44 6301
rect 8 6233 44 6267
rect 8 6199 9 6233
rect 43 6199 44 6233
rect 8 6165 44 6199
rect 8 6131 9 6165
rect 43 6131 44 6165
rect 8 6097 44 6131
rect 8 6063 9 6097
rect 43 6063 44 6097
rect 8 6029 44 6063
rect 8 5995 9 6029
rect 43 5995 44 6029
rect 8 5961 44 5995
rect 8 5927 9 5961
rect 43 5927 44 5961
rect 8 5893 44 5927
rect 8 5859 9 5893
rect 43 5859 44 5893
rect 8 5825 44 5859
rect 8 5791 9 5825
rect 43 5791 44 5825
rect 8 5757 44 5791
rect 8 5723 9 5757
rect 43 5723 44 5757
rect 8 5689 44 5723
rect 8 5655 9 5689
rect 43 5655 44 5689
rect 8 5621 44 5655
rect 8 5587 9 5621
rect 43 5587 44 5621
rect 8 5553 44 5587
rect 8 5519 9 5553
rect 43 5519 44 5553
rect 8 5485 44 5519
rect 8 5451 9 5485
rect 43 5451 44 5485
rect 8 5417 44 5451
rect 8 5383 9 5417
rect 43 5383 44 5417
rect 8 5349 44 5383
rect 8 5315 9 5349
rect 43 5315 44 5349
rect 8 5281 44 5315
rect 8 5247 9 5281
rect 43 5247 44 5281
rect 8 5213 44 5247
rect 8 5179 9 5213
rect 43 5179 44 5213
rect 8 5145 44 5179
rect 8 5111 9 5145
rect 43 5111 44 5145
rect 8 5077 44 5111
rect 8 5043 9 5077
rect 43 5043 44 5077
rect 8 5009 44 5043
rect 8 4975 9 5009
rect 43 4975 44 5009
rect 8 4941 44 4975
rect 8 4907 9 4941
rect 43 4907 44 4941
rect 8 4873 44 4907
rect 8 4839 9 4873
rect 43 4839 44 4873
rect 8 4805 44 4839
rect 8 4771 9 4805
rect 43 4771 44 4805
rect 8 4737 44 4771
rect 8 4703 9 4737
rect 43 4703 44 4737
rect 8 4669 44 4703
rect 8 4635 9 4669
rect 43 4635 44 4669
rect 8 4601 44 4635
rect 8 4567 9 4601
rect 43 4567 44 4601
rect 8 4533 44 4567
rect 8 4499 9 4533
rect 43 4499 44 4533
rect 8 4465 44 4499
rect 8 4431 9 4465
rect 43 4431 44 4465
rect 8 4397 44 4431
rect 8 4363 9 4397
rect 43 4363 44 4397
rect 8 4329 44 4363
rect 8 4295 9 4329
rect 43 4295 44 4329
rect 8 4261 44 4295
rect 8 4227 9 4261
rect 43 4227 44 4261
rect 8 4193 44 4227
rect 8 4159 9 4193
rect 43 4159 44 4193
rect 8 4125 44 4159
rect 8 4091 9 4125
rect 43 4091 44 4125
rect 8 4057 44 4091
rect 8 4023 9 4057
rect 43 4023 44 4057
rect 8 3989 44 4023
rect 8 3955 9 3989
rect 43 3955 44 3989
rect 8 3921 44 3955
rect 8 3887 9 3921
rect 43 3887 44 3921
rect 8 3853 44 3887
rect 8 3819 9 3853
rect 43 3819 44 3853
rect 8 3785 44 3819
rect 8 3751 9 3785
rect 43 3751 44 3785
rect 8 3717 44 3751
rect 8 3683 9 3717
rect 43 3683 44 3717
rect 8 3649 44 3683
rect 8 3615 9 3649
rect 43 3615 44 3649
rect 8 3581 44 3615
rect 8 3547 9 3581
rect 43 3547 44 3581
rect 8 3513 44 3547
rect 8 3479 9 3513
rect 43 3479 44 3513
rect 8 3445 44 3479
rect 8 3411 9 3445
rect 43 3411 44 3445
rect 8 3377 44 3411
rect 8 3343 9 3377
rect 43 3343 44 3377
rect 8 3309 44 3343
rect 8 3275 9 3309
rect 43 3275 44 3309
rect 8 3241 44 3275
rect 8 3207 9 3241
rect 43 3207 44 3241
rect 8 3173 44 3207
rect 8 3139 9 3173
rect 43 3139 44 3173
rect 8 3105 44 3139
rect 8 3071 9 3105
rect 43 3071 44 3105
rect 8 3037 44 3071
rect 8 3003 9 3037
rect 43 3003 44 3037
rect 8 2969 44 3003
rect 8 2935 9 2969
rect 43 2935 44 2969
rect 8 2901 44 2935
rect 8 2867 9 2901
rect 43 2867 44 2901
rect 8 2833 44 2867
rect 8 2799 9 2833
rect 43 2799 44 2833
rect 8 2765 44 2799
rect 8 2731 9 2765
rect 43 2731 44 2765
rect 8 2697 44 2731
rect 8 2663 9 2697
rect 43 2663 44 2697
rect 8 2629 44 2663
rect 8 2595 9 2629
rect 43 2595 44 2629
rect 8 2561 44 2595
rect 8 2527 9 2561
rect 43 2527 44 2561
rect 8 2493 44 2527
rect 8 2459 9 2493
rect 43 2459 44 2493
rect 8 2425 44 2459
rect 8 2391 9 2425
rect 43 2391 44 2425
rect 8 2357 44 2391
rect 8 2323 9 2357
rect 43 2323 44 2357
rect 8 2289 44 2323
rect 8 2255 9 2289
rect 43 2255 44 2289
rect 8 2221 44 2255
rect 8 2187 9 2221
rect 43 2187 44 2221
rect 8 2153 44 2187
rect 8 2119 9 2153
rect 43 2119 44 2153
rect 8 2085 44 2119
rect 8 2051 9 2085
rect 43 2051 44 2085
rect 8 2017 44 2051
rect 8 1983 9 2017
rect 43 1983 44 2017
rect 8 1949 44 1983
rect 8 1915 9 1949
rect 43 1915 44 1949
rect 8 1881 44 1915
rect 8 1847 9 1881
rect 43 1847 44 1881
rect 8 1813 44 1847
rect 8 1779 9 1813
rect 43 1779 44 1813
rect 8 1745 44 1779
rect 8 1711 9 1745
rect 43 1711 44 1745
rect 8 1677 44 1711
rect 8 1643 9 1677
rect 43 1643 44 1677
rect 8 1609 44 1643
rect 8 1575 9 1609
rect 43 1575 44 1609
rect 8 1541 44 1575
rect 8 1507 9 1541
rect 43 1507 44 1541
rect 8 1473 44 1507
rect 8 1439 9 1473
rect 43 1439 44 1473
rect 8 1405 44 1439
rect 8 1371 9 1405
rect 43 1371 44 1405
rect 8 1337 44 1371
rect 8 1303 9 1337
rect 43 1303 44 1337
rect 8 1269 44 1303
rect 8 1235 9 1269
rect 43 1235 44 1269
rect 8 1201 44 1235
rect 8 1167 9 1201
rect 43 1167 44 1201
rect 8 1133 44 1167
rect 8 1099 9 1133
rect 43 1099 44 1133
rect 8 1065 44 1099
rect 8 1031 9 1065
rect 43 1031 44 1065
rect 8 997 44 1031
rect 8 963 9 997
rect 43 963 44 997
rect 8 929 44 963
rect 8 895 9 929
rect 43 895 44 929
rect 8 861 44 895
rect 8 827 9 861
rect 43 827 44 861
rect 8 793 44 827
rect 8 759 9 793
rect 43 759 44 793
rect 8 725 44 759
rect 8 691 9 725
rect 43 691 44 725
rect 8 657 44 691
rect 8 623 9 657
rect 43 623 44 657
rect 8 589 44 623
rect 8 555 9 589
rect 43 555 44 589
rect 8 447 44 555
rect 1456 10675 1492 10709
rect 1456 10641 1457 10675
rect 1491 10641 1492 10675
rect 1456 10607 1492 10641
rect 1456 10573 1457 10607
rect 1491 10573 1492 10607
rect 1456 10539 1492 10573
rect 1456 10505 1457 10539
rect 1491 10505 1492 10539
rect 1456 10471 1492 10505
rect 1456 10437 1457 10471
rect 1491 10437 1492 10471
rect 1456 10403 1492 10437
rect 1456 10369 1457 10403
rect 1491 10369 1492 10403
rect 1456 10335 1492 10369
rect 1456 10301 1457 10335
rect 1491 10301 1492 10335
rect 1456 10267 1492 10301
rect 1456 10233 1457 10267
rect 1491 10233 1492 10267
rect 1456 10199 1492 10233
rect 1456 10165 1457 10199
rect 1491 10165 1492 10199
rect 1456 10131 1492 10165
rect 1456 10097 1457 10131
rect 1491 10097 1492 10131
rect 1456 10063 1492 10097
rect 1456 10029 1457 10063
rect 1491 10029 1492 10063
rect 1456 9995 1492 10029
rect 1456 9961 1457 9995
rect 1491 9961 1492 9995
rect 1456 9927 1492 9961
rect 1456 9893 1457 9927
rect 1491 9893 1492 9927
rect 1456 9859 1492 9893
rect 1456 9825 1457 9859
rect 1491 9825 1492 9859
rect 1456 9791 1492 9825
rect 1456 9757 1457 9791
rect 1491 9757 1492 9791
rect 1456 9723 1492 9757
rect 1456 9689 1457 9723
rect 1491 9689 1492 9723
rect 1456 9655 1492 9689
rect 1456 9621 1457 9655
rect 1491 9621 1492 9655
rect 1456 9587 1492 9621
rect 1456 9553 1457 9587
rect 1491 9553 1492 9587
rect 1456 9519 1492 9553
rect 1456 9485 1457 9519
rect 1491 9485 1492 9519
rect 1456 9451 1492 9485
rect 1456 9417 1457 9451
rect 1491 9417 1492 9451
rect 1456 9383 1492 9417
rect 1456 9349 1457 9383
rect 1491 9349 1492 9383
rect 1456 9315 1492 9349
rect 1456 9281 1457 9315
rect 1491 9281 1492 9315
rect 1456 9247 1492 9281
rect 1456 9213 1457 9247
rect 1491 9213 1492 9247
rect 1456 9179 1492 9213
rect 1456 9145 1457 9179
rect 1491 9145 1492 9179
rect 1456 9111 1492 9145
rect 1456 9077 1457 9111
rect 1491 9077 1492 9111
rect 1456 9043 1492 9077
rect 1456 9009 1457 9043
rect 1491 9009 1492 9043
rect 1456 8975 1492 9009
rect 1456 8941 1457 8975
rect 1491 8941 1492 8975
rect 1456 8907 1492 8941
rect 1456 8873 1457 8907
rect 1491 8873 1492 8907
rect 1456 8839 1492 8873
rect 1456 8805 1457 8839
rect 1491 8805 1492 8839
rect 1456 8771 1492 8805
rect 1456 8737 1457 8771
rect 1491 8737 1492 8771
rect 1456 8703 1492 8737
rect 1456 8669 1457 8703
rect 1491 8669 1492 8703
rect 1456 8635 1492 8669
rect 1456 8601 1457 8635
rect 1491 8601 1492 8635
rect 1456 8567 1492 8601
rect 1456 8533 1457 8567
rect 1491 8533 1492 8567
rect 1456 8499 1492 8533
rect 1456 8465 1457 8499
rect 1491 8465 1492 8499
rect 1456 8431 1492 8465
rect 1456 8397 1457 8431
rect 1491 8397 1492 8431
rect 1456 8363 1492 8397
rect 1456 8329 1457 8363
rect 1491 8329 1492 8363
rect 1456 8295 1492 8329
rect 1456 8261 1457 8295
rect 1491 8261 1492 8295
rect 1456 8227 1492 8261
rect 1456 8193 1457 8227
rect 1491 8193 1492 8227
rect 1456 8159 1492 8193
rect 1456 8125 1457 8159
rect 1491 8125 1492 8159
rect 1456 8091 1492 8125
rect 1456 8057 1457 8091
rect 1491 8057 1492 8091
rect 1456 8023 1492 8057
rect 1456 7989 1457 8023
rect 1491 7989 1492 8023
rect 1456 7955 1492 7989
rect 1456 7921 1457 7955
rect 1491 7921 1492 7955
rect 1456 7887 1492 7921
rect 1456 7853 1457 7887
rect 1491 7853 1492 7887
rect 1456 7819 1492 7853
rect 1456 7785 1457 7819
rect 1491 7785 1492 7819
rect 1456 7751 1492 7785
rect 1456 7717 1457 7751
rect 1491 7717 1492 7751
rect 1456 7683 1492 7717
rect 1456 7649 1457 7683
rect 1491 7649 1492 7683
rect 1456 7615 1492 7649
rect 1456 7581 1457 7615
rect 1491 7581 1492 7615
rect 1456 7547 1492 7581
rect 1456 7513 1457 7547
rect 1491 7513 1492 7547
rect 1456 7479 1492 7513
rect 1456 7445 1457 7479
rect 1491 7445 1492 7479
rect 8414 10717 8415 10751
rect 8449 10717 8450 10751
rect 8414 10683 8450 10717
rect 8414 10649 8415 10683
rect 8449 10649 8450 10683
rect 8414 10615 8450 10649
rect 8414 10581 8415 10615
rect 8449 10581 8450 10615
rect 8414 10547 8450 10581
rect 8414 10513 8415 10547
rect 8449 10513 8450 10547
rect 8414 10479 8450 10513
rect 8414 10445 8415 10479
rect 8449 10445 8450 10479
rect 8414 10411 8450 10445
rect 8414 10377 8415 10411
rect 8449 10377 8450 10411
rect 8414 10343 8450 10377
rect 8414 10309 8415 10343
rect 8449 10309 8450 10343
rect 8414 10275 8450 10309
rect 8414 10241 8415 10275
rect 8449 10241 8450 10275
rect 8414 10207 8450 10241
rect 8414 10173 8415 10207
rect 8449 10173 8450 10207
rect 8414 10139 8450 10173
rect 8414 10105 8415 10139
rect 8449 10105 8450 10139
rect 8414 10071 8450 10105
rect 8414 10037 8415 10071
rect 8449 10037 8450 10071
rect 8414 10003 8450 10037
rect 8414 9969 8415 10003
rect 8449 9969 8450 10003
rect 8414 9935 8450 9969
rect 8414 9901 8415 9935
rect 8449 9901 8450 9935
rect 8414 9867 8450 9901
rect 8414 9833 8415 9867
rect 8449 9833 8450 9867
rect 8414 9799 8450 9833
rect 8414 9765 8415 9799
rect 8449 9765 8450 9799
rect 8414 9731 8450 9765
rect 8414 9697 8415 9731
rect 8449 9697 8450 9731
rect 8414 9663 8450 9697
rect 8414 9629 8415 9663
rect 8449 9629 8450 9663
rect 8414 9595 8450 9629
rect 8414 9561 8415 9595
rect 8449 9561 8450 9595
rect 8414 9527 8450 9561
rect 8414 9493 8415 9527
rect 8449 9493 8450 9527
rect 8414 9459 8450 9493
rect 8414 9425 8415 9459
rect 8449 9425 8450 9459
rect 8414 9391 8450 9425
rect 8414 9357 8415 9391
rect 8449 9357 8450 9391
rect 8414 9323 8450 9357
rect 8414 9289 8415 9323
rect 8449 9289 8450 9323
rect 8414 9255 8450 9289
rect 8414 9221 8415 9255
rect 8449 9221 8450 9255
rect 8414 9187 8450 9221
rect 8414 9153 8415 9187
rect 8449 9153 8450 9187
rect 8414 9119 8450 9153
rect 8414 9085 8415 9119
rect 8449 9085 8450 9119
rect 8414 9051 8450 9085
rect 8414 9017 8415 9051
rect 8449 9017 8450 9051
rect 8414 8983 8450 9017
rect 8414 8949 8415 8983
rect 8449 8949 8450 8983
rect 8414 8915 8450 8949
rect 8414 8881 8415 8915
rect 8449 8881 8450 8915
rect 8414 8847 8450 8881
rect 8414 8813 8415 8847
rect 8449 8813 8450 8847
rect 8414 8779 8450 8813
rect 8414 8745 8415 8779
rect 8449 8745 8450 8779
rect 8414 8677 8450 8745
rect 8414 8643 8415 8677
rect 8449 8643 8450 8677
rect 8414 8553 8450 8643
rect 1456 7322 1492 7445
rect 1456 7321 4128 7322
rect 1456 7287 1490 7321
rect 1524 7287 1558 7321
rect 1592 7287 1626 7321
rect 1660 7287 1694 7321
rect 1728 7287 1762 7321
rect 1796 7287 1830 7321
rect 1864 7287 1898 7321
rect 1932 7287 1966 7321
rect 2000 7287 2034 7321
rect 2068 7287 2102 7321
rect 2136 7287 2170 7321
rect 2204 7287 2238 7321
rect 2272 7287 2306 7321
rect 2340 7287 2374 7321
rect 2408 7287 2442 7321
rect 2476 7287 2510 7321
rect 2544 7287 2578 7321
rect 2612 7287 2646 7321
rect 2680 7287 2714 7321
rect 2748 7287 2782 7321
rect 2816 7287 2850 7321
rect 2884 7287 2918 7321
rect 2952 7287 2986 7321
rect 3020 7287 3054 7321
rect 3088 7287 3122 7321
rect 3156 7287 3190 7321
rect 3224 7287 3258 7321
rect 3292 7287 3326 7321
rect 3360 7287 3394 7321
rect 3428 7287 3462 7321
rect 3496 7287 3530 7321
rect 3564 7287 3598 7321
rect 3632 7287 3666 7321
rect 3700 7287 3734 7321
rect 3768 7287 3802 7321
rect 3836 7287 3870 7321
rect 3904 7287 3938 7321
rect 3972 7287 4006 7321
rect 4040 7287 4128 7321
rect 1456 7286 4128 7287
rect 1456 7252 1492 7286
rect 1456 7218 1457 7252
rect 1491 7218 1492 7252
rect 1456 7184 1492 7218
rect 1456 7150 1457 7184
rect 1491 7150 1492 7184
rect 1456 7116 1492 7150
rect 1456 7082 1457 7116
rect 1491 7082 1492 7116
rect 4092 7226 4128 7286
rect 4092 7192 4093 7226
rect 4127 7192 4128 7226
rect 4092 7158 4128 7192
rect 4092 7124 4093 7158
rect 4127 7124 4128 7158
rect 1456 7048 1492 7082
rect 1456 7014 1457 7048
rect 1491 7014 1492 7048
rect 1456 6980 1492 7014
rect 1456 6946 1457 6980
rect 1491 6946 1492 6980
rect 1456 6912 1492 6946
rect 1456 6878 1457 6912
rect 1491 6878 1492 6912
rect 1456 6844 1492 6878
rect 1456 6810 1457 6844
rect 1491 6810 1492 6844
rect 1456 6776 1492 6810
rect 1456 6742 1457 6776
rect 1491 6742 1492 6776
rect 1456 6708 1492 6742
rect 1456 6674 1457 6708
rect 1491 6674 1492 6708
rect 1456 6640 1492 6674
rect 1456 6606 1457 6640
rect 1491 6606 1492 6640
rect 1456 6572 1492 6606
rect 1456 6538 1457 6572
rect 1491 6538 1492 6572
rect 1456 6504 1492 6538
rect 1456 6470 1457 6504
rect 1491 6470 1492 6504
rect 1456 6436 1492 6470
rect 1456 6402 1457 6436
rect 1491 6402 1492 6436
rect 1456 6368 1492 6402
rect 1456 6334 1457 6368
rect 1491 6334 1492 6368
rect 1456 6300 1492 6334
rect 1456 6266 1457 6300
rect 1491 6266 1492 6300
rect 1456 6232 1492 6266
rect 1456 6198 1457 6232
rect 1491 6198 1492 6232
rect 1456 6164 1492 6198
rect 1456 6130 1457 6164
rect 1491 6130 1492 6164
rect 1456 6096 1492 6130
rect 1456 6062 1457 6096
rect 1491 6062 1492 6096
rect 1456 6028 1492 6062
rect 1456 5994 1457 6028
rect 1491 5994 1492 6028
rect 1456 5960 1492 5994
rect 1456 5926 1457 5960
rect 1491 5926 1492 5960
rect 1456 5892 1492 5926
rect 1456 5858 1457 5892
rect 1491 5858 1492 5892
rect 1456 5824 1492 5858
rect 1456 5790 1457 5824
rect 1491 5790 1492 5824
rect 1456 5756 1492 5790
rect 1456 5722 1457 5756
rect 1491 5722 1492 5756
rect 1456 5688 1492 5722
rect 1456 5654 1457 5688
rect 1491 5654 1492 5688
rect 1456 5620 1492 5654
rect 1456 5586 1457 5620
rect 1491 5586 1492 5620
rect 1456 5552 1492 5586
rect 1456 5518 1457 5552
rect 1491 5518 1492 5552
rect 1456 5484 1492 5518
rect 1456 5450 1457 5484
rect 1491 5450 1492 5484
rect 1456 5416 1492 5450
rect 1456 5382 1457 5416
rect 1491 5382 1492 5416
rect 1456 5348 1492 5382
rect 1456 5314 1457 5348
rect 1491 5314 1492 5348
rect 1456 5280 1492 5314
rect 1456 5246 1457 5280
rect 1491 5246 1492 5280
rect 1456 5212 1492 5246
rect 1456 5178 1457 5212
rect 1491 5178 1492 5212
rect 1456 5144 1492 5178
rect 1456 5110 1457 5144
rect 1491 5110 1492 5144
rect 1456 5076 1492 5110
rect 1456 5042 1457 5076
rect 1491 5042 1492 5076
rect 1456 5008 1492 5042
rect 1456 4974 1457 5008
rect 1491 4974 1492 5008
rect 1456 4940 1492 4974
rect 1456 4906 1457 4940
rect 1491 4906 1492 4940
rect 1456 4872 1492 4906
rect 1456 4838 1457 4872
rect 1491 4838 1492 4872
rect 1456 4804 1492 4838
rect 1456 4770 1457 4804
rect 1491 4770 1492 4804
rect 1456 4736 1492 4770
rect 1456 4702 1457 4736
rect 1491 4702 1492 4736
rect 1456 4668 1492 4702
rect 1456 4634 1457 4668
rect 1491 4634 1492 4668
rect 1456 4600 1492 4634
rect 1456 4566 1457 4600
rect 1491 4566 1492 4600
rect 1456 4532 1492 4566
rect 1456 4498 1457 4532
rect 1491 4498 1492 4532
rect 1456 4464 1492 4498
rect 1456 4430 1457 4464
rect 1491 4430 1492 4464
rect 1456 4396 1492 4430
rect 1456 4362 1457 4396
rect 1491 4362 1492 4396
rect 1456 4328 1492 4362
rect 1456 4294 1457 4328
rect 1491 4294 1492 4328
rect 1456 4260 1492 4294
rect 1456 4226 1457 4260
rect 1491 4226 1492 4260
rect 1456 4192 1492 4226
rect 1456 4158 1457 4192
rect 1491 4158 1492 4192
rect 1456 4124 1492 4158
rect 1456 4090 1457 4124
rect 1491 4090 1492 4124
rect 1456 4056 1492 4090
rect 1456 4022 1457 4056
rect 1491 4022 1492 4056
rect 1456 3988 1492 4022
rect 1456 3954 1457 3988
rect 1491 3954 1492 3988
rect 1456 3920 1492 3954
rect 1456 3886 1457 3920
rect 1491 3886 1492 3920
rect 1456 3852 1492 3886
rect 1456 3818 1457 3852
rect 1491 3818 1492 3852
rect 1456 3784 1492 3818
rect 1456 3750 1457 3784
rect 1491 3750 1492 3784
rect 1456 3716 1492 3750
rect 1456 3682 1457 3716
rect 1491 3682 1492 3716
rect 1456 3648 1492 3682
rect 1456 3614 1457 3648
rect 1491 3614 1492 3648
rect 1456 3580 1492 3614
rect 1456 3546 1457 3580
rect 1491 3546 1492 3580
rect 1456 3512 1492 3546
rect 1456 3478 1457 3512
rect 1491 3478 1492 3512
rect 1456 3444 1492 3478
rect 1456 3410 1457 3444
rect 1491 3410 1492 3444
rect 1456 3376 1492 3410
rect 1456 3342 1457 3376
rect 1491 3342 1492 3376
rect 1456 3308 1492 3342
rect 1456 3274 1457 3308
rect 1491 3274 1492 3308
rect 1456 3240 1492 3274
rect 1456 3206 1457 3240
rect 1491 3206 1492 3240
rect 1456 3172 1492 3206
rect 1456 3138 1457 3172
rect 1491 3138 1492 3172
rect 1456 3104 1492 3138
rect 1456 3070 1457 3104
rect 1491 3070 1492 3104
rect 1456 3036 1492 3070
rect 1456 3002 1457 3036
rect 1491 3002 1492 3036
rect 1456 2968 1492 3002
rect 1456 2934 1457 2968
rect 1491 2934 1492 2968
rect 1456 2900 1492 2934
rect 1456 2866 1457 2900
rect 1491 2866 1492 2900
rect 1456 2832 1492 2866
rect 1456 2798 1457 2832
rect 1491 2798 1492 2832
rect 1456 2764 1492 2798
rect 1456 2730 1457 2764
rect 1491 2730 1492 2764
rect 1456 2696 1492 2730
rect 1456 2662 1457 2696
rect 1491 2662 1492 2696
rect 1456 2628 1492 2662
rect 1456 2594 1457 2628
rect 1491 2594 1492 2628
rect 1456 2560 1492 2594
rect 1456 2526 1457 2560
rect 1491 2526 1492 2560
rect 1456 2492 1492 2526
rect 1456 2458 1457 2492
rect 1491 2458 1492 2492
rect 1456 2424 1492 2458
rect 1456 2390 1457 2424
rect 1491 2390 1492 2424
rect 1456 2356 1492 2390
rect 1456 2322 1457 2356
rect 1491 2322 1492 2356
rect 1456 2288 1492 2322
rect 1456 2254 1457 2288
rect 1491 2254 1492 2288
rect 4092 7090 4128 7124
rect 4092 7056 4093 7090
rect 4127 7056 4128 7090
rect 4092 7022 4128 7056
rect 4092 6988 4093 7022
rect 4127 6988 4128 7022
rect 4092 6954 4128 6988
rect 4092 6920 4093 6954
rect 4127 6920 4128 6954
rect 4092 6886 4128 6920
rect 4092 6852 4093 6886
rect 4127 6852 4128 6886
rect 4092 6818 4128 6852
rect 4092 6784 4093 6818
rect 4127 6784 4128 6818
rect 4092 6750 4128 6784
rect 4092 6716 4093 6750
rect 4127 6716 4128 6750
rect 4092 6682 4128 6716
rect 4092 6648 4093 6682
rect 4127 6648 4128 6682
rect 4092 6614 4128 6648
rect 4092 6580 4093 6614
rect 4127 6580 4128 6614
rect 4092 6546 4128 6580
rect 4092 6512 4093 6546
rect 4127 6512 4128 6546
rect 4092 6478 4128 6512
rect 4092 6444 4093 6478
rect 4127 6444 4128 6478
rect 4092 6410 4128 6444
rect 4092 6376 4093 6410
rect 4127 6376 4128 6410
rect 4092 6342 4128 6376
rect 4092 6308 4093 6342
rect 4127 6308 4128 6342
rect 4092 6274 4128 6308
rect 4092 6240 4093 6274
rect 4127 6240 4128 6274
rect 4092 6206 4128 6240
rect 4092 6172 4093 6206
rect 4127 6172 4128 6206
rect 4092 6138 4128 6172
rect 4092 6104 4093 6138
rect 4127 6104 4128 6138
rect 4092 6070 4128 6104
rect 4092 6036 4093 6070
rect 4127 6036 4128 6070
rect 4092 6002 4128 6036
rect 4092 5968 4093 6002
rect 4127 5968 4128 6002
rect 4092 5934 4128 5968
rect 4092 5900 4093 5934
rect 4127 5900 4128 5934
rect 4092 5866 4128 5900
rect 4092 5832 4093 5866
rect 4127 5832 4128 5866
rect 4092 5798 4128 5832
rect 4092 5764 4093 5798
rect 4127 5764 4128 5798
rect 4092 5730 4128 5764
rect 4092 5696 4093 5730
rect 4127 5696 4128 5730
rect 4092 5662 4128 5696
rect 4092 5628 4093 5662
rect 4127 5628 4128 5662
rect 4092 5594 4128 5628
rect 4092 5560 4093 5594
rect 4127 5560 4128 5594
rect 4092 5526 4128 5560
rect 4092 5492 4093 5526
rect 4127 5492 4128 5526
rect 4092 5458 4128 5492
rect 4092 5424 4093 5458
rect 4127 5424 4128 5458
rect 4092 5390 4128 5424
rect 4092 5356 4093 5390
rect 4127 5356 4128 5390
rect 4092 5322 4128 5356
rect 4092 5288 4093 5322
rect 4127 5288 4128 5322
rect 4092 5254 4128 5288
rect 4092 5220 4093 5254
rect 4127 5220 4128 5254
rect 4092 5186 4128 5220
rect 4092 5152 4093 5186
rect 4127 5152 4128 5186
rect 4092 5118 4128 5152
rect 4092 5084 4093 5118
rect 4127 5084 4128 5118
rect 4092 5050 4128 5084
rect 4092 5016 4093 5050
rect 4127 5016 4128 5050
rect 4092 4982 4128 5016
rect 4092 4948 4093 4982
rect 4127 4948 4128 4982
rect 4092 4914 4128 4948
rect 4092 4880 4093 4914
rect 4127 4880 4128 4914
rect 4092 4846 4128 4880
rect 4092 4812 4093 4846
rect 4127 4812 4128 4846
rect 4092 4778 4128 4812
rect 4092 4744 4093 4778
rect 4127 4744 4128 4778
rect 4092 4710 4128 4744
rect 4092 4676 4093 4710
rect 4127 4676 4128 4710
rect 4092 4642 4128 4676
rect 4092 4608 4093 4642
rect 4127 4608 4128 4642
rect 4092 4574 4128 4608
rect 4092 4540 4093 4574
rect 4127 4540 4128 4574
rect 4092 4506 4128 4540
rect 4092 4472 4093 4506
rect 4127 4472 4128 4506
rect 4092 4438 4128 4472
rect 4092 4404 4093 4438
rect 4127 4404 4128 4438
rect 4092 4370 4128 4404
rect 4092 4336 4093 4370
rect 4127 4336 4128 4370
rect 4092 4302 4128 4336
rect 4092 4268 4093 4302
rect 4127 4268 4128 4302
rect 4092 4234 4128 4268
rect 4092 4200 4093 4234
rect 4127 4200 4128 4234
rect 4092 4166 4128 4200
rect 4092 4132 4093 4166
rect 4127 4132 4128 4166
rect 4092 4098 4128 4132
rect 4092 4064 4093 4098
rect 4127 4064 4128 4098
rect 4092 4030 4128 4064
rect 4092 3996 4093 4030
rect 4127 3996 4128 4030
rect 4092 3962 4128 3996
rect 4092 3928 4093 3962
rect 4127 3928 4128 3962
rect 4092 3894 4128 3928
rect 4092 3860 4093 3894
rect 4127 3860 4128 3894
rect 4092 3826 4128 3860
rect 4092 3792 4093 3826
rect 4127 3792 4128 3826
rect 4092 3758 4128 3792
rect 4092 3724 4093 3758
rect 4127 3724 4128 3758
rect 4092 3690 4128 3724
rect 4092 3656 4093 3690
rect 4127 3656 4128 3690
rect 4092 3622 4128 3656
rect 4092 3588 4093 3622
rect 4127 3588 4128 3622
rect 4092 3554 4128 3588
rect 4092 3520 4093 3554
rect 4127 3520 4128 3554
rect 4092 3486 4128 3520
rect 4092 3452 4093 3486
rect 4127 3452 4128 3486
rect 4092 3418 4128 3452
rect 4092 3384 4093 3418
rect 4127 3384 4128 3418
rect 4092 3350 4128 3384
rect 4092 3316 4093 3350
rect 4127 3316 4128 3350
rect 4092 3282 4128 3316
rect 4092 3248 4093 3282
rect 4127 3248 4128 3282
rect 4092 3214 4128 3248
rect 4092 3180 4093 3214
rect 4127 3180 4128 3214
rect 4092 3146 4128 3180
rect 4092 3112 4093 3146
rect 4127 3112 4128 3146
rect 4092 3078 4128 3112
rect 4092 3044 4093 3078
rect 4127 3044 4128 3078
rect 4092 3010 4128 3044
rect 4092 2976 4093 3010
rect 4127 2976 4128 3010
rect 4092 2942 4128 2976
rect 4092 2908 4093 2942
rect 4127 2908 4128 2942
rect 4092 2874 4128 2908
rect 4092 2840 4093 2874
rect 4127 2840 4128 2874
rect 4092 2806 4128 2840
rect 4092 2772 4093 2806
rect 4127 2772 4128 2806
rect 4092 2738 4128 2772
rect 4092 2704 4093 2738
rect 4127 2704 4128 2738
rect 4092 2670 4128 2704
rect 4092 2636 4093 2670
rect 4127 2636 4128 2670
rect 4092 2602 4128 2636
rect 4092 2568 4093 2602
rect 4127 2568 4128 2602
rect 4092 2534 4128 2568
rect 4092 2500 4093 2534
rect 4127 2500 4128 2534
rect 4092 2466 4128 2500
rect 4092 2432 4093 2466
rect 4127 2432 4128 2466
rect 4092 2398 4128 2432
rect 4092 2364 4093 2398
rect 4127 2364 4128 2398
rect 4092 2330 4128 2364
rect 4092 2296 4093 2330
rect 4127 2296 4128 2330
rect 4092 2262 4128 2296
rect 1456 2220 1492 2254
rect 1456 2186 1457 2220
rect 1491 2186 1492 2220
rect 1456 2152 1492 2186
rect 1456 2118 1457 2152
rect 1491 2118 1492 2152
rect 1456 2104 1492 2118
rect 4092 2228 4093 2262
rect 4127 2228 4128 2262
rect 4092 2194 4128 2228
rect 4092 2160 4093 2194
rect 4127 2160 4128 2194
rect 4092 2126 4128 2160
rect 4092 2104 4093 2126
rect 1456 2103 4093 2104
rect 1456 2069 1526 2103
rect 1560 2069 1594 2103
rect 1628 2069 1662 2103
rect 1696 2069 1730 2103
rect 1764 2069 1798 2103
rect 1832 2069 1866 2103
rect 1900 2069 1934 2103
rect 1968 2069 2002 2103
rect 2036 2069 2070 2103
rect 2104 2069 2138 2103
rect 2172 2069 2206 2103
rect 2240 2069 2274 2103
rect 2308 2069 2342 2103
rect 2376 2069 2410 2103
rect 2444 2069 2478 2103
rect 2512 2069 2546 2103
rect 2580 2069 2614 2103
rect 2648 2069 2682 2103
rect 2716 2069 2750 2103
rect 2784 2069 2818 2103
rect 2852 2069 2886 2103
rect 2920 2069 2954 2103
rect 2988 2069 3022 2103
rect 3056 2069 3090 2103
rect 3124 2069 3158 2103
rect 3192 2069 3226 2103
rect 3260 2069 3294 2103
rect 3328 2069 3362 2103
rect 3396 2069 3430 2103
rect 3464 2069 3498 2103
rect 3532 2069 3566 2103
rect 3600 2069 3634 2103
rect 3668 2069 3702 2103
rect 3736 2069 3770 2103
rect 3804 2069 3838 2103
rect 3872 2069 3906 2103
rect 3940 2069 3974 2103
rect 4008 2092 4093 2103
rect 4127 2092 4128 2126
rect 4008 2069 4128 2092
rect 1456 2068 4128 2069
rect 1456 1840 1492 2068
rect 4092 2058 4128 2068
rect 4092 2024 4093 2058
rect 4127 2024 4128 2058
rect 4092 1990 4128 2024
rect 1456 1806 1457 1840
rect 1491 1806 1492 1840
rect 1456 1772 1492 1806
rect 1456 1738 1457 1772
rect 1491 1738 1492 1772
rect 1456 1704 1492 1738
rect 1456 1670 1457 1704
rect 1491 1670 1492 1704
rect 1456 1636 1492 1670
rect 1456 1602 1457 1636
rect 1491 1602 1492 1636
rect 1456 1568 1492 1602
rect 1456 1534 1457 1568
rect 1491 1534 1492 1568
rect 1456 1500 1492 1534
rect 1456 1466 1457 1500
rect 1491 1466 1492 1500
rect 1456 1432 1492 1466
rect 1456 1398 1457 1432
rect 1491 1398 1492 1432
rect 1456 1364 1492 1398
rect 1456 1330 1457 1364
rect 1491 1330 1492 1364
rect 1456 1296 1492 1330
rect 1456 1262 1457 1296
rect 1491 1262 1492 1296
rect 1456 1228 1492 1262
rect 1456 1194 1457 1228
rect 1491 1194 1492 1228
rect 1456 1160 1492 1194
rect 1456 1126 1457 1160
rect 1491 1126 1492 1160
rect 1456 1092 1492 1126
rect 1456 1058 1457 1092
rect 1491 1058 1492 1092
rect 1456 1024 1492 1058
rect 1456 990 1457 1024
rect 1491 990 1492 1024
rect 1456 956 1492 990
rect 1456 922 1457 956
rect 1491 922 1492 956
rect 1456 888 1492 922
rect 1456 854 1457 888
rect 1491 854 1492 888
rect 1456 820 1492 854
rect 1456 786 1457 820
rect 1491 786 1492 820
rect 1456 752 1492 786
rect 1456 718 1457 752
rect 1491 718 1492 752
rect 1456 684 1492 718
rect 1456 650 1457 684
rect 1491 650 1492 684
rect 1456 616 1492 650
rect 1456 582 1457 616
rect 1491 582 1492 616
rect 1456 548 1492 582
rect 1456 514 1457 548
rect 1491 514 1492 548
rect 1456 462 1492 514
rect 4092 1956 4093 1990
rect 4127 1956 4128 1990
rect 4092 1922 4128 1956
rect 4092 1888 4093 1922
rect 4127 1888 4128 1922
rect 4092 1854 4128 1888
rect 4092 1820 4093 1854
rect 4127 1820 4128 1854
rect 4092 1786 4128 1820
rect 4092 1752 4093 1786
rect 4127 1752 4128 1786
rect 4092 1718 4128 1752
rect 4092 1684 4093 1718
rect 4127 1684 4128 1718
rect 4092 1650 4128 1684
rect 4092 1616 4093 1650
rect 4127 1616 4128 1650
rect 4092 1582 4128 1616
rect 4092 1548 4093 1582
rect 4127 1548 4128 1582
rect 4092 1514 4128 1548
rect 4092 1480 4093 1514
rect 4127 1480 4128 1514
rect 4092 1446 4128 1480
rect 4092 1412 4093 1446
rect 4127 1412 4128 1446
rect 4092 1378 4128 1412
rect 4092 1344 4093 1378
rect 4127 1344 4128 1378
rect 4092 1310 4128 1344
rect 4092 1276 4093 1310
rect 4127 1276 4128 1310
rect 4092 1242 4128 1276
rect 4092 1208 4093 1242
rect 4127 1208 4128 1242
rect 4092 1174 4128 1208
rect 4092 1140 4093 1174
rect 4127 1140 4128 1174
rect 4092 1106 4128 1140
rect 4092 1072 4093 1106
rect 4127 1072 4128 1106
rect 4092 1038 4128 1072
rect 4092 1004 4093 1038
rect 4127 1004 4128 1038
rect 4092 970 4128 1004
rect 4092 936 4093 970
rect 4127 936 4128 970
rect 4092 902 4128 936
rect 4092 868 4093 902
rect 4127 868 4128 902
rect 4092 834 4128 868
rect 4092 800 4093 834
rect 4127 800 4128 834
rect 4092 766 4128 800
rect 4092 732 4093 766
rect 4127 732 4128 766
rect 4092 698 4128 732
rect 4092 664 4093 698
rect 4127 664 4128 698
rect 4092 630 4128 664
rect 4092 596 4093 630
rect 4127 596 4128 630
rect 4092 562 4128 596
rect 4092 528 4093 562
rect 4127 528 4128 562
rect 4092 494 4128 528
rect 4092 462 4093 494
rect 8 413 9 447
rect 43 413 44 447
rect 8 312 44 413
rect 1266 461 4093 462
rect 1266 427 1300 461
rect 1334 427 1368 461
rect 1402 427 1490 461
rect 1524 427 1558 461
rect 1592 427 1626 461
rect 1660 427 1694 461
rect 1728 427 1762 461
rect 1796 427 1830 461
rect 1864 427 1898 461
rect 1932 427 1966 461
rect 2000 427 2034 461
rect 2068 427 2102 461
rect 2136 427 2170 461
rect 2204 427 2238 461
rect 2272 427 2306 461
rect 2340 427 2374 461
rect 2408 427 2442 461
rect 2476 427 2510 461
rect 2544 427 2578 461
rect 2612 427 2646 461
rect 2680 427 2714 461
rect 2748 427 2782 461
rect 2816 427 2850 461
rect 2884 427 2918 461
rect 2952 427 2986 461
rect 3020 427 3054 461
rect 3088 427 3122 461
rect 3156 427 3190 461
rect 3224 427 3258 461
rect 3292 427 3326 461
rect 3360 427 3394 461
rect 3428 427 3462 461
rect 3496 427 3530 461
rect 3564 427 3598 461
rect 3632 427 3666 461
rect 3700 427 3734 461
rect 3768 427 3802 461
rect 3836 427 3870 461
rect 3904 427 3938 461
rect 3972 427 4006 461
rect 4040 460 4093 461
rect 4127 460 4128 494
rect 4040 427 4128 460
rect 1266 426 4128 427
rect 1266 312 1302 426
rect 8 276 1302 312
<< mvpsubdiffcont >>
rect 198 10632 232 10666
rect 297 10665 331 10699
rect 365 10665 399 10699
rect 433 10665 467 10699
rect 501 10665 535 10699
rect 569 10665 603 10699
rect 637 10665 671 10699
rect 705 10665 739 10699
rect 773 10665 807 10699
rect 841 10665 875 10699
rect 909 10665 943 10699
rect 977 10665 1011 10699
rect 1045 10665 1079 10699
rect 198 10564 232 10598
rect 198 10496 232 10530
rect 1078 10563 1112 10597
rect 198 10428 232 10462
rect 198 10360 232 10394
rect 198 10292 232 10326
rect 198 10224 232 10258
rect 198 10156 232 10190
rect 198 10088 232 10122
rect 198 10020 232 10054
rect 198 9952 232 9986
rect 198 9884 232 9918
rect 198 9816 232 9850
rect 198 9748 232 9782
rect 198 9680 232 9714
rect 198 9612 232 9646
rect 198 9544 232 9578
rect 198 9476 232 9510
rect 198 9408 232 9442
rect 198 9340 232 9374
rect 198 9272 232 9306
rect 198 9204 232 9238
rect 198 9136 232 9170
rect 198 9068 232 9102
rect 198 9000 232 9034
rect 198 8932 232 8966
rect 198 8864 232 8898
rect 198 8796 232 8830
rect 198 8728 232 8762
rect 1078 10495 1112 10529
rect 1078 10427 1112 10461
rect 1078 10359 1112 10393
rect 1078 10291 1112 10325
rect 1078 10223 1112 10257
rect 1078 10155 1112 10189
rect 1078 10087 1112 10121
rect 1078 10019 1112 10053
rect 1078 9951 1112 9985
rect 1078 9883 1112 9917
rect 1078 9815 1112 9849
rect 1078 9747 1112 9781
rect 1078 9679 1112 9713
rect 1078 9611 1112 9645
rect 1078 9543 1112 9577
rect 1078 9475 1112 9509
rect 1078 9407 1112 9441
rect 1078 9339 1112 9373
rect 1078 9271 1112 9305
rect 1078 9203 1112 9237
rect 1078 9135 1112 9169
rect 1078 9067 1112 9101
rect 1078 8999 1112 9033
rect 1078 8931 1112 8965
rect 1078 8863 1112 8897
rect 1078 8795 1112 8829
rect 1078 8727 1112 8761
rect 198 8660 232 8694
rect 1078 8659 1112 8693
rect 198 8592 232 8626
rect 1078 8591 1112 8625
rect 198 8524 232 8558
rect 1078 8523 1112 8557
rect 198 8456 232 8490
rect 198 8388 232 8422
rect 198 8320 232 8354
rect 198 8252 232 8286
rect 198 8184 232 8218
rect 198 8116 232 8150
rect 198 8048 232 8082
rect 198 7980 232 8014
rect 198 7912 232 7946
rect 198 7844 232 7878
rect 198 7776 232 7810
rect 198 7708 232 7742
rect 198 7640 232 7674
rect 198 7572 232 7606
rect 198 7504 232 7538
rect 198 7436 232 7470
rect 198 7368 232 7402
rect 198 7300 232 7334
rect 198 7232 232 7266
rect 198 7164 232 7198
rect 198 7096 232 7130
rect 198 7028 232 7062
rect 198 6960 232 6994
rect 198 6892 232 6926
rect 198 6824 232 6858
rect 198 6756 232 6790
rect 198 6688 232 6722
rect 1078 8455 1112 8489
rect 1078 8387 1112 8421
rect 1078 8319 1112 8353
rect 1078 8251 1112 8285
rect 1078 8183 1112 8217
rect 1078 8115 1112 8149
rect 1078 8047 1112 8081
rect 1078 7979 1112 8013
rect 1078 7911 1112 7945
rect 1078 7843 1112 7877
rect 1078 7775 1112 7809
rect 1078 7707 1112 7741
rect 1078 7639 1112 7673
rect 1078 7571 1112 7605
rect 1078 7503 1112 7537
rect 1078 7435 1112 7469
rect 1078 7367 1112 7401
rect 1078 7299 1112 7333
rect 1078 7231 1112 7265
rect 1078 7163 1112 7197
rect 1078 7095 1112 7129
rect 1078 7027 1112 7061
rect 1078 6959 1112 6993
rect 1078 6891 1112 6925
rect 1078 6823 1112 6857
rect 1078 6755 1112 6789
rect 198 6620 232 6654
rect 1078 6687 1112 6721
rect 198 6552 232 6586
rect 1078 6619 1112 6653
rect 198 6484 232 6518
rect 1078 6551 1112 6585
rect 198 6416 232 6450
rect 198 6348 232 6382
rect 198 6280 232 6314
rect 198 6212 232 6246
rect 198 6144 232 6178
rect 198 6076 232 6110
rect 198 6008 232 6042
rect 198 5940 232 5974
rect 198 5872 232 5906
rect 198 5804 232 5838
rect 198 5736 232 5770
rect 198 5668 232 5702
rect 198 5600 232 5634
rect 198 5532 232 5566
rect 198 5464 232 5498
rect 198 5396 232 5430
rect 198 5328 232 5362
rect 198 5260 232 5294
rect 198 5192 232 5226
rect 198 5124 232 5158
rect 198 5056 232 5090
rect 198 4988 232 5022
rect 198 4920 232 4954
rect 198 4852 232 4886
rect 198 4784 232 4818
rect 198 4716 232 4750
rect 198 4648 232 4682
rect 1078 6483 1112 6517
rect 1078 6415 1112 6449
rect 1078 6347 1112 6381
rect 1078 6279 1112 6313
rect 1078 6211 1112 6245
rect 1078 6143 1112 6177
rect 1078 6075 1112 6109
rect 1078 6007 1112 6041
rect 1078 5939 1112 5973
rect 1078 5871 1112 5905
rect 1078 5803 1112 5837
rect 1078 5735 1112 5769
rect 1078 5667 1112 5701
rect 1078 5599 1112 5633
rect 1078 5531 1112 5565
rect 1078 5463 1112 5497
rect 1078 5395 1112 5429
rect 1078 5327 1112 5361
rect 1078 5259 1112 5293
rect 1078 5191 1112 5225
rect 1078 5123 1112 5157
rect 1078 5055 1112 5089
rect 1078 4987 1112 5021
rect 1078 4919 1112 4953
rect 1078 4851 1112 4885
rect 1078 4783 1112 4817
rect 1078 4715 1112 4749
rect 198 4580 232 4614
rect 1078 4647 1112 4681
rect 198 4512 232 4546
rect 1078 4579 1112 4613
rect 198 4444 232 4478
rect 1078 4511 1112 4545
rect 198 4376 232 4410
rect 198 4308 232 4342
rect 198 4240 232 4274
rect 198 4172 232 4206
rect 198 4104 232 4138
rect 198 4036 232 4070
rect 198 3968 232 4002
rect 198 3900 232 3934
rect 198 3832 232 3866
rect 198 3764 232 3798
rect 198 3696 232 3730
rect 198 3628 232 3662
rect 198 3560 232 3594
rect 198 3492 232 3526
rect 198 3424 232 3458
rect 198 3356 232 3390
rect 198 3288 232 3322
rect 198 3220 232 3254
rect 198 3152 232 3186
rect 198 3084 232 3118
rect 198 3016 232 3050
rect 198 2948 232 2982
rect 198 2880 232 2914
rect 198 2812 232 2846
rect 198 2744 232 2778
rect 198 2676 232 2710
rect 1078 4443 1112 4477
rect 1078 4375 1112 4409
rect 1078 4307 1112 4341
rect 1078 4239 1112 4273
rect 1078 4171 1112 4205
rect 1078 4103 1112 4137
rect 1078 4035 1112 4069
rect 1078 3967 1112 4001
rect 1078 3899 1112 3933
rect 1078 3831 1112 3865
rect 1078 3763 1112 3797
rect 1078 3695 1112 3729
rect 1078 3627 1112 3661
rect 1078 3559 1112 3593
rect 1078 3491 1112 3525
rect 1078 3423 1112 3457
rect 1078 3355 1112 3389
rect 1078 3287 1112 3321
rect 1078 3219 1112 3253
rect 1078 3151 1112 3185
rect 1078 3083 1112 3117
rect 1078 3015 1112 3049
rect 1078 2947 1112 2981
rect 1078 2879 1112 2913
rect 1078 2811 1112 2845
rect 1078 2743 1112 2777
rect 1078 2675 1112 2709
rect 198 2608 232 2642
rect 1078 2607 1112 2641
rect 198 2540 232 2574
rect 1078 2539 1112 2573
rect 198 2472 232 2506
rect 1078 2471 1112 2505
rect 198 2404 232 2438
rect 198 2336 232 2370
rect 198 2268 232 2302
rect 198 2200 232 2234
rect 198 2132 232 2166
rect 198 2064 232 2098
rect 198 1996 232 2030
rect 198 1928 232 1962
rect 198 1860 232 1894
rect 198 1792 232 1826
rect 198 1724 232 1758
rect 198 1656 232 1690
rect 198 1588 232 1622
rect 198 1520 232 1554
rect 198 1452 232 1486
rect 198 1384 232 1418
rect 198 1316 232 1350
rect 198 1248 232 1282
rect 198 1180 232 1214
rect 198 1112 232 1146
rect 198 1044 232 1078
rect 198 976 232 1010
rect 198 908 232 942
rect 198 840 232 874
rect 198 772 232 806
rect 198 704 232 738
rect 198 636 232 670
rect 1078 2403 1112 2437
rect 1078 2335 1112 2369
rect 1078 2267 1112 2301
rect 1078 2199 1112 2233
rect 1078 2131 1112 2165
rect 1078 2063 1112 2097
rect 1078 1995 1112 2029
rect 1078 1927 1112 1961
rect 1078 1859 1112 1893
rect 1078 1791 1112 1825
rect 1078 1723 1112 1757
rect 1078 1655 1112 1689
rect 1078 1587 1112 1621
rect 1078 1519 1112 1553
rect 1078 1451 1112 1485
rect 1078 1383 1112 1417
rect 1078 1315 1112 1349
rect 1078 1247 1112 1281
rect 1078 1179 1112 1213
rect 1078 1111 1112 1145
rect 1078 1043 1112 1077
rect 1078 975 1112 1009
rect 1078 907 1112 941
rect 1078 839 1112 873
rect 1078 771 1112 805
rect 1078 703 1112 737
rect 198 568 232 602
rect 1078 635 1112 669
rect 1078 567 1112 601
rect 231 466 265 500
rect 299 466 333 500
rect 367 466 401 500
rect 435 466 469 500
rect 503 466 537 500
rect 571 466 605 500
rect 639 466 673 500
rect 707 466 741 500
rect 775 466 809 500
rect 843 466 877 500
rect 911 466 945 500
rect 979 466 1013 500
rect 1078 499 1112 533
rect 1690 10656 1724 10690
rect 1801 10689 1835 10723
rect 1869 10689 1903 10723
rect 1937 10689 1971 10723
rect 2005 10689 2039 10723
rect 2073 10689 2107 10723
rect 2141 10689 2175 10723
rect 2209 10689 2243 10723
rect 2277 10689 2311 10723
rect 2345 10689 2379 10723
rect 2413 10689 2447 10723
rect 2481 10689 2515 10723
rect 2549 10689 2583 10723
rect 2617 10689 2651 10723
rect 2685 10689 2719 10723
rect 2753 10689 2787 10723
rect 2821 10689 2855 10723
rect 2889 10689 2923 10723
rect 2957 10689 2991 10723
rect 3025 10689 3059 10723
rect 3093 10689 3127 10723
rect 3161 10689 3195 10723
rect 3229 10689 3263 10723
rect 3297 10689 3331 10723
rect 3365 10689 3399 10723
rect 3433 10689 3467 10723
rect 3501 10689 3535 10723
rect 3569 10689 3603 10723
rect 3637 10689 3671 10723
rect 3705 10689 3739 10723
rect 3773 10689 3807 10723
rect 3841 10689 3875 10723
rect 3909 10689 3943 10723
rect 3977 10689 4011 10723
rect 4045 10689 4079 10723
rect 4113 10689 4147 10723
rect 4181 10689 4215 10723
rect 4249 10689 4283 10723
rect 4317 10689 4351 10723
rect 4385 10689 4419 10723
rect 4453 10689 4487 10723
rect 4521 10689 4555 10723
rect 4589 10689 4623 10723
rect 4657 10689 4691 10723
rect 4725 10689 4759 10723
rect 4793 10689 4827 10723
rect 4861 10689 4895 10723
rect 4929 10689 4963 10723
rect 4997 10689 5031 10723
rect 5065 10689 5099 10723
rect 5133 10689 5167 10723
rect 5201 10689 5235 10723
rect 5269 10689 5303 10723
rect 5337 10689 5371 10723
rect 5405 10689 5439 10723
rect 5473 10689 5507 10723
rect 5541 10689 5575 10723
rect 5609 10689 5643 10723
rect 5677 10689 5711 10723
rect 5745 10689 5779 10723
rect 5813 10689 5847 10723
rect 5881 10689 5915 10723
rect 5949 10689 5983 10723
rect 6017 10689 6051 10723
rect 6085 10689 6119 10723
rect 6153 10689 6187 10723
rect 6221 10689 6255 10723
rect 6289 10689 6323 10723
rect 6357 10689 6391 10723
rect 6425 10689 6459 10723
rect 6493 10689 6527 10723
rect 6561 10689 6595 10723
rect 6629 10689 6663 10723
rect 6697 10689 6731 10723
rect 6765 10689 6799 10723
rect 6833 10689 6867 10723
rect 6901 10689 6935 10723
rect 6969 10689 7003 10723
rect 7037 10689 7071 10723
rect 7105 10689 7139 10723
rect 7173 10689 7207 10723
rect 7241 10689 7275 10723
rect 7309 10689 7343 10723
rect 7377 10689 7411 10723
rect 7445 10689 7479 10723
rect 7513 10689 7547 10723
rect 7581 10689 7615 10723
rect 7649 10689 7683 10723
rect 7717 10689 7751 10723
rect 7785 10689 7819 10723
rect 7853 10689 7887 10723
rect 7921 10689 7955 10723
rect 7989 10689 8023 10723
rect 8057 10689 8091 10723
rect 8125 10689 8159 10723
rect 8193 10689 8227 10723
rect 1690 10588 1724 10622
rect 8226 10612 8260 10646
rect 1690 10520 1724 10554
rect 1690 10452 1724 10486
rect 1690 10384 1724 10418
rect 1690 10316 1724 10350
rect 1690 10248 1724 10282
rect 1690 10180 1724 10214
rect 1690 10112 1724 10146
rect 1690 10044 1724 10078
rect 1690 9976 1724 10010
rect 1690 9908 1724 9942
rect 1690 9840 1724 9874
rect 1690 9772 1724 9806
rect 8226 10544 8260 10578
rect 8226 10476 8260 10510
rect 8226 10408 8260 10442
rect 8226 10340 8260 10374
rect 8226 10272 8260 10306
rect 8226 10204 8260 10238
rect 8226 10136 8260 10170
rect 8226 10068 8260 10102
rect 8226 10000 8260 10034
rect 8226 9932 8260 9966
rect 8226 9864 8260 9898
rect 8226 9796 8260 9830
rect 1690 9704 1724 9738
rect 8226 9728 8260 9762
rect 1690 9636 1724 9670
rect 1690 9568 1724 9602
rect 1690 9500 1724 9534
rect 1690 9432 1724 9466
rect 1690 9364 1724 9398
rect 1690 9296 1724 9330
rect 1690 9228 1724 9262
rect 1690 9160 1724 9194
rect 1690 9092 1724 9126
rect 1690 9024 1724 9058
rect 1690 8956 1724 8990
rect 1690 8888 1724 8922
rect 8226 9660 8260 9694
rect 8226 9592 8260 9626
rect 8226 9524 8260 9558
rect 8226 9456 8260 9490
rect 8226 9388 8260 9422
rect 8226 9320 8260 9354
rect 8226 9252 8260 9286
rect 8226 9184 8260 9218
rect 8226 9116 8260 9150
rect 8226 9048 8260 9082
rect 8226 8980 8260 9014
rect 8226 8912 8260 8946
rect 8226 8844 8260 8878
rect 1646 8710 1680 8744
rect 1723 8743 1757 8777
rect 1791 8743 1825 8777
rect 1859 8743 1893 8777
rect 1927 8743 1961 8777
rect 1995 8743 2029 8777
rect 2063 8743 2097 8777
rect 2131 8743 2165 8777
rect 2199 8743 2233 8777
rect 2267 8743 2301 8777
rect 2335 8743 2369 8777
rect 2403 8743 2437 8777
rect 2471 8743 2505 8777
rect 2539 8743 2573 8777
rect 2607 8743 2641 8777
rect 2675 8743 2709 8777
rect 2743 8743 2777 8777
rect 2811 8743 2845 8777
rect 2879 8743 2913 8777
rect 2947 8743 2981 8777
rect 3015 8743 3049 8777
rect 3083 8743 3117 8777
rect 3151 8743 3185 8777
rect 3219 8743 3253 8777
rect 3287 8743 3321 8777
rect 3355 8743 3389 8777
rect 3423 8743 3457 8777
rect 3491 8743 3525 8777
rect 3559 8743 3593 8777
rect 3627 8743 3661 8777
rect 3695 8743 3729 8777
rect 3763 8743 3797 8777
rect 3831 8743 3865 8777
rect 3899 8743 3933 8777
rect 3967 8743 4001 8777
rect 4035 8743 4069 8777
rect 4103 8743 4137 8777
rect 4171 8743 4205 8777
rect 4239 8743 4273 8777
rect 4307 8743 4341 8777
rect 4375 8743 4409 8777
rect 4443 8743 4477 8777
rect 4511 8743 4545 8777
rect 4579 8743 4613 8777
rect 4647 8743 4681 8777
rect 4715 8743 4749 8777
rect 4783 8743 4817 8777
rect 4851 8743 4885 8777
rect 4919 8743 4953 8777
rect 4987 8743 5021 8777
rect 5055 8743 5089 8777
rect 5123 8743 5157 8777
rect 5191 8743 5225 8777
rect 5259 8743 5293 8777
rect 5327 8743 5361 8777
rect 5395 8743 5429 8777
rect 5463 8743 5497 8777
rect 5531 8743 5565 8777
rect 5599 8743 5633 8777
rect 5667 8743 5701 8777
rect 5735 8743 5769 8777
rect 5803 8743 5837 8777
rect 5871 8743 5905 8777
rect 5939 8743 5973 8777
rect 6007 8743 6041 8777
rect 6075 8743 6109 8777
rect 6143 8743 6177 8777
rect 6211 8743 6245 8777
rect 6279 8743 6313 8777
rect 6347 8743 6381 8777
rect 6415 8743 6449 8777
rect 6483 8743 6517 8777
rect 6551 8743 6585 8777
rect 6619 8743 6653 8777
rect 6687 8743 6721 8777
rect 6755 8743 6789 8777
rect 6823 8743 6857 8777
rect 6891 8743 6925 8777
rect 6959 8743 6993 8777
rect 7027 8743 7061 8777
rect 7095 8743 7129 8777
rect 7163 8743 7197 8777
rect 7231 8743 7265 8777
rect 7299 8743 7333 8777
rect 7367 8743 7401 8777
rect 7435 8743 7469 8777
rect 7503 8743 7537 8777
rect 7571 8743 7605 8777
rect 7639 8743 7673 8777
rect 7707 8743 7741 8777
rect 7775 8743 7809 8777
rect 7843 8743 7877 8777
rect 7911 8743 7945 8777
rect 7979 8743 8013 8777
rect 8047 8743 8081 8777
rect 8115 8743 8149 8777
rect 8226 8776 8260 8810
rect 1646 8642 1680 8676
rect 1646 8574 1680 8608
rect 1646 8506 1680 8540
rect 1646 8438 1680 8472
rect 1646 8370 1680 8404
rect 1646 8302 1680 8336
rect 1646 8234 1680 8268
rect 1646 8166 1680 8200
rect 1646 8098 1680 8132
rect 1646 8030 1680 8064
rect 1646 7962 1680 7996
rect 1646 7894 1680 7928
rect 1646 7826 1680 7860
rect 1646 7758 1680 7792
rect 1646 7690 1680 7724
rect 1646 7622 1680 7656
rect 1646 7554 1680 7588
rect 1679 7476 1713 7510
rect 1747 7476 1781 7510
rect 1815 7476 1849 7510
rect 1883 7476 1917 7510
rect 1951 7476 1985 7510
rect 2019 7476 2053 7510
rect 2087 7476 2121 7510
rect 2155 7476 2189 7510
rect 2223 7476 2257 7510
rect 2291 7476 2325 7510
rect 2359 7476 2393 7510
rect 2427 7476 2461 7510
rect 2495 7476 2529 7510
rect 2563 7476 2597 7510
rect 2631 7476 2665 7510
rect 2699 7476 2733 7510
rect 2767 7476 2801 7510
rect 2835 7476 2869 7510
rect 2903 7476 2937 7510
rect 2971 7476 3005 7510
rect 3039 7476 3073 7510
rect 3107 7476 3141 7510
rect 3175 7476 3209 7510
rect 3243 7476 3277 7510
rect 3311 7476 3345 7510
rect 3379 7476 3413 7510
rect 3447 7476 3481 7510
rect 3515 7476 3549 7510
rect 3583 7476 3617 7510
rect 3651 7476 3685 7510
rect 3719 7476 3753 7510
rect 3787 7476 3821 7510
rect 3855 7476 3889 7510
rect 3923 7476 3957 7510
rect 3991 7476 4025 7510
rect 4059 7476 4093 7510
rect 1646 7043 1680 7077
rect 1763 7076 1797 7110
rect 1831 7076 1865 7110
rect 1899 7076 1933 7110
rect 1967 7076 2001 7110
rect 2035 7076 2069 7110
rect 2103 7076 2137 7110
rect 2171 7076 2205 7110
rect 2239 7076 2273 7110
rect 2307 7076 2341 7110
rect 2375 7076 2409 7110
rect 2443 7076 2477 7110
rect 2511 7076 2545 7110
rect 2579 7076 2613 7110
rect 2647 7076 2681 7110
rect 2715 7076 2749 7110
rect 2783 7076 2817 7110
rect 2851 7076 2885 7110
rect 2919 7076 2953 7110
rect 2987 7076 3021 7110
rect 3055 7076 3089 7110
rect 3123 7076 3157 7110
rect 3191 7076 3225 7110
rect 3259 7076 3293 7110
rect 3327 7076 3361 7110
rect 3395 7076 3429 7110
rect 3463 7076 3497 7110
rect 3531 7076 3565 7110
rect 3599 7076 3633 7110
rect 3667 7076 3701 7110
rect 3735 7076 3769 7110
rect 3803 7076 3837 7110
rect 3871 7076 3905 7110
rect 1646 6975 1680 7009
rect 3904 7001 3938 7035
rect 1646 6907 1680 6941
rect 1646 6839 1680 6873
rect 1646 6771 1680 6805
rect 1646 6703 1680 6737
rect 1646 6635 1680 6669
rect 1646 6567 1680 6601
rect 1646 6499 1680 6533
rect 1646 6431 1680 6465
rect 1646 6363 1680 6397
rect 1646 6295 1680 6329
rect 1646 6227 1680 6261
rect 1646 6159 1680 6193
rect 1646 6091 1680 6125
rect 1646 6023 1680 6057
rect 1646 5955 1680 5989
rect 1646 5887 1680 5921
rect 3904 6933 3938 6967
rect 3904 6865 3938 6899
rect 3904 6797 3938 6831
rect 3904 6729 3938 6763
rect 3904 6661 3938 6695
rect 3904 6593 3938 6627
rect 3904 6525 3938 6559
rect 3904 6457 3938 6491
rect 3904 6389 3938 6423
rect 3904 6321 3938 6355
rect 3904 6253 3938 6287
rect 3904 6185 3938 6219
rect 3904 6117 3938 6151
rect 3904 6049 3938 6083
rect 3904 5981 3938 6015
rect 3904 5913 3938 5947
rect 1646 5819 1680 5853
rect 1646 5751 1680 5785
rect 3904 5845 3938 5879
rect 3904 5777 3938 5811
rect 1646 5683 1680 5717
rect 1646 5615 1680 5649
rect 1646 5547 1680 5581
rect 1646 5479 1680 5513
rect 1646 5411 1680 5445
rect 1646 5343 1680 5377
rect 1646 5275 1680 5309
rect 1646 5207 1680 5241
rect 1646 5139 1680 5173
rect 1646 5071 1680 5105
rect 1646 5003 1680 5037
rect 1646 4935 1680 4969
rect 1646 4867 1680 4901
rect 1646 4799 1680 4833
rect 1646 4731 1680 4765
rect 3904 5709 3938 5743
rect 3904 5641 3938 5675
rect 3904 5573 3938 5607
rect 3904 5505 3938 5539
rect 3904 5437 3938 5471
rect 3904 5369 3938 5403
rect 3904 5301 3938 5335
rect 3904 5233 3938 5267
rect 3904 5165 3938 5199
rect 3904 5097 3938 5131
rect 3904 5029 3938 5063
rect 3904 4961 3938 4995
rect 3904 4893 3938 4927
rect 3904 4825 3938 4859
rect 3904 4757 3938 4791
rect 1646 4663 1680 4697
rect 3904 4689 3938 4723
rect 1646 4595 1680 4629
rect 3904 4621 3938 4655
rect 1646 4527 1680 4561
rect 1646 4459 1680 4493
rect 1646 4391 1680 4425
rect 1646 4323 1680 4357
rect 1646 4255 1680 4289
rect 1646 4187 1680 4221
rect 1646 4119 1680 4153
rect 1646 4051 1680 4085
rect 1646 3983 1680 4017
rect 1646 3915 1680 3949
rect 1646 3847 1680 3881
rect 1646 3779 1680 3813
rect 1646 3711 1680 3745
rect 1646 3643 1680 3677
rect 1646 3575 1680 3609
rect 1646 3507 1680 3541
rect 3904 4553 3938 4587
rect 3904 4485 3938 4519
rect 3904 4417 3938 4451
rect 3904 4349 3938 4383
rect 3904 4281 3938 4315
rect 3904 4213 3938 4247
rect 3904 4145 3938 4179
rect 3904 4077 3938 4111
rect 3904 4009 3938 4043
rect 3904 3941 3938 3975
rect 3904 3873 3938 3907
rect 3904 3805 3938 3839
rect 3904 3737 3938 3771
rect 3904 3669 3938 3703
rect 3904 3601 3938 3635
rect 3904 3533 3938 3567
rect 1646 3439 1680 3473
rect 1646 3371 1680 3405
rect 1646 3303 1680 3337
rect 1646 3235 1680 3269
rect 1646 3167 1680 3201
rect 1646 3099 1680 3133
rect 1646 3031 1680 3065
rect 1646 2963 1680 2997
rect 1646 2895 1680 2929
rect 1646 2827 1680 2861
rect 1646 2759 1680 2793
rect 1646 2691 1680 2725
rect 1646 2623 1680 2657
rect 1646 2555 1680 2589
rect 1646 2487 1680 2521
rect 1646 2419 1680 2453
rect 3904 3243 3938 3277
rect 3904 3175 3938 3209
rect 3904 3107 3938 3141
rect 3904 3039 3938 3073
rect 3904 2971 3938 3005
rect 3904 2903 3938 2937
rect 3904 2835 3938 2869
rect 3904 2767 3938 2801
rect 3904 2699 3938 2733
rect 3904 2631 3938 2665
rect 3904 2563 3938 2597
rect 3904 2495 3938 2529
rect 3904 2427 3938 2461
rect 3904 2359 3938 2393
rect 1679 2258 1713 2292
rect 1747 2258 1781 2292
rect 1815 2258 1849 2292
rect 1883 2258 1917 2292
rect 1951 2258 1985 2292
rect 2019 2258 2053 2292
rect 2087 2258 2121 2292
rect 2155 2258 2189 2292
rect 2223 2258 2257 2292
rect 2291 2258 2325 2292
rect 2359 2258 2393 2292
rect 2427 2258 2461 2292
rect 2495 2258 2529 2292
rect 2563 2258 2597 2292
rect 2631 2258 2665 2292
rect 2699 2258 2733 2292
rect 2767 2258 2801 2292
rect 2835 2258 2869 2292
rect 2903 2258 2937 2292
rect 2971 2258 3005 2292
rect 3039 2258 3073 2292
rect 3107 2258 3141 2292
rect 3175 2258 3209 2292
rect 3243 2258 3277 2292
rect 3311 2258 3345 2292
rect 3379 2258 3413 2292
rect 3447 2258 3481 2292
rect 3515 2258 3549 2292
rect 3583 2258 3617 2292
rect 3651 2258 3685 2292
rect 3719 2258 3753 2292
rect 3787 2258 3821 2292
rect 3904 2291 3938 2325
<< mvnsubdiffcont >>
rect 42 10878 76 10912
rect 110 10878 144 10912
rect 178 10878 212 10912
rect 246 10878 280 10912
rect 314 10878 348 10912
rect 382 10878 416 10912
rect 450 10878 484 10912
rect 518 10878 552 10912
rect 586 10878 620 10912
rect 654 10878 688 10912
rect 722 10878 756 10912
rect 790 10878 824 10912
rect 858 10878 892 10912
rect 926 10878 960 10912
rect 994 10878 1028 10912
rect 1062 10878 1096 10912
rect 1130 10878 1164 10912
rect 1198 10878 1232 10912
rect 1266 10878 1300 10912
rect 1334 10878 1368 10912
rect 9 10755 43 10789
rect 9 10687 43 10721
rect 1457 10845 1491 10879
rect 1582 10878 1616 10912
rect 1650 10878 1684 10912
rect 1718 10878 1752 10912
rect 1786 10878 1820 10912
rect 1854 10878 1888 10912
rect 1922 10878 1956 10912
rect 1990 10878 2024 10912
rect 2058 10878 2092 10912
rect 2126 10878 2160 10912
rect 2194 10878 2228 10912
rect 2262 10878 2296 10912
rect 2330 10878 2364 10912
rect 2398 10878 2432 10912
rect 2466 10878 2500 10912
rect 2534 10878 2568 10912
rect 2602 10878 2636 10912
rect 2670 10878 2704 10912
rect 2738 10878 2772 10912
rect 2806 10878 2840 10912
rect 2874 10878 2908 10912
rect 2942 10878 2976 10912
rect 3010 10878 3044 10912
rect 3078 10878 3112 10912
rect 3146 10878 3180 10912
rect 3214 10878 3248 10912
rect 3282 10878 3316 10912
rect 3350 10878 3384 10912
rect 3418 10878 3452 10912
rect 3486 10878 3520 10912
rect 3554 10878 3588 10912
rect 3622 10878 3656 10912
rect 3690 10878 3724 10912
rect 3758 10878 3792 10912
rect 3826 10878 3860 10912
rect 3894 10878 3928 10912
rect 3962 10878 3996 10912
rect 4030 10878 4064 10912
rect 4098 10878 4132 10912
rect 4166 10878 4200 10912
rect 4234 10878 4268 10912
rect 4302 10878 4336 10912
rect 4370 10878 4404 10912
rect 4438 10878 4472 10912
rect 4506 10878 4540 10912
rect 4574 10878 4608 10912
rect 4642 10878 4676 10912
rect 4710 10878 4744 10912
rect 4778 10878 4812 10912
rect 4846 10878 4880 10912
rect 4914 10878 4948 10912
rect 4982 10878 5016 10912
rect 5050 10878 5084 10912
rect 5118 10878 5152 10912
rect 5186 10878 5220 10912
rect 5254 10878 5288 10912
rect 5322 10878 5356 10912
rect 5390 10878 5424 10912
rect 5458 10878 5492 10912
rect 5526 10878 5560 10912
rect 5594 10878 5628 10912
rect 5662 10878 5696 10912
rect 5730 10878 5764 10912
rect 5798 10878 5832 10912
rect 5866 10878 5900 10912
rect 5934 10878 5968 10912
rect 6002 10878 6036 10912
rect 6070 10878 6104 10912
rect 6138 10878 6172 10912
rect 6206 10878 6240 10912
rect 6274 10878 6308 10912
rect 6342 10878 6376 10912
rect 6410 10878 6444 10912
rect 6478 10878 6512 10912
rect 6546 10878 6580 10912
rect 6614 10878 6648 10912
rect 6682 10878 6716 10912
rect 6750 10878 6784 10912
rect 6818 10878 6852 10912
rect 6886 10878 6920 10912
rect 6954 10878 6988 10912
rect 7022 10878 7056 10912
rect 7090 10878 7124 10912
rect 7158 10878 7192 10912
rect 7226 10878 7260 10912
rect 7294 10878 7328 10912
rect 7362 10878 7396 10912
rect 7430 10878 7464 10912
rect 7498 10878 7532 10912
rect 7566 10878 7600 10912
rect 7634 10878 7668 10912
rect 7702 10878 7736 10912
rect 7770 10878 7804 10912
rect 7838 10878 7872 10912
rect 7906 10878 7940 10912
rect 7974 10878 8008 10912
rect 8042 10878 8076 10912
rect 8110 10878 8144 10912
rect 8178 10878 8212 10912
rect 8246 10878 8280 10912
rect 8314 10878 8348 10912
rect 8382 10878 8416 10912
rect 1457 10777 1491 10811
rect 1457 10709 1491 10743
rect 8415 10785 8449 10819
rect 9 10619 43 10653
rect 9 10551 43 10585
rect 9 10483 43 10517
rect 9 10415 43 10449
rect 9 10347 43 10381
rect 9 10279 43 10313
rect 9 10211 43 10245
rect 9 10143 43 10177
rect 9 10075 43 10109
rect 9 10007 43 10041
rect 9 9939 43 9973
rect 9 9871 43 9905
rect 9 9803 43 9837
rect 9 9735 43 9769
rect 9 9667 43 9701
rect 9 9599 43 9633
rect 9 9531 43 9565
rect 9 9463 43 9497
rect 9 9395 43 9429
rect 9 9327 43 9361
rect 9 9259 43 9293
rect 9 9191 43 9225
rect 9 9123 43 9157
rect 9 9055 43 9089
rect 9 8987 43 9021
rect 9 8919 43 8953
rect 9 8851 43 8885
rect 9 8783 43 8817
rect 9 8715 43 8749
rect 9 8647 43 8681
rect 9 8579 43 8613
rect 9 8511 43 8545
rect 9 8443 43 8477
rect 9 8375 43 8409
rect 9 8307 43 8341
rect 9 8239 43 8273
rect 9 8171 43 8205
rect 9 8103 43 8137
rect 9 8035 43 8069
rect 9 7967 43 8001
rect 9 7899 43 7933
rect 9 7831 43 7865
rect 9 7763 43 7797
rect 9 7695 43 7729
rect 9 7627 43 7661
rect 9 7559 43 7593
rect 9 7491 43 7525
rect 9 7423 43 7457
rect 9 7355 43 7389
rect 9 7287 43 7321
rect 9 7219 43 7253
rect 9 7151 43 7185
rect 9 7083 43 7117
rect 9 7015 43 7049
rect 9 6947 43 6981
rect 9 6879 43 6913
rect 9 6811 43 6845
rect 9 6743 43 6777
rect 9 6675 43 6709
rect 9 6607 43 6641
rect 9 6539 43 6573
rect 9 6471 43 6505
rect 9 6403 43 6437
rect 9 6335 43 6369
rect 9 6267 43 6301
rect 9 6199 43 6233
rect 9 6131 43 6165
rect 9 6063 43 6097
rect 9 5995 43 6029
rect 9 5927 43 5961
rect 9 5859 43 5893
rect 9 5791 43 5825
rect 9 5723 43 5757
rect 9 5655 43 5689
rect 9 5587 43 5621
rect 9 5519 43 5553
rect 9 5451 43 5485
rect 9 5383 43 5417
rect 9 5315 43 5349
rect 9 5247 43 5281
rect 9 5179 43 5213
rect 9 5111 43 5145
rect 9 5043 43 5077
rect 9 4975 43 5009
rect 9 4907 43 4941
rect 9 4839 43 4873
rect 9 4771 43 4805
rect 9 4703 43 4737
rect 9 4635 43 4669
rect 9 4567 43 4601
rect 9 4499 43 4533
rect 9 4431 43 4465
rect 9 4363 43 4397
rect 9 4295 43 4329
rect 9 4227 43 4261
rect 9 4159 43 4193
rect 9 4091 43 4125
rect 9 4023 43 4057
rect 9 3955 43 3989
rect 9 3887 43 3921
rect 9 3819 43 3853
rect 9 3751 43 3785
rect 9 3683 43 3717
rect 9 3615 43 3649
rect 9 3547 43 3581
rect 9 3479 43 3513
rect 9 3411 43 3445
rect 9 3343 43 3377
rect 9 3275 43 3309
rect 9 3207 43 3241
rect 9 3139 43 3173
rect 9 3071 43 3105
rect 9 3003 43 3037
rect 9 2935 43 2969
rect 9 2867 43 2901
rect 9 2799 43 2833
rect 9 2731 43 2765
rect 9 2663 43 2697
rect 9 2595 43 2629
rect 9 2527 43 2561
rect 9 2459 43 2493
rect 9 2391 43 2425
rect 9 2323 43 2357
rect 9 2255 43 2289
rect 9 2187 43 2221
rect 9 2119 43 2153
rect 9 2051 43 2085
rect 9 1983 43 2017
rect 9 1915 43 1949
rect 9 1847 43 1881
rect 9 1779 43 1813
rect 9 1711 43 1745
rect 9 1643 43 1677
rect 9 1575 43 1609
rect 9 1507 43 1541
rect 9 1439 43 1473
rect 9 1371 43 1405
rect 9 1303 43 1337
rect 9 1235 43 1269
rect 9 1167 43 1201
rect 9 1099 43 1133
rect 9 1031 43 1065
rect 9 963 43 997
rect 9 895 43 929
rect 9 827 43 861
rect 9 759 43 793
rect 9 691 43 725
rect 9 623 43 657
rect 9 555 43 589
rect 1457 10641 1491 10675
rect 1457 10573 1491 10607
rect 1457 10505 1491 10539
rect 1457 10437 1491 10471
rect 1457 10369 1491 10403
rect 1457 10301 1491 10335
rect 1457 10233 1491 10267
rect 1457 10165 1491 10199
rect 1457 10097 1491 10131
rect 1457 10029 1491 10063
rect 1457 9961 1491 9995
rect 1457 9893 1491 9927
rect 1457 9825 1491 9859
rect 1457 9757 1491 9791
rect 1457 9689 1491 9723
rect 1457 9621 1491 9655
rect 1457 9553 1491 9587
rect 1457 9485 1491 9519
rect 1457 9417 1491 9451
rect 1457 9349 1491 9383
rect 1457 9281 1491 9315
rect 1457 9213 1491 9247
rect 1457 9145 1491 9179
rect 1457 9077 1491 9111
rect 1457 9009 1491 9043
rect 1457 8941 1491 8975
rect 1457 8873 1491 8907
rect 1457 8805 1491 8839
rect 1457 8737 1491 8771
rect 1457 8669 1491 8703
rect 1457 8601 1491 8635
rect 1457 8533 1491 8567
rect 1457 8465 1491 8499
rect 1457 8397 1491 8431
rect 1457 8329 1491 8363
rect 1457 8261 1491 8295
rect 1457 8193 1491 8227
rect 1457 8125 1491 8159
rect 1457 8057 1491 8091
rect 1457 7989 1491 8023
rect 1457 7921 1491 7955
rect 1457 7853 1491 7887
rect 1457 7785 1491 7819
rect 1457 7717 1491 7751
rect 1457 7649 1491 7683
rect 1457 7581 1491 7615
rect 1457 7513 1491 7547
rect 1457 7445 1491 7479
rect 8415 10717 8449 10751
rect 8415 10649 8449 10683
rect 8415 10581 8449 10615
rect 8415 10513 8449 10547
rect 8415 10445 8449 10479
rect 8415 10377 8449 10411
rect 8415 10309 8449 10343
rect 8415 10241 8449 10275
rect 8415 10173 8449 10207
rect 8415 10105 8449 10139
rect 8415 10037 8449 10071
rect 8415 9969 8449 10003
rect 8415 9901 8449 9935
rect 8415 9833 8449 9867
rect 8415 9765 8449 9799
rect 8415 9697 8449 9731
rect 8415 9629 8449 9663
rect 8415 9561 8449 9595
rect 8415 9493 8449 9527
rect 8415 9425 8449 9459
rect 8415 9357 8449 9391
rect 8415 9289 8449 9323
rect 8415 9221 8449 9255
rect 8415 9153 8449 9187
rect 8415 9085 8449 9119
rect 8415 9017 8449 9051
rect 8415 8949 8449 8983
rect 8415 8881 8449 8915
rect 8415 8813 8449 8847
rect 8415 8745 8449 8779
rect 8415 8643 8449 8677
rect 1490 7287 1524 7321
rect 1558 7287 1592 7321
rect 1626 7287 1660 7321
rect 1694 7287 1728 7321
rect 1762 7287 1796 7321
rect 1830 7287 1864 7321
rect 1898 7287 1932 7321
rect 1966 7287 2000 7321
rect 2034 7287 2068 7321
rect 2102 7287 2136 7321
rect 2170 7287 2204 7321
rect 2238 7287 2272 7321
rect 2306 7287 2340 7321
rect 2374 7287 2408 7321
rect 2442 7287 2476 7321
rect 2510 7287 2544 7321
rect 2578 7287 2612 7321
rect 2646 7287 2680 7321
rect 2714 7287 2748 7321
rect 2782 7287 2816 7321
rect 2850 7287 2884 7321
rect 2918 7287 2952 7321
rect 2986 7287 3020 7321
rect 3054 7287 3088 7321
rect 3122 7287 3156 7321
rect 3190 7287 3224 7321
rect 3258 7287 3292 7321
rect 3326 7287 3360 7321
rect 3394 7287 3428 7321
rect 3462 7287 3496 7321
rect 3530 7287 3564 7321
rect 3598 7287 3632 7321
rect 3666 7287 3700 7321
rect 3734 7287 3768 7321
rect 3802 7287 3836 7321
rect 3870 7287 3904 7321
rect 3938 7287 3972 7321
rect 4006 7287 4040 7321
rect 1457 7218 1491 7252
rect 1457 7150 1491 7184
rect 1457 7082 1491 7116
rect 4093 7192 4127 7226
rect 4093 7124 4127 7158
rect 1457 7014 1491 7048
rect 1457 6946 1491 6980
rect 1457 6878 1491 6912
rect 1457 6810 1491 6844
rect 1457 6742 1491 6776
rect 1457 6674 1491 6708
rect 1457 6606 1491 6640
rect 1457 6538 1491 6572
rect 1457 6470 1491 6504
rect 1457 6402 1491 6436
rect 1457 6334 1491 6368
rect 1457 6266 1491 6300
rect 1457 6198 1491 6232
rect 1457 6130 1491 6164
rect 1457 6062 1491 6096
rect 1457 5994 1491 6028
rect 1457 5926 1491 5960
rect 1457 5858 1491 5892
rect 1457 5790 1491 5824
rect 1457 5722 1491 5756
rect 1457 5654 1491 5688
rect 1457 5586 1491 5620
rect 1457 5518 1491 5552
rect 1457 5450 1491 5484
rect 1457 5382 1491 5416
rect 1457 5314 1491 5348
rect 1457 5246 1491 5280
rect 1457 5178 1491 5212
rect 1457 5110 1491 5144
rect 1457 5042 1491 5076
rect 1457 4974 1491 5008
rect 1457 4906 1491 4940
rect 1457 4838 1491 4872
rect 1457 4770 1491 4804
rect 1457 4702 1491 4736
rect 1457 4634 1491 4668
rect 1457 4566 1491 4600
rect 1457 4498 1491 4532
rect 1457 4430 1491 4464
rect 1457 4362 1491 4396
rect 1457 4294 1491 4328
rect 1457 4226 1491 4260
rect 1457 4158 1491 4192
rect 1457 4090 1491 4124
rect 1457 4022 1491 4056
rect 1457 3954 1491 3988
rect 1457 3886 1491 3920
rect 1457 3818 1491 3852
rect 1457 3750 1491 3784
rect 1457 3682 1491 3716
rect 1457 3614 1491 3648
rect 1457 3546 1491 3580
rect 1457 3478 1491 3512
rect 1457 3410 1491 3444
rect 1457 3342 1491 3376
rect 1457 3274 1491 3308
rect 1457 3206 1491 3240
rect 1457 3138 1491 3172
rect 1457 3070 1491 3104
rect 1457 3002 1491 3036
rect 1457 2934 1491 2968
rect 1457 2866 1491 2900
rect 1457 2798 1491 2832
rect 1457 2730 1491 2764
rect 1457 2662 1491 2696
rect 1457 2594 1491 2628
rect 1457 2526 1491 2560
rect 1457 2458 1491 2492
rect 1457 2390 1491 2424
rect 1457 2322 1491 2356
rect 1457 2254 1491 2288
rect 4093 7056 4127 7090
rect 4093 6988 4127 7022
rect 4093 6920 4127 6954
rect 4093 6852 4127 6886
rect 4093 6784 4127 6818
rect 4093 6716 4127 6750
rect 4093 6648 4127 6682
rect 4093 6580 4127 6614
rect 4093 6512 4127 6546
rect 4093 6444 4127 6478
rect 4093 6376 4127 6410
rect 4093 6308 4127 6342
rect 4093 6240 4127 6274
rect 4093 6172 4127 6206
rect 4093 6104 4127 6138
rect 4093 6036 4127 6070
rect 4093 5968 4127 6002
rect 4093 5900 4127 5934
rect 4093 5832 4127 5866
rect 4093 5764 4127 5798
rect 4093 5696 4127 5730
rect 4093 5628 4127 5662
rect 4093 5560 4127 5594
rect 4093 5492 4127 5526
rect 4093 5424 4127 5458
rect 4093 5356 4127 5390
rect 4093 5288 4127 5322
rect 4093 5220 4127 5254
rect 4093 5152 4127 5186
rect 4093 5084 4127 5118
rect 4093 5016 4127 5050
rect 4093 4948 4127 4982
rect 4093 4880 4127 4914
rect 4093 4812 4127 4846
rect 4093 4744 4127 4778
rect 4093 4676 4127 4710
rect 4093 4608 4127 4642
rect 4093 4540 4127 4574
rect 4093 4472 4127 4506
rect 4093 4404 4127 4438
rect 4093 4336 4127 4370
rect 4093 4268 4127 4302
rect 4093 4200 4127 4234
rect 4093 4132 4127 4166
rect 4093 4064 4127 4098
rect 4093 3996 4127 4030
rect 4093 3928 4127 3962
rect 4093 3860 4127 3894
rect 4093 3792 4127 3826
rect 4093 3724 4127 3758
rect 4093 3656 4127 3690
rect 4093 3588 4127 3622
rect 4093 3520 4127 3554
rect 4093 3452 4127 3486
rect 4093 3384 4127 3418
rect 4093 3316 4127 3350
rect 4093 3248 4127 3282
rect 4093 3180 4127 3214
rect 4093 3112 4127 3146
rect 4093 3044 4127 3078
rect 4093 2976 4127 3010
rect 4093 2908 4127 2942
rect 4093 2840 4127 2874
rect 4093 2772 4127 2806
rect 4093 2704 4127 2738
rect 4093 2636 4127 2670
rect 4093 2568 4127 2602
rect 4093 2500 4127 2534
rect 4093 2432 4127 2466
rect 4093 2364 4127 2398
rect 4093 2296 4127 2330
rect 1457 2186 1491 2220
rect 1457 2118 1491 2152
rect 4093 2228 4127 2262
rect 4093 2160 4127 2194
rect 1526 2069 1560 2103
rect 1594 2069 1628 2103
rect 1662 2069 1696 2103
rect 1730 2069 1764 2103
rect 1798 2069 1832 2103
rect 1866 2069 1900 2103
rect 1934 2069 1968 2103
rect 2002 2069 2036 2103
rect 2070 2069 2104 2103
rect 2138 2069 2172 2103
rect 2206 2069 2240 2103
rect 2274 2069 2308 2103
rect 2342 2069 2376 2103
rect 2410 2069 2444 2103
rect 2478 2069 2512 2103
rect 2546 2069 2580 2103
rect 2614 2069 2648 2103
rect 2682 2069 2716 2103
rect 2750 2069 2784 2103
rect 2818 2069 2852 2103
rect 2886 2069 2920 2103
rect 2954 2069 2988 2103
rect 3022 2069 3056 2103
rect 3090 2069 3124 2103
rect 3158 2069 3192 2103
rect 3226 2069 3260 2103
rect 3294 2069 3328 2103
rect 3362 2069 3396 2103
rect 3430 2069 3464 2103
rect 3498 2069 3532 2103
rect 3566 2069 3600 2103
rect 3634 2069 3668 2103
rect 3702 2069 3736 2103
rect 3770 2069 3804 2103
rect 3838 2069 3872 2103
rect 3906 2069 3940 2103
rect 3974 2069 4008 2103
rect 4093 2092 4127 2126
rect 4093 2024 4127 2058
rect 1457 1806 1491 1840
rect 1457 1738 1491 1772
rect 1457 1670 1491 1704
rect 1457 1602 1491 1636
rect 1457 1534 1491 1568
rect 1457 1466 1491 1500
rect 1457 1398 1491 1432
rect 1457 1330 1491 1364
rect 1457 1262 1491 1296
rect 1457 1194 1491 1228
rect 1457 1126 1491 1160
rect 1457 1058 1491 1092
rect 1457 990 1491 1024
rect 1457 922 1491 956
rect 1457 854 1491 888
rect 1457 786 1491 820
rect 1457 718 1491 752
rect 1457 650 1491 684
rect 1457 582 1491 616
rect 1457 514 1491 548
rect 4093 1956 4127 1990
rect 4093 1888 4127 1922
rect 4093 1820 4127 1854
rect 4093 1752 4127 1786
rect 4093 1684 4127 1718
rect 4093 1616 4127 1650
rect 4093 1548 4127 1582
rect 4093 1480 4127 1514
rect 4093 1412 4127 1446
rect 4093 1344 4127 1378
rect 4093 1276 4127 1310
rect 4093 1208 4127 1242
rect 4093 1140 4127 1174
rect 4093 1072 4127 1106
rect 4093 1004 4127 1038
rect 4093 936 4127 970
rect 4093 868 4127 902
rect 4093 800 4127 834
rect 4093 732 4127 766
rect 4093 664 4127 698
rect 4093 596 4127 630
rect 4093 528 4127 562
rect 9 413 43 447
rect 1300 427 1334 461
rect 1368 427 1402 461
rect 1490 427 1524 461
rect 1558 427 1592 461
rect 1626 427 1660 461
rect 1694 427 1728 461
rect 1762 427 1796 461
rect 1830 427 1864 461
rect 1898 427 1932 461
rect 1966 427 2000 461
rect 2034 427 2068 461
rect 2102 427 2136 461
rect 2170 427 2204 461
rect 2238 427 2272 461
rect 2306 427 2340 461
rect 2374 427 2408 461
rect 2442 427 2476 461
rect 2510 427 2544 461
rect 2578 427 2612 461
rect 2646 427 2680 461
rect 2714 427 2748 461
rect 2782 427 2816 461
rect 2850 427 2884 461
rect 2918 427 2952 461
rect 2986 427 3020 461
rect 3054 427 3088 461
rect 3122 427 3156 461
rect 3190 427 3224 461
rect 3258 427 3292 461
rect 3326 427 3360 461
rect 3394 427 3428 461
rect 3462 427 3496 461
rect 3530 427 3564 461
rect 3598 427 3632 461
rect 3666 427 3700 461
rect 3734 427 3768 461
rect 3802 427 3836 461
rect 3870 427 3904 461
rect 3938 427 3972 461
rect 4006 427 4040 461
rect 4093 460 4127 494
<< poly >>
rect 1757 9761 1821 10561
rect 3871 9761 3949 10561
rect 6001 9761 6079 10561
rect 8131 9761 8193 10561
rect 1757 8905 1821 9705
rect 6001 8905 6079 9705
rect 8131 8905 8193 9705
rect 1808 8692 2104 8708
rect 1808 8658 1824 8692
rect 1858 8658 1892 8692
rect 1926 8658 1986 8692
rect 2020 8658 2054 8692
rect 2088 8658 2104 8692
rect 1808 8642 2104 8658
rect 2160 8692 2360 8708
rect 2160 8658 2209 8692
rect 2243 8658 2277 8692
rect 2311 8658 2360 8692
rect 2160 8636 2360 8658
rect 2416 8692 2616 8708
rect 2416 8658 2465 8692
rect 2499 8658 2533 8692
rect 2567 8658 2616 8692
rect 2416 8636 2616 8658
rect 2672 8692 2872 8708
rect 2672 8658 2721 8692
rect 2755 8658 2789 8692
rect 2823 8658 2872 8692
rect 2672 8636 2872 8658
rect 2928 8692 3128 8708
rect 2928 8658 2977 8692
rect 3011 8658 3045 8692
rect 3079 8658 3128 8692
rect 2928 8636 3128 8658
rect 3184 8692 3384 8708
rect 3184 8658 3233 8692
rect 3267 8658 3301 8692
rect 3335 8658 3384 8692
rect 3184 8636 3384 8658
rect 3440 8692 3640 8708
rect 3440 8658 3489 8692
rect 3523 8658 3557 8692
rect 3591 8658 3640 8692
rect 3440 8636 3640 8658
rect 3696 8692 3896 8708
rect 3696 8658 3745 8692
rect 3779 8658 3813 8692
rect 3847 8658 3896 8692
rect 3696 8636 3896 8658
rect 3952 8692 4152 8708
rect 3952 8658 4001 8692
rect 4035 8658 4069 8692
rect 4103 8658 4152 8692
rect 4208 8692 4328 8708
rect 4208 8662 4251 8692
rect 3952 8636 4152 8658
rect 4235 8658 4251 8662
rect 4285 8662 4328 8692
rect 4285 8658 4301 8662
rect 4235 8642 4301 8658
rect 1774 7025 1908 7041
rect 1774 6991 1790 7025
rect 1824 6991 1858 7025
rect 1892 6991 1908 7025
rect 1774 6975 1908 6991
rect 1964 6969 2764 7041
rect 2820 6969 3620 7041
rect 3676 7025 3810 7041
rect 3676 6991 3692 7025
rect 3726 6991 3760 7025
rect 3794 6991 3810 7025
rect 3676 6975 3810 6991
rect 1808 5849 1908 5891
rect 3676 5849 3776 5891
rect 1774 5833 1908 5849
rect 1774 5799 1790 5833
rect 1824 5799 1858 5833
rect 1892 5799 1908 5833
rect 1774 5783 1908 5799
rect 1964 5777 2764 5849
rect 2820 5777 3620 5849
rect 3676 5833 3810 5849
rect 3676 5799 3692 5833
rect 3726 5799 3760 5833
rect 3794 5799 3810 5833
rect 3676 5783 3810 5799
rect 1808 4657 1908 4699
rect 3676 4657 3776 4699
rect 1774 4641 1908 4657
rect 1774 4607 1790 4641
rect 1824 4607 1858 4641
rect 1892 4607 1908 4641
rect 1774 4591 1908 4607
rect 1964 4585 2764 4657
rect 2820 4585 3620 4657
rect 3676 4641 3810 4657
rect 3676 4607 3692 4641
rect 3726 4607 3760 4641
rect 3794 4607 3810 4641
rect 3676 4591 3810 4607
rect 1808 3465 1908 3507
rect 1774 3449 1908 3465
rect 1774 3415 1790 3449
rect 1824 3415 1858 3449
rect 1892 3415 1908 3449
rect 1774 3399 1908 3415
rect 1964 3393 2764 3465
rect 2820 3393 3620 3465
rect 3676 3449 3810 3465
rect 3676 3415 3692 3449
rect 3726 3415 3760 3449
rect 3794 3415 3810 3449
rect 3676 3399 3810 3415
rect 1652 2018 1852 2034
rect 1652 1984 1668 2018
rect 1702 1984 1736 2018
rect 1770 1984 1852 2018
rect 1652 1968 1852 1984
rect 1908 2018 2308 2034
rect 1908 1984 1955 2018
rect 1989 1984 2023 2018
rect 2057 1984 2091 2018
rect 2125 1984 2159 2018
rect 2193 1984 2227 2018
rect 2261 1984 2308 2018
rect 1908 1968 2308 1984
rect 2364 2018 2764 2034
rect 2364 1984 2411 2018
rect 2445 1984 2479 2018
rect 2513 1984 2547 2018
rect 2581 1984 2615 2018
rect 2649 1984 2683 2018
rect 2717 1984 2764 2018
rect 2364 1968 2764 1984
rect 2820 2018 3220 2034
rect 2820 1984 2867 2018
rect 2901 1984 2935 2018
rect 2969 1984 3003 2018
rect 3037 1984 3071 2018
rect 3105 1984 3139 2018
rect 3173 1984 3220 2018
rect 2820 1968 3220 1984
rect 3276 2018 3676 2034
rect 3276 1984 3323 2018
rect 3357 1984 3391 2018
rect 3425 1984 3459 2018
rect 3493 1984 3527 2018
rect 3561 1984 3595 2018
rect 3629 1984 3676 2018
rect 3276 1968 3676 1984
rect 3732 2018 3932 2034
rect 3732 1984 3814 2018
rect 3848 1984 3882 2018
rect 3916 1984 3932 2018
rect 3732 1968 3932 1984
<< polycont >>
rect 1824 8658 1858 8692
rect 1892 8658 1926 8692
rect 1986 8658 2020 8692
rect 2054 8658 2088 8692
rect 2209 8658 2243 8692
rect 2277 8658 2311 8692
rect 2465 8658 2499 8692
rect 2533 8658 2567 8692
rect 2721 8658 2755 8692
rect 2789 8658 2823 8692
rect 2977 8658 3011 8692
rect 3045 8658 3079 8692
rect 3233 8658 3267 8692
rect 3301 8658 3335 8692
rect 3489 8658 3523 8692
rect 3557 8658 3591 8692
rect 3745 8658 3779 8692
rect 3813 8658 3847 8692
rect 4001 8658 4035 8692
rect 4069 8658 4103 8692
rect 4251 8658 4285 8692
rect 1790 6991 1824 7025
rect 1858 6991 1892 7025
rect 3692 6991 3726 7025
rect 3760 6991 3794 7025
rect 1790 5799 1824 5833
rect 1858 5799 1892 5833
rect 3692 5799 3726 5833
rect 3760 5799 3794 5833
rect 1790 4607 1824 4641
rect 1858 4607 1892 4641
rect 3692 4607 3726 4641
rect 3760 4607 3794 4641
rect 1790 3415 1824 3449
rect 1858 3415 1892 3449
rect 3692 3415 3726 3449
rect 3760 3415 3794 3449
rect 1668 1984 1702 2018
rect 1736 1984 1770 2018
rect 1955 1984 1989 2018
rect 2023 1984 2057 2018
rect 2091 1984 2125 2018
rect 2159 1984 2193 2018
rect 2227 1984 2261 2018
rect 2411 1984 2445 2018
rect 2479 1984 2513 2018
rect 2547 1984 2581 2018
rect 2615 1984 2649 2018
rect 2683 1984 2717 2018
rect 2867 1984 2901 2018
rect 2935 1984 2969 2018
rect 3003 1984 3037 2018
rect 3071 1984 3105 2018
rect 3139 1984 3173 2018
rect 3323 1984 3357 2018
rect 3391 1984 3425 2018
rect 3459 1984 3493 2018
rect 3527 1984 3561 2018
rect 3595 1984 3629 2018
rect 3814 1984 3848 2018
rect 3882 1984 3916 2018
<< locali >>
rect 8 10912 8450 10913
rect 8 10878 42 10912
rect 76 10878 110 10912
rect 144 10878 178 10912
rect 212 10878 246 10912
rect 280 10878 314 10912
rect 348 10878 382 10912
rect 416 10878 450 10912
rect 484 10878 518 10912
rect 552 10878 586 10912
rect 620 10878 654 10912
rect 688 10878 722 10912
rect 756 10878 790 10912
rect 824 10878 858 10912
rect 892 10878 926 10912
rect 960 10878 994 10912
rect 1028 10878 1062 10912
rect 1096 10878 1130 10912
rect 1164 10878 1198 10912
rect 1232 10878 1266 10912
rect 1300 10878 1334 10912
rect 1368 10879 1582 10912
rect 1368 10878 1457 10879
rect 8 10877 1457 10878
rect 8 10872 61 10877
rect 1391 10872 1457 10877
rect 8 10789 44 10872
rect 8 10755 9 10789
rect 43 10755 44 10789
rect 8 10721 44 10755
rect 1456 10845 1457 10872
rect 1491 10878 1582 10879
rect 1616 10878 1650 10912
rect 1684 10878 1718 10912
rect 1752 10878 1786 10912
rect 1820 10878 1854 10912
rect 1888 10878 1922 10912
rect 1956 10878 1990 10912
rect 2024 10878 2058 10912
rect 2092 10878 2126 10912
rect 2160 10878 2194 10912
rect 2228 10878 2262 10912
rect 2296 10878 2330 10912
rect 2364 10878 2398 10912
rect 2432 10878 2466 10912
rect 2500 10878 2534 10912
rect 2568 10878 2602 10912
rect 2636 10878 2670 10912
rect 2704 10878 2738 10912
rect 2772 10878 2806 10912
rect 2840 10878 2874 10912
rect 2908 10878 2942 10912
rect 2976 10878 3010 10912
rect 3044 10878 3078 10912
rect 3112 10878 3146 10912
rect 3180 10878 3214 10912
rect 3248 10878 3282 10912
rect 3316 10878 3350 10912
rect 3384 10878 3418 10912
rect 3452 10878 3486 10912
rect 3520 10878 3554 10912
rect 3588 10878 3622 10912
rect 3656 10878 3690 10912
rect 3724 10878 3758 10912
rect 3792 10878 3826 10912
rect 3860 10878 3894 10912
rect 3928 10878 3962 10912
rect 3996 10878 4030 10912
rect 4064 10878 4098 10912
rect 4132 10878 4166 10912
rect 4200 10878 4234 10912
rect 4268 10878 4302 10912
rect 4336 10878 4370 10912
rect 4404 10878 4438 10912
rect 4472 10878 4506 10912
rect 4540 10878 4574 10912
rect 4608 10878 4642 10912
rect 4676 10878 4710 10912
rect 4744 10878 4778 10912
rect 4812 10878 4846 10912
rect 4880 10878 4914 10912
rect 4948 10878 4982 10912
rect 5016 10878 5050 10912
rect 5084 10878 5118 10912
rect 5152 10878 5186 10912
rect 5220 10878 5254 10912
rect 5288 10878 5322 10912
rect 5356 10878 5390 10912
rect 5424 10878 5458 10912
rect 5492 10878 5526 10912
rect 5560 10878 5594 10912
rect 5628 10878 5662 10912
rect 5696 10878 5730 10912
rect 5764 10878 5798 10912
rect 5832 10878 5866 10912
rect 5900 10878 5934 10912
rect 5968 10878 6002 10912
rect 6036 10878 6070 10912
rect 6104 10878 6138 10912
rect 6172 10878 6206 10912
rect 6240 10878 6274 10912
rect 6308 10878 6342 10912
rect 6376 10878 6410 10912
rect 6444 10878 6478 10912
rect 6512 10878 6546 10912
rect 6580 10878 6614 10912
rect 6648 10878 6682 10912
rect 6716 10878 6750 10912
rect 6784 10878 6818 10912
rect 6852 10878 6886 10912
rect 6920 10878 6954 10912
rect 6988 10878 7022 10912
rect 7056 10878 7090 10912
rect 7124 10878 7158 10912
rect 7192 10878 7226 10912
rect 7260 10878 7294 10912
rect 7328 10878 7362 10912
rect 7396 10878 7430 10912
rect 7464 10878 7498 10912
rect 7532 10878 7566 10912
rect 7600 10878 7634 10912
rect 7668 10878 7702 10912
rect 7736 10878 7770 10912
rect 7804 10878 7838 10912
rect 7872 10878 7906 10912
rect 7940 10878 7974 10912
rect 8008 10878 8042 10912
rect 8076 10878 8110 10912
rect 8144 10878 8178 10912
rect 8212 10878 8246 10912
rect 8280 10878 8314 10912
rect 8348 10878 8382 10912
rect 8416 10878 8450 10912
rect 1491 10877 8450 10878
rect 1491 10872 1557 10877
rect 8376 10872 8450 10877
rect 1491 10845 1502 10872
rect 1456 10811 1502 10845
rect 1456 10777 1457 10811
rect 1491 10800 1502 10811
rect 8414 10819 8450 10872
rect 1491 10777 1492 10800
rect 1456 10743 1492 10777
rect 8 10687 9 10721
rect 43 10687 44 10721
rect 8 10653 44 10687
rect 8 10619 9 10653
rect 43 10619 44 10653
rect 8 10585 44 10619
rect 8 10551 9 10585
rect 43 10551 44 10585
rect 8 10517 44 10551
rect 8 10483 9 10517
rect 43 10483 44 10517
rect 8 10449 44 10483
rect 8 10415 9 10449
rect 43 10415 44 10449
rect 8 10381 44 10415
rect 8 10347 9 10381
rect 43 10347 44 10381
rect 8 10313 44 10347
rect 8 10279 9 10313
rect 43 10279 44 10313
rect 8 10245 44 10279
rect 8 10211 9 10245
rect 43 10211 44 10245
rect 8 10177 44 10211
rect 8 10143 9 10177
rect 43 10143 44 10177
rect 8 10109 44 10143
rect 8 10075 9 10109
rect 43 10075 44 10109
rect 8 10041 44 10075
rect 8 10007 9 10041
rect 43 10007 44 10041
rect 8 9973 44 10007
rect 8 9939 9 9973
rect 43 9939 44 9973
rect 8 9905 44 9939
rect 8 9871 9 9905
rect 43 9871 44 9905
rect 8 9837 44 9871
rect 8 9803 9 9837
rect 43 9803 44 9837
rect 8 9769 44 9803
rect 8 9735 9 9769
rect 43 9735 44 9769
rect 8 9701 44 9735
rect 8 9667 9 9701
rect 43 9667 44 9701
rect 8 9633 44 9667
rect 8 9599 9 9633
rect 43 9599 44 9633
rect 8 9565 44 9599
rect 8 9531 9 9565
rect 43 9531 44 9565
rect 8 9497 44 9531
rect 8 9463 9 9497
rect 43 9463 44 9497
rect 8 9429 44 9463
rect 8 9395 9 9429
rect 43 9395 44 9429
rect 8 9361 44 9395
rect 8 9327 9 9361
rect 43 9327 44 9361
rect 8 9293 44 9327
rect 8 9259 9 9293
rect 43 9259 44 9293
rect 8 9225 44 9259
rect 8 9191 9 9225
rect 43 9191 44 9225
rect 8 9157 44 9191
rect 8 9123 9 9157
rect 43 9123 44 9157
rect 8 9089 44 9123
rect 8 9055 9 9089
rect 43 9055 44 9089
rect 8 9021 44 9055
rect 8 8987 9 9021
rect 43 8987 44 9021
rect 8 8953 44 8987
rect 8 8919 9 8953
rect 43 8919 44 8953
rect 8 8885 44 8919
rect 8 8851 9 8885
rect 43 8851 44 8885
rect 8 8817 44 8851
rect 8 8783 9 8817
rect 43 8783 44 8817
rect 8 8749 44 8783
rect 8 8715 9 8749
rect 43 8715 44 8749
rect 8 8681 44 8715
rect 8 8647 9 8681
rect 43 8647 44 8681
rect 8 8613 44 8647
rect 8 8579 9 8613
rect 43 8579 44 8613
rect 8 8545 44 8579
rect 8 8511 9 8545
rect 43 8511 44 8545
rect 8 8477 44 8511
rect 8 8443 9 8477
rect 43 8443 44 8477
rect 8 8409 44 8443
rect 8 8375 9 8409
rect 43 8375 44 8409
rect 8 8341 44 8375
rect 8 8307 9 8341
rect 43 8307 44 8341
rect 8 8273 44 8307
rect 8 8239 9 8273
rect 43 8239 44 8273
rect 8 8205 44 8239
rect 8 8171 9 8205
rect 43 8171 44 8205
rect 8 8137 44 8171
rect 8 8103 9 8137
rect 43 8103 44 8137
rect 8 8069 44 8103
rect 8 8035 9 8069
rect 43 8035 44 8069
rect 8 8001 44 8035
rect 8 7967 9 8001
rect 43 7967 44 8001
rect 8 7933 44 7967
rect 8 7899 9 7933
rect 43 7899 44 7933
rect 8 7865 44 7899
rect 8 7831 9 7865
rect 43 7831 44 7865
rect 8 7797 44 7831
rect 8 7763 9 7797
rect 43 7763 44 7797
rect 8 7729 44 7763
rect 8 7695 9 7729
rect 43 7695 44 7729
rect 8 7661 44 7695
rect 8 7627 9 7661
rect 43 7627 44 7661
rect 8 7593 44 7627
rect 8 7559 9 7593
rect 43 7559 44 7593
rect 8 7525 44 7559
rect 8 7491 9 7525
rect 43 7491 44 7525
rect 8 7457 44 7491
rect 8 7423 9 7457
rect 43 7423 44 7457
rect 8 7389 44 7423
rect 8 7355 9 7389
rect 43 7355 44 7389
rect 8 7321 44 7355
rect 8 7287 9 7321
rect 43 7287 44 7321
rect 8 7253 44 7287
rect 8 7219 9 7253
rect 43 7219 44 7253
rect 8 7185 44 7219
rect 8 7151 9 7185
rect 43 7151 44 7185
rect 8 7117 44 7151
rect 8 7083 9 7117
rect 43 7083 44 7117
rect 8 7049 44 7083
rect 8 7015 9 7049
rect 43 7015 44 7049
rect 8 6981 44 7015
rect 8 6947 9 6981
rect 43 6947 44 6981
rect 8 6913 44 6947
rect 8 6879 9 6913
rect 43 6879 44 6913
rect 8 6845 44 6879
rect 8 6811 9 6845
rect 43 6811 44 6845
rect 8 6777 44 6811
rect 8 6743 9 6777
rect 43 6743 44 6777
rect 8 6709 44 6743
rect 8 6675 9 6709
rect 43 6675 44 6709
rect 8 6641 44 6675
rect 8 6607 9 6641
rect 43 6607 44 6641
rect 8 6573 44 6607
rect 8 6539 9 6573
rect 43 6539 44 6573
rect 8 6505 44 6539
rect 8 6471 9 6505
rect 43 6471 44 6505
rect 8 6437 44 6471
rect 8 6403 9 6437
rect 43 6403 44 6437
rect 8 6369 44 6403
rect 8 6335 9 6369
rect 43 6335 44 6369
rect 8 6301 44 6335
rect 8 6267 9 6301
rect 43 6267 44 6301
rect 8 6233 44 6267
rect 8 6199 9 6233
rect 43 6199 44 6233
rect 8 6165 44 6199
rect 8 6131 9 6165
rect 43 6131 44 6165
rect 8 6097 44 6131
rect 8 6063 9 6097
rect 43 6063 44 6097
rect 8 6029 44 6063
rect 8 5995 9 6029
rect 43 5995 44 6029
rect 8 5961 44 5995
rect 8 5927 9 5961
rect 43 5927 44 5961
rect 8 5893 44 5927
rect 8 5859 9 5893
rect 43 5859 44 5893
rect 8 5825 44 5859
rect 8 5791 9 5825
rect 43 5791 44 5825
rect 8 5757 44 5791
rect 8 5723 9 5757
rect 43 5723 44 5757
rect 8 5689 44 5723
rect 8 5655 9 5689
rect 43 5655 44 5689
rect 8 5621 44 5655
rect 8 5587 9 5621
rect 43 5587 44 5621
rect 8 5553 44 5587
rect 8 5519 9 5553
rect 43 5519 44 5553
rect 8 5485 44 5519
rect 8 5451 9 5485
rect 43 5451 44 5485
rect 8 5417 44 5451
rect 8 5383 9 5417
rect 43 5383 44 5417
rect 8 5349 44 5383
rect 8 5315 9 5349
rect 43 5315 44 5349
rect 8 5281 44 5315
rect 8 5247 9 5281
rect 43 5247 44 5281
rect 8 5213 44 5247
rect 8 5179 9 5213
rect 43 5179 44 5213
rect 8 5145 44 5179
rect 8 5111 9 5145
rect 43 5111 44 5145
rect 8 5077 44 5111
rect 8 5043 9 5077
rect 43 5043 44 5077
rect 8 5009 44 5043
rect 8 4975 9 5009
rect 43 4975 44 5009
rect 8 4941 44 4975
rect 8 4907 9 4941
rect 43 4907 44 4941
rect 8 4873 44 4907
rect 8 4839 9 4873
rect 43 4839 44 4873
rect 8 4805 44 4839
rect 8 4771 9 4805
rect 43 4771 44 4805
rect 8 4737 44 4771
rect 8 4703 9 4737
rect 43 4703 44 4737
rect 8 4669 44 4703
rect 8 4635 9 4669
rect 43 4635 44 4669
rect 8 4601 44 4635
rect 8 4567 9 4601
rect 43 4567 44 4601
rect 8 4533 44 4567
rect 8 4499 9 4533
rect 43 4499 44 4533
rect 8 4465 44 4499
rect 8 4431 9 4465
rect 43 4431 44 4465
rect 8 4397 44 4431
rect 8 4363 9 4397
rect 43 4363 44 4397
rect 8 4329 44 4363
rect 8 4295 9 4329
rect 43 4295 44 4329
rect 8 4261 44 4295
rect 8 4227 9 4261
rect 43 4227 44 4261
rect 8 4193 44 4227
rect 8 4159 9 4193
rect 43 4159 44 4193
rect 8 4125 44 4159
rect 8 4091 9 4125
rect 43 4091 44 4125
rect 8 4057 44 4091
rect 8 4023 9 4057
rect 43 4023 44 4057
rect 8 3989 44 4023
rect 8 3955 9 3989
rect 43 3955 44 3989
rect 8 3921 44 3955
rect 8 3887 9 3921
rect 43 3887 44 3921
rect 8 3853 44 3887
rect 8 3819 9 3853
rect 43 3819 44 3853
rect 8 3785 44 3819
rect 8 3751 9 3785
rect 43 3751 44 3785
rect 8 3717 44 3751
rect 8 3683 9 3717
rect 43 3683 44 3717
rect 8 3649 44 3683
rect 8 3615 9 3649
rect 43 3615 44 3649
rect 8 3581 44 3615
rect 8 3547 9 3581
rect 43 3547 44 3581
rect 8 3513 44 3547
rect 8 3479 9 3513
rect 43 3479 44 3513
rect 8 3445 44 3479
rect 8 3411 9 3445
rect 43 3411 44 3445
rect 8 3377 44 3411
rect 8 3343 9 3377
rect 43 3343 44 3377
rect 8 3309 44 3343
rect 8 3275 9 3309
rect 43 3275 44 3309
rect 8 3241 44 3275
rect 8 3207 9 3241
rect 43 3207 44 3241
rect 8 3173 44 3207
rect 8 3139 9 3173
rect 43 3139 44 3173
rect 8 3105 44 3139
rect 8 3071 9 3105
rect 43 3071 44 3105
rect 8 3037 44 3071
rect 8 3003 9 3037
rect 43 3003 44 3037
rect 8 2969 44 3003
rect 8 2935 9 2969
rect 43 2935 44 2969
rect 8 2901 44 2935
rect 8 2867 9 2901
rect 43 2867 44 2901
rect 8 2833 44 2867
rect 8 2799 9 2833
rect 43 2799 44 2833
rect 8 2765 44 2799
rect 8 2731 9 2765
rect 43 2731 44 2765
rect 8 2697 44 2731
rect 8 2663 9 2697
rect 43 2663 44 2697
rect 8 2629 44 2663
rect 8 2595 9 2629
rect 43 2595 44 2629
rect 8 2561 44 2595
rect 8 2527 9 2561
rect 43 2527 44 2561
rect 8 2493 44 2527
rect 8 2459 9 2493
rect 43 2459 44 2493
rect 8 2425 44 2459
rect 8 2391 9 2425
rect 43 2391 44 2425
rect 8 2357 44 2391
rect 8 2323 9 2357
rect 43 2323 44 2357
rect 8 2289 44 2323
rect 8 2255 9 2289
rect 43 2255 44 2289
rect 8 2221 44 2255
rect 8 2187 9 2221
rect 43 2187 44 2221
rect 8 2153 44 2187
rect 8 2119 9 2153
rect 43 2119 44 2153
rect 8 2085 44 2119
rect 8 2051 9 2085
rect 43 2051 44 2085
rect 8 2017 44 2051
rect 8 1983 9 2017
rect 43 1983 44 2017
rect 8 1949 44 1983
rect 8 1915 9 1949
rect 43 1915 44 1949
rect 8 1881 44 1915
rect 8 1847 9 1881
rect 43 1847 44 1881
rect 8 1813 44 1847
rect 8 1779 9 1813
rect 43 1779 44 1813
rect 8 1745 44 1779
rect 8 1711 9 1745
rect 43 1711 44 1745
rect 8 1677 44 1711
rect 8 1643 9 1677
rect 43 1643 44 1677
rect 8 1609 44 1643
rect 8 1575 9 1609
rect 43 1575 44 1609
rect 8 1541 44 1575
rect 8 1507 9 1541
rect 43 1507 44 1541
rect 8 1473 44 1507
rect 8 1439 9 1473
rect 43 1439 44 1473
rect 8 1405 44 1439
rect 8 1371 9 1405
rect 43 1371 44 1405
rect 8 1337 44 1371
rect 8 1303 9 1337
rect 43 1303 44 1337
rect 8 1269 44 1303
rect 8 1235 9 1269
rect 43 1235 44 1269
rect 8 1201 44 1235
rect 8 1167 9 1201
rect 43 1167 44 1201
rect 8 1133 44 1167
rect 8 1099 9 1133
rect 43 1099 44 1133
rect 8 1065 44 1099
rect 8 1031 9 1065
rect 43 1031 44 1065
rect 8 997 44 1031
rect 8 963 9 997
rect 43 963 44 997
rect 8 929 44 963
rect 8 895 9 929
rect 43 895 44 929
rect 8 861 44 895
rect 8 827 9 861
rect 43 827 44 861
rect 8 793 44 827
rect 8 759 9 793
rect 43 759 44 793
rect 8 725 44 759
rect 8 691 9 725
rect 43 691 44 725
rect 8 657 44 691
rect 8 623 9 657
rect 43 623 44 657
rect 8 589 44 623
rect 8 555 9 589
rect 43 555 44 589
rect 8 447 44 555
rect 8 413 9 447
rect 43 413 44 447
rect 197 10700 278 10724
rect 1032 10700 1113 10724
rect 197 10699 1113 10700
rect 197 10666 297 10699
rect 197 10632 198 10666
rect 232 10665 297 10666
rect 331 10665 365 10699
rect 399 10665 433 10699
rect 467 10665 501 10699
rect 535 10665 569 10699
rect 603 10665 637 10699
rect 671 10665 705 10699
rect 739 10665 773 10699
rect 807 10665 841 10699
rect 875 10665 909 10699
rect 943 10665 977 10699
rect 1011 10665 1045 10699
rect 1079 10665 1113 10699
rect 232 10664 1113 10665
rect 232 10632 233 10664
rect 197 10598 233 10632
rect 197 10564 198 10598
rect 232 10564 233 10598
rect 1077 10597 1113 10664
rect 197 10530 233 10564
rect 197 10496 198 10530
rect 232 10496 233 10530
rect 307 10536 323 10582
rect 357 10536 373 10582
rect 307 10514 373 10536
rect 433 10536 449 10582
rect 483 10536 499 10582
rect 433 10514 499 10536
rect 559 10536 575 10582
rect 609 10536 625 10582
rect 559 10514 625 10536
rect 685 10536 701 10582
rect 735 10536 751 10582
rect 685 10514 751 10536
rect 811 10536 827 10582
rect 861 10536 877 10582
rect 811 10514 877 10536
rect 937 10536 953 10582
rect 987 10536 1003 10582
rect 937 10514 1003 10536
rect 1077 10563 1078 10597
rect 1112 10563 1113 10597
rect 1077 10529 1113 10563
rect 197 10462 233 10496
rect 323 10498 357 10514
rect 197 10428 198 10462
rect 232 10428 233 10462
rect 307 10464 323 10480
rect 449 10498 483 10514
rect 357 10464 373 10480
rect 307 10452 373 10464
rect 433 10464 449 10480
rect 575 10498 609 10514
rect 483 10464 499 10480
rect 433 10452 499 10464
rect 559 10464 575 10480
rect 701 10498 735 10514
rect 609 10464 625 10480
rect 559 10452 625 10464
rect 685 10464 701 10480
rect 827 10498 861 10514
rect 735 10464 751 10480
rect 685 10452 751 10464
rect 811 10464 827 10480
rect 953 10498 987 10514
rect 861 10464 877 10480
rect 811 10452 877 10464
rect 937 10464 953 10480
rect 1077 10495 1078 10529
rect 1112 10495 1113 10529
rect 987 10464 1003 10480
rect 937 10452 1003 10464
rect 1077 10461 1113 10495
rect 197 10394 233 10428
rect 197 10360 198 10394
rect 232 10360 233 10394
rect 197 10326 233 10360
rect 197 10292 198 10326
rect 232 10292 233 10326
rect 197 10258 233 10292
rect 197 10224 198 10258
rect 232 10224 233 10258
rect 197 10190 233 10224
rect 197 10156 198 10190
rect 232 10156 233 10190
rect 197 10122 233 10156
rect 197 10088 198 10122
rect 232 10088 233 10122
rect 197 10054 233 10088
rect 197 10020 198 10054
rect 232 10020 233 10054
rect 197 9986 233 10020
rect 197 9952 198 9986
rect 232 9952 233 9986
rect 197 9918 233 9952
rect 197 9884 198 9918
rect 232 9884 233 9918
rect 197 9850 233 9884
rect 197 9816 198 9850
rect 232 9816 233 9850
rect 197 9782 233 9816
rect 197 9748 198 9782
rect 232 9748 233 9782
rect 197 9714 233 9748
rect 197 9680 198 9714
rect 232 9680 233 9714
rect 197 9646 233 9680
rect 197 9612 198 9646
rect 232 9612 233 9646
rect 197 9578 233 9612
rect 197 9544 198 9578
rect 232 9544 233 9578
rect 197 9510 233 9544
rect 197 9476 198 9510
rect 232 9476 233 9510
rect 197 9442 233 9476
rect 197 9408 198 9442
rect 232 9408 233 9442
rect 197 9374 233 9408
rect 197 9340 198 9374
rect 232 9340 233 9374
rect 197 9306 233 9340
rect 197 9272 198 9306
rect 232 9272 233 9306
rect 197 9238 233 9272
rect 197 9204 198 9238
rect 232 9204 233 9238
rect 197 9170 233 9204
rect 197 9136 198 9170
rect 232 9136 233 9170
rect 197 9102 233 9136
rect 197 9068 198 9102
rect 232 9068 233 9102
rect 197 9034 233 9068
rect 197 9000 198 9034
rect 232 9000 233 9034
rect 197 8966 233 9000
rect 197 8932 198 8966
rect 232 8932 233 8966
rect 197 8898 233 8932
rect 197 8864 198 8898
rect 232 8864 233 8898
rect 197 8830 233 8864
rect 197 8796 198 8830
rect 232 8796 233 8830
rect 197 8762 233 8796
rect 1077 10427 1078 10461
rect 1112 10427 1113 10461
rect 1077 10393 1113 10427
rect 1077 10359 1078 10393
rect 1112 10359 1113 10393
rect 1077 10325 1113 10359
rect 1077 10291 1078 10325
rect 1112 10291 1113 10325
rect 1077 10257 1113 10291
rect 1077 10223 1078 10257
rect 1112 10223 1113 10257
rect 1077 10189 1113 10223
rect 1077 10155 1078 10189
rect 1112 10155 1113 10189
rect 1077 10121 1113 10155
rect 1077 10087 1078 10121
rect 1112 10087 1113 10121
rect 1077 10053 1113 10087
rect 1077 10019 1078 10053
rect 1112 10019 1113 10053
rect 1077 9985 1113 10019
rect 1077 9951 1078 9985
rect 1112 9951 1113 9985
rect 1077 9917 1113 9951
rect 1077 9883 1078 9917
rect 1112 9883 1113 9917
rect 1077 9849 1113 9883
rect 1077 9815 1078 9849
rect 1112 9815 1113 9849
rect 1077 9781 1113 9815
rect 1077 9747 1078 9781
rect 1112 9747 1113 9781
rect 1077 9713 1113 9747
rect 1077 9679 1078 9713
rect 1112 9679 1113 9713
rect 1077 9645 1113 9679
rect 1077 9611 1078 9645
rect 1112 9611 1113 9645
rect 1077 9577 1113 9611
rect 1077 9543 1078 9577
rect 1112 9543 1113 9577
rect 1077 9509 1113 9543
rect 1077 9475 1078 9509
rect 1112 9475 1113 9509
rect 1077 9441 1113 9475
rect 1077 9407 1078 9441
rect 1112 9407 1113 9441
rect 1077 9373 1113 9407
rect 1077 9339 1078 9373
rect 1112 9339 1113 9373
rect 1077 9305 1113 9339
rect 1077 9271 1078 9305
rect 1112 9271 1113 9305
rect 1077 9237 1113 9271
rect 1077 9203 1078 9237
rect 1112 9203 1113 9237
rect 1077 9169 1113 9203
rect 1077 9135 1078 9169
rect 1112 9135 1113 9169
rect 1077 9101 1113 9135
rect 1077 9067 1078 9101
rect 1112 9067 1113 9101
rect 1077 9033 1113 9067
rect 1077 8999 1078 9033
rect 1112 8999 1113 9033
rect 1077 8965 1113 8999
rect 1077 8931 1078 8965
rect 1112 8931 1113 8965
rect 1077 8897 1113 8931
rect 1077 8863 1078 8897
rect 1112 8863 1113 8897
rect 1077 8829 1113 8863
rect 1077 8795 1078 8829
rect 1112 8795 1113 8829
rect 197 8728 198 8762
rect 232 8728 233 8762
rect 307 8761 373 8773
rect 307 8745 323 8761
rect 197 8694 233 8728
rect 357 8745 373 8761
rect 433 8761 499 8773
rect 433 8745 449 8761
rect 323 8711 357 8727
rect 483 8745 499 8761
rect 559 8761 625 8773
rect 559 8745 575 8761
rect 449 8711 483 8727
rect 609 8745 625 8761
rect 685 8761 751 8773
rect 685 8745 701 8761
rect 575 8711 609 8727
rect 735 8745 751 8761
rect 811 8761 877 8773
rect 811 8745 827 8761
rect 701 8711 735 8727
rect 861 8745 877 8761
rect 937 8761 1003 8773
rect 937 8745 953 8761
rect 827 8711 861 8727
rect 987 8745 1003 8761
rect 1077 8761 1113 8795
rect 953 8711 987 8727
rect 1077 8727 1078 8761
rect 1112 8727 1113 8761
rect 197 8660 198 8694
rect 232 8660 233 8694
rect 197 8626 233 8660
rect 307 8689 373 8711
rect 307 8643 323 8689
rect 357 8643 373 8689
rect 433 8689 499 8711
rect 433 8643 449 8689
rect 483 8643 499 8689
rect 559 8689 625 8711
rect 559 8643 575 8689
rect 609 8643 625 8689
rect 685 8689 751 8711
rect 685 8643 701 8689
rect 735 8643 751 8689
rect 811 8689 877 8711
rect 811 8643 827 8689
rect 861 8643 877 8689
rect 937 8689 1003 8711
rect 937 8643 953 8689
rect 987 8643 1003 8689
rect 1077 8693 1113 8727
rect 1077 8659 1078 8693
rect 1112 8659 1113 8693
rect 197 8592 198 8626
rect 232 8592 233 8626
rect 197 8558 233 8592
rect 1077 8625 1113 8659
rect 1077 8591 1078 8625
rect 1112 8591 1113 8625
rect 197 8524 198 8558
rect 232 8524 233 8558
rect 197 8490 233 8524
rect 307 8521 323 8567
rect 357 8521 373 8567
rect 307 8499 373 8521
rect 433 8521 449 8567
rect 483 8521 499 8567
rect 433 8499 499 8521
rect 559 8521 575 8567
rect 609 8521 625 8567
rect 559 8499 625 8521
rect 685 8521 701 8567
rect 735 8521 751 8567
rect 685 8499 751 8521
rect 811 8521 827 8567
rect 861 8521 877 8567
rect 811 8499 877 8521
rect 937 8521 953 8567
rect 987 8521 1003 8567
rect 937 8499 1003 8521
rect 1077 8557 1113 8591
rect 1077 8523 1078 8557
rect 1112 8523 1113 8557
rect 197 8456 198 8490
rect 232 8456 233 8490
rect 323 8483 357 8499
rect 197 8422 233 8456
rect 307 8449 323 8465
rect 449 8483 483 8499
rect 357 8449 373 8465
rect 307 8437 373 8449
rect 433 8449 449 8465
rect 575 8483 609 8499
rect 483 8449 499 8465
rect 433 8437 499 8449
rect 559 8449 575 8465
rect 701 8483 735 8499
rect 609 8449 625 8465
rect 559 8437 625 8449
rect 685 8449 701 8465
rect 827 8483 861 8499
rect 735 8449 751 8465
rect 685 8437 751 8449
rect 811 8449 827 8465
rect 953 8483 987 8499
rect 861 8449 877 8465
rect 811 8437 877 8449
rect 937 8449 953 8465
rect 1077 8489 1113 8523
rect 987 8449 1003 8465
rect 937 8437 1003 8449
rect 1077 8455 1078 8489
rect 1112 8455 1113 8489
rect 197 8388 198 8422
rect 232 8388 233 8422
rect 197 8354 233 8388
rect 197 8320 198 8354
rect 232 8320 233 8354
rect 197 8286 233 8320
rect 197 8252 198 8286
rect 232 8252 233 8286
rect 197 8218 233 8252
rect 197 8184 198 8218
rect 232 8184 233 8218
rect 197 8150 233 8184
rect 197 8116 198 8150
rect 232 8116 233 8150
rect 197 8082 233 8116
rect 197 8048 198 8082
rect 232 8048 233 8082
rect 197 8014 233 8048
rect 197 7980 198 8014
rect 232 7980 233 8014
rect 197 7946 233 7980
rect 197 7912 198 7946
rect 232 7912 233 7946
rect 197 7878 233 7912
rect 197 7844 198 7878
rect 232 7844 233 7878
rect 197 7810 233 7844
rect 197 7776 198 7810
rect 232 7776 233 7810
rect 197 7742 233 7776
rect 197 7708 198 7742
rect 232 7708 233 7742
rect 197 7674 233 7708
rect 197 7640 198 7674
rect 232 7640 233 7674
rect 197 7606 233 7640
rect 197 7572 198 7606
rect 232 7572 233 7606
rect 197 7538 233 7572
rect 197 7504 198 7538
rect 232 7504 233 7538
rect 197 7470 233 7504
rect 197 7436 198 7470
rect 232 7436 233 7470
rect 197 7402 233 7436
rect 197 7368 198 7402
rect 232 7368 233 7402
rect 197 7334 233 7368
rect 197 7300 198 7334
rect 232 7300 233 7334
rect 197 7266 233 7300
rect 197 7232 198 7266
rect 232 7232 233 7266
rect 197 7198 233 7232
rect 197 7164 198 7198
rect 232 7164 233 7198
rect 197 7130 233 7164
rect 197 7096 198 7130
rect 232 7096 233 7130
rect 197 7062 233 7096
rect 197 7028 198 7062
rect 232 7028 233 7062
rect 197 6994 233 7028
rect 197 6960 198 6994
rect 232 6960 233 6994
rect 197 6926 233 6960
rect 197 6892 198 6926
rect 232 6892 233 6926
rect 197 6858 233 6892
rect 197 6824 198 6858
rect 232 6824 233 6858
rect 197 6790 233 6824
rect 197 6756 198 6790
rect 232 6756 233 6790
rect 1077 8421 1113 8455
rect 1077 8387 1078 8421
rect 1112 8387 1113 8421
rect 1077 8353 1113 8387
rect 1077 8319 1078 8353
rect 1112 8319 1113 8353
rect 1077 8285 1113 8319
rect 1077 8251 1078 8285
rect 1112 8251 1113 8285
rect 1077 8217 1113 8251
rect 1077 8183 1078 8217
rect 1112 8183 1113 8217
rect 1077 8149 1113 8183
rect 1077 8115 1078 8149
rect 1112 8115 1113 8149
rect 1077 8081 1113 8115
rect 1077 8047 1078 8081
rect 1112 8047 1113 8081
rect 1077 8013 1113 8047
rect 1077 7979 1078 8013
rect 1112 7979 1113 8013
rect 1077 7945 1113 7979
rect 1077 7911 1078 7945
rect 1112 7911 1113 7945
rect 1077 7877 1113 7911
rect 1077 7843 1078 7877
rect 1112 7843 1113 7877
rect 1077 7809 1113 7843
rect 1077 7775 1078 7809
rect 1112 7775 1113 7809
rect 1077 7741 1113 7775
rect 1077 7707 1078 7741
rect 1112 7707 1113 7741
rect 1077 7673 1113 7707
rect 1077 7639 1078 7673
rect 1112 7639 1113 7673
rect 1077 7605 1113 7639
rect 1077 7571 1078 7605
rect 1112 7571 1113 7605
rect 1077 7537 1113 7571
rect 1077 7503 1078 7537
rect 1112 7503 1113 7537
rect 1077 7469 1113 7503
rect 1077 7435 1078 7469
rect 1112 7435 1113 7469
rect 1077 7401 1113 7435
rect 1077 7367 1078 7401
rect 1112 7367 1113 7401
rect 1077 7333 1113 7367
rect 1077 7299 1078 7333
rect 1112 7299 1113 7333
rect 1077 7265 1113 7299
rect 1077 7231 1078 7265
rect 1112 7231 1113 7265
rect 1077 7197 1113 7231
rect 1077 7163 1078 7197
rect 1112 7163 1113 7197
rect 1077 7129 1113 7163
rect 1077 7095 1078 7129
rect 1112 7095 1113 7129
rect 1077 7061 1113 7095
rect 1077 7027 1078 7061
rect 1112 7027 1113 7061
rect 1077 6993 1113 7027
rect 1077 6959 1078 6993
rect 1112 6959 1113 6993
rect 1077 6925 1113 6959
rect 1077 6891 1078 6925
rect 1112 6891 1113 6925
rect 1077 6857 1113 6891
rect 1077 6823 1078 6857
rect 1112 6823 1113 6857
rect 1077 6789 1113 6823
rect 197 6722 233 6756
rect 307 6746 373 6758
rect 307 6730 323 6746
rect 197 6688 198 6722
rect 232 6688 233 6722
rect 357 6730 373 6746
rect 433 6746 499 6758
rect 433 6730 449 6746
rect 323 6696 357 6712
rect 483 6730 499 6746
rect 559 6746 625 6758
rect 559 6730 575 6746
rect 449 6696 483 6712
rect 609 6730 625 6746
rect 685 6746 751 6758
rect 685 6730 701 6746
rect 575 6696 609 6712
rect 735 6730 751 6746
rect 811 6746 877 6758
rect 811 6730 827 6746
rect 701 6696 735 6712
rect 861 6730 877 6746
rect 937 6746 1003 6758
rect 937 6730 953 6746
rect 827 6696 861 6712
rect 987 6730 1003 6746
rect 1077 6755 1078 6789
rect 1112 6755 1113 6789
rect 953 6696 987 6712
rect 1077 6721 1113 6755
rect 197 6654 233 6688
rect 197 6620 198 6654
rect 232 6620 233 6654
rect 307 6674 373 6696
rect 307 6628 323 6674
rect 357 6628 373 6674
rect 433 6674 499 6696
rect 433 6628 449 6674
rect 483 6628 499 6674
rect 559 6674 625 6696
rect 559 6628 575 6674
rect 609 6628 625 6674
rect 685 6674 751 6696
rect 685 6628 701 6674
rect 735 6628 751 6674
rect 811 6674 877 6696
rect 811 6628 827 6674
rect 861 6628 877 6674
rect 937 6674 1003 6696
rect 937 6628 953 6674
rect 987 6628 1003 6674
rect 1077 6681 1078 6721
rect 1112 6681 1113 6721
rect 1077 6653 1113 6681
rect 197 6586 233 6620
rect 197 6552 198 6586
rect 232 6552 233 6586
rect 1077 6609 1078 6653
rect 1112 6609 1113 6653
rect 1077 6585 1113 6609
rect 197 6518 233 6552
rect 197 6484 198 6518
rect 232 6484 233 6518
rect 307 6506 323 6552
rect 357 6506 373 6552
rect 307 6484 373 6506
rect 433 6506 449 6552
rect 483 6506 499 6552
rect 433 6484 499 6506
rect 559 6506 575 6552
rect 609 6506 625 6552
rect 559 6484 625 6506
rect 685 6506 701 6552
rect 735 6506 751 6552
rect 685 6484 751 6506
rect 811 6506 827 6552
rect 861 6506 877 6552
rect 811 6484 877 6506
rect 937 6506 953 6552
rect 987 6506 1003 6552
rect 937 6484 1003 6506
rect 1077 6537 1078 6585
rect 1112 6537 1113 6585
rect 1077 6517 1113 6537
rect 197 6450 233 6484
rect 323 6468 357 6484
rect 197 6416 198 6450
rect 232 6416 233 6450
rect 307 6434 323 6450
rect 449 6468 483 6484
rect 357 6434 373 6450
rect 307 6422 373 6434
rect 433 6434 449 6450
rect 575 6468 609 6484
rect 483 6434 499 6450
rect 433 6422 499 6434
rect 559 6434 575 6450
rect 701 6468 735 6484
rect 609 6434 625 6450
rect 559 6422 625 6434
rect 685 6434 701 6450
rect 827 6468 861 6484
rect 735 6434 751 6450
rect 685 6422 751 6434
rect 811 6434 827 6450
rect 953 6468 987 6484
rect 861 6434 877 6450
rect 811 6422 877 6434
rect 937 6434 953 6450
rect 1077 6465 1078 6517
rect 1112 6465 1113 6517
rect 987 6434 1003 6450
rect 937 6422 1003 6434
rect 1077 6449 1113 6465
rect 197 6382 233 6416
rect 197 6348 198 6382
rect 232 6348 233 6382
rect 197 6314 233 6348
rect 197 6280 198 6314
rect 232 6280 233 6314
rect 197 6246 233 6280
rect 197 6212 198 6246
rect 232 6212 233 6246
rect 197 6178 233 6212
rect 197 6144 198 6178
rect 232 6144 233 6178
rect 197 6110 233 6144
rect 197 6076 198 6110
rect 232 6076 233 6110
rect 197 6042 233 6076
rect 197 6008 198 6042
rect 232 6008 233 6042
rect 197 5974 233 6008
rect 197 5940 198 5974
rect 232 5940 233 5974
rect 197 5906 233 5940
rect 197 5872 198 5906
rect 232 5872 233 5906
rect 197 5838 233 5872
rect 197 5804 198 5838
rect 232 5804 233 5838
rect 197 5770 233 5804
rect 197 5736 198 5770
rect 232 5736 233 5770
rect 197 5702 233 5736
rect 197 5668 198 5702
rect 232 5668 233 5702
rect 197 5634 233 5668
rect 197 5600 198 5634
rect 232 5600 233 5634
rect 197 5566 233 5600
rect 197 5532 198 5566
rect 232 5532 233 5566
rect 197 5498 233 5532
rect 197 5464 198 5498
rect 232 5464 233 5498
rect 197 5430 233 5464
rect 197 5396 198 5430
rect 232 5396 233 5430
rect 197 5362 233 5396
rect 197 5328 198 5362
rect 232 5328 233 5362
rect 197 5294 233 5328
rect 197 5260 198 5294
rect 232 5260 233 5294
rect 197 5226 233 5260
rect 197 5192 198 5226
rect 232 5192 233 5226
rect 197 5158 233 5192
rect 197 5124 198 5158
rect 232 5124 233 5158
rect 197 5090 233 5124
rect 197 5056 198 5090
rect 232 5056 233 5090
rect 197 5022 233 5056
rect 197 4988 198 5022
rect 232 4988 233 5022
rect 197 4954 233 4988
rect 197 4920 198 4954
rect 232 4920 233 4954
rect 197 4886 233 4920
rect 197 4852 198 4886
rect 232 4852 233 4886
rect 197 4818 233 4852
rect 197 4784 198 4818
rect 232 4784 233 4818
rect 197 4750 233 4784
rect 197 4716 198 4750
rect 232 4716 233 4750
rect 1077 6415 1078 6449
rect 1112 6415 1113 6449
rect 1077 6381 1113 6415
rect 1077 6347 1078 6381
rect 1112 6347 1113 6381
rect 1077 6313 1113 6347
rect 1077 6279 1078 6313
rect 1112 6279 1113 6313
rect 1077 6245 1113 6279
rect 1077 6211 1078 6245
rect 1112 6211 1113 6245
rect 1077 6177 1113 6211
rect 1077 6143 1078 6177
rect 1112 6143 1113 6177
rect 1077 6109 1113 6143
rect 1077 6075 1078 6109
rect 1112 6075 1113 6109
rect 1077 6041 1113 6075
rect 1077 6007 1078 6041
rect 1112 6007 1113 6041
rect 1077 5973 1113 6007
rect 1077 5939 1078 5973
rect 1112 5939 1113 5973
rect 1077 5905 1113 5939
rect 1077 5871 1078 5905
rect 1112 5871 1113 5905
rect 1077 5837 1113 5871
rect 1077 5803 1078 5837
rect 1112 5803 1113 5837
rect 1077 5769 1113 5803
rect 1077 5735 1078 5769
rect 1112 5735 1113 5769
rect 1077 5701 1113 5735
rect 1077 5667 1078 5701
rect 1112 5667 1113 5701
rect 1077 5633 1113 5667
rect 1077 5599 1078 5633
rect 1112 5599 1113 5633
rect 1077 5565 1113 5599
rect 1077 5531 1078 5565
rect 1112 5531 1113 5565
rect 1077 5497 1113 5531
rect 1077 5463 1078 5497
rect 1112 5463 1113 5497
rect 1077 5429 1113 5463
rect 1077 5395 1078 5429
rect 1112 5395 1113 5429
rect 1077 5361 1113 5395
rect 1077 5327 1078 5361
rect 1112 5327 1113 5361
rect 1077 5293 1113 5327
rect 1077 5259 1078 5293
rect 1112 5259 1113 5293
rect 1077 5225 1113 5259
rect 1077 5191 1078 5225
rect 1112 5191 1113 5225
rect 1077 5157 1113 5191
rect 1077 5123 1078 5157
rect 1112 5123 1113 5157
rect 1077 5089 1113 5123
rect 1077 5055 1078 5089
rect 1112 5055 1113 5089
rect 1077 5021 1113 5055
rect 1077 4987 1078 5021
rect 1112 4987 1113 5021
rect 1077 4953 1113 4987
rect 1077 4919 1078 4953
rect 1112 4919 1113 4953
rect 1077 4885 1113 4919
rect 1077 4851 1078 4885
rect 1112 4851 1113 4885
rect 1077 4817 1113 4851
rect 1077 4783 1078 4817
rect 1112 4783 1113 4817
rect 1077 4749 1113 4783
rect 197 4682 233 4716
rect 307 4731 373 4743
rect 307 4715 323 4731
rect 197 4648 198 4682
rect 232 4648 233 4682
rect 357 4715 373 4731
rect 433 4731 499 4743
rect 433 4715 449 4731
rect 323 4681 357 4697
rect 483 4715 499 4731
rect 559 4731 625 4743
rect 559 4715 575 4731
rect 449 4681 483 4697
rect 609 4715 625 4731
rect 685 4731 751 4743
rect 685 4715 701 4731
rect 575 4681 609 4697
rect 735 4715 751 4731
rect 811 4731 877 4743
rect 811 4715 827 4731
rect 701 4681 735 4697
rect 861 4715 877 4731
rect 937 4731 1003 4743
rect 937 4715 953 4731
rect 827 4681 861 4697
rect 987 4715 1003 4731
rect 1077 4715 1078 4749
rect 1112 4715 1113 4749
rect 953 4681 987 4697
rect 1077 4681 1113 4715
rect 197 4614 233 4648
rect 197 4580 198 4614
rect 232 4580 233 4614
rect 307 4659 373 4681
rect 307 4613 323 4659
rect 357 4613 373 4659
rect 433 4659 499 4681
rect 433 4613 449 4659
rect 483 4613 499 4659
rect 559 4659 625 4681
rect 559 4613 575 4659
rect 609 4613 625 4659
rect 685 4659 751 4681
rect 685 4613 701 4659
rect 735 4613 751 4659
rect 811 4659 877 4681
rect 811 4613 827 4659
rect 861 4613 877 4659
rect 937 4659 1003 4681
rect 937 4613 953 4659
rect 987 4613 1003 4659
rect 1077 4647 1078 4681
rect 1112 4647 1113 4681
rect 1077 4613 1113 4647
rect 197 4546 233 4580
rect 197 4512 198 4546
rect 232 4512 233 4546
rect 1077 4579 1078 4613
rect 1112 4579 1113 4613
rect 1077 4545 1113 4579
rect 197 4478 233 4512
rect 197 4444 198 4478
rect 232 4444 233 4478
rect 307 4491 323 4537
rect 357 4491 373 4537
rect 307 4469 373 4491
rect 433 4491 449 4537
rect 483 4491 499 4537
rect 433 4469 499 4491
rect 559 4491 575 4537
rect 609 4491 625 4537
rect 559 4469 625 4491
rect 685 4491 701 4537
rect 735 4491 751 4537
rect 685 4469 751 4491
rect 811 4491 827 4537
rect 861 4491 877 4537
rect 811 4469 877 4491
rect 937 4491 953 4537
rect 987 4491 1003 4537
rect 937 4469 1003 4491
rect 1077 4511 1078 4545
rect 1112 4511 1113 4545
rect 1077 4477 1113 4511
rect 197 4410 233 4444
rect 323 4453 357 4469
rect 197 4376 198 4410
rect 232 4376 233 4410
rect 307 4419 323 4435
rect 449 4453 483 4469
rect 357 4419 373 4435
rect 307 4407 373 4419
rect 433 4419 449 4435
rect 575 4453 609 4469
rect 483 4419 499 4435
rect 433 4407 499 4419
rect 559 4419 575 4435
rect 701 4453 735 4469
rect 609 4419 625 4435
rect 559 4407 625 4419
rect 685 4419 701 4435
rect 827 4453 861 4469
rect 735 4419 751 4435
rect 685 4407 751 4419
rect 811 4419 827 4435
rect 953 4453 987 4469
rect 861 4419 877 4435
rect 811 4407 877 4419
rect 937 4419 953 4435
rect 1077 4443 1078 4477
rect 1112 4443 1113 4477
rect 987 4419 1003 4435
rect 937 4407 1003 4419
rect 1077 4409 1113 4443
rect 197 4342 233 4376
rect 197 4308 198 4342
rect 232 4308 233 4342
rect 197 4274 233 4308
rect 197 4240 198 4274
rect 232 4240 233 4274
rect 197 4206 233 4240
rect 197 4172 198 4206
rect 232 4172 233 4206
rect 197 4138 233 4172
rect 197 4104 198 4138
rect 232 4104 233 4138
rect 197 4070 233 4104
rect 197 4036 198 4070
rect 232 4036 233 4070
rect 197 4002 233 4036
rect 197 3968 198 4002
rect 232 3968 233 4002
rect 197 3934 233 3968
rect 197 3900 198 3934
rect 232 3900 233 3934
rect 197 3866 233 3900
rect 197 3832 198 3866
rect 232 3832 233 3866
rect 197 3798 233 3832
rect 197 3764 198 3798
rect 232 3764 233 3798
rect 197 3730 233 3764
rect 197 3696 198 3730
rect 232 3696 233 3730
rect 197 3662 233 3696
rect 197 3628 198 3662
rect 232 3628 233 3662
rect 197 3594 233 3628
rect 197 3560 198 3594
rect 232 3560 233 3594
rect 197 3526 233 3560
rect 197 3492 198 3526
rect 232 3492 233 3526
rect 197 3458 233 3492
rect 197 3424 198 3458
rect 232 3424 233 3458
rect 197 3390 233 3424
rect 197 3356 198 3390
rect 232 3356 233 3390
rect 197 3322 233 3356
rect 197 3288 198 3322
rect 232 3288 233 3322
rect 197 3254 233 3288
rect 197 3220 198 3254
rect 232 3220 233 3254
rect 197 3186 233 3220
rect 197 3152 198 3186
rect 232 3152 233 3186
rect 197 3118 233 3152
rect 197 3084 198 3118
rect 232 3084 233 3118
rect 197 3050 233 3084
rect 197 3016 198 3050
rect 232 3016 233 3050
rect 197 2982 233 3016
rect 197 2948 198 2982
rect 232 2948 233 2982
rect 197 2914 233 2948
rect 197 2880 198 2914
rect 232 2880 233 2914
rect 197 2846 233 2880
rect 197 2812 198 2846
rect 232 2812 233 2846
rect 197 2778 233 2812
rect 197 2744 198 2778
rect 232 2744 233 2778
rect 197 2710 233 2744
rect 1077 4375 1078 4409
rect 1112 4375 1113 4409
rect 1077 4341 1113 4375
rect 1077 4307 1078 4341
rect 1112 4307 1113 4341
rect 1077 4273 1113 4307
rect 1077 4239 1078 4273
rect 1112 4239 1113 4273
rect 1077 4205 1113 4239
rect 1077 4171 1078 4205
rect 1112 4171 1113 4205
rect 1077 4137 1113 4171
rect 1077 4103 1078 4137
rect 1112 4103 1113 4137
rect 1077 4069 1113 4103
rect 1077 4035 1078 4069
rect 1112 4035 1113 4069
rect 1077 4001 1113 4035
rect 1077 3967 1078 4001
rect 1112 3967 1113 4001
rect 1077 3933 1113 3967
rect 1077 3899 1078 3933
rect 1112 3899 1113 3933
rect 1077 3865 1113 3899
rect 1077 3831 1078 3865
rect 1112 3831 1113 3865
rect 1077 3797 1113 3831
rect 1077 3763 1078 3797
rect 1112 3763 1113 3797
rect 1077 3729 1113 3763
rect 1077 3695 1078 3729
rect 1112 3695 1113 3729
rect 1077 3661 1113 3695
rect 1077 3627 1078 3661
rect 1112 3627 1113 3661
rect 1077 3593 1113 3627
rect 1077 3559 1078 3593
rect 1112 3559 1113 3593
rect 1077 3525 1113 3559
rect 1077 3491 1078 3525
rect 1112 3491 1113 3525
rect 1077 3457 1113 3491
rect 1077 3423 1078 3457
rect 1112 3423 1113 3457
rect 1077 3389 1113 3423
rect 1077 3355 1078 3389
rect 1112 3355 1113 3389
rect 1077 3321 1113 3355
rect 1077 3287 1078 3321
rect 1112 3287 1113 3321
rect 1077 3253 1113 3287
rect 1077 3219 1078 3253
rect 1112 3219 1113 3253
rect 1077 3185 1113 3219
rect 1077 3151 1078 3185
rect 1112 3151 1113 3185
rect 1077 3117 1113 3151
rect 1077 3083 1078 3117
rect 1112 3083 1113 3117
rect 1077 3049 1113 3083
rect 1077 3015 1078 3049
rect 1112 3015 1113 3049
rect 1077 2981 1113 3015
rect 1077 2947 1078 2981
rect 1112 2947 1113 2981
rect 1077 2913 1113 2947
rect 1077 2879 1078 2913
rect 1112 2879 1113 2913
rect 1077 2845 1113 2879
rect 1077 2811 1078 2845
rect 1112 2811 1113 2845
rect 1077 2777 1113 2811
rect 1077 2743 1078 2777
rect 1112 2743 1113 2777
rect 197 2676 198 2710
rect 232 2676 233 2710
rect 307 2716 373 2728
rect 307 2700 323 2716
rect 197 2642 233 2676
rect 357 2700 373 2716
rect 433 2716 499 2728
rect 433 2700 449 2716
rect 323 2666 357 2682
rect 483 2700 499 2716
rect 559 2716 625 2728
rect 559 2700 575 2716
rect 449 2666 483 2682
rect 609 2700 625 2716
rect 685 2716 751 2728
rect 685 2700 701 2716
rect 575 2666 609 2682
rect 735 2700 751 2716
rect 811 2716 877 2728
rect 811 2700 827 2716
rect 701 2666 735 2682
rect 861 2700 877 2716
rect 937 2716 1003 2728
rect 937 2700 953 2716
rect 827 2666 861 2682
rect 987 2700 1003 2716
rect 1077 2709 1113 2743
rect 953 2666 987 2682
rect 1077 2675 1078 2709
rect 1112 2675 1113 2709
rect 197 2608 198 2642
rect 232 2608 233 2642
rect 197 2574 233 2608
rect 307 2644 373 2666
rect 307 2598 323 2644
rect 357 2598 373 2644
rect 433 2644 499 2666
rect 433 2598 449 2644
rect 483 2598 499 2644
rect 559 2644 625 2666
rect 559 2598 575 2644
rect 609 2598 625 2644
rect 685 2644 751 2666
rect 685 2598 701 2644
rect 735 2598 751 2644
rect 811 2644 877 2666
rect 811 2598 827 2644
rect 861 2598 877 2644
rect 937 2644 1003 2666
rect 937 2598 953 2644
rect 987 2598 1003 2644
rect 1077 2641 1113 2675
rect 1077 2607 1078 2641
rect 1112 2607 1113 2641
rect 197 2540 198 2574
rect 232 2540 233 2574
rect 197 2506 233 2540
rect 1077 2573 1113 2607
rect 1077 2539 1078 2573
rect 1112 2539 1113 2573
rect 197 2472 198 2506
rect 232 2472 233 2506
rect 197 2438 233 2472
rect 307 2476 323 2522
rect 357 2476 373 2522
rect 307 2454 373 2476
rect 433 2476 449 2522
rect 483 2476 499 2522
rect 433 2454 499 2476
rect 559 2476 575 2522
rect 609 2476 625 2522
rect 559 2454 625 2476
rect 685 2476 701 2522
rect 735 2476 751 2522
rect 685 2454 751 2476
rect 811 2476 827 2522
rect 861 2476 877 2522
rect 811 2454 877 2476
rect 937 2476 953 2522
rect 987 2476 1003 2522
rect 937 2454 1003 2476
rect 1077 2505 1113 2539
rect 1077 2471 1078 2505
rect 1112 2471 1113 2505
rect 197 2404 198 2438
rect 232 2404 233 2438
rect 323 2438 357 2454
rect 197 2370 233 2404
rect 307 2404 323 2420
rect 449 2438 483 2454
rect 357 2404 373 2420
rect 307 2392 373 2404
rect 433 2404 449 2420
rect 575 2438 609 2454
rect 483 2404 499 2420
rect 433 2392 499 2404
rect 559 2404 575 2420
rect 701 2438 735 2454
rect 609 2404 625 2420
rect 559 2392 625 2404
rect 685 2404 701 2420
rect 827 2438 861 2454
rect 735 2404 751 2420
rect 685 2392 751 2404
rect 811 2404 827 2420
rect 953 2438 987 2454
rect 861 2404 877 2420
rect 811 2392 877 2404
rect 937 2404 953 2420
rect 1077 2437 1113 2471
rect 987 2404 1003 2420
rect 937 2392 1003 2404
rect 1077 2403 1078 2437
rect 1112 2403 1113 2437
rect 197 2336 198 2370
rect 232 2336 233 2370
rect 197 2302 233 2336
rect 197 2268 198 2302
rect 232 2268 233 2302
rect 197 2234 233 2268
rect 197 2200 198 2234
rect 232 2200 233 2234
rect 197 2166 233 2200
rect 197 2132 198 2166
rect 232 2132 233 2166
rect 197 2098 233 2132
rect 197 2064 198 2098
rect 232 2064 233 2098
rect 197 2030 233 2064
rect 197 1996 198 2030
rect 232 1996 233 2030
rect 197 1962 233 1996
rect 197 1928 198 1962
rect 232 1928 233 1962
rect 197 1894 233 1928
rect 197 1860 198 1894
rect 232 1860 233 1894
rect 197 1826 233 1860
rect 197 1792 198 1826
rect 232 1792 233 1826
rect 197 1758 233 1792
rect 197 1724 198 1758
rect 232 1724 233 1758
rect 197 1690 233 1724
rect 197 1656 198 1690
rect 232 1656 233 1690
rect 197 1622 233 1656
rect 197 1588 198 1622
rect 232 1588 233 1622
rect 197 1554 233 1588
rect 197 1520 198 1554
rect 232 1520 233 1554
rect 197 1486 233 1520
rect 197 1452 198 1486
rect 232 1452 233 1486
rect 197 1418 233 1452
rect 197 1384 198 1418
rect 232 1384 233 1418
rect 197 1350 233 1384
rect 197 1316 198 1350
rect 232 1316 233 1350
rect 197 1282 233 1316
rect 197 1248 198 1282
rect 232 1248 233 1282
rect 197 1214 233 1248
rect 197 1180 198 1214
rect 232 1180 233 1214
rect 197 1146 233 1180
rect 197 1112 198 1146
rect 232 1112 233 1146
rect 197 1078 233 1112
rect 197 1044 198 1078
rect 232 1044 233 1078
rect 197 1010 233 1044
rect 197 976 198 1010
rect 232 976 233 1010
rect 197 942 233 976
rect 197 908 198 942
rect 232 908 233 942
rect 197 874 233 908
rect 197 840 198 874
rect 232 840 233 874
rect 197 806 233 840
rect 197 772 198 806
rect 232 772 233 806
rect 197 738 233 772
rect 197 704 198 738
rect 232 704 233 738
rect 1077 2369 1113 2403
rect 1077 2335 1078 2369
rect 1112 2335 1113 2369
rect 1077 2301 1113 2335
rect 1077 2267 1078 2301
rect 1112 2267 1113 2301
rect 1077 2233 1113 2267
rect 1077 2199 1078 2233
rect 1112 2199 1113 2233
rect 1077 2165 1113 2199
rect 1077 2131 1078 2165
rect 1112 2131 1113 2165
rect 1077 2097 1113 2131
rect 1077 2063 1078 2097
rect 1112 2063 1113 2097
rect 1456 10706 1457 10743
rect 1491 10706 1492 10743
rect 8414 10785 8415 10819
rect 8449 10785 8450 10819
rect 8414 10751 8450 10785
rect 1456 10675 1492 10706
rect 1456 10634 1457 10675
rect 1491 10634 1492 10675
rect 1456 10607 1492 10634
rect 1456 10562 1457 10607
rect 1491 10562 1492 10607
rect 1456 10539 1492 10562
rect 1456 10490 1457 10539
rect 1491 10490 1492 10539
rect 1456 10471 1492 10490
rect 1456 10437 1457 10471
rect 1491 10437 1492 10471
rect 1456 10403 1492 10437
rect 1456 10369 1457 10403
rect 1491 10369 1492 10403
rect 1456 10335 1492 10369
rect 1456 10301 1457 10335
rect 1491 10301 1492 10335
rect 1456 10267 1492 10301
rect 1456 10233 1457 10267
rect 1491 10233 1492 10267
rect 1456 10199 1492 10233
rect 1456 10165 1457 10199
rect 1491 10165 1492 10199
rect 1456 10131 1492 10165
rect 1456 10097 1457 10131
rect 1491 10097 1492 10131
rect 1456 10063 1492 10097
rect 1456 10029 1457 10063
rect 1491 10029 1492 10063
rect 1456 9995 1492 10029
rect 1456 9961 1457 9995
rect 1491 9961 1492 9995
rect 1456 9927 1492 9961
rect 1456 9893 1457 9927
rect 1491 9893 1492 9927
rect 1456 9859 1492 9893
rect 1456 9825 1457 9859
rect 1491 9825 1492 9859
rect 1456 9822 1492 9825
rect 1490 9791 1492 9822
rect 1456 9757 1457 9788
rect 1491 9757 1492 9791
rect 1456 9750 1492 9757
rect 1490 9723 1492 9750
rect 1456 9689 1457 9716
rect 1491 9689 1492 9723
rect 1456 9678 1492 9689
rect 1490 9655 1492 9678
rect 1456 9621 1457 9644
rect 1491 9621 1492 9655
rect 1456 9587 1492 9621
rect 1456 9553 1457 9587
rect 1491 9553 1492 9587
rect 1456 9519 1492 9553
rect 1456 9485 1457 9519
rect 1491 9485 1492 9519
rect 1456 9451 1492 9485
rect 1456 9417 1457 9451
rect 1491 9417 1492 9451
rect 1456 9383 1492 9417
rect 1456 9349 1457 9383
rect 1491 9349 1492 9383
rect 1456 9315 1492 9349
rect 1456 9281 1457 9315
rect 1491 9281 1492 9315
rect 1456 9247 1492 9281
rect 1456 9213 1457 9247
rect 1491 9213 1492 9247
rect 1456 9179 1492 9213
rect 1456 9145 1457 9179
rect 1491 9145 1492 9179
rect 1456 9111 1492 9145
rect 1456 9077 1457 9111
rect 1491 9077 1492 9111
rect 1456 9043 1492 9077
rect 1456 9009 1457 9043
rect 1491 9009 1492 9043
rect 1456 8975 1492 9009
rect 1456 8941 1457 8975
rect 1491 8941 1492 8975
rect 1456 8919 1492 8941
rect 1490 8907 1492 8919
rect 1456 8873 1457 8885
rect 1491 8873 1492 8907
rect 1456 8847 1492 8873
rect 1490 8839 1492 8847
rect 1456 8805 1457 8813
rect 1491 8805 1492 8839
rect 1456 8775 1492 8805
rect 1689 10690 1691 10724
rect 1725 10723 8261 10724
rect 1725 10690 1801 10723
rect 1689 10656 1690 10690
rect 1724 10689 1801 10690
rect 1835 10689 1869 10723
rect 1903 10689 1937 10723
rect 1971 10689 2005 10723
rect 2039 10689 2073 10723
rect 2107 10689 2141 10723
rect 2175 10689 2209 10723
rect 2243 10689 2277 10723
rect 2311 10689 2345 10723
rect 2379 10689 2413 10723
rect 2447 10689 2481 10723
rect 2515 10689 2549 10723
rect 2583 10689 2617 10723
rect 2651 10689 2685 10723
rect 2719 10689 2753 10723
rect 2787 10689 2821 10723
rect 2855 10689 2889 10723
rect 2923 10689 2957 10723
rect 2991 10689 3025 10723
rect 3059 10689 3093 10723
rect 3127 10689 3161 10723
rect 3195 10689 3229 10723
rect 3263 10689 3297 10723
rect 3331 10689 3365 10723
rect 3399 10689 3433 10723
rect 3467 10689 3501 10723
rect 3535 10689 3569 10723
rect 3603 10689 3637 10723
rect 3671 10689 3705 10723
rect 3739 10689 3773 10723
rect 3807 10689 3841 10723
rect 3875 10689 3909 10723
rect 3943 10689 3977 10723
rect 4011 10689 4045 10723
rect 4079 10689 4113 10723
rect 4147 10689 4181 10723
rect 4215 10689 4249 10723
rect 4283 10689 4317 10723
rect 4351 10689 4385 10723
rect 4419 10689 4453 10723
rect 4487 10689 4521 10723
rect 4555 10689 4589 10723
rect 4623 10689 4657 10723
rect 4691 10689 4725 10723
rect 4759 10689 4793 10723
rect 4827 10689 4861 10723
rect 4895 10689 4929 10723
rect 4963 10689 4997 10723
rect 5031 10689 5065 10723
rect 5099 10689 5133 10723
rect 5167 10689 5201 10723
rect 5235 10689 5269 10723
rect 5303 10689 5337 10723
rect 5371 10689 5405 10723
rect 5439 10689 5473 10723
rect 5507 10689 5541 10723
rect 5575 10689 5609 10723
rect 5643 10689 5677 10723
rect 5711 10689 5745 10723
rect 5779 10689 5813 10723
rect 5847 10689 5881 10723
rect 5915 10689 5949 10723
rect 5983 10689 6017 10723
rect 6051 10689 6085 10723
rect 6119 10689 6153 10723
rect 6187 10689 6221 10723
rect 6255 10689 6289 10723
rect 6323 10689 6357 10723
rect 6391 10689 6425 10723
rect 6459 10689 6493 10723
rect 6527 10689 6561 10723
rect 6595 10689 6629 10723
rect 6663 10689 6697 10723
rect 6731 10689 6765 10723
rect 6799 10689 6833 10723
rect 6867 10689 6901 10723
rect 6935 10689 6969 10723
rect 7003 10689 7037 10723
rect 7071 10689 7105 10723
rect 7139 10689 7173 10723
rect 7207 10689 7241 10723
rect 7275 10689 7309 10723
rect 7343 10689 7377 10723
rect 7411 10689 7445 10723
rect 7479 10689 7513 10723
rect 7547 10689 7581 10723
rect 7615 10689 7649 10723
rect 7683 10689 7717 10723
rect 7751 10689 7785 10723
rect 7819 10689 7853 10723
rect 7887 10689 7921 10723
rect 7955 10689 7989 10723
rect 8023 10689 8057 10723
rect 8091 10689 8125 10723
rect 8159 10689 8193 10723
rect 8227 10689 8261 10723
rect 1724 10688 8261 10689
rect 1724 10656 1725 10688
rect 1689 10652 1725 10656
rect 1689 10622 1691 10652
rect 1689 10588 1690 10622
rect 1724 10588 1725 10618
rect 1689 10580 1725 10588
rect 1689 10554 1691 10580
rect 1689 10520 1690 10554
rect 1724 10520 1725 10546
rect 8225 10646 8261 10688
rect 8225 10612 8226 10646
rect 8260 10612 8261 10646
rect 8225 10578 8261 10612
rect 8225 10544 8226 10578
rect 8260 10544 8261 10578
rect 1689 10486 1725 10520
rect 1689 10452 1690 10486
rect 1724 10452 1725 10486
rect 1689 10418 1725 10452
rect 1689 10384 1690 10418
rect 1724 10384 1725 10418
rect 1689 10350 1725 10384
rect 1689 10316 1690 10350
rect 1724 10316 1725 10350
rect 1689 10282 1725 10316
rect 1689 10248 1690 10282
rect 1724 10248 1725 10282
rect 1689 10214 1725 10248
rect 1689 10180 1690 10214
rect 1724 10180 1725 10214
rect 1689 10146 1725 10180
rect 1689 10112 1690 10146
rect 1724 10112 1725 10146
rect 1689 10078 1725 10112
rect 1689 10044 1690 10078
rect 1724 10044 1725 10078
rect 1689 10010 1725 10044
rect 1689 9976 1690 10010
rect 1724 9976 1725 10010
rect 1689 9942 1725 9976
rect 1689 9908 1690 9942
rect 1724 9908 1725 9942
rect 1689 9874 1725 9908
rect 1689 9840 1690 9874
rect 1724 9840 1725 9874
rect 1689 9822 1725 9840
rect 1689 9772 1690 9822
rect 1724 9772 1725 9822
rect 1799 10418 1840 10534
rect 8112 10418 8153 10534
rect 1799 10384 1806 10418
rect 1799 10346 1840 10384
rect 1799 10312 1806 10346
rect 1799 10274 1840 10312
rect 1799 10240 1806 10274
rect 1799 10202 1840 10240
rect 1799 10168 1806 10202
rect 1799 10130 1840 10168
rect 1799 10096 1806 10130
rect 1799 10058 1840 10096
rect 1799 10024 1806 10058
rect 1799 9986 1840 10024
rect 1799 9952 1806 9986
rect 3893 10346 3927 10384
rect 3893 10274 3927 10312
rect 3893 10202 3927 10240
rect 3893 10130 3927 10168
rect 3893 10058 3927 10096
rect 3893 9986 3927 10024
rect 6023 10346 6057 10384
rect 6023 10274 6057 10312
rect 6023 10202 6057 10240
rect 6023 10130 6057 10168
rect 6023 10058 6057 10096
rect 6023 9986 6057 10024
rect 8146 10384 8153 10418
rect 8112 10346 8153 10384
rect 8146 10312 8153 10346
rect 8112 10274 8153 10312
rect 8146 10240 8153 10274
rect 8112 10202 8153 10240
rect 8146 10168 8153 10202
rect 8112 10130 8153 10168
rect 8146 10096 8153 10130
rect 8112 10058 8153 10096
rect 8146 10024 8153 10058
rect 8112 9986 8153 10024
rect 8146 9952 8153 9986
rect 1799 9788 1840 9952
rect 8112 9788 8153 9952
rect 8225 10510 8261 10544
rect 8225 10476 8226 10510
rect 8260 10476 8261 10510
rect 8225 10442 8261 10476
rect 8225 10408 8226 10442
rect 8260 10408 8261 10442
rect 8225 10374 8261 10408
rect 8225 10340 8226 10374
rect 8260 10340 8261 10374
rect 8225 10306 8261 10340
rect 8225 10272 8226 10306
rect 8260 10272 8261 10306
rect 8225 10238 8261 10272
rect 8225 10204 8226 10238
rect 8260 10204 8261 10238
rect 8225 10170 8261 10204
rect 8225 10136 8226 10170
rect 8260 10136 8261 10170
rect 8225 10102 8261 10136
rect 8225 10068 8226 10102
rect 8260 10068 8261 10102
rect 8225 10034 8261 10068
rect 8225 10000 8226 10034
rect 8260 10000 8261 10034
rect 8225 9966 8261 10000
rect 8225 9932 8226 9966
rect 8260 9932 8261 9966
rect 8225 9898 8261 9932
rect 8225 9864 8226 9898
rect 8260 9864 8261 9898
rect 8225 9830 8261 9864
rect 8225 9796 8226 9830
rect 8260 9796 8261 9830
rect 1689 9750 1725 9772
rect 1689 9704 1690 9750
rect 1724 9704 1725 9750
rect 1689 9678 1725 9704
rect 8225 9762 8261 9796
rect 8225 9728 8226 9762
rect 8260 9728 8261 9762
rect 8225 9694 8261 9728
rect 1689 9636 1690 9678
rect 1724 9636 1725 9678
rect 1689 9602 1725 9636
rect 1689 9568 1690 9602
rect 1724 9568 1725 9602
rect 1689 9534 1725 9568
rect 1689 9500 1690 9534
rect 1724 9500 1725 9534
rect 1689 9466 1725 9500
rect 1689 9432 1690 9466
rect 1724 9432 1725 9466
rect 1689 9398 1725 9432
rect 1689 9364 1690 9398
rect 1724 9364 1725 9398
rect 1689 9330 1725 9364
rect 1689 9296 1690 9330
rect 1724 9296 1725 9330
rect 1799 9310 1840 9678
rect 8112 9514 8153 9678
rect 1689 9262 1725 9296
rect 1689 9228 1690 9262
rect 1724 9228 1725 9262
rect 1689 9194 1725 9228
rect 1689 9160 1690 9194
rect 1724 9160 1725 9194
rect 1689 9126 1725 9160
rect 1689 9092 1690 9126
rect 1724 9092 1725 9126
rect 1689 9058 1725 9092
rect 1689 9024 1690 9058
rect 1724 9024 1725 9058
rect 1689 8990 1725 9024
rect 1689 8956 1690 8990
rect 1724 8956 1725 8990
rect 1807 9276 1840 9310
rect 1773 9238 1840 9276
rect 1807 9204 1840 9238
rect 1773 9166 1840 9204
rect 1807 9132 1840 9166
rect 1773 9094 1840 9132
rect 1807 9060 1840 9094
rect 1773 9022 1840 9060
rect 6023 9442 6057 9480
rect 6023 9370 6057 9408
rect 6023 9298 6057 9336
rect 6023 9226 6057 9264
rect 6023 9154 6057 9192
rect 6023 9082 6057 9120
rect 8146 9480 8153 9514
rect 8112 9442 8153 9480
rect 8146 9408 8153 9442
rect 8112 9370 8153 9408
rect 8146 9336 8153 9370
rect 8112 9298 8153 9336
rect 8146 9264 8153 9298
rect 8112 9226 8153 9264
rect 8146 9192 8153 9226
rect 8112 9154 8153 9192
rect 8146 9120 8153 9154
rect 8112 9082 8153 9120
rect 8146 9048 8153 9082
rect 1807 8988 1840 9022
rect 1689 8922 1725 8956
rect 1799 8932 1840 8988
rect 8112 8932 8153 9048
rect 8225 9660 8226 9694
rect 8260 9660 8261 9694
rect 8225 9626 8261 9660
rect 8225 9592 8226 9626
rect 8260 9592 8261 9626
rect 8225 9558 8261 9592
rect 8225 9524 8226 9558
rect 8260 9524 8261 9558
rect 8225 9490 8261 9524
rect 8225 9456 8226 9490
rect 8260 9456 8261 9490
rect 8225 9422 8261 9456
rect 8225 9388 8226 9422
rect 8260 9388 8261 9422
rect 8225 9354 8261 9388
rect 8225 9320 8226 9354
rect 8260 9320 8261 9354
rect 8225 9286 8261 9320
rect 8225 9252 8226 9286
rect 8260 9252 8261 9286
rect 8225 9218 8261 9252
rect 8225 9184 8226 9218
rect 8260 9184 8261 9218
rect 8225 9150 8261 9184
rect 8225 9116 8226 9150
rect 8260 9116 8261 9150
rect 8225 9082 8261 9116
rect 8225 9048 8226 9082
rect 8260 9048 8261 9082
rect 8225 9014 8261 9048
rect 8225 8980 8226 9014
rect 8260 8980 8261 9014
rect 8225 8946 8261 8980
rect 1689 8886 1690 8922
rect 1724 8886 1725 8922
rect 1689 8848 1725 8886
rect 1689 8814 1690 8848
rect 1724 8814 1725 8848
rect 1689 8778 1725 8814
rect 8225 8912 8226 8946
rect 8260 8912 8261 8946
rect 8225 8878 8261 8912
rect 8225 8844 8226 8878
rect 8260 8844 8261 8878
rect 8225 8810 8261 8844
rect 8225 8778 8226 8810
rect 1490 8771 1492 8775
rect 1456 8737 1457 8741
rect 1491 8737 1492 8771
rect 1456 8703 1492 8737
rect 1456 8669 1457 8703
rect 1491 8669 1492 8703
rect 1456 8635 1492 8669
rect 1456 8601 1457 8635
rect 1491 8601 1492 8635
rect 1456 8567 1492 8601
rect 1456 8533 1457 8567
rect 1491 8533 1492 8567
rect 1456 8499 1492 8533
rect 1456 8465 1457 8499
rect 1491 8465 1492 8499
rect 1456 8431 1492 8465
rect 1456 8397 1457 8431
rect 1491 8397 1492 8431
rect 1456 8363 1492 8397
rect 1456 8329 1457 8363
rect 1491 8329 1492 8363
rect 1456 8295 1492 8329
rect 1456 8261 1457 8295
rect 1491 8261 1492 8295
rect 1456 8227 1492 8261
rect 1456 8193 1457 8227
rect 1491 8193 1492 8227
rect 1456 8159 1492 8193
rect 1456 8125 1457 8159
rect 1491 8125 1492 8159
rect 1456 8091 1492 8125
rect 1456 8057 1457 8091
rect 1491 8057 1492 8091
rect 1456 8023 1492 8057
rect 1456 7989 1457 8023
rect 1491 7989 1492 8023
rect 1456 7955 1492 7989
rect 1456 7921 1457 7955
rect 1491 7921 1492 7955
rect 1456 7887 1492 7921
rect 1456 7853 1457 7887
rect 1491 7853 1492 7887
rect 1456 7819 1492 7853
rect 1456 7785 1457 7819
rect 1491 7785 1492 7819
rect 1456 7751 1492 7785
rect 1456 7717 1457 7751
rect 1491 7717 1492 7751
rect 1456 7683 1492 7717
rect 1456 7649 1457 7683
rect 1491 7649 1492 7683
rect 1456 7615 1492 7649
rect 1456 7581 1457 7615
rect 1491 7581 1492 7615
rect 1456 7547 1492 7581
rect 1456 7513 1457 7547
rect 1491 7513 1492 7547
rect 1456 7479 1492 7513
rect 1456 7445 1457 7479
rect 1491 7445 1492 7479
rect 1645 8777 8226 8778
rect 1645 8744 1723 8777
rect 1645 8710 1646 8744
rect 1680 8743 1723 8744
rect 1757 8743 1791 8777
rect 1825 8743 1859 8777
rect 1893 8743 1927 8777
rect 1961 8743 1995 8777
rect 2029 8743 2063 8777
rect 2097 8743 2131 8777
rect 2165 8743 2199 8777
rect 2233 8743 2267 8777
rect 2301 8743 2335 8777
rect 2369 8743 2403 8777
rect 2437 8743 2471 8777
rect 2505 8743 2539 8777
rect 2573 8743 2607 8777
rect 2641 8743 2675 8777
rect 2709 8743 2743 8777
rect 2777 8743 2811 8777
rect 2845 8743 2879 8777
rect 2913 8743 2947 8777
rect 2981 8743 3015 8777
rect 3049 8743 3083 8777
rect 3117 8743 3151 8777
rect 3185 8743 3219 8777
rect 3253 8743 3287 8777
rect 3321 8743 3355 8777
rect 3389 8743 3423 8777
rect 3457 8743 3491 8777
rect 3525 8743 3559 8777
rect 3593 8743 3627 8777
rect 3661 8743 3695 8777
rect 3729 8743 3763 8777
rect 3797 8743 3831 8777
rect 3865 8743 3899 8777
rect 3933 8743 3967 8777
rect 4001 8743 4035 8777
rect 4069 8743 4103 8777
rect 4137 8743 4171 8777
rect 4205 8743 4239 8777
rect 4273 8743 4307 8777
rect 4341 8743 4375 8777
rect 4409 8743 4443 8777
rect 4477 8743 4511 8777
rect 4545 8743 4579 8777
rect 4613 8743 4647 8777
rect 4681 8743 4715 8777
rect 4749 8743 4783 8777
rect 4817 8743 4851 8777
rect 4885 8743 4919 8777
rect 4953 8743 4987 8777
rect 5021 8743 5055 8777
rect 5089 8743 5123 8777
rect 5157 8743 5191 8777
rect 5225 8743 5259 8777
rect 5293 8743 5327 8777
rect 5361 8743 5395 8777
rect 5429 8743 5463 8777
rect 5497 8743 5531 8777
rect 5565 8743 5599 8777
rect 5633 8743 5667 8777
rect 5701 8743 5735 8777
rect 5769 8743 5803 8777
rect 5837 8743 5871 8777
rect 5905 8743 5939 8777
rect 5973 8743 6007 8777
rect 6041 8743 6075 8777
rect 6109 8743 6143 8777
rect 6177 8743 6211 8777
rect 6245 8743 6279 8777
rect 6313 8743 6347 8777
rect 6381 8743 6415 8777
rect 6449 8743 6483 8777
rect 6517 8743 6551 8777
rect 6585 8743 6619 8777
rect 6653 8743 6687 8777
rect 6721 8743 6755 8777
rect 6789 8743 6823 8777
rect 6857 8743 6891 8777
rect 6925 8743 6959 8777
rect 6993 8743 7027 8777
rect 7061 8743 7095 8777
rect 7129 8743 7163 8777
rect 7197 8743 7231 8777
rect 7265 8743 7299 8777
rect 7333 8743 7367 8777
rect 7401 8743 7435 8777
rect 7469 8743 7503 8777
rect 7537 8743 7571 8777
rect 7605 8743 7639 8777
rect 7673 8743 7707 8777
rect 7741 8743 7775 8777
rect 7809 8743 7843 8777
rect 7877 8743 7911 8777
rect 7945 8743 7979 8777
rect 8013 8743 8047 8777
rect 8081 8743 8115 8777
rect 8149 8776 8226 8777
rect 8260 8776 8261 8810
rect 8149 8743 8261 8776
rect 1680 8742 8261 8743
rect 8414 10717 8415 10751
rect 8449 10717 8450 10751
rect 8414 10683 8450 10717
rect 8414 10649 8415 10683
rect 8449 10649 8450 10683
rect 8414 10615 8450 10649
rect 8414 10581 8415 10615
rect 8449 10581 8450 10615
rect 8414 10547 8450 10581
rect 8414 10513 8415 10547
rect 8449 10513 8450 10547
rect 8414 10479 8450 10513
rect 8414 10445 8415 10479
rect 8449 10445 8450 10479
rect 8414 10411 8450 10445
rect 8414 10377 8415 10411
rect 8449 10377 8450 10411
rect 8414 10343 8450 10377
rect 8414 10309 8415 10343
rect 8449 10309 8450 10343
rect 8414 10275 8450 10309
rect 8414 10241 8415 10275
rect 8449 10241 8450 10275
rect 8414 10207 8450 10241
rect 8414 10173 8415 10207
rect 8449 10173 8450 10207
rect 8414 10139 8450 10173
rect 8414 10105 8415 10139
rect 8449 10105 8450 10139
rect 8414 10071 8450 10105
rect 8414 10037 8415 10071
rect 8449 10037 8450 10071
rect 8414 10003 8450 10037
rect 8414 9969 8415 10003
rect 8449 9969 8450 10003
rect 8414 9935 8450 9969
rect 8414 9901 8415 9935
rect 8449 9901 8450 9935
rect 8414 9867 8450 9901
rect 8414 9833 8415 9867
rect 8449 9833 8450 9867
rect 8414 9799 8450 9833
rect 8414 9765 8415 9799
rect 8449 9765 8450 9799
rect 8414 9731 8450 9765
rect 8414 9697 8415 9731
rect 8449 9697 8450 9731
rect 8414 9663 8450 9697
rect 8414 9629 8415 9663
rect 8449 9629 8450 9663
rect 8414 9595 8450 9629
rect 8414 9561 8415 9595
rect 8449 9561 8450 9595
rect 8414 9527 8450 9561
rect 8414 9493 8415 9527
rect 8449 9493 8450 9527
rect 8414 9459 8450 9493
rect 8414 9425 8415 9459
rect 8449 9425 8450 9459
rect 8414 9391 8450 9425
rect 8414 9357 8415 9391
rect 8449 9357 8450 9391
rect 8414 9323 8450 9357
rect 8414 9289 8415 9323
rect 8449 9289 8450 9323
rect 8414 9255 8450 9289
rect 8414 9221 8415 9255
rect 8449 9221 8450 9255
rect 8414 9187 8450 9221
rect 8414 9153 8415 9187
rect 8449 9153 8450 9187
rect 8414 9119 8450 9153
rect 8414 9085 8415 9119
rect 8449 9085 8450 9119
rect 8414 9051 8450 9085
rect 8414 9017 8415 9051
rect 8449 9017 8450 9051
rect 8414 8983 8450 9017
rect 8414 8949 8415 8983
rect 8449 8949 8450 8983
rect 8414 8915 8450 8949
rect 8414 8881 8415 8915
rect 8449 8881 8450 8915
rect 8414 8847 8450 8881
rect 8414 8813 8415 8847
rect 8449 8813 8450 8847
rect 8414 8779 8450 8813
rect 8414 8745 8415 8779
rect 8449 8745 8450 8779
rect 1680 8710 1681 8742
rect 1645 8676 1681 8710
rect 1645 8642 1646 8676
rect 1680 8642 1681 8676
rect 1808 8658 1824 8692
rect 1858 8658 1892 8692
rect 1926 8658 1986 8692
rect 2020 8658 2054 8692
rect 2088 8658 2104 8692
rect 2193 8658 2209 8692
rect 2243 8658 2277 8692
rect 2311 8658 2327 8692
rect 2449 8658 2465 8692
rect 2499 8658 2533 8692
rect 2567 8658 2583 8692
rect 2705 8658 2721 8692
rect 2755 8658 2789 8692
rect 2823 8658 2839 8692
rect 2961 8658 2977 8692
rect 3011 8658 3045 8692
rect 3079 8658 3095 8692
rect 3217 8658 3233 8692
rect 3267 8658 3301 8692
rect 3335 8658 3351 8692
rect 3473 8658 3489 8692
rect 3523 8658 3557 8692
rect 3591 8658 3607 8692
rect 3729 8658 3745 8692
rect 3779 8658 3813 8692
rect 3847 8658 3863 8692
rect 3985 8658 4001 8692
rect 4035 8658 4069 8692
rect 4103 8658 4119 8692
rect 4235 8658 4251 8692
rect 4285 8658 4301 8692
rect 8414 8677 8450 8745
rect 1645 8608 1681 8642
rect 1645 8574 1646 8608
rect 1680 8574 1681 8608
rect 1905 8624 2011 8658
rect 1939 8590 1977 8624
rect 4251 8612 4285 8658
rect 1645 8540 1681 8574
rect 1645 8506 1646 8540
rect 1680 8506 1681 8540
rect 4251 8540 4285 8578
rect 8414 8643 8415 8677
rect 8449 8643 8450 8677
rect 8414 8553 8450 8643
rect 1645 8472 1681 8506
rect 1645 8438 1646 8472
rect 1680 8438 1681 8472
rect 1645 8404 1681 8438
rect 1645 8370 1646 8404
rect 1680 8370 1681 8404
rect 1645 8336 1681 8370
rect 1645 8302 1646 8336
rect 1680 8302 1681 8336
rect 1645 8268 1681 8302
rect 1645 8234 1646 8268
rect 1680 8234 1681 8268
rect 1645 8200 1681 8234
rect 1645 8166 1646 8200
rect 1680 8166 1681 8200
rect 1645 8132 1681 8166
rect 1645 8098 1646 8132
rect 1680 8098 1681 8132
rect 1645 8064 1681 8098
rect 1645 8030 1646 8064
rect 1680 8030 1681 8064
rect 1645 7996 1681 8030
rect 1645 7962 1646 7996
rect 1680 7962 1681 7996
rect 1645 7928 1681 7962
rect 1645 7894 1646 7928
rect 1680 7894 1681 7928
rect 1645 7860 1681 7894
rect 1645 7826 1646 7860
rect 1680 7826 1681 7860
rect 1645 7792 1681 7826
rect 1645 7758 1646 7792
rect 1680 7758 1681 7792
rect 1645 7724 1681 7758
rect 1645 7690 1646 7724
rect 1680 7690 1681 7724
rect 1645 7656 1681 7690
rect 1645 7622 1646 7656
rect 1680 7622 1681 7656
rect 1645 7588 1681 7622
rect 1645 7554 1646 7588
rect 1680 7554 1681 7588
rect 1645 7511 1681 7554
rect 1645 7510 4139 7511
rect 1645 7476 1679 7510
rect 1713 7476 1747 7510
rect 1781 7476 1815 7510
rect 1849 7476 1883 7510
rect 1917 7476 1951 7510
rect 1985 7476 2019 7510
rect 2053 7476 2087 7510
rect 2121 7476 2155 7510
rect 2189 7476 2223 7510
rect 2257 7476 2291 7510
rect 2325 7476 2359 7510
rect 2393 7476 2427 7510
rect 2461 7476 2495 7510
rect 2529 7476 2563 7510
rect 2597 7476 2631 7510
rect 2665 7476 2699 7510
rect 2733 7476 2767 7510
rect 2801 7476 2835 7510
rect 2869 7476 2903 7510
rect 2937 7476 2971 7510
rect 3005 7476 3039 7510
rect 3073 7476 3107 7510
rect 3141 7476 3175 7510
rect 3209 7476 3243 7510
rect 3277 7476 3311 7510
rect 3345 7476 3379 7510
rect 3413 7476 3447 7510
rect 3481 7476 3515 7510
rect 3549 7476 3583 7510
rect 3617 7476 3651 7510
rect 3685 7476 3719 7510
rect 3753 7476 3787 7510
rect 3821 7476 3855 7510
rect 3889 7476 3923 7510
rect 3957 7476 3991 7510
rect 4025 7476 4059 7510
rect 4093 7476 4139 7510
rect 1645 7475 4139 7476
rect 1456 7322 1492 7445
rect 1456 7321 4128 7322
rect 1456 7287 1490 7321
rect 1524 7287 1558 7321
rect 1592 7287 1626 7321
rect 1660 7287 1694 7321
rect 1728 7287 1762 7321
rect 1796 7287 1830 7321
rect 1864 7287 1898 7321
rect 1932 7287 1966 7321
rect 2000 7287 2034 7321
rect 2068 7287 2102 7321
rect 2136 7287 2170 7321
rect 2204 7287 2238 7321
rect 2272 7287 2306 7321
rect 2340 7287 2374 7321
rect 2408 7287 2442 7321
rect 2476 7287 2510 7321
rect 2544 7287 2578 7321
rect 2612 7287 2646 7321
rect 2680 7287 2714 7321
rect 2748 7287 2782 7321
rect 2816 7287 2850 7321
rect 2884 7287 2918 7321
rect 2952 7287 2986 7321
rect 3020 7287 3054 7321
rect 3088 7287 3122 7321
rect 3156 7287 3190 7321
rect 3224 7287 3258 7321
rect 3292 7287 3326 7321
rect 3360 7287 3394 7321
rect 3428 7287 3462 7321
rect 3496 7287 3530 7321
rect 3564 7287 3598 7321
rect 3632 7287 3666 7321
rect 3700 7287 3734 7321
rect 3768 7287 3802 7321
rect 3836 7287 3870 7321
rect 3904 7287 3938 7321
rect 3972 7287 4006 7321
rect 4040 7287 4128 7321
rect 1456 7286 4128 7287
rect 1456 7252 1492 7286
rect 1456 7218 1457 7252
rect 1491 7218 1492 7252
rect 1456 7184 1492 7218
rect 1456 7150 1457 7184
rect 1491 7150 1492 7184
rect 1456 7116 1492 7150
rect 1456 7082 1457 7116
rect 1491 7082 1492 7116
rect 4092 7226 4128 7286
rect 4092 7192 4093 7226
rect 4127 7192 4128 7226
rect 4092 7158 4128 7192
rect 4092 7124 4093 7158
rect 4127 7124 4128 7158
rect 1456 7048 1492 7082
rect 1456 7014 1457 7048
rect 1491 7014 1492 7048
rect 1456 6980 1492 7014
rect 1456 6946 1457 6980
rect 1491 6946 1492 6980
rect 1456 6912 1492 6946
rect 1456 6878 1457 6912
rect 1491 6878 1492 6912
rect 1456 6844 1492 6878
rect 1456 6810 1457 6844
rect 1491 6810 1492 6844
rect 1456 6776 1492 6810
rect 1456 6742 1457 6776
rect 1491 6742 1492 6776
rect 1456 6708 1492 6742
rect 1456 6674 1457 6708
rect 1491 6674 1492 6708
rect 1456 6640 1492 6674
rect 1456 6606 1457 6640
rect 1491 6606 1492 6640
rect 1456 6572 1492 6606
rect 1456 6538 1457 6572
rect 1491 6538 1492 6572
rect 1456 6504 1492 6538
rect 1456 6470 1457 6504
rect 1491 6470 1492 6504
rect 1456 6436 1492 6470
rect 1456 6402 1457 6436
rect 1491 6402 1492 6436
rect 1456 6368 1492 6402
rect 1456 6334 1457 6368
rect 1491 6334 1492 6368
rect 1456 6300 1492 6334
rect 1456 6266 1457 6300
rect 1491 6266 1492 6300
rect 1456 6232 1492 6266
rect 1456 6198 1457 6232
rect 1491 6198 1492 6232
rect 1456 6164 1492 6198
rect 1456 6130 1457 6164
rect 1491 6130 1492 6164
rect 1456 6096 1492 6130
rect 1456 6062 1457 6096
rect 1491 6062 1492 6096
rect 1456 6028 1492 6062
rect 1456 5994 1457 6028
rect 1491 5994 1492 6028
rect 1456 5960 1492 5994
rect 1456 5926 1457 5960
rect 1491 5926 1492 5960
rect 1456 5892 1492 5926
rect 1456 5858 1457 5892
rect 1491 5858 1492 5892
rect 1456 5824 1492 5858
rect 1456 5790 1457 5824
rect 1491 5790 1492 5824
rect 1456 5756 1492 5790
rect 1456 5722 1457 5756
rect 1491 5722 1492 5756
rect 1456 5688 1492 5722
rect 1456 5654 1457 5688
rect 1491 5654 1492 5688
rect 1456 5620 1492 5654
rect 1456 5586 1457 5620
rect 1491 5586 1492 5620
rect 1456 5552 1492 5586
rect 1456 5518 1457 5552
rect 1491 5518 1492 5552
rect 1456 5484 1492 5518
rect 1456 5450 1457 5484
rect 1491 5450 1492 5484
rect 1456 5416 1492 5450
rect 1456 5382 1457 5416
rect 1491 5382 1492 5416
rect 1456 5348 1492 5382
rect 1456 5314 1457 5348
rect 1491 5314 1492 5348
rect 1456 5280 1492 5314
rect 1456 5246 1457 5280
rect 1491 5246 1492 5280
rect 1456 5212 1492 5246
rect 1456 5178 1457 5212
rect 1491 5178 1492 5212
rect 1456 5144 1492 5178
rect 1456 5110 1457 5144
rect 1491 5110 1492 5144
rect 1456 5076 1492 5110
rect 1456 5042 1457 5076
rect 1491 5042 1492 5076
rect 1456 5008 1492 5042
rect 1456 4974 1457 5008
rect 1491 4974 1492 5008
rect 1456 4940 1492 4974
rect 1456 4906 1457 4940
rect 1491 4906 1492 4940
rect 1456 4872 1492 4906
rect 1456 4838 1457 4872
rect 1491 4838 1492 4872
rect 1456 4804 1492 4838
rect 1456 4770 1457 4804
rect 1491 4770 1492 4804
rect 1456 4736 1492 4770
rect 1456 4702 1457 4736
rect 1491 4702 1492 4736
rect 1456 4668 1492 4702
rect 1456 4634 1457 4668
rect 1491 4634 1492 4668
rect 1456 4600 1492 4634
rect 1456 4566 1457 4600
rect 1491 4566 1492 4600
rect 1456 4532 1492 4566
rect 1456 4498 1457 4532
rect 1491 4498 1492 4532
rect 1456 4464 1492 4498
rect 1456 4430 1457 4464
rect 1491 4430 1492 4464
rect 1456 4396 1492 4430
rect 1456 4362 1457 4396
rect 1491 4362 1492 4396
rect 1456 4328 1492 4362
rect 1456 4294 1457 4328
rect 1491 4294 1492 4328
rect 1456 4260 1492 4294
rect 1456 4226 1457 4260
rect 1491 4226 1492 4260
rect 1456 4192 1492 4226
rect 1456 4158 1457 4192
rect 1491 4158 1492 4192
rect 1456 4124 1492 4158
rect 1456 4090 1457 4124
rect 1491 4090 1492 4124
rect 1456 4056 1492 4090
rect 1456 4022 1457 4056
rect 1491 4022 1492 4056
rect 1456 3988 1492 4022
rect 1456 3954 1457 3988
rect 1491 3954 1492 3988
rect 1456 3920 1492 3954
rect 1456 3886 1457 3920
rect 1491 3886 1492 3920
rect 1456 3852 1492 3886
rect 1456 3818 1457 3852
rect 1491 3818 1492 3852
rect 1456 3784 1492 3818
rect 1456 3750 1457 3784
rect 1491 3750 1492 3784
rect 1456 3716 1492 3750
rect 1456 3682 1457 3716
rect 1491 3682 1492 3716
rect 1456 3648 1492 3682
rect 1456 3614 1457 3648
rect 1491 3614 1492 3648
rect 1456 3580 1492 3614
rect 1456 3546 1457 3580
rect 1491 3546 1492 3580
rect 1456 3512 1492 3546
rect 1456 3478 1457 3512
rect 1491 3478 1492 3512
rect 1456 3444 1492 3478
rect 1456 3410 1457 3444
rect 1491 3410 1492 3444
rect 1456 3376 1492 3410
rect 1456 3342 1457 3376
rect 1491 3342 1492 3376
rect 1456 3308 1492 3342
rect 1456 3274 1457 3308
rect 1491 3274 1492 3308
rect 1456 3240 1492 3274
rect 1456 3206 1457 3240
rect 1491 3206 1492 3240
rect 1456 3172 1492 3206
rect 1456 3138 1457 3172
rect 1491 3138 1492 3172
rect 1456 3104 1492 3138
rect 1456 3070 1457 3104
rect 1491 3070 1492 3104
rect 1456 3036 1492 3070
rect 1456 3002 1457 3036
rect 1491 3002 1492 3036
rect 1456 2968 1492 3002
rect 1456 2934 1457 2968
rect 1491 2934 1492 2968
rect 1456 2900 1492 2934
rect 1456 2866 1457 2900
rect 1491 2866 1492 2900
rect 1456 2832 1492 2866
rect 1456 2798 1457 2832
rect 1491 2798 1492 2832
rect 1456 2764 1492 2798
rect 1456 2730 1457 2764
rect 1491 2730 1492 2764
rect 1456 2696 1492 2730
rect 1456 2662 1457 2696
rect 1491 2662 1492 2696
rect 1456 2628 1492 2662
rect 1456 2594 1457 2628
rect 1491 2594 1492 2628
rect 1456 2560 1492 2594
rect 1456 2526 1457 2560
rect 1491 2526 1492 2560
rect 1456 2492 1492 2526
rect 1456 2458 1457 2492
rect 1491 2458 1492 2492
rect 1456 2424 1492 2458
rect 1456 2390 1457 2424
rect 1491 2390 1492 2424
rect 1456 2356 1492 2390
rect 1456 2322 1457 2356
rect 1491 2322 1492 2356
rect 1456 2288 1492 2322
rect 1456 2254 1457 2288
rect 1491 2254 1492 2288
rect 1645 7110 3939 7111
rect 1645 7077 1763 7110
rect 1645 7043 1646 7077
rect 1680 7076 1763 7077
rect 1797 7076 1831 7110
rect 1865 7076 1899 7110
rect 1933 7076 1967 7110
rect 2001 7076 2035 7110
rect 2069 7076 2103 7110
rect 2137 7076 2171 7110
rect 2205 7076 2239 7110
rect 2273 7076 2307 7110
rect 2341 7076 2375 7110
rect 2409 7076 2443 7110
rect 2477 7076 2511 7110
rect 2545 7076 2579 7110
rect 2613 7076 2647 7110
rect 2681 7076 2715 7110
rect 2749 7076 2783 7110
rect 2817 7076 2851 7110
rect 2885 7076 2919 7110
rect 2953 7076 2987 7110
rect 3021 7076 3055 7110
rect 3089 7076 3123 7110
rect 3157 7076 3191 7110
rect 3225 7076 3259 7110
rect 3293 7076 3327 7110
rect 3361 7076 3395 7110
rect 3429 7076 3463 7110
rect 3497 7076 3531 7110
rect 3565 7076 3599 7110
rect 3633 7076 3667 7110
rect 3701 7076 3735 7110
rect 3769 7076 3803 7110
rect 3837 7076 3871 7110
rect 3905 7076 3939 7110
rect 1680 7075 3939 7076
rect 1680 7043 1681 7075
rect 1645 7009 1681 7043
rect 1645 6975 1646 7009
rect 1680 6975 1681 7009
rect 1742 7025 1892 7041
rect 1742 7005 1790 7025
rect 1645 6941 1681 6975
rect 1645 6907 1646 6941
rect 1680 6907 1681 6941
rect 1645 6873 1681 6907
rect 1763 6991 1790 7005
rect 1824 6991 1858 7025
rect 1763 6975 1892 6991
rect 3692 7025 3842 7041
rect 3726 6991 3760 7025
rect 3794 7005 3842 7025
rect 3903 7035 3939 7075
rect 3794 6991 3821 7005
rect 3692 6975 3821 6991
rect 1763 6889 1797 6975
rect 3787 6889 3821 6975
rect 3903 7001 3904 7035
rect 3938 7001 3939 7035
rect 3903 6967 3939 7001
rect 3903 6933 3904 6967
rect 3938 6933 3939 6967
rect 3903 6899 3939 6933
rect 1645 6839 1646 6873
rect 1680 6839 1681 6873
rect 1645 6805 1681 6839
rect 1645 6771 1646 6805
rect 1680 6771 1681 6805
rect 1645 6737 1681 6771
rect 1645 6703 1646 6737
rect 1680 6703 1681 6737
rect 1645 6669 1681 6703
rect 1645 6635 1646 6669
rect 1680 6635 1681 6669
rect 1645 6601 1681 6635
rect 1645 6567 1646 6601
rect 1680 6567 1681 6601
rect 1645 6533 1681 6567
rect 1645 6499 1646 6533
rect 1680 6499 1681 6533
rect 1645 6465 1681 6499
rect 1645 6431 1646 6465
rect 1680 6431 1681 6465
rect 1645 6397 1681 6431
rect 1645 6363 1646 6397
rect 1680 6363 1681 6397
rect 1645 6329 1681 6363
rect 1645 6295 1646 6329
rect 1680 6295 1681 6329
rect 1645 6261 1681 6295
rect 1645 6227 1646 6261
rect 1680 6227 1681 6261
rect 1645 6193 1681 6227
rect 1645 6159 1646 6193
rect 1680 6159 1681 6193
rect 1645 6125 1681 6159
rect 1645 6091 1646 6125
rect 1680 6091 1681 6125
rect 1645 6057 1681 6091
rect 1645 6023 1646 6057
rect 1680 6023 1681 6057
rect 1645 5989 1681 6023
rect 1645 5955 1646 5989
rect 1680 5955 1681 5989
rect 1645 5921 1681 5955
rect 3903 6865 3904 6899
rect 3938 6865 3939 6899
rect 3903 6831 3939 6865
rect 3903 6797 3904 6831
rect 3938 6797 3939 6831
rect 3903 6763 3939 6797
rect 3903 6729 3904 6763
rect 3938 6729 3939 6763
rect 3903 6695 3939 6729
rect 3903 6661 3904 6695
rect 3938 6661 3939 6695
rect 3903 6627 3939 6661
rect 3903 6593 3904 6627
rect 3938 6593 3939 6627
rect 3903 6559 3939 6593
rect 3903 6525 3904 6559
rect 3938 6525 3939 6559
rect 3903 6491 3939 6525
rect 3903 6457 3904 6491
rect 3938 6457 3939 6491
rect 3903 6423 3939 6457
rect 3903 6389 3904 6423
rect 3938 6389 3939 6423
rect 3903 6355 3939 6389
rect 3903 6321 3904 6355
rect 3938 6321 3939 6355
rect 3903 6287 3939 6321
rect 3903 6253 3904 6287
rect 3938 6253 3939 6287
rect 3903 6219 3939 6253
rect 3903 6185 3904 6219
rect 3938 6185 3939 6219
rect 3903 6151 3939 6185
rect 3903 6117 3904 6151
rect 3938 6117 3939 6151
rect 3903 6083 3939 6117
rect 3903 6049 3904 6083
rect 3938 6049 3939 6083
rect 3903 6015 3939 6049
rect 3903 5981 3904 6015
rect 3938 5981 3939 6015
rect 3903 5947 3939 5981
rect 1645 5887 1646 5921
rect 1680 5887 1681 5921
rect 1645 5853 1681 5887
rect 1645 5819 1646 5853
rect 1680 5819 1681 5853
rect 1645 5785 1681 5819
rect 1645 5751 1646 5785
rect 1680 5751 1681 5785
rect 1645 5717 1681 5751
rect 1645 5683 1646 5717
rect 1680 5683 1681 5717
rect 1763 5849 1797 5939
rect 3787 5849 3821 5939
rect 1763 5833 1892 5849
rect 1763 5799 1790 5833
rect 1824 5799 1858 5833
rect 1763 5783 1892 5799
rect 3692 5833 3821 5849
rect 3726 5799 3760 5833
rect 3794 5799 3821 5833
rect 3692 5783 3821 5799
rect 1763 5697 1797 5783
rect 3787 5697 3821 5783
rect 3903 5913 3904 5947
rect 3938 5913 3939 5947
rect 3903 5879 3939 5913
rect 3903 5845 3904 5879
rect 3938 5845 3939 5879
rect 3903 5811 3939 5845
rect 3903 5777 3904 5811
rect 3938 5777 3939 5811
rect 3903 5743 3939 5777
rect 3903 5709 3904 5743
rect 3938 5709 3939 5743
rect 1645 5649 1681 5683
rect 1645 5615 1646 5649
rect 1680 5615 1681 5649
rect 1645 5581 1681 5615
rect 1645 5547 1646 5581
rect 1680 5547 1681 5581
rect 1645 5513 1681 5547
rect 1645 5479 1646 5513
rect 1680 5479 1681 5513
rect 1645 5445 1681 5479
rect 1645 5411 1646 5445
rect 1680 5411 1681 5445
rect 1645 5377 1681 5411
rect 1645 5343 1646 5377
rect 1680 5343 1681 5377
rect 1645 5309 1681 5343
rect 1645 5275 1646 5309
rect 1680 5275 1681 5309
rect 1645 5241 1681 5275
rect 1645 5207 1646 5241
rect 1680 5207 1681 5241
rect 1645 5173 1681 5207
rect 1645 5139 1646 5173
rect 1680 5139 1681 5173
rect 1645 5105 1681 5139
rect 1645 5071 1646 5105
rect 1680 5071 1681 5105
rect 1645 5037 1681 5071
rect 1645 5003 1646 5037
rect 1680 5003 1681 5037
rect 1645 4969 1681 5003
rect 1645 4935 1646 4969
rect 1680 4935 1681 4969
rect 1645 4901 1681 4935
rect 1645 4867 1646 4901
rect 1680 4867 1681 4901
rect 1645 4833 1681 4867
rect 1645 4799 1646 4833
rect 1680 4799 1681 4833
rect 1645 4765 1681 4799
rect 1645 4731 1646 4765
rect 1680 4731 1681 4765
rect 3903 5675 3939 5709
rect 3903 5641 3904 5675
rect 3938 5641 3939 5675
rect 3903 5607 3939 5641
rect 3903 5573 3904 5607
rect 3938 5573 3939 5607
rect 3903 5539 3939 5573
rect 3903 5505 3904 5539
rect 3938 5505 3939 5539
rect 3903 5471 3939 5505
rect 3903 5437 3904 5471
rect 3938 5437 3939 5471
rect 3903 5403 3939 5437
rect 3903 5369 3904 5403
rect 3938 5369 3939 5403
rect 3903 5335 3939 5369
rect 3903 5301 3904 5335
rect 3938 5301 3939 5335
rect 3903 5267 3939 5301
rect 3903 5233 3904 5267
rect 3938 5233 3939 5267
rect 3903 5199 3939 5233
rect 3903 5165 3904 5199
rect 3938 5165 3939 5199
rect 3903 5131 3939 5165
rect 3903 5097 3904 5131
rect 3938 5097 3939 5131
rect 3903 5063 3939 5097
rect 3903 5029 3904 5063
rect 3938 5029 3939 5063
rect 3903 4995 3939 5029
rect 3903 4961 3904 4995
rect 3938 4961 3939 4995
rect 3903 4927 3939 4961
rect 3903 4893 3904 4927
rect 3938 4893 3939 4927
rect 3903 4859 3939 4893
rect 3903 4825 3904 4859
rect 3938 4825 3939 4859
rect 3903 4791 3939 4825
rect 3903 4757 3904 4791
rect 3938 4757 3939 4791
rect 1645 4697 1681 4731
rect 1645 4663 1646 4697
rect 1680 4663 1681 4697
rect 1645 4629 1681 4663
rect 1645 4595 1646 4629
rect 1680 4595 1681 4629
rect 1645 4561 1681 4595
rect 1645 4527 1646 4561
rect 1680 4527 1681 4561
rect 1645 4493 1681 4527
rect 1763 4657 1797 4747
rect 3787 4657 3821 4747
rect 1763 4641 1892 4657
rect 1763 4607 1790 4641
rect 1824 4607 1858 4641
rect 1763 4591 1892 4607
rect 3692 4641 3821 4657
rect 3726 4607 3760 4641
rect 3794 4607 3821 4641
rect 3692 4591 3821 4607
rect 1763 4505 1797 4591
rect 3787 4505 3821 4591
rect 3903 4723 3939 4757
rect 3903 4689 3904 4723
rect 3938 4689 3939 4723
rect 3903 4655 3939 4689
rect 3903 4621 3904 4655
rect 3938 4621 3939 4655
rect 3903 4587 3939 4621
rect 3903 4553 3904 4587
rect 3938 4553 3939 4587
rect 3903 4519 3939 4553
rect 1645 4459 1646 4493
rect 1680 4459 1681 4493
rect 1645 4425 1681 4459
rect 1645 4391 1646 4425
rect 1680 4391 1681 4425
rect 1645 4357 1681 4391
rect 1645 4323 1646 4357
rect 1680 4323 1681 4357
rect 1645 4289 1681 4323
rect 1645 4255 1646 4289
rect 1680 4255 1681 4289
rect 1645 4221 1681 4255
rect 1645 4187 1646 4221
rect 1680 4187 1681 4221
rect 1645 4153 1681 4187
rect 1645 4119 1646 4153
rect 1680 4119 1681 4153
rect 1645 4085 1681 4119
rect 1645 4051 1646 4085
rect 1680 4051 1681 4085
rect 1645 4017 1681 4051
rect 1645 3983 1646 4017
rect 1680 3983 1681 4017
rect 1645 3949 1681 3983
rect 1645 3915 1646 3949
rect 1680 3915 1681 3949
rect 1645 3881 1681 3915
rect 1645 3847 1646 3881
rect 1680 3847 1681 3881
rect 1645 3813 1681 3847
rect 1645 3779 1646 3813
rect 1680 3779 1681 3813
rect 1645 3745 1681 3779
rect 1645 3711 1646 3745
rect 1680 3711 1681 3745
rect 1645 3677 1681 3711
rect 1645 3643 1646 3677
rect 1680 3643 1681 3677
rect 1645 3609 1681 3643
rect 1645 3575 1646 3609
rect 1680 3575 1681 3609
rect 1645 3541 1681 3575
rect 3903 4485 3904 4519
rect 3938 4485 3939 4519
rect 3903 4451 3939 4485
rect 3903 4417 3904 4451
rect 3938 4417 3939 4451
rect 3903 4383 3939 4417
rect 3903 4349 3904 4383
rect 3938 4349 3939 4383
rect 3903 4315 3939 4349
rect 3903 4281 3904 4315
rect 3938 4281 3939 4315
rect 3903 4247 3939 4281
rect 3903 4213 3904 4247
rect 3938 4213 3939 4247
rect 3903 4179 3939 4213
rect 3903 4145 3904 4179
rect 3938 4145 3939 4179
rect 3903 4111 3939 4145
rect 3903 4077 3904 4111
rect 3938 4077 3939 4111
rect 3903 4043 3939 4077
rect 3903 4009 3904 4043
rect 3938 4009 3939 4043
rect 3903 3975 3939 4009
rect 3903 3941 3904 3975
rect 3938 3941 3939 3975
rect 3903 3907 3939 3941
rect 3903 3873 3904 3907
rect 3938 3873 3939 3907
rect 3903 3839 3939 3873
rect 3903 3805 3904 3839
rect 3938 3805 3939 3839
rect 3903 3771 3939 3805
rect 3903 3737 3904 3771
rect 3938 3737 3939 3771
rect 3903 3703 3939 3737
rect 3903 3669 3904 3703
rect 3938 3669 3939 3703
rect 3903 3635 3939 3669
rect 3903 3601 3904 3635
rect 3938 3601 3939 3635
rect 3903 3567 3939 3601
rect 1645 3507 1646 3541
rect 1680 3507 1681 3541
rect 1645 3473 1681 3507
rect 1645 3439 1646 3473
rect 1680 3439 1681 3473
rect 1645 3405 1681 3439
rect 1645 3371 1646 3405
rect 1680 3371 1681 3405
rect 1645 3337 1681 3371
rect 1645 3303 1646 3337
rect 1680 3303 1681 3337
rect 1763 3465 1797 3555
rect 3787 3518 3821 3555
rect 3903 3533 3904 3567
rect 3938 3533 3939 3567
rect 3903 3499 3939 3533
rect 4092 7090 4128 7124
rect 4092 7056 4093 7090
rect 4127 7056 4128 7090
rect 4092 7022 4128 7056
rect 4092 6988 4093 7022
rect 4127 6988 4128 7022
rect 4092 6954 4128 6988
rect 4092 6920 4093 6954
rect 4127 6920 4128 6954
rect 4092 6886 4128 6920
rect 4092 6852 4093 6886
rect 4127 6852 4128 6886
rect 4092 6818 4128 6852
rect 4092 6784 4093 6818
rect 4127 6784 4128 6818
rect 4092 6750 4128 6784
rect 4092 6716 4093 6750
rect 4127 6716 4128 6750
rect 4092 6682 4128 6716
rect 4092 6648 4093 6682
rect 4127 6648 4128 6682
rect 4092 6614 4128 6648
rect 4092 6580 4093 6614
rect 4127 6580 4128 6614
rect 4092 6546 4128 6580
rect 4092 6512 4093 6546
rect 4127 6512 4128 6546
rect 4092 6478 4128 6512
rect 4092 6444 4093 6478
rect 4127 6444 4128 6478
rect 4092 6410 4128 6444
rect 4092 6376 4093 6410
rect 4127 6376 4128 6410
rect 4092 6342 4128 6376
rect 4092 6308 4093 6342
rect 4127 6308 4128 6342
rect 4092 6274 4128 6308
rect 4092 6240 4093 6274
rect 4127 6240 4128 6274
rect 4092 6206 4128 6240
rect 4092 6172 4093 6206
rect 4127 6172 4128 6206
rect 4092 6138 4128 6172
rect 4092 6104 4093 6138
rect 4127 6104 4128 6138
rect 4092 6070 4128 6104
rect 4092 6036 4093 6070
rect 4127 6036 4128 6070
rect 4092 6002 4128 6036
rect 4092 5968 4093 6002
rect 4127 5968 4128 6002
rect 4092 5934 4128 5968
rect 4092 5900 4093 5934
rect 4127 5900 4128 5934
rect 4092 5866 4128 5900
rect 4092 5832 4093 5866
rect 4127 5832 4128 5866
rect 4092 5798 4128 5832
rect 4092 5764 4093 5798
rect 4127 5764 4128 5798
rect 4092 5730 4128 5764
rect 4092 5696 4093 5730
rect 4127 5696 4128 5730
rect 4092 5662 4128 5696
rect 4092 5628 4093 5662
rect 4127 5628 4128 5662
rect 4092 5594 4128 5628
rect 4092 5560 4093 5594
rect 4127 5560 4128 5594
rect 4092 5526 4128 5560
rect 4092 5492 4093 5526
rect 4127 5492 4128 5526
rect 4092 5458 4128 5492
rect 4092 5424 4093 5458
rect 4127 5424 4128 5458
rect 4092 5390 4128 5424
rect 4092 5356 4093 5390
rect 4127 5356 4128 5390
rect 4092 5322 4128 5356
rect 4092 5288 4093 5322
rect 4127 5288 4128 5322
rect 4092 5254 4128 5288
rect 4092 5220 4093 5254
rect 4127 5220 4128 5254
rect 4092 5186 4128 5220
rect 4092 5152 4093 5186
rect 4127 5152 4128 5186
rect 4092 5118 4128 5152
rect 4092 5084 4093 5118
rect 4127 5084 4128 5118
rect 4092 5050 4128 5084
rect 4092 5016 4093 5050
rect 4127 5016 4128 5050
rect 4092 4982 4128 5016
rect 4092 4948 4093 4982
rect 4127 4948 4128 4982
rect 4092 4914 4128 4948
rect 4092 4880 4093 4914
rect 4127 4880 4128 4914
rect 4092 4846 4128 4880
rect 4092 4812 4093 4846
rect 4127 4812 4128 4846
rect 4092 4778 4128 4812
rect 4092 4744 4093 4778
rect 4127 4744 4128 4778
rect 4092 4710 4128 4744
rect 4092 4676 4093 4710
rect 4127 4676 4128 4710
rect 4092 4642 4128 4676
rect 4092 4608 4093 4642
rect 4127 4608 4128 4642
rect 4092 4574 4128 4608
rect 4092 4540 4093 4574
rect 4127 4540 4128 4574
rect 4092 4506 4128 4540
rect 4092 4472 4093 4506
rect 4127 4472 4128 4506
rect 4092 4438 4128 4472
rect 4092 4404 4093 4438
rect 4127 4404 4128 4438
rect 4092 4370 4128 4404
rect 4092 4336 4093 4370
rect 4127 4336 4128 4370
rect 4092 4302 4128 4336
rect 4092 4268 4093 4302
rect 4127 4268 4128 4302
rect 4092 4234 4128 4268
rect 4092 4200 4093 4234
rect 4127 4200 4128 4234
rect 4092 4166 4128 4200
rect 4092 4132 4093 4166
rect 4127 4132 4128 4166
rect 4092 4098 4128 4132
rect 4092 4064 4093 4098
rect 4127 4064 4128 4098
rect 4092 4030 4128 4064
rect 4092 3996 4093 4030
rect 4127 3996 4128 4030
rect 4092 3962 4128 3996
rect 4092 3928 4093 3962
rect 4127 3928 4128 3962
rect 4092 3894 4128 3928
rect 4092 3860 4093 3894
rect 4127 3860 4128 3894
rect 4092 3826 4128 3860
rect 4092 3792 4093 3826
rect 4127 3792 4128 3826
rect 4092 3758 4128 3792
rect 4092 3724 4093 3758
rect 4127 3724 4128 3758
rect 4092 3690 4128 3724
rect 4092 3656 4093 3690
rect 4127 3656 4128 3690
rect 4092 3622 4128 3656
rect 4092 3588 4093 3622
rect 4127 3588 4128 3622
rect 4092 3554 4128 3588
rect 4092 3520 4093 3554
rect 4127 3520 4128 3554
rect 4092 3486 4128 3520
rect 1763 3449 1892 3465
rect 1763 3415 1790 3449
rect 1824 3415 1858 3449
rect 1763 3399 1892 3415
rect 3692 3453 4033 3465
rect 3692 3449 3999 3453
rect 3726 3415 3760 3449
rect 3794 3419 3999 3449
rect 3794 3415 4033 3419
rect 3692 3399 4033 3415
rect 1763 3313 1797 3399
rect 3999 3381 4033 3399
rect 3787 3313 3821 3333
rect 1645 3269 1681 3303
rect 1645 3235 1646 3269
rect 1680 3235 1681 3269
rect 1645 3201 1681 3235
rect 1645 3167 1646 3201
rect 1680 3167 1681 3201
rect 1645 3133 1681 3167
rect 1645 3099 1646 3133
rect 1680 3099 1681 3133
rect 1645 3065 1681 3099
rect 1645 3031 1646 3065
rect 1680 3031 1681 3065
rect 1645 2997 1681 3031
rect 1645 2963 1646 2997
rect 1680 2963 1681 2997
rect 1645 2929 1681 2963
rect 1645 2895 1646 2929
rect 1680 2895 1681 2929
rect 1645 2861 1681 2895
rect 1645 2827 1646 2861
rect 1680 2827 1681 2861
rect 1645 2793 1681 2827
rect 1645 2759 1646 2793
rect 1680 2759 1681 2793
rect 1645 2725 1681 2759
rect 1645 2691 1646 2725
rect 1680 2691 1681 2725
rect 1645 2657 1681 2691
rect 1645 2623 1646 2657
rect 1680 2623 1681 2657
rect 1645 2589 1681 2623
rect 1645 2555 1646 2589
rect 1680 2555 1681 2589
rect 1645 2521 1681 2555
rect 1645 2487 1646 2521
rect 1680 2487 1681 2521
rect 1645 2453 1681 2487
rect 1645 2419 1646 2453
rect 1680 2419 1681 2453
rect 1645 2293 1681 2419
rect 3903 3277 3939 3348
rect 4092 3452 4093 3486
rect 4127 3452 4128 3486
rect 4092 3418 4128 3452
rect 4092 3384 4093 3418
rect 4127 3384 4128 3418
rect 4092 3350 4128 3384
rect 3903 3243 3904 3277
rect 3938 3243 3939 3277
rect 3903 3209 3939 3243
rect 3903 3175 3904 3209
rect 3938 3175 3939 3209
rect 3903 3141 3939 3175
rect 3903 3107 3904 3141
rect 3938 3107 3939 3141
rect 3903 3073 3939 3107
rect 3903 3039 3904 3073
rect 3938 3039 3939 3073
rect 3903 3005 3939 3039
rect 3903 2971 3904 3005
rect 3938 2971 3939 3005
rect 3903 2937 3939 2971
rect 3903 2903 3904 2937
rect 3938 2903 3939 2937
rect 3903 2869 3939 2903
rect 3903 2835 3904 2869
rect 3938 2835 3939 2869
rect 3903 2801 3939 2835
rect 3903 2767 3904 2801
rect 3938 2767 3939 2801
rect 3903 2733 3939 2767
rect 3903 2699 3904 2733
rect 3938 2699 3939 2733
rect 3903 2665 3939 2699
rect 3903 2631 3904 2665
rect 3938 2631 3939 2665
rect 3903 2597 3939 2631
rect 3903 2563 3904 2597
rect 3938 2563 3939 2597
rect 3903 2529 3939 2563
rect 3903 2495 3904 2529
rect 3938 2495 3939 2529
rect 3903 2461 3939 2495
rect 3903 2427 3904 2461
rect 3938 2427 3939 2461
rect 3903 2393 3939 2427
rect 3903 2359 3904 2393
rect 3938 2359 3939 2393
rect 3903 2325 3939 2359
rect 3903 2293 3904 2325
rect 1645 2292 3904 2293
rect 1645 2258 1679 2292
rect 1713 2258 1747 2292
rect 1793 2258 1815 2292
rect 1865 2258 1883 2292
rect 1917 2258 1951 2292
rect 1985 2258 2019 2292
rect 2053 2258 2087 2292
rect 2121 2258 2155 2292
rect 2189 2258 2223 2292
rect 2257 2258 2291 2292
rect 2325 2258 2359 2292
rect 2393 2258 2427 2292
rect 2461 2258 2495 2292
rect 2529 2258 2563 2292
rect 2597 2258 2631 2292
rect 2665 2258 2699 2292
rect 2733 2258 2767 2292
rect 2801 2258 2835 2292
rect 2869 2258 2903 2292
rect 2937 2258 2971 2292
rect 3005 2258 3039 2292
rect 3073 2258 3107 2292
rect 3141 2258 3175 2292
rect 3209 2258 3243 2292
rect 3277 2258 3311 2292
rect 3345 2258 3379 2292
rect 3413 2258 3447 2292
rect 3481 2258 3515 2292
rect 3549 2258 3583 2292
rect 3617 2258 3651 2292
rect 3685 2258 3719 2292
rect 3753 2258 3787 2292
rect 3825 2291 3904 2292
rect 3938 2291 3939 2325
rect 3825 2258 3939 2291
rect 1645 2257 3939 2258
rect 4092 3316 4093 3350
rect 4127 3316 4128 3350
rect 4092 3282 4128 3316
rect 4092 3248 4093 3282
rect 4127 3248 4128 3282
rect 4092 3214 4128 3248
rect 4092 3180 4093 3214
rect 4127 3180 4128 3214
rect 4092 3146 4128 3180
rect 4092 3112 4093 3146
rect 4127 3112 4128 3146
rect 4092 3078 4128 3112
rect 4092 3044 4093 3078
rect 4127 3044 4128 3078
rect 4092 3010 4128 3044
rect 4092 2976 4093 3010
rect 4127 2976 4128 3010
rect 4092 2942 4128 2976
rect 4092 2908 4093 2942
rect 4127 2908 4128 2942
rect 4092 2874 4128 2908
rect 4092 2840 4093 2874
rect 4127 2840 4128 2874
rect 4092 2806 4128 2840
rect 4092 2772 4093 2806
rect 4127 2772 4128 2806
rect 4092 2738 4128 2772
rect 4092 2704 4093 2738
rect 4127 2704 4128 2738
rect 4092 2670 4128 2704
rect 4092 2636 4093 2670
rect 4127 2636 4128 2670
rect 4092 2602 4128 2636
rect 4092 2568 4093 2602
rect 4127 2568 4128 2602
rect 4092 2534 4128 2568
rect 4092 2500 4093 2534
rect 4127 2500 4128 2534
rect 4092 2466 4128 2500
rect 4092 2432 4093 2466
rect 4127 2432 4128 2466
rect 4092 2398 4128 2432
rect 4092 2364 4093 2398
rect 4127 2364 4128 2398
rect 4092 2330 4128 2364
rect 4092 2296 4093 2330
rect 4127 2296 4128 2330
rect 4092 2262 4128 2296
rect 1456 2220 1492 2254
rect 1456 2186 1457 2220
rect 1491 2186 1492 2220
rect 1456 2152 1492 2186
rect 1456 2118 1457 2152
rect 1491 2118 1492 2152
rect 1456 2104 1492 2118
rect 4092 2228 4093 2262
rect 4127 2228 4128 2262
rect 4092 2194 4128 2228
rect 4092 2160 4093 2194
rect 4127 2160 4128 2194
rect 4092 2126 4128 2160
rect 4092 2104 4093 2126
rect 1456 2103 4093 2104
rect 1456 2069 1526 2103
rect 1560 2069 1594 2103
rect 1628 2069 1662 2103
rect 1696 2069 1730 2103
rect 1764 2069 1798 2103
rect 1836 2069 1866 2103
rect 1908 2069 1934 2103
rect 1980 2069 2002 2103
rect 2052 2069 2070 2103
rect 2104 2069 2138 2103
rect 2172 2069 2206 2103
rect 2240 2069 2274 2103
rect 2308 2069 2342 2103
rect 2376 2069 2410 2103
rect 2444 2069 2478 2103
rect 2512 2069 2546 2103
rect 2604 2069 2614 2103
rect 2676 2069 2682 2103
rect 2748 2069 2750 2103
rect 2784 2069 2786 2103
rect 2852 2069 2858 2103
rect 2920 2069 2930 2103
rect 2988 2069 3022 2103
rect 3056 2069 3090 2103
rect 3124 2069 3158 2103
rect 3192 2069 3226 2103
rect 3260 2069 3294 2103
rect 3328 2069 3362 2103
rect 3396 2069 3430 2103
rect 3464 2069 3498 2103
rect 3532 2069 3566 2103
rect 3600 2069 3629 2103
rect 3668 2069 3701 2103
rect 3736 2069 3770 2103
rect 3807 2069 3838 2103
rect 3879 2069 3906 2103
rect 3951 2069 3974 2103
rect 4023 2092 4093 2103
rect 4127 2092 4128 2126
rect 4023 2069 4128 2092
rect 1456 2068 4128 2069
rect 1077 2029 1113 2063
rect 4092 2058 4128 2068
rect 1077 1995 1078 2029
rect 1112 1995 1113 2029
rect 1077 1961 1113 1995
rect 1077 1927 1078 1961
rect 1112 1927 1113 1961
rect 1077 1893 1113 1927
rect 1349 2022 1770 2034
rect 1383 2018 1770 2022
rect 1383 1988 1668 2018
rect 1349 1984 1668 1988
rect 1702 1984 1736 2018
rect 1349 1968 1770 1984
rect 1955 2018 2261 2034
rect 1989 1984 2023 2018
rect 2057 1984 2091 2018
rect 2125 1984 2149 2018
rect 2193 1984 2221 2018
rect 1955 1968 2261 1984
rect 2411 2018 2717 2034
rect 2451 1984 2479 2018
rect 2523 1984 2547 2018
rect 2581 1984 2615 2018
rect 2649 1984 2683 2018
rect 2411 1968 2717 1984
rect 2867 2018 3173 2034
rect 2901 1984 2935 2018
rect 2969 1984 3003 2018
rect 3037 1984 3061 2018
rect 3105 1984 3133 2018
rect 2867 1968 3173 1984
rect 3323 2018 3629 2034
rect 3363 1984 3391 2018
rect 3435 1984 3459 2018
rect 3493 1984 3527 2018
rect 3561 1984 3595 2018
rect 3323 1968 3629 1984
rect 3814 2018 3977 2034
rect 3848 1984 3882 2018
rect 3916 1984 3977 2018
rect 3814 1968 3977 1984
rect 1349 1950 1383 1968
rect 3943 1930 3977 1968
rect 4092 2024 4093 2058
rect 4127 2024 4128 2058
rect 4092 1990 4128 2024
rect 4092 1956 4093 1990
rect 4127 1956 4128 1990
rect 4092 1922 4128 1956
rect 1077 1859 1078 1893
rect 1112 1859 1113 1893
rect 4092 1888 4093 1922
rect 4127 1888 4128 1922
rect 1077 1825 1113 1859
rect 1077 1791 1078 1825
rect 1112 1791 1113 1825
rect 1077 1757 1113 1791
rect 1077 1723 1078 1757
rect 1112 1723 1113 1757
rect 1077 1689 1113 1723
rect 1077 1655 1078 1689
rect 1112 1655 1113 1689
rect 1077 1621 1113 1655
rect 1077 1587 1078 1621
rect 1112 1587 1113 1621
rect 1077 1553 1113 1587
rect 1077 1519 1078 1553
rect 1112 1519 1113 1553
rect 1077 1485 1113 1519
rect 1077 1451 1078 1485
rect 1112 1451 1113 1485
rect 1077 1417 1113 1451
rect 1077 1383 1078 1417
rect 1112 1383 1113 1417
rect 1077 1349 1113 1383
rect 1077 1315 1078 1349
rect 1112 1315 1113 1349
rect 1077 1281 1113 1315
rect 1077 1247 1078 1281
rect 1112 1247 1113 1281
rect 1077 1213 1113 1247
rect 1077 1179 1078 1213
rect 1112 1179 1113 1213
rect 1077 1145 1113 1179
rect 1077 1111 1078 1145
rect 1112 1111 1113 1145
rect 1077 1077 1113 1111
rect 1077 1043 1078 1077
rect 1112 1043 1113 1077
rect 1077 1009 1113 1043
rect 1077 975 1078 1009
rect 1112 975 1113 1009
rect 1077 941 1113 975
rect 1077 907 1078 941
rect 1112 907 1113 941
rect 1077 873 1113 907
rect 1077 839 1078 873
rect 1112 839 1113 873
rect 1077 805 1113 839
rect 1077 771 1078 805
rect 1112 771 1113 805
rect 1077 737 1113 771
rect 197 670 233 704
rect 307 701 373 713
rect 307 685 323 701
rect 197 636 198 670
rect 232 636 233 670
rect 357 685 373 701
rect 433 701 499 713
rect 433 685 449 701
rect 323 651 357 667
rect 483 685 499 701
rect 559 701 625 713
rect 559 685 575 701
rect 449 651 483 667
rect 609 685 625 701
rect 685 701 751 713
rect 685 685 701 701
rect 575 651 609 667
rect 735 685 751 701
rect 811 701 877 713
rect 811 685 827 701
rect 701 651 735 667
rect 861 685 877 701
rect 937 701 1003 713
rect 937 685 953 701
rect 827 651 861 667
rect 987 685 1003 701
rect 1077 703 1078 737
rect 1112 703 1113 737
rect 953 651 987 667
rect 1077 669 1113 703
rect 197 602 233 636
rect 197 568 198 602
rect 232 568 233 602
rect 307 629 373 651
rect 307 583 323 629
rect 357 583 373 629
rect 433 629 499 651
rect 433 583 449 629
rect 483 583 499 629
rect 559 629 625 651
rect 559 583 575 629
rect 609 583 625 629
rect 685 629 751 651
rect 685 583 701 629
rect 735 583 751 629
rect 811 629 877 651
rect 811 583 827 629
rect 861 583 877 629
rect 937 629 1003 651
rect 937 583 953 629
rect 987 583 1003 629
rect 1077 635 1078 669
rect 1112 635 1113 669
rect 1077 601 1113 635
rect 197 501 233 568
rect 1077 567 1078 601
rect 1112 567 1113 601
rect 1077 533 1113 567
rect 1077 501 1078 533
rect 197 500 1078 501
rect 197 466 231 500
rect 265 466 299 500
rect 333 466 367 500
rect 401 466 435 500
rect 469 466 503 500
rect 537 466 571 500
rect 605 466 639 500
rect 673 466 707 500
rect 741 466 775 500
rect 809 466 843 500
rect 877 466 911 500
rect 945 466 979 500
rect 1013 499 1078 500
rect 1112 499 1113 533
rect 1013 466 1113 499
rect 197 429 1113 466
rect 1456 1840 1492 1874
rect 1456 1806 1457 1840
rect 1491 1806 1492 1840
rect 1456 1772 1492 1806
rect 1456 1738 1457 1772
rect 1491 1738 1492 1772
rect 1456 1704 1492 1738
rect 1456 1670 1457 1704
rect 1491 1670 1492 1704
rect 1456 1636 1492 1670
rect 1456 1602 1457 1636
rect 1491 1602 1492 1636
rect 1456 1568 1492 1602
rect 1456 1534 1457 1568
rect 1491 1534 1492 1568
rect 1456 1500 1492 1534
rect 1456 1466 1457 1500
rect 1491 1466 1492 1500
rect 1456 1432 1492 1466
rect 1456 1398 1457 1432
rect 1491 1398 1492 1432
rect 1456 1364 1492 1398
rect 1456 1330 1457 1364
rect 1491 1330 1492 1364
rect 1456 1296 1492 1330
rect 1456 1262 1457 1296
rect 1491 1262 1492 1296
rect 1456 1228 1492 1262
rect 1456 1194 1457 1228
rect 1491 1194 1492 1228
rect 1456 1160 1492 1194
rect 1456 1126 1457 1160
rect 1491 1126 1492 1160
rect 1456 1092 1492 1126
rect 1456 1058 1457 1092
rect 1491 1058 1492 1092
rect 1456 1024 1492 1058
rect 1456 990 1457 1024
rect 1491 990 1492 1024
rect 1456 956 1492 990
rect 1456 922 1457 956
rect 1491 922 1492 956
rect 1456 888 1492 922
rect 1456 854 1457 888
rect 1491 854 1492 888
rect 1456 820 1492 854
rect 1456 786 1457 820
rect 1491 786 1492 820
rect 1456 752 1492 786
rect 1456 718 1457 752
rect 1491 718 1492 752
rect 1456 684 1492 718
rect 1456 650 1457 684
rect 1491 650 1492 684
rect 1456 616 1492 650
rect 1456 582 1457 616
rect 1491 582 1492 616
rect 1456 548 1492 582
rect 1456 514 1457 548
rect 1491 514 1492 548
rect 1456 462 1492 514
rect 4092 1854 4128 1888
rect 4092 1820 4093 1854
rect 4127 1820 4128 1854
rect 4092 1786 4128 1820
rect 4092 1752 4093 1786
rect 4127 1752 4128 1786
rect 4092 1718 4128 1752
rect 4092 1684 4093 1718
rect 4127 1684 4128 1718
rect 4092 1650 4128 1684
rect 4092 1616 4093 1650
rect 4127 1616 4128 1650
rect 4092 1582 4128 1616
rect 4092 1548 4093 1582
rect 4127 1548 4128 1582
rect 4092 1514 4128 1548
rect 4092 1480 4093 1514
rect 4127 1480 4128 1514
rect 4092 1446 4128 1480
rect 4092 1412 4093 1446
rect 4127 1412 4128 1446
rect 4092 1378 4128 1412
rect 4092 1344 4093 1378
rect 4127 1344 4128 1378
rect 4092 1310 4128 1344
rect 4092 1276 4093 1310
rect 4127 1276 4128 1310
rect 4092 1242 4128 1276
rect 4092 1208 4093 1242
rect 4127 1208 4128 1242
rect 4092 1174 4128 1208
rect 4092 1140 4093 1174
rect 4127 1140 4128 1174
rect 4092 1106 4128 1140
rect 4092 1072 4093 1106
rect 4127 1072 4128 1106
rect 4092 1038 4128 1072
rect 4092 1004 4093 1038
rect 4127 1004 4128 1038
rect 4092 970 4128 1004
rect 4092 936 4093 970
rect 4127 936 4128 970
rect 4092 902 4128 936
rect 4092 868 4093 902
rect 4127 868 4128 902
rect 4092 834 4128 868
rect 4092 800 4093 834
rect 4127 800 4128 834
rect 4092 766 4128 800
rect 4092 732 4093 766
rect 4127 732 4128 766
rect 4092 698 4128 732
rect 4092 664 4093 698
rect 4127 664 4128 698
rect 4092 630 4128 664
rect 4092 596 4093 630
rect 4127 596 4128 630
rect 4092 562 4128 596
rect 4092 528 4093 562
rect 4127 528 4128 562
rect 4092 494 4128 528
rect 4092 462 4093 494
rect 1266 461 4093 462
rect 8 294 44 413
rect 1266 427 1299 461
rect 1334 427 1368 461
rect 1405 427 1443 461
rect 1477 427 1490 461
rect 1524 427 1558 461
rect 1592 427 1626 461
rect 1660 427 1694 461
rect 1728 427 1762 461
rect 1796 427 1830 461
rect 1864 427 1898 461
rect 1932 427 1966 461
rect 2000 427 2034 461
rect 2068 427 2102 461
rect 2136 427 2170 461
rect 2204 427 2238 461
rect 2272 427 2306 461
rect 2340 427 2374 461
rect 2408 427 2442 461
rect 2476 427 2510 461
rect 2544 427 2578 461
rect 2612 427 2646 461
rect 2680 427 2714 461
rect 2748 427 2782 461
rect 2816 427 2850 461
rect 2884 427 2918 461
rect 2952 427 2986 461
rect 3020 427 3054 461
rect 3088 427 3122 461
rect 3156 427 3190 461
rect 3224 427 3258 461
rect 3292 427 3326 461
rect 3360 427 3394 461
rect 3428 427 3462 461
rect 3496 427 3530 461
rect 3564 427 3598 461
rect 3632 427 3666 461
rect 3700 427 3734 461
rect 3768 427 3802 461
rect 3836 427 3870 461
rect 3904 427 3938 461
rect 3972 427 4006 461
rect 4040 460 4093 461
rect 4127 460 4128 494
rect 4040 427 4128 460
rect 1266 426 4128 427
rect 1266 381 1302 426
rect 1266 347 1267 381
rect 1301 347 1302 381
rect 1266 311 1302 347
rect 1247 277 1302 311
<< viali >>
rect 323 10548 357 10570
rect 323 10536 357 10548
rect 449 10548 483 10570
rect 449 10536 483 10548
rect 575 10548 609 10570
rect 575 10536 609 10548
rect 701 10548 735 10570
rect 701 10536 735 10548
rect 827 10548 861 10570
rect 827 10536 861 10548
rect 953 10548 987 10570
rect 953 10536 987 10548
rect 323 10464 357 10498
rect 449 10464 483 10498
rect 575 10464 609 10498
rect 701 10464 735 10498
rect 827 10464 861 10498
rect 953 10464 987 10498
rect 323 8727 357 8761
rect 449 8727 483 8761
rect 575 8727 609 8761
rect 701 8727 735 8761
rect 827 8727 861 8761
rect 953 8727 987 8761
rect 323 8677 357 8689
rect 323 8655 357 8677
rect 449 8677 483 8689
rect 449 8655 483 8677
rect 575 8677 609 8689
rect 575 8655 609 8677
rect 701 8677 735 8689
rect 701 8655 735 8677
rect 827 8677 861 8689
rect 827 8655 861 8677
rect 953 8677 987 8689
rect 953 8655 987 8677
rect 323 8533 357 8555
rect 323 8521 357 8533
rect 449 8533 483 8555
rect 449 8521 483 8533
rect 575 8533 609 8555
rect 575 8521 609 8533
rect 701 8533 735 8555
rect 701 8521 735 8533
rect 827 8533 861 8555
rect 827 8521 861 8533
rect 953 8533 987 8555
rect 953 8521 987 8533
rect 323 8449 357 8483
rect 449 8449 483 8483
rect 575 8449 609 8483
rect 701 8449 735 8483
rect 827 8449 861 8483
rect 953 8449 987 8483
rect 323 6712 357 6746
rect 449 6712 483 6746
rect 575 6712 609 6746
rect 701 6712 735 6746
rect 827 6712 861 6746
rect 953 6712 987 6746
rect 323 6662 357 6674
rect 323 6640 357 6662
rect 449 6662 483 6674
rect 449 6640 483 6662
rect 575 6662 609 6674
rect 575 6640 609 6662
rect 701 6662 735 6674
rect 701 6640 735 6662
rect 827 6662 861 6674
rect 827 6640 861 6662
rect 953 6662 987 6674
rect 953 6640 987 6662
rect 1078 6687 1112 6715
rect 1078 6681 1112 6687
rect 1078 6619 1112 6643
rect 1078 6609 1112 6619
rect 323 6518 357 6540
rect 323 6506 357 6518
rect 449 6518 483 6540
rect 449 6506 483 6518
rect 575 6518 609 6540
rect 575 6506 609 6518
rect 701 6518 735 6540
rect 701 6506 735 6518
rect 827 6518 861 6540
rect 827 6506 861 6518
rect 953 6518 987 6540
rect 953 6506 987 6518
rect 1078 6551 1112 6571
rect 1078 6537 1112 6551
rect 323 6434 357 6468
rect 449 6434 483 6468
rect 575 6434 609 6468
rect 701 6434 735 6468
rect 827 6434 861 6468
rect 953 6434 987 6468
rect 1078 6483 1112 6499
rect 1078 6465 1112 6483
rect 323 4697 357 4731
rect 449 4697 483 4731
rect 575 4697 609 4731
rect 701 4697 735 4731
rect 827 4697 861 4731
rect 953 4697 987 4731
rect 323 4647 357 4659
rect 323 4625 357 4647
rect 449 4647 483 4659
rect 449 4625 483 4647
rect 575 4647 609 4659
rect 575 4625 609 4647
rect 701 4647 735 4659
rect 701 4625 735 4647
rect 827 4647 861 4659
rect 827 4625 861 4647
rect 953 4647 987 4659
rect 953 4625 987 4647
rect 323 4503 357 4525
rect 323 4491 357 4503
rect 449 4503 483 4525
rect 449 4491 483 4503
rect 575 4503 609 4525
rect 575 4491 609 4503
rect 701 4503 735 4525
rect 701 4491 735 4503
rect 827 4503 861 4525
rect 827 4491 861 4503
rect 953 4503 987 4525
rect 953 4491 987 4503
rect 323 4419 357 4453
rect 449 4419 483 4453
rect 575 4419 609 4453
rect 701 4419 735 4453
rect 827 4419 861 4453
rect 953 4419 987 4453
rect 323 2682 357 2716
rect 449 2682 483 2716
rect 575 2682 609 2716
rect 701 2682 735 2716
rect 827 2682 861 2716
rect 953 2682 987 2716
rect 323 2632 357 2644
rect 323 2610 357 2632
rect 449 2632 483 2644
rect 449 2610 483 2632
rect 575 2632 609 2644
rect 575 2610 609 2632
rect 701 2632 735 2644
rect 701 2610 735 2632
rect 827 2632 861 2644
rect 827 2610 861 2632
rect 953 2632 987 2644
rect 953 2610 987 2632
rect 323 2488 357 2510
rect 323 2476 357 2488
rect 449 2488 483 2510
rect 449 2476 483 2488
rect 575 2488 609 2510
rect 575 2476 609 2488
rect 701 2488 735 2510
rect 701 2476 735 2488
rect 827 2488 861 2510
rect 827 2476 861 2488
rect 953 2488 987 2510
rect 953 2476 987 2488
rect 323 2404 357 2438
rect 449 2404 483 2438
rect 575 2404 609 2438
rect 701 2404 735 2438
rect 827 2404 861 2438
rect 953 2404 987 2438
rect 1457 10709 1491 10740
rect 1457 10706 1491 10709
rect 1457 10641 1491 10668
rect 1457 10634 1491 10641
rect 1457 10573 1491 10596
rect 1457 10562 1491 10573
rect 1457 10505 1491 10524
rect 1457 10490 1491 10505
rect 1456 9791 1490 9822
rect 1456 9788 1457 9791
rect 1457 9788 1490 9791
rect 1456 9723 1490 9750
rect 1456 9716 1457 9723
rect 1457 9716 1490 9723
rect 1456 9655 1490 9678
rect 1456 9644 1457 9655
rect 1457 9644 1490 9655
rect 1456 8907 1490 8919
rect 1456 8885 1457 8907
rect 1457 8885 1490 8907
rect 1456 8839 1490 8847
rect 1456 8813 1457 8839
rect 1457 8813 1490 8839
rect 1691 10690 1725 10724
rect 1691 10622 1725 10652
rect 1691 10618 1724 10622
rect 1724 10618 1725 10622
rect 1691 10554 1725 10580
rect 1691 10546 1724 10554
rect 1724 10546 1725 10554
rect 1690 9806 1724 9822
rect 1690 9788 1724 9806
rect 1806 10384 1840 10418
rect 1806 10312 1840 10346
rect 1806 10240 1840 10274
rect 1806 10168 1840 10202
rect 1806 10096 1840 10130
rect 1806 10024 1840 10058
rect 1806 9952 1840 9986
rect 3893 10384 3927 10418
rect 3893 10312 3927 10346
rect 3893 10240 3927 10274
rect 3893 10168 3927 10202
rect 3893 10096 3927 10130
rect 3893 10024 3927 10058
rect 3893 9952 3927 9986
rect 6023 10384 6057 10418
rect 6023 10312 6057 10346
rect 6023 10240 6057 10274
rect 6023 10168 6057 10202
rect 6023 10096 6057 10130
rect 6023 10024 6057 10058
rect 6023 9952 6057 9986
rect 8112 10384 8146 10418
rect 8112 10312 8146 10346
rect 8112 10240 8146 10274
rect 8112 10168 8146 10202
rect 8112 10096 8146 10130
rect 8112 10024 8146 10058
rect 8112 9952 8146 9986
rect 1690 9738 1724 9750
rect 1690 9716 1724 9738
rect 1690 9670 1724 9678
rect 1690 9644 1724 9670
rect 1773 9276 1807 9310
rect 1773 9204 1807 9238
rect 1773 9132 1807 9166
rect 1773 9060 1807 9094
rect 6023 9480 6057 9514
rect 6023 9408 6057 9442
rect 6023 9336 6057 9370
rect 6023 9264 6057 9298
rect 6023 9192 6057 9226
rect 6023 9120 6057 9154
rect 6023 9048 6057 9082
rect 8112 9480 8146 9514
rect 8112 9408 8146 9442
rect 8112 9336 8146 9370
rect 8112 9264 8146 9298
rect 8112 9192 8146 9226
rect 8112 9120 8146 9154
rect 8112 9048 8146 9082
rect 1773 8988 1807 9022
rect 1690 8888 1724 8920
rect 1690 8886 1724 8888
rect 1690 8814 1724 8848
rect 1456 8771 1490 8775
rect 1456 8741 1457 8771
rect 1457 8741 1490 8771
rect 1905 8590 1939 8624
rect 1977 8590 2011 8624
rect 4251 8578 4285 8612
rect 4251 8506 4285 8540
rect 3999 3419 4033 3453
rect 3999 3347 4033 3381
rect 1759 2258 1781 2292
rect 1781 2258 1793 2292
rect 1831 2258 1849 2292
rect 1849 2258 1865 2292
rect 3719 2258 3753 2292
rect 3791 2258 3821 2292
rect 3821 2258 3825 2292
rect 1730 2069 1764 2103
rect 1802 2069 1832 2103
rect 1832 2069 1836 2103
rect 1874 2069 1900 2103
rect 1900 2069 1908 2103
rect 1946 2069 1968 2103
rect 1968 2069 1980 2103
rect 2018 2069 2036 2103
rect 2036 2069 2052 2103
rect 2570 2069 2580 2103
rect 2580 2069 2604 2103
rect 2642 2069 2648 2103
rect 2648 2069 2676 2103
rect 2714 2069 2716 2103
rect 2716 2069 2748 2103
rect 2786 2069 2818 2103
rect 2818 2069 2820 2103
rect 2858 2069 2886 2103
rect 2886 2069 2892 2103
rect 2930 2069 2954 2103
rect 2954 2069 2964 2103
rect 3629 2069 3634 2103
rect 3634 2069 3663 2103
rect 3701 2069 3702 2103
rect 3702 2069 3735 2103
rect 3773 2069 3804 2103
rect 3804 2069 3807 2103
rect 3845 2069 3872 2103
rect 3872 2069 3879 2103
rect 3917 2069 3940 2103
rect 3940 2069 3951 2103
rect 3989 2069 4008 2103
rect 4008 2069 4023 2103
rect 1349 1988 1383 2022
rect 2149 1984 2159 2018
rect 2159 1984 2183 2018
rect 2221 1984 2227 2018
rect 2227 1984 2255 2018
rect 2417 1984 2445 2018
rect 2445 1984 2451 2018
rect 2489 1984 2513 2018
rect 2513 1984 2523 2018
rect 3061 1984 3071 2018
rect 3071 1984 3095 2018
rect 3133 1984 3139 2018
rect 3139 1984 3167 2018
rect 3329 1984 3357 2018
rect 3357 1984 3363 2018
rect 3401 1984 3425 2018
rect 3425 1984 3435 2018
rect 1349 1916 1383 1950
rect 323 667 357 701
rect 449 667 483 701
rect 575 667 609 701
rect 701 667 735 701
rect 827 667 861 701
rect 953 667 987 701
rect 323 617 357 629
rect 323 595 357 617
rect 449 617 483 629
rect 449 595 483 617
rect 575 617 609 629
rect 575 595 609 617
rect 701 617 735 629
rect 701 595 735 617
rect 827 617 861 629
rect 827 595 861 617
rect 953 617 987 629
rect 953 595 987 617
rect 1299 427 1300 461
rect 1300 427 1333 461
rect 1371 427 1402 461
rect 1402 427 1405 461
rect 1443 427 1477 461
rect 1267 347 1301 381
<< metal1 >>
rect -3 11100 2702 11152
rect 2754 11100 2766 11152
rect 2818 11100 2830 11152
rect 2882 11100 4796 11152
rect 4848 11100 4860 11152
rect 4912 11100 4924 11152
rect 4976 11100 4988 11152
rect 5040 11100 5052 11152
rect 5104 11100 7167 11152
rect 7219 11100 7231 11152
rect 7283 11100 7295 11152
rect 7347 11100 7359 11152
rect 7411 11100 8522 11152
rect -3 11020 7757 11072
rect 7809 11020 7821 11072
rect 7873 11020 7885 11072
rect 7937 11020 7949 11072
rect 8001 11020 8013 11072
rect 8065 11020 8522 11072
rect -3 10940 2702 10992
rect 2754 10940 2766 10992
rect 2818 10940 2830 10992
rect 2882 10940 4796 10992
rect 4848 10940 4860 10992
rect 4912 10940 4924 10992
rect 4976 10940 4988 10992
rect 5040 10940 5052 10992
rect 5104 10940 7167 10992
rect 7219 10940 7231 10992
rect 7283 10940 7295 10992
rect 7347 10940 7359 10992
rect 7411 10940 8522 10992
rect 1403 10881 1503 10912
rect 8388 10911 8522 10912
rect 1403 10866 1449 10881
tri 1418 10839 1445 10866 ne
rect 1445 10829 1449 10866
rect 1501 10866 1503 10881
rect 1549 10866 1555 10911
rect 1501 10859 1555 10866
rect 1607 10859 1619 10911
rect 1671 10859 1677 10911
tri 1677 10859 1684 10866 nw
tri 8125 10859 8132 10866 ne
rect 8132 10859 8138 10911
rect 8190 10859 8202 10911
rect 8254 10859 8266 10911
rect 8318 10859 8330 10911
rect 8382 10859 8522 10911
rect 1501 10829 1503 10859
rect -3 10821 1204 10827
rect -3 10781 1152 10821
tri 1127 10756 1152 10781 ne
rect 1152 10757 1204 10769
tri 213 10706 243 10736 se
rect 243 10706 272 10736
rect 1038 10733 1121 10736
tri 197 10690 213 10706 se
rect 213 10690 272 10706
tri 186 10679 197 10690 se
rect 197 10679 272 10690
rect 993 10681 999 10733
rect 1051 10681 1063 10733
rect 1115 10681 1121 10733
rect 1152 10699 1204 10705
rect 1445 10817 1503 10829
rect 1445 10765 1449 10817
rect 1501 10765 1503 10817
tri 1503 10813 1549 10859 nw
tri 8357 10838 8378 10859 ne
rect 8378 10838 8522 10859
rect 2971 10786 2977 10838
rect 3029 10786 3041 10838
rect 3093 10786 3105 10838
rect 3157 10786 4517 10838
rect 4569 10786 4581 10838
rect 4633 10786 4645 10838
rect 4697 10786 5473 10838
rect 5525 10786 5537 10838
rect 5589 10786 5601 10838
rect 5653 10786 5659 10838
tri 8378 10813 8403 10838 ne
rect 8403 10788 8522 10838
rect 1445 10753 1503 10765
rect 1445 10701 1449 10753
rect 1501 10701 1503 10753
rect 186 10678 272 10679
rect 1038 10678 1121 10681
rect 1445 10689 1503 10701
rect 186 10668 259 10678
tri 259 10668 269 10678 nw
rect 186 10646 244 10668
tri 244 10653 259 10668 nw
tri 344 10646 348 10650 se
rect 348 10646 1253 10650
tri 332 10634 344 10646 se
rect 344 10634 1253 10646
tri 1253 10634 1269 10650 sw
rect 1445 10637 1449 10689
rect 1501 10637 1503 10689
rect 1445 10634 1457 10637
rect 1491 10634 1503 10637
tri 316 10618 332 10634 se
rect 332 10619 1269 10634
tri 1269 10619 1284 10634 sw
rect 332 10618 1284 10619
tri 311 10613 316 10618 se
rect 316 10613 1284 10618
rect 311 10610 1284 10613
rect 311 10596 380 10610
tri 380 10596 394 10610 nw
tri 916 10596 930 10610 ne
rect 930 10596 1010 10610
tri 1010 10596 1024 10610 nw
tri 1207 10596 1221 10610 ne
rect 1221 10604 1284 10610
rect 1221 10596 1232 10604
rect 311 10570 369 10596
tri 369 10585 380 10596 nw
tri 930 10585 941 10596 ne
rect 311 10536 323 10570
rect 357 10536 369 10570
rect 311 10498 369 10536
rect 311 10464 323 10498
rect 357 10464 369 10498
rect 311 8761 369 10464
rect 437 10570 621 10582
rect 437 10536 449 10570
rect 483 10536 575 10570
rect 609 10536 621 10570
rect 437 10498 621 10536
rect 437 10464 449 10498
rect 483 10464 575 10498
rect 609 10464 621 10498
rect 437 10452 621 10464
rect 689 10570 873 10582
rect 689 10536 701 10570
rect 735 10536 827 10570
rect 861 10536 873 10570
rect 689 10498 873 10536
rect 689 10464 701 10498
rect 735 10464 827 10498
rect 861 10464 873 10498
rect 689 10452 873 10464
rect 941 10570 999 10596
tri 999 10585 1010 10596 nw
tri 1221 10585 1232 10596 ne
rect 941 10536 953 10570
rect 987 10536 999 10570
rect 941 10498 999 10536
rect 941 10464 953 10498
rect 987 10464 999 10498
rect 311 8727 323 8761
rect 357 8727 369 8761
rect 311 8689 369 8727
rect 311 8655 323 8689
rect 357 8655 369 8689
rect 311 8555 369 8655
rect 311 8521 323 8555
rect 357 8521 369 8555
rect 311 8483 369 8521
rect 311 8449 323 8483
rect 357 8449 369 8483
rect 311 6746 369 8449
rect 437 8761 495 8773
rect 437 8727 449 8761
rect 483 8727 495 8761
rect 437 8689 495 8727
rect 437 8655 449 8689
rect 483 8655 495 8689
rect 437 8555 495 8655
rect 437 8521 449 8555
rect 483 8521 495 8555
rect 437 8483 495 8521
rect 437 8449 449 8483
rect 483 8449 495 8483
rect 437 8437 495 8449
rect 563 8761 621 8773
rect 563 8727 575 8761
rect 609 8727 621 8761
rect 563 8689 621 8727
rect 563 8655 575 8689
rect 609 8655 621 8689
rect 563 8555 621 8655
rect 563 8521 575 8555
rect 609 8521 621 8555
rect 563 8483 621 8521
rect 563 8449 575 8483
rect 609 8449 621 8483
rect 563 8437 621 8449
rect 689 8761 747 8773
rect 689 8727 701 8761
rect 735 8727 747 8761
rect 689 8689 747 8727
rect 689 8655 701 8689
rect 735 8655 747 8689
rect 689 8555 747 8655
rect 689 8521 701 8555
rect 735 8521 747 8555
rect 689 8483 747 8521
rect 689 8449 701 8483
rect 735 8449 747 8483
rect 689 8437 747 8449
rect 815 8761 873 8773
rect 815 8727 827 8761
rect 861 8727 873 8761
rect 815 8689 873 8727
rect 815 8655 827 8689
rect 861 8655 873 8689
rect 815 8555 873 8655
rect 815 8521 827 8555
rect 861 8521 873 8555
rect 815 8483 873 8521
rect 815 8449 827 8483
rect 861 8449 873 8483
rect 815 8437 873 8449
rect 941 8761 999 10464
rect 1232 10540 1284 10552
rect 1232 10476 1284 10488
rect 1445 10625 1503 10634
rect 1445 10573 1449 10625
rect 1501 10573 1503 10625
rect 1445 10562 1457 10573
rect 1491 10562 1503 10573
rect 1445 10524 1503 10562
rect 1679 10726 8272 10732
rect 1679 10724 2015 10726
rect 1679 10690 1691 10724
rect 1725 10690 2015 10724
rect 1679 10674 2015 10690
rect 2067 10674 3517 10726
rect 3569 10674 4651 10726
rect 4703 10674 7822 10726
rect 1679 10662 7822 10674
rect 1679 10652 2015 10662
rect 1679 10618 1691 10652
rect 1725 10618 2015 10652
rect 1679 10610 2015 10618
rect 2067 10610 3517 10662
rect 3569 10610 4651 10662
rect 4703 10610 7822 10662
rect 1679 10598 7822 10610
rect 1679 10580 2015 10598
rect 1679 10546 1691 10580
rect 1725 10546 2015 10580
rect 2067 10546 3517 10598
rect 3569 10546 4651 10598
rect 4703 10546 7822 10598
rect 7938 10546 8272 10726
rect 1679 10540 8272 10546
rect 1445 10490 1457 10524
rect 1491 10490 1503 10524
tri 8189 10515 8214 10540 ne
rect 1445 10484 1503 10490
rect 1232 10418 1284 10424
rect 1340 9941 1415 10428
rect 1416 9942 1417 10427
rect 1453 9942 1454 10427
rect 1455 10418 8158 10428
rect 1455 10384 1806 10418
rect 1840 10384 3893 10418
rect 3927 10384 6023 10418
rect 6057 10384 8112 10418
rect 8146 10384 8158 10418
rect 1455 10346 8158 10384
rect 1455 10312 1806 10346
rect 1840 10312 3893 10346
rect 3927 10312 6023 10346
rect 6057 10312 8112 10346
rect 8146 10312 8158 10346
rect 1455 10274 8158 10312
rect 1455 10240 1806 10274
rect 1840 10240 3893 10274
rect 3927 10240 6023 10274
rect 6057 10240 8112 10274
rect 8146 10240 8158 10274
rect 1455 10202 8158 10240
rect 1455 10168 1806 10202
rect 1840 10168 3893 10202
rect 3927 10168 6023 10202
rect 6057 10168 8112 10202
rect 8146 10168 8158 10202
rect 1455 10130 8158 10168
rect 1455 10096 1806 10130
rect 1840 10096 3893 10130
rect 3927 10096 6023 10130
rect 6057 10096 8112 10130
rect 8146 10096 8158 10130
rect 1455 10058 8158 10096
rect 1455 10024 1806 10058
rect 1840 10024 3893 10058
rect 3927 10024 6023 10058
rect 6057 10024 8112 10058
rect 8146 10024 8158 10058
rect 1455 9986 8158 10024
rect 1455 9952 1806 9986
rect 1840 9952 3893 9986
rect 3927 9952 6023 9986
rect 6057 9952 8112 9986
rect 8146 9952 8158 9986
rect 1455 9941 8158 9952
tri 1392 9916 1417 9941 nw
tri 1512 9916 1537 9941 ne
rect 1537 9916 1617 9941
tri 1537 9890 1563 9916 ne
rect 1563 9892 1617 9916
tri 1617 9892 1666 9941 nw
rect 1615 9891 1616 9892
tri 1616 9891 1617 9892 nw
rect 1564 9890 1614 9891
tri 1615 9890 1616 9891 nw
rect 1563 9854 1615 9890
tri 1538 9829 1563 9854 se
rect 1564 9853 1614 9854
tri 1615 9853 1616 9854 sw
tri 8213 9853 8214 9854 se
rect 1615 9852 1616 9853
tri 1616 9852 1617 9853 sw
tri 8212 9852 8213 9853 se
rect 8213 9852 8214 9853
rect 1563 9829 1617 9852
tri 1617 9829 1640 9852 sw
tri 8189 9829 8212 9852 se
rect 8212 9829 8214 9852
rect 1444 9823 1502 9829
rect 1444 9771 1449 9823
rect 1501 9771 1502 9823
rect 1444 9759 1502 9771
rect 1444 9707 1449 9759
rect 1501 9707 1502 9759
rect 1444 9695 1502 9707
rect 1444 9643 1449 9695
rect 1501 9643 1502 9695
rect 1444 9637 1502 9643
rect 1538 9823 8214 9829
rect 1538 9822 2015 9823
rect 1538 9788 1690 9822
rect 1724 9788 2015 9822
rect 1538 9771 2015 9788
rect 2067 9771 3517 9823
rect 3569 9771 4651 9823
rect 4703 9771 7822 9823
rect 1538 9759 7822 9771
rect 1538 9750 2015 9759
rect 1538 9716 1690 9750
rect 1724 9716 2015 9750
rect 1538 9707 2015 9716
rect 2067 9707 3517 9759
rect 3569 9707 4651 9759
rect 4703 9707 7822 9759
rect 1538 9695 7822 9707
rect 1538 9678 2015 9695
rect 1538 9644 1690 9678
rect 1724 9644 2015 9678
rect 1538 9643 2015 9644
rect 2067 9643 3517 9695
rect 3569 9643 4651 9695
rect 4703 9643 7822 9695
rect 7938 9643 8214 9823
rect 1538 9637 8214 9643
tri 1538 9612 1563 9637 ne
rect 1563 9614 1617 9637
tri 1617 9614 1640 9637 nw
tri 8189 9614 8212 9637 ne
rect 8212 9614 8214 9637
rect 1615 9613 1616 9614
tri 1616 9613 1617 9614 nw
tri 8212 9613 8213 9614 ne
rect 8213 9613 8214 9614
rect 1564 9612 1614 9613
tri 1615 9612 1616 9613 nw
tri 8213 9612 8214 9613 ne
rect 1563 9576 1615 9612
tri 1392 9551 1417 9576 sw
tri 1538 9551 1563 9576 se
rect 1564 9575 1614 9576
tri 1615 9575 1616 9576 sw
rect 1615 9574 1616 9575
tri 1616 9574 1617 9575 sw
rect 1563 9551 1617 9574
tri 1617 9551 1640 9574 sw
rect 1363 9411 1415 9551
rect 1416 9412 1417 9550
rect 1453 9412 1454 9550
rect 1455 9514 8158 9551
rect 1455 9480 6023 9514
rect 6057 9480 8112 9514
rect 8146 9480 8158 9514
rect 1455 9442 8158 9480
rect 1455 9411 6023 9442
rect 1392 9408 1414 9411
tri 1414 9408 1417 9411 nw
tri 5986 9408 5989 9411 ne
rect 5989 9408 6023 9411
rect 6057 9411 8112 9442
rect 6057 9408 6091 9411
tri 6091 9408 6094 9411 nw
tri 8075 9408 8078 9411 ne
rect 8078 9408 8112 9411
rect 8146 9408 8158 9442
tri 1392 9386 1414 9408 nw
tri 5989 9386 6011 9408 ne
rect 6011 9370 6069 9408
tri 6069 9386 6091 9408 nw
tri 8078 9386 8100 9408 ne
rect 6011 9336 6023 9370
rect 6057 9336 6069 9370
rect 1761 9310 1819 9316
rect 1761 9276 1773 9310
rect 1807 9276 1819 9310
rect 1761 9238 1819 9276
tri 1392 9204 1395 9207 sw
tri 1758 9204 1761 9207 se
rect 1761 9204 1773 9238
rect 1807 9204 1819 9238
rect 1392 9192 1395 9204
tri 1395 9192 1407 9204 sw
tri 1746 9192 1758 9204 se
rect 1758 9192 1819 9204
rect 1392 9182 1407 9192
tri 1407 9182 1417 9192 sw
tri 1736 9182 1746 9192 se
rect 1746 9182 1819 9192
rect 1363 9012 1415 9182
rect 1417 9181 1453 9182
rect 1416 9013 1454 9181
rect 1455 9166 1819 9182
rect 1455 9132 1773 9166
rect 1807 9132 1819 9166
rect 1455 9094 1819 9132
rect 1455 9060 1773 9094
rect 1807 9060 1819 9094
rect 1455 9022 1819 9060
rect 6011 9298 6069 9336
rect 6011 9264 6023 9298
rect 6057 9264 6069 9298
rect 6011 9226 6069 9264
rect 6011 9192 6023 9226
rect 6057 9192 6069 9226
rect 6011 9154 6069 9192
rect 6011 9120 6023 9154
rect 6057 9120 6069 9154
rect 6011 9082 6069 9120
rect 6011 9048 6023 9082
rect 6057 9048 6069 9082
rect 6011 9042 6069 9048
rect 8100 9370 8158 9408
rect 8100 9336 8112 9370
rect 8146 9336 8158 9370
rect 8100 9298 8158 9336
rect 8100 9264 8112 9298
rect 8146 9264 8158 9298
rect 8100 9226 8158 9264
rect 8100 9192 8112 9226
rect 8146 9192 8158 9226
rect 8100 9154 8158 9192
rect 8100 9120 8112 9154
rect 8146 9120 8158 9154
rect 8100 9082 8158 9120
rect 8100 9048 8112 9082
rect 8146 9048 8158 9082
rect 8100 9042 8158 9048
rect 1417 9012 1453 9013
rect 1455 9012 1773 9022
tri 1538 8988 1562 9012 ne
rect 1562 8989 1617 9012
tri 1617 8989 1640 9012 nw
tri 1731 8989 1754 9012 ne
rect 1754 8989 1773 9012
rect 1562 8988 1563 8989
rect 1615 8988 1616 8989
tri 1616 8988 1617 8989 nw
tri 1754 8988 1755 8989 ne
rect 1755 8988 1773 8989
rect 1807 8988 1819 9022
tri 1562 8987 1563 8988 ne
rect 1564 8987 1614 8988
tri 1615 8987 1616 8988 nw
tri 1755 8987 1756 8988 ne
rect 1756 8987 1819 8988
tri 1756 8982 1761 8987 ne
rect 1761 8982 1819 8987
tri 1538 8926 1563 8951 se
rect 1564 8950 1614 8951
tri 1615 8950 1616 8951 sw
tri 8213 8950 8214 8951 se
rect 1615 8949 1616 8950
tri 1616 8949 1617 8950 sw
tri 8212 8949 8213 8950 se
rect 8213 8949 8214 8950
rect 1563 8926 1617 8949
tri 1617 8926 1640 8949 sw
tri 8189 8926 8212 8949 se
rect 8212 8926 8214 8949
rect 1444 8920 1502 8926
rect 1444 8868 1449 8920
rect 1501 8868 1502 8920
rect 1444 8856 1502 8868
rect 941 8727 953 8761
rect 987 8727 999 8761
rect 941 8689 999 8727
rect 941 8655 953 8689
rect 987 8655 999 8689
rect 941 8555 999 8655
rect 1152 8838 1204 8844
rect 1152 8774 1204 8786
rect 1444 8804 1449 8856
rect 1501 8804 1502 8856
rect 1444 8792 1502 8804
rect 1444 8740 1449 8792
rect 1501 8740 1502 8792
rect 1444 8734 1502 8740
rect 1538 8920 8272 8926
rect 1538 8886 1690 8920
rect 1724 8886 2015 8920
rect 1538 8868 2015 8886
rect 2067 8868 3517 8920
rect 3569 8868 4651 8920
rect 4703 8868 7822 8920
rect 1538 8856 7822 8868
rect 1538 8848 2015 8856
rect 1538 8814 1690 8848
rect 1724 8814 2015 8848
rect 1538 8804 2015 8814
rect 2067 8804 3517 8856
rect 3569 8804 4651 8856
rect 4703 8804 7822 8856
rect 1538 8792 7822 8804
rect 1538 8740 2015 8792
rect 2067 8740 3517 8792
rect 3569 8740 4651 8792
rect 4703 8740 7822 8792
rect 7938 8740 8272 8920
rect 1538 8734 8272 8740
rect 1152 8710 1204 8722
tri 1204 8698 1229 8723 sw
rect 1204 8658 4385 8698
rect 1152 8652 1868 8658
tri 1868 8652 1874 8658 nw
tri 2051 8652 2057 8658 ne
rect 2057 8652 4385 8658
tri 1887 8624 1893 8630 se
rect 1893 8624 2023 8630
tri 2023 8624 2029 8630 sw
rect 941 8521 953 8555
rect 987 8521 999 8555
rect 941 8483 999 8521
rect 941 8449 953 8483
rect 987 8449 999 8483
rect 941 6936 999 8449
rect 1152 8618 1905 8624
rect 1204 8596 1905 8618
rect 1204 8590 1223 8596
tri 1223 8590 1229 8596 nw
tri 1881 8590 1887 8596 ne
rect 1887 8590 1905 8596
rect 1939 8590 1977 8624
rect 2011 8612 4291 8624
rect 2011 8596 4251 8612
rect 2011 8590 2023 8596
rect 1204 8578 1211 8590
tri 1211 8578 1223 8590 nw
tri 1887 8584 1893 8590 ne
rect 1893 8584 2023 8590
tri 2023 8584 2035 8596 nw
tri 4220 8584 4232 8596 ne
rect 4232 8584 4251 8596
tri 4232 8578 4238 8584 ne
rect 4238 8578 4251 8584
rect 4285 8578 4291 8612
tri 1204 8571 1211 8578 nw
tri 4238 8571 4245 8578 ne
rect 1152 8554 1204 8566
rect 1751 8556 1865 8568
tri 1865 8556 1877 8568 sw
tri 2039 8556 2051 8568 se
rect 2051 8556 2260 8568
rect 2262 8567 2298 8568
rect 1445 8509 1503 8519
rect 1152 8490 1204 8502
rect 1152 8432 1204 8438
rect 1751 8404 2260 8556
rect 2261 8405 2299 8567
rect 2262 8404 2298 8405
rect 2300 8404 4015 8568
rect 4017 8567 4053 8568
rect 4016 8405 4054 8567
rect 4055 8564 4205 8568
tri 4205 8564 4209 8568 sw
rect 4017 8404 4053 8405
rect 4055 8404 4209 8564
rect 4245 8540 4291 8578
rect 4245 8506 4251 8540
rect 4285 8506 4291 8540
rect 4245 8494 4291 8506
tri 1809 8379 1834 8404 nw
tri 2078 8379 2103 8404 ne
rect 2103 8369 2161 8404
tri 2161 8379 2186 8404 nw
tri 2590 8379 2615 8404 ne
tri 2673 8379 2698 8404 nw
tri 3102 8379 3127 8404 ne
tri 3185 8379 3210 8404 nw
tri 3614 8379 3639 8404 ne
tri 3697 8379 3722 8404 nw
tri 4126 8379 4151 8404 ne
rect 4151 8369 4209 8404
rect 2359 7720 2417 7772
rect 2360 7718 2416 7719
rect 2360 7681 2416 7682
rect 2359 7655 2417 7680
tri 2417 7655 2442 7680 sw
tri 2846 7655 2871 7680 se
rect 2871 7655 2929 7766
rect 3383 7720 3441 7772
rect 3384 7718 3440 7719
rect 3895 7720 3953 7772
rect 3896 7718 3952 7719
rect 3384 7681 3440 7682
rect 3896 7681 3952 7682
tri 2929 7655 2954 7680 sw
tri 3358 7655 3383 7680 se
rect 3383 7655 3441 7680
tri 3441 7655 3466 7680 sw
tri 3870 7655 3895 7680 se
rect 3895 7655 3953 7680
rect 2359 7628 3953 7655
tri 2359 7603 2384 7628 ne
rect 2384 7603 3928 7628
tri 3928 7603 3953 7628 nw
tri 1692 7516 1717 7541 sw
tri 1902 7516 1927 7541 se
rect 1927 7516 1985 7603
tri 2738 7578 2763 7603 ne
tri 1985 7516 2010 7541 sw
rect 1634 7508 2721 7516
rect 1634 7392 1756 7508
rect 1936 7456 2015 7508
rect 2067 7456 2669 7508
rect 1936 7444 2721 7456
rect 1936 7392 2015 7444
rect 2067 7392 2669 7444
rect 1634 7383 2721 7392
tri 1500 7327 1537 7364 sw
rect 1500 7275 1555 7327
rect 1607 7275 1619 7327
rect 1671 7275 1677 7327
tri 1677 7275 1702 7300 nw
rect 1500 7239 1503 7275
tri 1503 7239 1539 7275 nw
rect 1340 7202 1417 7208
rect 1392 7150 1417 7202
rect 1340 7144 1417 7150
rect 1445 7202 2641 7208
rect 1445 7150 2525 7202
rect 2577 7150 2589 7202
rect 1445 7144 2641 7150
rect 1340 7138 1392 7144
rect 1232 7122 1284 7128
rect 1232 7058 1284 7070
rect 1232 6994 1284 7006
tri 999 6936 1024 6961 sw
tri 1207 6936 1232 6961 se
rect 1232 6936 1284 6942
rect 941 6927 1284 6936
tri 941 6896 972 6927 ne
rect 972 6896 1253 6927
tri 1253 6896 1284 6927 nw
tri 1392 7119 1417 7144 nw
rect 1340 7074 1392 7086
tri 1634 7090 1660 7116 se
rect 1660 7090 1741 7116
rect 1634 7083 1741 7090
rect 1692 7070 1741 7083
rect 1340 7010 1392 7022
rect 1340 6946 1392 6958
tri 1315 6868 1340 6893 se
rect 1340 6882 1392 6894
tri 815 6809 874 6868 se
rect 874 6830 1340 6868
rect 874 6810 1392 6830
rect 874 6809 897 6810
tri 897 6809 898 6810 nw
rect 311 6712 323 6746
rect 357 6712 369 6746
rect 311 6674 369 6712
rect 311 6640 323 6674
rect 357 6640 369 6674
rect 311 6540 369 6640
rect 311 6506 323 6540
rect 357 6506 369 6540
rect 311 6468 369 6506
rect 311 6434 323 6468
rect 357 6434 369 6468
rect 311 4731 369 6434
rect 437 6746 495 6758
rect 437 6712 449 6746
rect 483 6712 495 6746
rect 437 6674 495 6712
rect 437 6640 449 6674
rect 483 6640 495 6674
rect 437 6540 495 6640
rect 563 6746 747 6758
rect 563 6712 575 6746
rect 609 6712 701 6746
rect 735 6712 747 6746
rect 563 6674 747 6712
rect 563 6640 575 6674
rect 609 6640 701 6674
rect 735 6640 747 6674
rect 563 6628 747 6640
rect 815 6746 873 6809
tri 873 6785 897 6809 nw
rect 815 6712 827 6746
rect 861 6712 873 6746
rect 815 6674 873 6712
rect 815 6640 827 6674
rect 861 6640 873 6674
rect 815 6610 873 6640
rect 816 6608 872 6609
rect 815 6572 873 6608
rect 816 6571 872 6572
rect 437 6506 449 6540
rect 483 6506 495 6540
rect 437 6468 495 6506
rect 437 6434 449 6468
rect 483 6434 495 6468
rect 437 6422 495 6434
rect 563 6540 747 6552
rect 563 6506 575 6540
rect 609 6506 701 6540
rect 735 6506 747 6540
rect 563 6468 747 6506
rect 563 6434 575 6468
rect 609 6434 701 6468
rect 735 6434 747 6468
rect 563 6422 747 6434
rect 815 6540 873 6570
rect 815 6506 827 6540
rect 861 6506 873 6540
rect 815 6468 873 6506
rect 815 6434 827 6468
rect 861 6434 873 6468
rect 815 6364 873 6434
tri 941 6758 965 6782 se
rect 965 6758 1260 6782
tri 1260 6758 1284 6782 sw
rect 941 6749 1284 6758
rect 941 6746 999 6749
rect 941 6712 953 6746
rect 987 6712 999 6746
tri 999 6724 1024 6749 nw
tri 1207 6724 1232 6749 ne
rect 1232 6744 1284 6749
rect 941 6674 999 6712
rect 941 6640 953 6674
rect 987 6640 999 6674
rect 941 6540 999 6640
rect 941 6506 953 6540
rect 987 6506 999 6540
rect 941 6468 999 6506
rect 941 6434 953 6468
rect 987 6434 999 6468
rect 1066 6715 1124 6721
rect 1066 6712 1078 6715
rect 1112 6712 1124 6715
rect 1066 6660 1069 6712
rect 1121 6660 1124 6712
rect 1066 6648 1124 6660
rect 1066 6596 1069 6648
rect 1121 6596 1124 6648
rect 1066 6584 1124 6596
rect 1066 6532 1069 6584
rect 1121 6532 1124 6584
rect 1066 6520 1124 6532
rect 1066 6468 1069 6520
rect 1121 6468 1124 6520
rect 1066 6465 1078 6468
rect 1112 6465 1124 6468
rect 1066 6459 1124 6465
rect 1232 6680 1284 6692
rect 1232 6616 1284 6628
rect 1232 6552 1284 6564
rect 1232 6488 1284 6500
rect 941 6431 999 6434
tri 999 6431 1024 6456 sw
tri 1207 6431 1232 6456 se
rect 1232 6431 1284 6436
rect 941 6422 1284 6431
tri 941 6391 972 6422 ne
rect 972 6391 1253 6422
tri 1253 6391 1284 6422 nw
rect 1448 6401 1500 6403
rect 1634 6395 1785 7070
tri 1785 7045 1810 7070 nw
rect 2561 7031 2613 7037
tri 2535 6953 2561 6979 ne
rect 2561 6967 2613 6979
tri 2613 6953 2639 6979 nw
rect 2561 6909 2613 6915
tri 1912 6388 1913 6389 se
tri 815 6306 873 6364 ne
tri 873 6363 898 6388 sw
tri 1887 6363 1912 6388 se
rect 1912 6363 1913 6388
rect 873 6306 1913 6363
tri 873 6305 874 6306 ne
rect 874 6305 1913 6306
tri 1887 6279 1913 6305 ne
tri 941 6246 972 6277 se
rect 972 6246 1253 6277
tri 1253 6246 1284 6277 sw
rect 941 6237 1284 6246
rect 311 4697 323 4731
rect 357 4697 369 4731
rect 311 4659 369 4697
rect 311 4625 323 4659
rect 357 4625 369 4659
rect 311 4525 369 4625
rect 311 4491 323 4525
rect 357 4491 369 4525
rect 311 4453 369 4491
rect 311 4419 323 4453
rect 357 4419 369 4453
rect 311 2716 369 4419
rect 437 4731 495 4743
rect 437 4697 449 4731
rect 483 4697 495 4731
rect 437 4659 495 4697
rect 437 4625 449 4659
rect 483 4625 495 4659
rect 437 4525 495 4625
rect 437 4491 449 4525
rect 483 4491 495 4525
rect 437 4453 495 4491
rect 437 4419 449 4453
rect 483 4419 495 4453
rect 437 4407 495 4419
rect 563 4731 621 4743
rect 563 4697 575 4731
rect 609 4697 621 4731
rect 563 4659 621 4697
rect 563 4625 575 4659
rect 609 4625 621 4659
rect 563 4525 621 4625
rect 563 4491 575 4525
rect 609 4491 621 4525
rect 563 4453 621 4491
rect 563 4419 575 4453
rect 609 4419 621 4453
rect 563 4407 621 4419
rect 689 4731 747 4743
rect 689 4697 701 4731
rect 735 4697 747 4731
rect 689 4659 747 4697
rect 689 4625 701 4659
rect 735 4625 747 4659
rect 689 4525 747 4625
rect 689 4491 701 4525
rect 735 4491 747 4525
rect 689 4453 747 4491
rect 689 4419 701 4453
rect 735 4419 747 4453
rect 689 4407 747 4419
rect 815 4731 873 4743
rect 815 4697 827 4731
rect 861 4697 873 4731
rect 815 4659 873 4697
rect 815 4625 827 4659
rect 861 4625 873 4659
rect 815 4525 873 4625
rect 815 4491 827 4525
rect 861 4491 873 4525
rect 815 4453 873 4491
rect 815 4419 827 4453
rect 861 4419 873 4453
rect 815 4407 873 4419
rect 941 4731 999 6237
tri 999 6212 1024 6237 nw
tri 1207 6212 1232 6237 ne
rect 1232 6231 1284 6237
rect 1232 6167 1284 6179
rect 1232 6103 1284 6115
rect 1232 6045 1284 6051
rect 941 4697 953 4731
rect 987 4697 999 4731
rect 941 4659 999 4697
rect 941 4625 953 4659
rect 987 4625 999 4659
rect 941 4525 999 4625
rect 941 4491 953 4525
rect 987 4491 999 4525
rect 941 4453 999 4491
rect 941 4419 953 4453
rect 987 4419 999 4453
rect 311 2682 323 2716
rect 357 2682 369 2716
rect 311 2644 369 2682
rect 311 2610 323 2644
rect 357 2610 369 2644
rect 311 2510 369 2610
rect 311 2476 323 2510
rect 357 2476 369 2510
rect 311 2438 369 2476
rect 311 2404 323 2438
rect 357 2404 369 2438
rect 311 701 369 2404
rect 437 2716 495 2728
rect 437 2682 449 2716
rect 483 2682 495 2716
rect 437 2644 495 2682
rect 437 2610 449 2644
rect 483 2610 495 2644
rect 437 2510 495 2610
rect 437 2476 449 2510
rect 483 2476 495 2510
rect 437 2438 495 2476
rect 437 2404 449 2438
rect 483 2404 495 2438
rect 437 2392 495 2404
rect 563 2716 621 2728
rect 563 2682 575 2716
rect 609 2682 621 2716
rect 563 2644 621 2682
rect 563 2610 575 2644
rect 609 2610 621 2644
rect 563 2510 621 2610
rect 563 2476 575 2510
rect 609 2476 621 2510
rect 563 2438 621 2476
rect 563 2404 575 2438
rect 609 2404 621 2438
rect 563 2392 621 2404
rect 689 2716 747 2728
rect 689 2682 701 2716
rect 735 2682 747 2716
rect 689 2644 747 2682
rect 689 2610 701 2644
rect 735 2610 747 2644
rect 689 2510 747 2610
rect 689 2476 701 2510
rect 735 2476 747 2510
rect 689 2438 747 2476
rect 689 2404 701 2438
rect 735 2404 747 2438
rect 689 2392 747 2404
rect 815 2716 873 2728
rect 815 2682 827 2716
rect 861 2682 873 2716
rect 815 2644 873 2682
rect 815 2610 827 2644
rect 861 2610 873 2644
rect 815 2510 873 2610
rect 815 2476 827 2510
rect 861 2476 873 2510
rect 815 2438 873 2476
rect 815 2404 827 2438
rect 861 2404 873 2438
rect 815 2392 873 2404
rect 941 2716 999 4419
rect 941 2682 953 2716
rect 987 2682 999 2716
rect 941 2644 999 2682
rect 941 2610 953 2644
rect 987 2610 999 2644
rect 941 2510 999 2610
rect 941 2476 953 2510
rect 987 2476 999 2510
rect 941 2438 999 2476
rect 941 2404 953 2438
rect 987 2404 999 2438
rect 311 667 323 701
rect 357 667 369 701
rect 311 629 369 667
rect 311 595 323 629
rect 357 595 369 629
rect 311 555 369 595
rect 437 701 621 713
rect 437 667 449 701
rect 483 667 575 701
rect 609 667 621 701
rect 437 629 621 667
rect 437 595 449 629
rect 483 595 575 629
rect 609 595 621 629
rect 437 583 621 595
rect 689 701 873 713
rect 689 667 701 701
rect 735 667 827 701
rect 861 667 873 701
rect 689 629 873 667
rect 689 595 701 629
rect 735 595 827 629
rect 861 595 873 629
rect 689 583 873 595
rect 941 701 999 2404
rect 1634 2298 1785 6226
rect 1913 5907 1959 5927
tri 1913 5861 1959 5907 ne
tri 1959 5891 1995 5927 sw
rect 2669 5909 2721 5915
rect 1959 5861 1995 5891
tri 1959 5825 1995 5861 ne
tri 1995 5825 2061 5891 sw
tri 2643 5845 2669 5871 se
rect 2669 5845 2721 5857
tri 1995 5805 2015 5825 ne
tri 1893 4715 1959 4781 se
tri 1873 4695 1893 4715 se
rect 1893 4695 1939 4715
tri 1939 4695 1959 4715 nw
tri 1827 4649 1873 4695 se
rect 1827 3431 1873 4649
tri 1873 4629 1939 4695 nw
tri 1985 4629 2015 4659 se
rect 2015 4639 2061 5825
rect 2669 5787 2721 5793
rect 2453 5590 2721 5596
rect 2505 5538 2669 5590
rect 2453 5526 2721 5538
rect 2505 5474 2669 5526
rect 2453 5468 2721 5474
tri 1949 4593 1985 4629 se
rect 1985 4593 2015 4629
tri 2015 4593 2061 4639 nw
rect 2561 4647 2613 4653
tri 2535 4593 2537 4595 ne
rect 2537 4593 2613 4595
tri 1913 4557 1949 4593 se
rect 1949 4557 1959 4593
rect 1913 4537 1959 4557
tri 1959 4537 2015 4593 nw
tri 2537 4569 2561 4593 ne
rect 2561 4583 2613 4593
tri 2613 4569 2639 4595 nw
rect 2561 4525 2613 4531
rect 2453 3774 2721 3780
rect 2505 3722 2669 3774
rect 2453 3710 2721 3722
rect 2505 3658 2669 3710
rect 2453 3652 2721 3658
rect 1913 3523 1959 3543
tri 1913 3477 1959 3523 ne
tri 1959 3507 1995 3543 sw
rect 2669 3525 2721 3531
rect 1959 3477 1995 3507
tri 1959 3453 1983 3477 ne
rect 1983 3453 1995 3477
tri 1995 3453 2049 3507 sw
tri 2643 3461 2669 3487 se
rect 2669 3461 2721 3473
tri 1983 3451 1985 3453 ne
rect 1985 3451 2049 3453
tri 1873 3431 1893 3451 sw
tri 1985 3441 1995 3451 ne
rect 1995 3441 2049 3451
tri 2049 3441 2061 3453 sw
tri 1995 3431 2005 3441 ne
rect 2005 3431 2061 3441
tri 1827 3419 1839 3431 ne
rect 1839 3419 1893 3431
tri 1893 3419 1905 3431 sw
tri 2005 3421 2015 3431 ne
tri 1839 3381 1877 3419 ne
rect 1877 3381 1905 3419
tri 1905 3381 1943 3419 sw
tri 1877 3365 1893 3381 ne
rect 1893 3365 1943 3381
tri 1943 3365 1959 3381 sw
tri 1893 3347 1911 3365 ne
rect 1911 3347 1959 3365
tri 1911 3299 1959 3347 ne
rect 2015 2425 2061 3431
rect 2669 3403 2721 3409
tri 2061 2425 2067 2431 sw
rect 2015 2419 2067 2425
tri 1785 2298 1810 2323 sw
rect 1692 2292 1877 2298
rect 1692 2285 1759 2292
rect 1634 2278 1759 2285
tri 1634 2258 1654 2278 ne
rect 1654 2258 1759 2278
rect 1793 2258 1831 2292
rect 1865 2258 1877 2292
tri 1654 2252 1660 2258 ne
rect 1660 2252 1877 2258
tri 1886 2166 1913 2193 se
rect 1913 2166 1959 2359
rect 2015 2355 2067 2367
rect 2763 2351 2821 7603
tri 2821 7578 2846 7603 nw
tri 4302 7516 4327 7541 se
rect 4327 7516 4385 7603
tri 4385 7516 4410 7541 sw
rect 2863 7508 4410 7516
rect 2915 7456 3517 7508
rect 3569 7456 3648 7508
rect 2863 7444 3648 7456
rect 2915 7392 3517 7444
rect 3569 7392 3648 7444
rect 3828 7392 3924 7508
rect 4104 7392 4410 7508
rect 2863 7383 4410 7392
tri 3882 7275 3907 7300 ne
rect 3907 7275 3913 7327
rect 3965 7275 3977 7327
rect 4029 7275 4139 7327
tri 4047 7241 4081 7275 ne
rect 4081 7236 4139 7275
rect 3843 7090 3924 7116
tri 3924 7090 3950 7116 sw
rect 3843 7083 3950 7090
rect 3843 7070 3892 7083
tri 3774 7045 3799 7070 ne
rect 2971 7031 3023 7037
tri 2945 6953 2971 6979 ne
rect 2971 6967 3023 6979
tri 3023 6953 3049 6979 nw
rect 2971 6909 3023 6915
tri 3569 5871 3625 5927 se
rect 3625 5907 3671 5927
rect 3625 5871 3635 5907
tri 3635 5871 3671 5907 nw
tri 3543 5845 3569 5871 se
rect 2863 5839 2915 5845
tri 3523 5825 3543 5845 se
rect 3543 5825 3569 5845
rect 2863 5775 2915 5787
tri 2915 5761 2941 5787 nw
rect 2863 5717 2915 5723
rect 2863 5590 3131 5596
rect 2915 5538 3079 5590
rect 2863 5526 3131 5538
rect 2915 5474 3079 5526
rect 2863 5468 3131 5474
rect 2971 4647 3023 4653
rect 3523 4639 3569 5825
tri 3569 5805 3635 5871 nw
tri 3625 4715 3691 4781 sw
tri 3625 4659 3681 4715 ne
rect 3681 4659 3691 4715
tri 3523 4595 3567 4639 ne
rect 3567 4623 3569 4639
tri 3569 4623 3605 4659 sw
tri 3681 4649 3691 4659 ne
tri 3691 4649 3757 4715 sw
tri 3691 4629 3711 4649 ne
rect 3567 4595 3605 4623
tri 2945 4569 2971 4595 ne
rect 2971 4583 3023 4595
tri 3023 4569 3049 4595 nw
tri 3567 4593 3569 4595 ne
rect 3569 4593 3605 4595
tri 3569 4569 3593 4593 ne
rect 3593 4569 3605 4593
tri 3593 4557 3605 4569 ne
tri 3605 4557 3671 4623 sw
tri 3605 4537 3625 4557 ne
rect 3625 4537 3671 4557
rect 2971 4525 3023 4531
rect 2863 3774 3131 3780
rect 2915 3722 3079 3774
rect 2863 3710 3131 3722
rect 2915 3658 3079 3710
rect 2863 3652 3131 3658
tri 3559 3477 3625 3543 se
rect 3625 3523 3671 3543
tri 3625 3477 3671 3523 nw
tri 3543 3461 3559 3477 se
rect 3559 3461 3601 3477
rect 2863 3455 2915 3461
tri 3535 3453 3543 3461 se
rect 3543 3453 3601 3461
tri 3601 3453 3625 3477 nw
tri 3523 3441 3535 3453 se
rect 3535 3441 3569 3453
rect 2863 3391 2919 3403
rect 2915 3381 2919 3391
tri 2919 3381 2941 3403 nw
tri 2915 3377 2919 3381 nw
rect 2863 3333 2915 3339
tri 3517 2425 3523 2431 se
rect 3523 2425 3569 3441
tri 3569 3421 3601 3453 nw
tri 3681 3421 3711 3451 se
rect 3711 3431 3757 4649
rect 3711 3421 3745 3431
tri 3679 3419 3681 3421 se
rect 3681 3419 3745 3421
tri 3745 3419 3757 3431 nw
tri 3645 3385 3679 3419 se
rect 3679 3385 3711 3419
tri 3711 3385 3745 3419 nw
tri 3641 3381 3645 3385 se
rect 3645 3381 3707 3385
tri 3707 3381 3711 3385 nw
tri 3625 3365 3641 3381 se
rect 3641 3365 3691 3381
tri 3691 3365 3707 3381 nw
rect 3625 3347 3673 3365
tri 3673 3347 3691 3365 nw
tri 3625 3299 3673 3347 nw
rect 3517 2419 3569 2425
rect 3517 2355 3569 2367
rect 2015 2224 2067 2303
tri 2722 2298 2728 2304 se
rect 2728 2298 2734 2304
rect 2677 2252 2734 2298
rect 2786 2252 2798 2304
rect 2850 2298 2856 2304
tri 2856 2298 2862 2304 sw
rect 2850 2252 2907 2298
rect 3517 2297 3569 2303
tri 2067 2224 2092 2249 sw
tri 3600 2224 3625 2249 se
rect 3625 2224 3671 2359
tri 3774 2298 3799 2323 se
rect 3799 2298 3950 7070
rect 3707 2292 3950 2298
rect 3707 2258 3719 2292
rect 3753 2258 3791 2292
rect 3825 2278 3950 2292
rect 3825 2258 3924 2278
rect 3707 2252 3924 2258
tri 3924 2252 3950 2278 nw
rect 3993 3453 4039 3465
rect 3993 3419 3999 3453
rect 4033 3419 4039 3453
rect 3993 3381 4039 3419
rect 3993 3347 3999 3381
rect 4033 3347 4039 3381
rect 2015 2221 3671 2224
tri 2015 2195 2041 2221 ne
rect 2041 2195 3645 2221
tri 3645 2195 3671 2221 nw
tri 1959 2166 1986 2193 sw
rect 3993 2192 4039 3347
rect 4081 2220 4139 2222
tri 4039 2192 4064 2217 sw
rect 1595 2140 3543 2166
tri 3543 2140 3569 2166 sw
rect 3993 2146 4154 2192
rect 1595 2137 3569 2140
rect 1152 2028 1392 2034
rect 1204 1976 1340 2028
rect 1152 1964 1392 1976
rect 1204 1912 1340 1964
rect 1445 1936 1503 2099
rect 1595 1936 1653 2137
tri 1653 2110 1680 2137 nw
tri 2142 2110 2169 2137 ne
rect 2169 2110 2231 2137
tri 2169 2109 2170 2110 ne
rect 2170 2109 2231 2110
rect 1718 2103 2064 2109
tri 2170 2106 2173 2109 ne
rect 2173 2106 2231 2109
tri 2231 2106 2262 2137 nw
tri 2410 2106 2441 2137 ne
rect 2174 2104 2230 2105
rect 1718 2069 1730 2103
rect 1764 2069 1802 2103
rect 1836 2069 1874 2103
rect 1908 2069 1946 2103
rect 1980 2069 2018 2103
rect 2052 2069 2064 2103
rect 1718 2063 2064 2069
rect 2174 2067 2230 2068
tri 2170 2063 2173 2066 se
rect 2173 2063 2231 2066
tri 1819 2031 1851 2063 ne
rect 1851 1936 1909 2063
tri 1909 2031 1941 2063 nw
tri 2006 2031 2038 2063 ne
rect 2038 2031 2064 2063
tri 2038 2024 2045 2031 ne
rect 2045 2030 2064 2031
tri 2064 2030 2097 2063 sw
tri 2137 2030 2170 2063 se
rect 2170 2036 2231 2063
tri 2231 2036 2261 2066 sw
rect 2170 2030 2261 2036
rect 2045 1972 2097 2030
rect 2099 2029 2135 2030
rect 2098 1973 2136 2029
rect 2137 2018 2261 2030
rect 2137 1984 2149 2018
rect 2183 1984 2221 2018
rect 2255 1984 2261 2018
rect 2099 1972 2135 1973
rect 2137 1972 2261 1984
tri 2411 2036 2441 2066 se
rect 2441 2036 2499 2137
tri 2499 2106 2530 2137 nw
tri 3054 2109 3082 2137 ne
rect 3082 2109 3143 2137
rect 2558 2103 2976 2109
tri 3082 2106 3085 2109 ne
rect 3085 2106 3143 2109
tri 3143 2106 3174 2137 nw
tri 3322 2106 3353 2137 ne
rect 3086 2104 3142 2105
rect 2558 2069 2570 2103
rect 2604 2069 2642 2103
rect 2676 2069 2714 2103
rect 2748 2069 2786 2103
rect 2820 2069 2858 2103
rect 2892 2069 2930 2103
rect 2964 2069 2976 2103
tri 2499 2036 2529 2066 sw
rect 2558 2063 2976 2069
rect 3086 2067 3142 2068
tri 3082 2063 3085 2066 se
rect 3085 2063 3143 2066
rect 2411 2018 2529 2036
tri 2731 2031 2763 2063 ne
rect 2411 1984 2417 2018
rect 2451 1984 2489 2018
rect 2523 1984 2529 2018
rect 2411 1972 2529 1984
rect 2763 1936 2821 2063
tri 2821 2031 2853 2063 nw
tri 2918 2031 2950 2063 ne
rect 2950 2031 2976 2063
tri 2950 2024 2957 2031 ne
rect 2957 2030 2976 2031
tri 2976 2030 3009 2063 sw
tri 3049 2030 3082 2063 se
rect 3082 2036 3143 2063
tri 3143 2036 3173 2066 sw
rect 3082 2030 3173 2036
rect 2957 1972 3009 2030
rect 3011 2029 3047 2030
rect 3010 1973 3048 2029
rect 3049 2018 3173 2030
rect 3049 1984 3061 2018
rect 3095 1984 3133 2018
rect 3167 1984 3173 2018
rect 3011 1972 3047 1973
rect 3049 1972 3173 1984
tri 3323 2036 3353 2066 se
rect 3353 2036 3411 2137
tri 3411 2106 3442 2137 nw
tri 3491 2111 3517 2137 ne
tri 3411 2036 3441 2066 sw
rect 3323 2018 3441 2036
rect 3323 1984 3329 2018
rect 3363 1984 3401 2018
rect 3435 1984 3441 2018
rect 3323 1972 3441 1984
tri 3490 1936 3517 1963 se
rect 3517 1936 3569 2137
rect 3617 2103 4139 2109
rect 3617 2069 3629 2103
rect 3663 2069 3701 2103
rect 3735 2069 3773 2103
rect 3807 2069 3845 2103
rect 3879 2069 3917 2103
rect 3951 2069 3989 2103
rect 4023 2069 4139 2103
rect 3617 2063 4139 2069
tri 3643 2031 3675 2063 ne
rect 3675 1936 3733 2063
tri 3733 2031 3765 2063 nw
tri 3899 2031 3931 2063 ne
rect 1152 1904 1392 1912
rect 2015 1930 2307 1936
rect 2067 1884 2307 1930
rect 2015 1866 2067 1878
tri 2067 1857 2094 1884 nw
tri 2280 1857 2307 1884 ne
rect 3277 1930 3569 1936
rect 3277 1884 3517 1930
tri 3277 1857 3304 1884 nw
tri 3490 1857 3517 1884 ne
rect 3517 1866 3569 1878
rect 2015 1808 2067 1814
rect 3517 1808 3569 1814
tri 1500 754 1535 789 sw
tri 1819 754 1851 786 se
tri 1909 754 1941 786 sw
tri 2731 754 2763 786 se
tri 2821 754 2853 786 sw
tri 3643 754 3675 786 se
tri 3733 754 3765 786 sw
tri 3899 754 3931 786 se
rect 3931 754 4139 2063
rect 941 667 953 701
rect 987 667 999 701
rect 941 629 999 667
rect 941 595 953 629
rect 987 595 999 629
tri 369 555 396 582 sw
tri 914 555 941 582 se
rect 941 555 999 595
rect 1232 743 1284 749
rect 1232 679 1284 691
rect 1232 615 1284 627
tri 999 555 1026 582 sw
tri 1205 555 1232 582 se
rect 1232 555 1284 563
rect 311 554 1284 555
tri 311 520 345 554 ne
rect 345 548 1284 554
rect 345 520 1239 548
rect 186 486 244 520
tri 345 512 353 520 ne
rect 353 512 1239 520
tri 244 486 270 512 sw
tri 353 503 362 512 ne
rect 362 503 1239 512
tri 1239 503 1284 548 nw
rect 1500 522 4139 754
tri 1426 503 1445 522 se
rect 1445 503 4139 522
tri 1409 486 1426 503 se
rect 1426 486 4139 503
tri 186 461 211 486 ne
rect 211 475 270 486
tri 270 475 281 486 sw
tri 1398 475 1409 486 se
rect 1409 475 4139 486
rect 211 461 272 475
tri 211 427 245 461 ne
rect 245 427 272 461
tri 245 417 255 427 ne
rect 255 417 272 427
rect 993 423 999 475
rect 1051 423 1063 475
rect 1115 423 1121 475
tri 1396 473 1398 475 se
rect 1398 473 4139 475
tri 1281 461 1293 473 se
rect 1293 467 4139 473
rect 1293 461 1503 467
rect 1038 417 1121 423
tri 1261 441 1281 461 se
rect 1281 441 1299 461
rect 1261 427 1299 441
rect 1333 427 1371 461
rect 1405 427 1443 461
rect 1477 427 1503 461
rect 4009 448 4139 467
tri 1503 435 1508 440 nw
rect 1261 421 1503 427
rect 4009 421 4112 448
tri 4112 421 4139 448 nw
rect 1261 415 1483 421
tri 1483 415 1489 421 nw
rect 1261 381 1307 415
tri 1307 390 1332 415 nw
tri 1259 354 1261 356 se
rect 1261 354 1267 381
rect -3 347 55 354
tri 1253 348 1259 354 se
rect 1259 348 1267 354
tri 55 347 56 348 sw
tri 1252 347 1253 348 se
rect 1253 347 1267 348
rect 1301 347 1307 381
rect -3 322 56 347
tri -3 271 48 322 ne
rect 48 317 56 322
tri 56 317 86 347 sw
tri 1222 317 1252 347 se
rect 1252 317 1307 347
rect 48 271 121 317
rect 1259 301 1307 317
rect 1259 271 1277 301
tri 1277 271 1307 301 nw
<< rmetal1 >>
rect 1415 10427 1417 10428
rect 1415 9942 1416 10427
rect 1415 9941 1417 9942
rect 1453 10427 1455 10428
rect 1454 9942 1455 10427
rect 1453 9941 1455 9942
rect 1563 9891 1615 9892
rect 1563 9890 1564 9891
rect 1614 9890 1615 9891
rect 1563 9853 1564 9854
rect 1614 9853 1615 9854
rect 1563 9852 1615 9853
rect 1563 9613 1615 9614
rect 1563 9612 1564 9613
rect 1614 9612 1615 9613
rect 1563 9575 1564 9576
rect 1614 9575 1615 9576
rect 1563 9574 1615 9575
rect 1415 9550 1417 9551
rect 1415 9412 1416 9550
rect 1415 9411 1417 9412
rect 1453 9550 1455 9551
rect 1454 9412 1455 9550
rect 1453 9411 1455 9412
rect 1415 9181 1417 9182
rect 1453 9181 1455 9182
rect 1415 9013 1416 9181
rect 1454 9013 1455 9181
rect 1415 9012 1417 9013
rect 1453 9012 1455 9013
rect 1563 8988 1615 8989
rect 1563 8987 1564 8988
rect 1614 8987 1615 8988
rect 1563 8950 1564 8951
rect 1614 8950 1615 8951
rect 1563 8949 1615 8950
rect 2260 8567 2262 8568
rect 2298 8567 2300 8568
rect 2260 8405 2261 8567
rect 2299 8405 2300 8567
rect 2260 8404 2262 8405
rect 2298 8404 2300 8405
rect 4015 8567 4017 8568
rect 4053 8567 4055 8568
rect 4015 8405 4016 8567
rect 4054 8405 4055 8567
rect 4015 8404 4017 8405
rect 4053 8404 4055 8405
rect 2359 7719 2417 7720
rect 2359 7718 2360 7719
rect 2416 7718 2417 7719
rect 2359 7681 2360 7682
rect 2416 7681 2417 7682
rect 2359 7680 2417 7681
rect 3383 7719 3441 7720
rect 3383 7718 3384 7719
rect 3440 7718 3441 7719
rect 3895 7719 3953 7720
rect 3895 7718 3896 7719
rect 3952 7718 3953 7719
rect 3383 7681 3384 7682
rect 3440 7681 3441 7682
rect 3383 7680 3441 7681
rect 3895 7681 3896 7682
rect 3952 7681 3953 7682
rect 3895 7680 3953 7681
rect 815 6609 873 6610
rect 815 6608 816 6609
rect 872 6608 873 6609
rect 815 6571 816 6572
rect 872 6571 873 6572
rect 815 6570 873 6571
rect 2173 2105 2231 2106
rect 2173 2104 2174 2105
rect 2230 2104 2231 2105
rect 2173 2067 2174 2068
rect 2230 2067 2231 2068
rect 2173 2066 2231 2067
rect 2097 2029 2099 2030
rect 2135 2029 2137 2030
rect 2097 1973 2098 2029
rect 2136 1973 2137 2029
rect 2097 1972 2099 1973
rect 2135 1972 2137 1973
rect 3085 2105 3143 2106
rect 3085 2104 3086 2105
rect 3142 2104 3143 2105
rect 3085 2067 3086 2068
rect 3142 2067 3143 2068
rect 3085 2066 3143 2067
rect 3009 2029 3011 2030
rect 3047 2029 3049 2030
rect 3009 1973 3010 2029
rect 3048 1973 3049 2029
rect 3009 1972 3011 1973
rect 3047 1972 3049 1973
<< via1 >>
rect 2702 11100 2754 11152
rect 2766 11100 2818 11152
rect 2830 11100 2882 11152
rect 4796 11100 4848 11152
rect 4860 11100 4912 11152
rect 4924 11100 4976 11152
rect 4988 11100 5040 11152
rect 5052 11100 5104 11152
rect 7167 11100 7219 11152
rect 7231 11100 7283 11152
rect 7295 11100 7347 11152
rect 7359 11100 7411 11152
rect 7757 11020 7809 11072
rect 7821 11020 7873 11072
rect 7885 11020 7937 11072
rect 7949 11020 8001 11072
rect 8013 11020 8065 11072
rect 2702 10940 2754 10992
rect 2766 10940 2818 10992
rect 2830 10940 2882 10992
rect 4796 10940 4848 10992
rect 4860 10940 4912 10992
rect 4924 10940 4976 10992
rect 4988 10940 5040 10992
rect 5052 10940 5104 10992
rect 7167 10940 7219 10992
rect 7231 10940 7283 10992
rect 7295 10940 7347 10992
rect 7359 10940 7411 10992
rect 1449 10829 1501 10881
rect 1555 10859 1607 10911
rect 1619 10859 1671 10911
rect 8138 10859 8190 10911
rect 8202 10859 8254 10911
rect 8266 10859 8318 10911
rect 8330 10859 8382 10911
rect 1152 10769 1204 10821
rect 999 10681 1051 10733
rect 1063 10681 1115 10733
rect 1152 10705 1204 10757
rect 1449 10765 1501 10817
rect 2977 10786 3029 10838
rect 3041 10786 3093 10838
rect 3105 10786 3157 10838
rect 4517 10786 4569 10838
rect 4581 10786 4633 10838
rect 4645 10786 4697 10838
rect 5473 10786 5525 10838
rect 5537 10786 5589 10838
rect 5601 10786 5653 10838
rect 1449 10740 1501 10753
rect 1449 10706 1457 10740
rect 1457 10706 1491 10740
rect 1491 10706 1501 10740
rect 1449 10701 1501 10706
rect 1449 10668 1501 10689
rect 1449 10637 1457 10668
rect 1457 10637 1491 10668
rect 1491 10637 1501 10668
rect 1232 10552 1284 10604
rect 1232 10488 1284 10540
rect 1449 10596 1501 10625
rect 1449 10573 1457 10596
rect 1457 10573 1491 10596
rect 1491 10573 1501 10596
rect 2015 10674 2067 10726
rect 3517 10674 3569 10726
rect 4651 10674 4703 10726
rect 2015 10610 2067 10662
rect 3517 10610 3569 10662
rect 4651 10610 4703 10662
rect 2015 10546 2067 10598
rect 3517 10546 3569 10598
rect 4651 10546 4703 10598
rect 7822 10546 7938 10726
rect 1232 10424 1284 10476
rect 1449 9822 1501 9823
rect 1449 9788 1456 9822
rect 1456 9788 1490 9822
rect 1490 9788 1501 9822
rect 1449 9771 1501 9788
rect 1449 9750 1501 9759
rect 1449 9716 1456 9750
rect 1456 9716 1490 9750
rect 1490 9716 1501 9750
rect 1449 9707 1501 9716
rect 1449 9678 1501 9695
rect 1449 9644 1456 9678
rect 1456 9644 1490 9678
rect 1490 9644 1501 9678
rect 1449 9643 1501 9644
rect 2015 9771 2067 9823
rect 3517 9771 3569 9823
rect 4651 9771 4703 9823
rect 2015 9707 2067 9759
rect 3517 9707 3569 9759
rect 4651 9707 4703 9759
rect 2015 9643 2067 9695
rect 3517 9643 3569 9695
rect 4651 9643 4703 9695
rect 7822 9643 7938 9823
rect 1449 8919 1501 8920
rect 1449 8885 1456 8919
rect 1456 8885 1490 8919
rect 1490 8885 1501 8919
rect 1449 8868 1501 8885
rect 1152 8786 1204 8838
rect 1152 8722 1204 8774
rect 1449 8847 1501 8856
rect 1449 8813 1456 8847
rect 1456 8813 1490 8847
rect 1490 8813 1501 8847
rect 1449 8804 1501 8813
rect 1449 8775 1501 8792
rect 1449 8741 1456 8775
rect 1456 8741 1490 8775
rect 1490 8741 1501 8775
rect 1449 8740 1501 8741
rect 2015 8868 2067 8920
rect 3517 8868 3569 8920
rect 4651 8868 4703 8920
rect 2015 8804 2067 8856
rect 3517 8804 3569 8856
rect 4651 8804 4703 8856
rect 2015 8740 2067 8792
rect 3517 8740 3569 8792
rect 4651 8740 4703 8792
rect 7822 8740 7938 8920
rect 1152 8658 1204 8710
rect 1152 8566 1204 8618
rect 1152 8502 1204 8554
rect 1152 8438 1204 8490
rect 1756 7392 1936 7508
rect 2015 7456 2067 7508
rect 2669 7456 2721 7508
rect 2015 7392 2067 7444
rect 2669 7392 2721 7444
rect 1555 7275 1607 7327
rect 1619 7275 1671 7327
rect 1340 7150 1392 7202
rect 2525 7150 2577 7202
rect 2589 7150 2641 7202
rect 1232 7070 1284 7122
rect 1232 7006 1284 7058
rect 1232 6942 1284 6994
rect 1340 7086 1392 7138
rect 1340 7022 1392 7074
rect 1340 6958 1392 7010
rect 1340 6894 1392 6946
rect 1340 6830 1392 6882
rect 1069 6681 1078 6712
rect 1078 6681 1112 6712
rect 1112 6681 1121 6712
rect 1069 6660 1121 6681
rect 1069 6643 1121 6648
rect 1069 6609 1078 6643
rect 1078 6609 1112 6643
rect 1112 6609 1121 6643
rect 1069 6596 1121 6609
rect 1069 6571 1121 6584
rect 1069 6537 1078 6571
rect 1078 6537 1112 6571
rect 1112 6537 1121 6571
rect 1069 6532 1121 6537
rect 1069 6499 1121 6520
rect 1069 6468 1078 6499
rect 1078 6468 1112 6499
rect 1112 6468 1121 6499
rect 1232 6692 1284 6744
rect 1232 6628 1284 6680
rect 1232 6564 1284 6616
rect 1232 6500 1284 6552
rect 1232 6436 1284 6488
rect 2561 6979 2613 7031
rect 2561 6915 2613 6967
rect 1232 6179 1284 6231
rect 1232 6115 1284 6167
rect 1232 6051 1284 6103
rect 2669 5857 2721 5909
rect 2669 5793 2721 5845
rect 2453 5538 2505 5590
rect 2669 5538 2721 5590
rect 2453 5474 2505 5526
rect 2669 5474 2721 5526
rect 2561 4595 2613 4647
rect 2561 4531 2613 4583
rect 2453 3722 2505 3774
rect 2669 3722 2721 3774
rect 2453 3658 2505 3710
rect 2669 3658 2721 3710
rect 2669 3473 2721 3525
rect 2669 3409 2721 3461
rect 2015 2367 2067 2419
rect 2015 2303 2067 2355
rect 2863 7456 2915 7508
rect 3517 7456 3569 7508
rect 2863 7392 2915 7444
rect 3517 7392 3569 7444
rect 3648 7392 3828 7508
rect 3924 7392 4104 7508
rect 3913 7275 3965 7327
rect 3977 7275 4029 7327
rect 2971 6979 3023 7031
rect 2971 6915 3023 6967
rect 2863 5787 2915 5839
rect 2863 5723 2915 5775
rect 2863 5538 2915 5590
rect 3079 5538 3131 5590
rect 2863 5474 2915 5526
rect 3079 5474 3131 5526
rect 2971 4595 3023 4647
rect 2971 4531 3023 4583
rect 2863 3722 2915 3774
rect 3079 3722 3131 3774
rect 2863 3658 2915 3710
rect 3079 3658 3131 3710
rect 2863 3403 2915 3455
rect 2863 3339 2915 3391
rect 3517 2367 3569 2419
rect 2734 2252 2786 2304
rect 2798 2252 2850 2304
rect 3517 2303 3569 2355
rect 1152 1976 1204 2028
rect 1340 2022 1392 2028
rect 1340 1988 1349 2022
rect 1349 1988 1383 2022
rect 1383 1988 1392 2022
rect 1340 1976 1392 1988
rect 1152 1912 1204 1964
rect 1340 1950 1392 1964
rect 1340 1916 1349 1950
rect 1349 1916 1383 1950
rect 1383 1916 1392 1950
rect 1340 1912 1392 1916
rect 2015 1878 2067 1930
rect 2015 1814 2067 1866
rect 3517 1878 3569 1930
rect 3517 1814 3569 1866
rect 1232 691 1284 743
rect 1232 627 1284 679
rect 1232 563 1284 615
rect 999 423 1051 475
rect 1063 423 1115 475
<< metal2 >>
rect 2669 11100 2702 11152
rect 2754 11100 2766 11152
rect 2818 11100 2830 11152
rect 2882 11100 2915 11152
rect 2669 10992 2915 11100
rect 2669 10940 2702 10992
rect 2754 10940 2766 10992
rect 2818 10940 2830 10992
rect 2882 10940 2915 10992
tri -82 475 0 557 se
rect 0 475 133 10912
rect 1448 10911 1677 10912
rect 1448 10881 1555 10911
rect 1448 10829 1449 10881
rect 1501 10859 1555 10881
rect 1607 10859 1619 10911
rect 1671 10859 1677 10911
rect 1501 10829 1677 10859
rect 1152 10821 1204 10827
rect 1152 10757 1204 10769
tri -134 423 -82 475 se
rect -82 423 133 475
tri -286 271 -134 423 se
rect -134 271 133 423
rect -286 226 133 271
rect 189 226 317 10733
rect 373 226 937 10733
rect 993 10681 999 10733
rect 1051 10681 1063 10733
rect 1115 10681 1121 10733
rect 993 6712 1121 10681
rect 1152 8838 1204 10705
rect 1448 10817 1677 10829
rect 1448 10765 1449 10817
rect 1501 10765 1677 10817
rect 1448 10753 1677 10765
rect 1448 10701 1449 10753
rect 1501 10701 1677 10753
rect 1448 10689 1677 10701
rect 1448 10637 1449 10689
rect 1501 10637 1677 10689
rect 1448 10625 1677 10637
rect 1152 8774 1204 8786
rect 1152 8710 1204 8722
rect 1152 8652 1204 8658
rect 1232 10604 1284 10610
rect 1232 10540 1284 10552
rect 1232 10476 1284 10488
rect 993 6660 1069 6712
rect 993 6648 1121 6660
rect 993 6596 1069 6648
rect 993 6584 1121 6596
rect 993 6532 1069 6584
rect 993 6520 1121 6532
rect 993 6468 1069 6520
rect 993 475 1121 6468
rect 1152 8618 1204 8624
rect 1152 8554 1204 8566
rect 1152 8490 1204 8502
rect 1152 2028 1204 8438
rect 1152 1964 1204 1976
rect 1152 1906 1204 1912
rect 1232 7122 1284 10424
rect 1448 10573 1449 10625
rect 1501 10573 1677 10625
rect 1448 9823 1677 10573
rect 1448 9771 1449 9823
rect 1501 9771 1677 9823
rect 1448 9759 1677 9771
rect 1448 9707 1449 9759
rect 1501 9707 1677 9759
rect 1448 9695 1677 9707
rect 1448 9643 1449 9695
rect 1501 9643 1677 9695
rect 1232 7058 1284 7070
rect 1232 6994 1284 7006
rect 1232 6744 1284 6942
rect 1340 7202 1392 9012
rect 1340 7138 1392 7150
rect 1340 7074 1392 7086
rect 1340 7010 1392 7022
rect 1340 6946 1392 6958
rect 1340 6882 1392 6894
rect 1340 6824 1392 6830
rect 1448 8920 1677 9643
rect 1448 8868 1449 8920
rect 1501 8868 1677 8920
rect 1448 8856 1677 8868
rect 1448 8804 1449 8856
rect 1501 8804 1677 8856
rect 1448 8792 1677 8804
rect 1448 8740 1449 8792
rect 1501 8740 1677 8792
rect 1448 7327 1677 8740
rect 1448 7275 1555 7327
rect 1607 7275 1619 7327
rect 1671 7275 1677 7327
rect 1232 6680 1284 6692
rect 1232 6616 1284 6628
rect 1232 6552 1284 6564
rect 1232 6488 1284 6500
rect 1232 6231 1284 6436
rect 1232 6167 1284 6179
rect 1232 6103 1284 6115
rect 1232 743 1284 6051
rect 1232 679 1284 691
rect 1232 615 1284 627
rect 1232 557 1284 563
rect 1340 2028 1392 2034
rect 1340 1964 1392 1976
rect 993 423 999 475
rect 1051 423 1063 475
rect 1115 423 1121 475
rect 993 260 1121 423
rect 1340 400 1392 1912
rect 1448 715 1677 7275
rect 1733 7508 1959 10732
rect 1733 7392 1756 7508
rect 1936 7392 1959 7508
rect 1733 1130 1959 7392
rect 2015 10726 2067 10732
rect 2015 10662 2067 10674
rect 2015 10598 2067 10610
rect 2015 9823 2067 10546
rect 2015 9759 2067 9771
rect 2015 9695 2067 9707
rect 2015 8920 2067 9643
rect 2015 8856 2067 8868
rect 2015 8792 2067 8804
rect 2015 7508 2067 8740
rect 2015 7444 2067 7456
rect 2015 2473 2067 7392
rect 2123 7284 2505 10732
rect 2123 7068 2497 7284
tri 2497 7276 2505 7284 nw
tri 2525 7208 2561 7244 se
rect 2561 7216 2613 10732
rect 2669 7508 2915 10940
tri 4647 10859 4651 10863 se
rect 4651 10859 4703 11152
tri 4626 10838 4647 10859 se
rect 4647 10838 4703 10859
rect 2721 7456 2863 7508
rect 2669 7444 2915 7456
rect 2721 7392 2863 7444
tri 2613 7216 2641 7244 sw
rect 2561 7208 2641 7216
rect 2525 7202 2641 7208
rect 2577 7150 2589 7202
rect 2525 7144 2641 7150
tri 2525 7108 2561 7144 ne
rect 2561 7136 2641 7144
tri 2497 7068 2505 7076 sw
rect 2123 5590 2505 7068
rect 2123 5538 2453 5590
rect 2123 5526 2505 5538
rect 2123 5474 2453 5526
rect 2123 3774 2505 5474
rect 2123 3722 2453 3774
rect 2123 3710 2505 3722
rect 2123 3658 2453 3710
rect 2015 2419 2067 2425
rect 2015 2355 2067 2367
rect 2015 1930 2067 2303
rect 2015 1866 2067 1878
rect 2015 1808 2067 1814
rect 2123 1387 2505 3658
tri 2123 1204 2306 1387 ne
rect 1733 862 1916 1130
tri 1916 1087 1959 1130 nw
tri 2188 887 2306 1005 se
rect 2306 887 2505 1387
tri 1916 862 1941 887 sw
tri 2163 862 2188 887 se
rect 2188 862 2505 887
rect 1733 839 2505 862
tri 1733 801 1771 839 ne
rect 1771 801 2505 839
tri 1677 715 1763 801 sw
tri 1771 715 1857 801 ne
rect 1857 715 2505 801
rect 1448 621 1763 715
tri 1763 621 1857 715 sw
tri 1857 621 1951 715 ne
rect 1951 621 2505 715
rect 1448 602 1857 621
tri 1392 400 1398 406 sw
rect 1448 400 1571 602
tri 1571 577 1596 602 nw
tri 1630 577 1655 602 ne
rect 1655 577 1857 602
tri 1655 452 1780 577 ne
rect 1780 563 1857 577
tri 1857 563 1915 621 sw
tri 1951 563 2009 621 ne
rect 2009 563 2505 621
rect 1780 469 1915 563
tri 1915 469 2009 563 sw
rect 1780 400 2009 469
tri 2009 449 2123 563 ne
rect 2123 400 2505 563
rect 2561 7031 2613 7136
tri 2613 7108 2641 7136 nw
rect 2561 6967 2613 6979
rect 2561 5731 2613 6915
rect 2669 6036 2915 7392
tri 2669 6009 2696 6036 ne
rect 2696 6009 2888 6036
tri 2888 6009 2915 6036 nw
rect 2971 10786 2977 10838
rect 3029 10786 3041 10838
rect 3093 10786 3105 10838
rect 3157 10786 3163 10838
rect 4511 10786 4517 10838
rect 4569 10786 4581 10838
rect 4633 10786 4645 10838
rect 4697 10786 4703 10838
rect 4759 11100 4796 11152
rect 4848 11100 4860 11152
rect 4912 11100 4924 11152
rect 4976 11100 4988 11152
rect 5040 11100 5052 11152
rect 5104 11100 5141 11152
rect 4759 10992 5141 11100
rect 4759 10940 4796 10992
rect 4848 10940 4860 10992
rect 4912 10940 4924 10992
rect 4976 10940 4988 10992
rect 5040 10940 5052 10992
rect 5104 10940 5141 10992
rect 2971 7031 3023 10786
tri 3023 10761 3048 10786 nw
rect 2971 6967 3023 6979
tri 2944 5953 2971 5980 se
rect 2971 5953 3023 6915
tri 2669 5915 2707 5953 se
rect 2707 5915 3023 5953
rect 2669 5909 3023 5915
rect 2721 5901 3023 5909
tri 2721 5874 2748 5901 nw
tri 2944 5874 2971 5901 ne
rect 2669 5845 2721 5857
rect 2669 5787 2721 5793
rect 2863 5839 2915 5845
rect 2863 5775 2915 5787
tri 2613 5731 2640 5758 sw
tri 2836 5731 2863 5758 se
rect 2561 5723 2863 5731
rect 2561 5717 2915 5723
rect 2561 5679 2877 5717
tri 2877 5679 2915 5717 nw
rect 2561 4647 2613 5679
tri 2613 5652 2640 5679 nw
rect 2561 4583 2613 4595
rect 2561 3347 2613 4531
tri 2669 5596 2696 5623 se
rect 2696 5596 2888 5623
tri 2888 5596 2915 5623 sw
rect 2669 5590 2915 5596
rect 2721 5538 2863 5590
rect 2669 5526 2915 5538
rect 2721 5474 2863 5526
rect 2669 3774 2915 5474
rect 2721 3722 2863 3774
rect 2669 3710 2915 3722
rect 2721 3658 2863 3710
rect 2669 3652 2915 3658
tri 2669 3625 2696 3652 ne
rect 2696 3625 2888 3652
tri 2888 3625 2915 3652 nw
rect 2971 4647 3023 5901
rect 2971 4583 3023 4595
tri 2944 3569 2971 3596 se
rect 2971 3569 3023 4531
tri 2669 3531 2707 3569 se
rect 2707 3531 3023 3569
rect 2669 3525 3023 3531
rect 2721 3517 3023 3525
tri 2721 3490 2748 3517 nw
tri 2944 3490 2971 3517 ne
rect 2669 3461 2721 3473
rect 2669 3403 2721 3409
rect 2863 3455 2915 3461
rect 2863 3391 2915 3403
tri 2613 3347 2640 3374 sw
tri 2836 3347 2863 3374 se
rect 2561 3339 2863 3347
rect 2561 3333 2915 3339
rect 2561 3295 2877 3333
tri 2877 3295 2915 3333 nw
rect 2561 400 2613 3295
tri 2613 3268 2640 3295 nw
tri 2669 3212 2696 3239 se
rect 2696 3212 2888 3239
tri 2888 3212 2915 3239 sw
rect 2669 2304 2915 3212
rect 2669 2252 2734 2304
rect 2786 2252 2798 2304
rect 2850 2252 2915 2304
rect 2669 400 2915 2252
rect 2971 400 3023 3517
rect 3079 5590 3461 10732
rect 3131 5538 3461 5590
rect 3079 5526 3461 5538
rect 3131 5474 3461 5526
rect 3079 3774 3461 5474
rect 3131 3722 3461 3774
rect 3079 3710 3461 3722
rect 3131 3658 3461 3710
rect 3079 400 3461 3658
rect 3517 10726 3569 10732
rect 3517 10662 3569 10674
rect 3517 10598 3569 10610
rect 3517 9823 3569 10546
rect 3517 9759 3569 9771
rect 3517 9695 3569 9707
rect 3517 8920 3569 9643
rect 3517 8856 3569 8868
rect 3517 8792 3569 8804
rect 3517 7508 3569 8740
rect 3517 7444 3569 7456
rect 3517 2473 3569 7392
rect 3625 7508 3851 10732
rect 3625 7392 3648 7508
rect 3828 7392 3851 7508
rect 3517 2419 3569 2425
rect 3517 2355 3569 2367
rect 3517 1930 3569 2303
rect 3517 1866 3569 1878
rect 3517 1808 3569 1814
tri 3517 1676 3625 1784 se
rect 3625 1676 3851 7392
rect 3907 7508 4313 10732
rect 4369 8734 4595 10732
rect 4651 10726 4703 10732
rect 4651 10662 4703 10674
rect 4651 10598 4703 10610
rect 4651 9823 4703 10546
rect 4651 9759 4703 9771
rect 4651 9695 4703 9707
rect 4651 8920 4703 9643
rect 4651 8856 4703 8868
rect 4651 8792 4703 8804
rect 4651 8734 4703 8740
rect 4759 8734 5141 10940
rect 7155 11100 7167 11152
rect 7219 11100 7231 11152
rect 7283 11100 7295 11152
rect 7347 11100 7359 11152
rect 7411 11100 7423 11152
rect 7155 10992 7423 11100
rect 7751 11020 7757 11072
rect 7809 11020 7821 11072
rect 7873 11020 7885 11072
rect 7937 11020 7949 11072
rect 8001 11020 8013 11072
rect 8065 11020 8071 11072
tri 7994 10995 8019 11020 ne
rect 7155 10940 7167 10992
rect 7219 10940 7231 10992
rect 7283 10940 7295 10992
rect 7347 10940 7359 10992
rect 7411 10940 7423 10992
rect 5467 10786 5473 10838
rect 5525 10786 5537 10838
rect 5589 10786 5601 10838
rect 5653 10786 5659 10838
tri 5582 10761 5607 10786 ne
rect 5197 8734 5249 10732
rect 5305 8734 5551 10732
rect 5607 8734 5659 10786
rect 5715 8734 6097 10732
rect 6153 8734 6205 10732
rect 6261 8734 6487 10732
rect 6543 8734 6772 10732
rect 6831 8734 7099 10732
rect 7155 8734 7423 10940
rect 7479 8734 7747 10732
rect 7803 10726 7957 10732
rect 7803 10546 7822 10726
rect 7938 10546 7957 10726
rect 7803 9823 7957 10546
rect 7803 9643 7822 9823
rect 7938 9643 7957 9823
rect 7803 8920 7957 9643
rect 7803 8740 7822 8920
rect 7938 8740 7957 8920
rect 8019 8786 8071 11020
rect 8132 10911 8522 10912
rect 8132 10859 8138 10911
rect 8190 10859 8202 10911
rect 8254 10859 8266 10911
rect 8318 10859 8330 10911
rect 8382 10859 8522 10911
tri 8229 10763 8325 10859 ne
rect 7803 8734 7957 8740
rect 8127 8734 8272 10732
rect 8325 8734 8522 10859
rect 3907 7392 3924 7508
rect 4104 7392 4313 7508
rect 3907 7386 4313 7392
rect 3517 400 3851 1676
rect 3907 7275 3913 7327
rect 3965 7275 3977 7327
rect 4029 7275 4136 7327
rect 3907 508 4136 7275
tri 3907 400 4015 508 ne
rect 4015 400 4136 508
tri 1121 260 1132 271 sw
rect 993 226 1132 260
rect 1340 266 1398 400
tri 1398 266 1532 400 sw
tri 4015 372 4043 400 ne
rect 4043 372 4136 400
rect 1340 226 1532 266
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_0
timestamp 1704896540
transform 0 -1 369 -1 0 2530
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_1
timestamp 1704896540
transform 0 -1 495 -1 0 2530
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_2
timestamp 1704896540
transform 0 -1 621 -1 0 2530
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_3
timestamp 1704896540
transform 0 -1 747 -1 0 2530
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_4
timestamp 1704896540
transform 0 -1 873 -1 0 2530
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_5
timestamp 1704896540
transform 0 -1 999 -1 0 2530
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_6
timestamp 1704896540
transform 0 -1 999 -1 0 4545
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_7
timestamp 1704896540
transform 0 -1 873 -1 0 4545
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_8
timestamp 1704896540
transform 0 -1 747 -1 0 4545
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_9
timestamp 1704896540
transform 0 -1 621 -1 0 4545
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_10
timestamp 1704896540
transform 0 -1 495 -1 0 4545
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_11
timestamp 1704896540
transform 0 -1 369 -1 0 4545
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_12
timestamp 1704896540
transform 0 -1 369 -1 0 6560
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_13
timestamp 1704896540
transform 0 -1 495 -1 0 6560
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_14
timestamp 1704896540
transform 0 -1 621 -1 0 6560
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_15
timestamp 1704896540
transform 0 -1 747 -1 0 6560
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_16
timestamp 1704896540
transform 0 -1 873 -1 0 6560
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_17
timestamp 1704896540
transform 0 -1 999 -1 0 6560
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_18
timestamp 1704896540
transform 0 -1 999 -1 0 8575
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_19
timestamp 1704896540
transform 0 -1 873 -1 0 8575
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_20
timestamp 1704896540
transform 0 -1 747 -1 0 8575
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_21
timestamp 1704896540
transform 0 -1 621 -1 0 8575
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_22
timestamp 1704896540
transform 0 -1 495 -1 0 8575
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_23
timestamp 1704896540
transform 0 -1 369 -1 0 8575
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_24
timestamp 1704896540
transform 0 -1 999 -1 0 10590
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_25
timestamp 1704896540
transform 0 -1 873 -1 0 10590
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_26
timestamp 1704896540
transform 0 -1 747 -1 0 10590
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_27
timestamp 1704896540
transform 0 -1 621 -1 0 10590
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_28
timestamp 1704896540
transform 0 -1 495 -1 0 10590
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_29
timestamp 1704896540
transform 0 -1 369 -1 0 10590
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_30
timestamp 1704896540
transform 0 -1 999 1 0 575
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_31
timestamp 1704896540
transform 0 -1 873 1 0 575
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_32
timestamp 1704896540
transform 0 -1 747 1 0 575
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_33
timestamp 1704896540
transform 0 -1 621 1 0 575
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_34
timestamp 1704896540
transform 0 -1 495 1 0 575
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_35
timestamp 1704896540
transform 0 -1 369 1 0 575
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_36
timestamp 1704896540
transform 0 -1 369 1 0 2590
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_37
timestamp 1704896540
transform 0 -1 495 1 0 2590
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_38
timestamp 1704896540
transform 0 -1 621 1 0 2590
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_39
timestamp 1704896540
transform 0 -1 747 1 0 2590
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_40
timestamp 1704896540
transform 0 -1 873 1 0 2590
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_41
timestamp 1704896540
transform 0 -1 999 1 0 2590
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_42
timestamp 1704896540
transform 0 -1 999 1 0 4605
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_43
timestamp 1704896540
transform 0 -1 873 1 0 4605
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_44
timestamp 1704896540
transform 0 -1 747 1 0 4605
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_45
timestamp 1704896540
transform 0 -1 621 1 0 4605
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_46
timestamp 1704896540
transform 0 -1 495 1 0 4605
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_47
timestamp 1704896540
transform 0 -1 369 1 0 4605
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_48
timestamp 1704896540
transform 0 -1 369 1 0 6620
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_49
timestamp 1704896540
transform 0 -1 495 1 0 6620
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_50
timestamp 1704896540
transform 0 -1 621 1 0 6620
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_51
timestamp 1704896540
transform 0 -1 747 1 0 6620
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_52
timestamp 1704896540
transform 0 -1 873 1 0 6620
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_53
timestamp 1704896540
transform 0 -1 999 1 0 6620
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_54
timestamp 1704896540
transform 0 -1 999 1 0 8635
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_55
timestamp 1704896540
transform 0 -1 873 1 0 8635
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_56
timestamp 1704896540
transform 0 -1 747 1 0 8635
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_57
timestamp 1704896540
transform 0 -1 621 1 0 8635
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_58
timestamp 1704896540
transform 0 -1 495 1 0 8635
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_59
timestamp 1704896540
transform 0 -1 369 1 0 8635
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_0
timestamp 1704896540
transform -1 0 987 0 1 8449
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_1
timestamp 1704896540
transform -1 0 861 0 1 8449
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_2
timestamp 1704896540
transform -1 0 861 0 1 10464
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_3
timestamp 1704896540
transform -1 0 735 0 1 10464
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_4
timestamp 1704896540
transform -1 0 609 0 1 10464
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_5
timestamp 1704896540
transform -1 0 483 0 1 10464
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_6
timestamp 1704896540
transform -1 0 357 0 1 10464
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_7
timestamp 1704896540
transform -1 0 357 0 1 8449
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_8
timestamp 1704896540
transform -1 0 483 0 1 8449
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_9
timestamp 1704896540
transform -1 0 609 0 1 8449
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_10
timestamp 1704896540
transform -1 0 735 0 1 8449
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_11
timestamp 1704896540
transform -1 0 987 0 1 10464
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_12
timestamp 1704896540
transform -1 0 357 0 1 6434
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_13
timestamp 1704896540
transform -1 0 483 0 1 6434
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_14
timestamp 1704896540
transform -1 0 609 0 1 6434
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_15
timestamp 1704896540
transform -1 0 735 0 1 6434
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_16
timestamp 1704896540
transform -1 0 861 0 1 6434
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_17
timestamp 1704896540
transform -1 0 987 0 1 6434
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_18
timestamp 1704896540
transform -1 0 357 0 1 4419
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_19
timestamp 1704896540
transform -1 0 483 0 1 4419
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_20
timestamp 1704896540
transform -1 0 609 0 1 4419
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_21
timestamp 1704896540
transform -1 0 735 0 1 4419
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_22
timestamp 1704896540
transform -1 0 861 0 1 4419
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_23
timestamp 1704896540
transform -1 0 987 0 1 4419
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_24
timestamp 1704896540
transform -1 0 357 0 1 2404
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_25
timestamp 1704896540
transform -1 0 483 0 1 2404
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_26
timestamp 1704896540
transform -1 0 609 0 1 2404
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_27
timestamp 1704896540
transform -1 0 735 0 1 2404
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_28
timestamp 1704896540
transform -1 0 861 0 1 2404
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_29
timestamp 1704896540
transform -1 0 987 0 1 2404
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_30
timestamp 1704896540
transform -1 0 357 0 -1 8761
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_31
timestamp 1704896540
transform -1 0 483 0 -1 8761
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_32
timestamp 1704896540
transform -1 0 609 0 -1 8761
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_33
timestamp 1704896540
transform -1 0 735 0 -1 8761
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_34
timestamp 1704896540
transform -1 0 861 0 -1 8761
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_35
timestamp 1704896540
transform -1 0 987 0 -1 8761
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_36
timestamp 1704896540
transform -1 0 357 0 -1 6746
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_37
timestamp 1704896540
transform -1 0 483 0 -1 6746
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_38
timestamp 1704896540
transform -1 0 609 0 -1 6746
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_39
timestamp 1704896540
transform -1 0 735 0 -1 6746
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_40
timestamp 1704896540
transform -1 0 861 0 -1 6746
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_41
timestamp 1704896540
transform -1 0 987 0 -1 6746
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_42
timestamp 1704896540
transform -1 0 357 0 -1 4731
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_43
timestamp 1704896540
transform -1 0 483 0 -1 4731
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_44
timestamp 1704896540
transform -1 0 609 0 -1 4731
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_45
timestamp 1704896540
transform -1 0 735 0 -1 4731
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_46
timestamp 1704896540
transform -1 0 861 0 -1 4731
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_47
timestamp 1704896540
transform -1 0 987 0 -1 4731
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_48
timestamp 1704896540
transform -1 0 357 0 -1 2716
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_49
timestamp 1704896540
transform -1 0 483 0 -1 2716
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_50
timestamp 1704896540
transform -1 0 609 0 -1 2716
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_51
timestamp 1704896540
transform -1 0 735 0 -1 2716
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_52
timestamp 1704896540
transform -1 0 861 0 -1 2716
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_53
timestamp 1704896540
transform -1 0 987 0 -1 2716
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_54
timestamp 1704896540
transform -1 0 357 0 -1 701
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_55
timestamp 1704896540
transform -1 0 483 0 -1 701
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_56
timestamp 1704896540
transform -1 0 609 0 -1 701
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_57
timestamp 1704896540
transform -1 0 735 0 -1 701
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_58
timestamp 1704896540
transform -1 0 861 0 -1 701
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_59
timestamp 1704896540
transform -1 0 987 0 -1 701
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_60
timestamp 1704896540
transform 0 1 2417 1 0 1984
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_61
timestamp 1704896540
transform 0 1 3329 1 0 1984
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_62
timestamp 1704896540
transform 0 -1 2255 1 0 1984
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_63
timestamp 1704896540
transform 0 -1 3167 1 0 1984
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_64
timestamp 1704896540
transform 1 0 1690 0 -1 8920
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1704896540
transform 0 1 3999 -1 0 3453
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1704896540
transform -1 0 2011 0 1 8590
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1704896540
transform -1 0 3825 0 1 2258
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1704896540
transform 0 1 4251 1 0 8506
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_4
timestamp 1704896540
transform 0 -1 1383 1 0 1916
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_5
timestamp 1704896540
transform 1 0 1759 0 1 2258
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_0
timestamp 1704896540
transform 0 1 1299 1 0 427
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_1
timestamp 1704896540
transform 1 0 1456 0 -1 8919
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_2
timestamp 1704896540
transform 1 0 1456 0 -1 9822
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_3
timestamp 1704896540
transform 1 0 1691 0 1 10546
box 0 0 1 1
use L1M1_CDNS_52468879185192  L1M1_CDNS_52468879185192_4
timestamp 1704896540
transform 1 0 1690 0 1 9644
box 0 0 1 1
use L1M1_CDNS_52468879185193  L1M1_CDNS_52468879185193_0
timestamp 1704896540
transform -1 0 2052 0 1 2069
box 0 0 1 1
use L1M1_CDNS_52468879185195  L1M1_CDNS_52468879185195_0
timestamp 1704896540
transform -1 0 3457 0 1 2258
box -12 -6 550 40
use L1M1_CDNS_52468879185195  L1M1_CDNS_52468879185195_1
timestamp 1704896540
transform 1 0 2127 0 1 2258
box -12 -6 550 40
use L1M1_CDNS_52468879185308  L1M1_CDNS_52468879185308_0
timestamp 1704896540
transform -1 0 4023 0 1 2069
box 0 0 1 1
use L1M1_CDNS_52468879185308  L1M1_CDNS_52468879185308_1
timestamp 1704896540
transform -1 0 2964 0 1 2069
box 0 0 1 1
use L1M1_CDNS_52468879185316  L1M1_CDNS_52468879185316_0
timestamp 1704896540
transform 0 -1 1776 -1 0 7017
box -12 -6 622 40
use L1M1_CDNS_52468879185326  L1M1_CDNS_52468879185326_0
timestamp 1704896540
transform 0 -1 1491 1 0 6413
box -12 -6 694 40
use L1M1_CDNS_52468879185335  L1M1_CDNS_52468879185335_0
timestamp 1704896540
transform 1 0 133 0 -1 311
box -12 -6 1126 40
use L1M1_CDNS_52468879185381  L1M1_CDNS_52468879185381_0
timestamp 1704896540
transform 1 0 1797 0 1 7476
box -12 -6 910 40
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_0
timestamp 1704896540
transform 0 1 1267 -1 0 381
box 0 0 1 1
use L1M1_CDNS_52468879185955  L1M1_CDNS_52468879185955_0
timestamp 1704896540
transform 0 1 3805 -1 0 3333
box -12 -6 982 40
use L1M1_CDNS_52468879185955  L1M1_CDNS_52468879185955_1
timestamp 1704896540
transform -1 0 2723 0 1 7076
box -12 -6 982 40
use L1M1_CDNS_52468879185955  L1M1_CDNS_52468879185955_2
timestamp 1704896540
transform 1 0 2861 0 1 7076
box -12 -6 982 40
use L1M1_CDNS_52468879185956  L1M1_CDNS_52468879185956_0
timestamp 1704896540
transform 1 0 1515 0 1 427
box -12 -6 2494 40
use L1M1_CDNS_524688791851011  L1M1_CDNS_524688791851011_0
timestamp 1704896540
transform -1 0 4047 0 1 7287
box -12 -6 1198 40
use L1M1_CDNS_524688791851011  L1M1_CDNS_524688791851011_1
timestamp 1704896540
transform -1 0 4075 0 1 7476
box -12 -6 1198 40
use L1M1_CDNS_524688791851011  L1M1_CDNS_524688791851011_2
timestamp 1704896540
transform 1 0 1537 0 1 7287
box -12 -6 1198 40
use L1M1_CDNS_524688791851014  L1M1_CDNS_524688791851014_0
timestamp 1704896540
transform 0 1 278 1 0 429
box -12 -6 46 760
use L1M1_CDNS_524688791851014  L1M1_CDNS_524688791851014_1
timestamp 1704896540
transform 0 1 278 1 0 10690
box -12 -6 46 760
use L1M1_CDNS_524688791851014  L1M1_CDNS_524688791851014_2
timestamp 1704896540
transform 1 0 1939 0 -1 8363
box -12 -6 46 760
use L1M1_CDNS_524688791851015  L1M1_CDNS_524688791851015_0
timestamp 1704896540
transform 1 0 4339 0 1 7609
box -12 -6 46 904
use L1M1_CDNS_524688791851015  L1M1_CDNS_524688791851015_1
timestamp 1704896540
transform 1 0 2115 0 1 7660
box -12 -6 46 904
use L1M1_CDNS_524688791851015  L1M1_CDNS_524688791851015_2
timestamp 1704896540
transform 1 0 1763 0 1 7660
box -12 -6 46 904
use L1M1_CDNS_524688791851015  L1M1_CDNS_524688791851015_3
timestamp 1704896540
transform 1 0 4163 0 1 7660
box -12 -6 46 904
use L1M1_CDNS_524688791851016  L1M1_CDNS_524688791851016_0
timestamp 1704896540
transform 0 1 2869 1 0 6991
box -12 -6 46 616
use L1M1_CDNS_524688791851016  L1M1_CDNS_524688791851016_1
timestamp 1704896540
transform 0 1 2869 1 0 3415
box -12 -6 46 616
use L1M1_CDNS_524688791851016  L1M1_CDNS_524688791851016_2
timestamp 1704896540
transform 0 1 2869 1 0 5799
box -12 -6 46 616
use L1M1_CDNS_524688791851016  L1M1_CDNS_524688791851016_3
timestamp 1704896540
transform 0 1 2869 1 0 4607
box -12 -6 46 616
use L1M1_CDNS_524688791851016  L1M1_CDNS_524688791851016_4
timestamp 1704896540
transform 0 -1 2715 1 0 6991
box -12 -6 46 616
use L1M1_CDNS_524688791851016  L1M1_CDNS_524688791851016_5
timestamp 1704896540
transform 0 -1 2715 1 0 4607
box -12 -6 46 616
use L1M1_CDNS_524688791851016  L1M1_CDNS_524688791851016_6
timestamp 1704896540
transform 0 -1 2715 1 0 3415
box -12 -6 46 616
use L1M1_CDNS_524688791851016  L1M1_CDNS_524688791851016_7
timestamp 1704896540
transform 0 -1 2715 1 0 5799
box -12 -6 46 616
use L1M1_CDNS_524688791851016  L1M1_CDNS_524688791851016_8
timestamp 1704896540
transform 1 0 2883 0 -1 8342
box -12 -6 46 616
use L1M1_CDNS_524688791851016  L1M1_CDNS_524688791851016_9
timestamp 1704896540
transform 1 0 2371 0 -1 8342
box -12 -6 46 616
use L1M1_CDNS_524688791851016  L1M1_CDNS_524688791851016_10
timestamp 1704896540
transform 1 0 3395 0 -1 8342
box -12 -6 46 616
use L1M1_CDNS_524688791851016  L1M1_CDNS_524688791851016_11
timestamp 1704896540
transform 1 0 3907 0 -1 8342
box -12 -6 46 616
use L1M1_CDNS_524688791851017  L1M1_CDNS_524688791851017_0
timestamp 1704896540
transform 1 0 2173 0 1 8658
box -12 -6 1918 40
use L1M1_CDNS_524688791851018  L1M1_CDNS_524688791851018_0
timestamp 1704896540
transform 1 0 3139 0 1 7732
box -12 -6 46 832
use L1M1_CDNS_524688791851018  L1M1_CDNS_524688791851018_1
timestamp 1704896540
transform 1 0 2627 0 1 7732
box -12 -6 46 832
use L1M1_CDNS_524688791851018  L1M1_CDNS_524688791851018_2
timestamp 1704896540
transform 1 0 3651 0 1 7732
box -12 -6 46 832
use L1M1_CDNS_524688791851042  L1M1_CDNS_524688791851042_0
timestamp 1704896540
transform -1 0 1391 0 1 10872
box -12 -6 1342 40
use L1M1_CDNS_524688791851044  L1M1_CDNS_524688791851044_0
timestamp 1704896540
transform 1 0 4093 0 -1 7230
box -12 -6 46 5008
use L1M1_CDNS_524688791851053  L1M1_CDNS_524688791851053_0
timestamp 1704896540
transform 1 0 1779 0 1 8743
box -12 -6 6454 40
use L1M1_CDNS_524688791851053  L1M1_CDNS_524688791851053_1
timestamp 1704896540
transform 1 0 1779 0 1 10689
box -12 -6 6454 40
use L1M1_CDNS_524688791851054  L1M1_CDNS_524688791851054_0
timestamp 1704896540
transform 1 0 3687 0 -1 1930
box -12 -6 46 1408
use L1M1_CDNS_524688791851054  L1M1_CDNS_524688791851054_1
timestamp 1704896540
transform 1 0 2775 0 -1 1930
box -12 -6 46 1408
use L1M1_CDNS_524688791851054  L1M1_CDNS_524688791851054_2
timestamp 1704896540
transform 1 0 1863 0 -1 1930
box -12 -6 46 1408
use L1M1_CDNS_524688791851054  L1M1_CDNS_524688791851054_3
timestamp 1704896540
transform 1 0 3943 0 -1 1930
box -12 -6 46 1408
use L1M1_CDNS_524688791851054  L1M1_CDNS_524688791851054_4
timestamp 1704896540
transform 1 0 1457 0 -1 1930
box -12 -6 46 1408
use L1M1_CDNS_524688791851055  L1M1_CDNS_524688791851055_0
timestamp 1704896540
transform 1 0 2319 0 -1 1930
box -12 -6 46 1120
use L1M1_CDNS_524688791851055  L1M1_CDNS_524688791851055_1
timestamp 1704896540
transform 1 0 3231 0 -1 1930
box -12 -6 46 1120
use L1M1_CDNS_524688791851055  L1M1_CDNS_524688791851055_2
timestamp 1704896540
transform 1 0 1607 0 -1 1930
box -12 -6 46 1120
use L1M1_CDNS_524688791851056  L1M1_CDNS_524688791851056_0
timestamp 1704896540
transform 1 0 198 0 1 526
box -12 -6 46 10120
use L1M1_CDNS_524688791851057  L1M1_CDNS_524688791851057_0
timestamp 1704896540
transform 1 0 1078 0 -1 6715
box 0 0 1 1
use L1M1_CDNS_524688791851057  L1M1_CDNS_524688791851057_1
timestamp 1704896540
transform 1 0 1457 0 1 10490
box 0 0 1 1
use L1M1_CDNS_524688791851058  L1M1_CDNS_524688791851058_0
timestamp 1704896540
transform 1 0 1078 0 -1 6203
box -12 -6 46 5584
use L1M1_CDNS_524688791851059  L1M1_CDNS_524688791851059_0
timestamp 1704896540
transform 1 0 3904 0 -1 7077
box -12 -6 46 3568
use L1M1_CDNS_524688791851059  L1M1_CDNS_524688791851059_1
timestamp 1704896540
transform 1 0 1078 0 1 6979
box -12 -6 46 3568
use L1M1_CDNS_524688791851060  L1M1_CDNS_524688791851060_0
timestamp 1704896540
transform 1 0 1646 0 -1 8551
box -12 -6 46 1048
use L1M1_CDNS_524688791851061  L1M1_CDNS_524688791851061_0
timestamp 1704896540
transform -1 0 7985 0 1 10572
box -12 -6 6094 40
use L1M1_CDNS_524688791851061  L1M1_CDNS_524688791851061_1
timestamp 1704896540
transform -1 0 7985 0 1 9716
box -12 -6 6094 40
use L1M1_CDNS_524688791851061  L1M1_CDNS_524688791851061_2
timestamp 1704896540
transform -1 0 7985 0 1 8860
box -12 -6 6094 40
use L1M1_CDNS_524688791851062  L1M1_CDNS_524688791851062_0
timestamp 1704896540
transform -1 0 1840 0 -1 10418
box 0 0 1 1
use L1M1_CDNS_524688791851062  L1M1_CDNS_524688791851062_1
timestamp 1704896540
transform 1 0 8112 0 -1 9514
box 0 0 1 1
use L1M1_CDNS_524688791851062  L1M1_CDNS_524688791851062_2
timestamp 1704896540
transform 1 0 6023 0 -1 10418
box 0 0 1 1
use L1M1_CDNS_524688791851062  L1M1_CDNS_524688791851062_3
timestamp 1704896540
transform 1 0 3893 0 -1 10418
box 0 0 1 1
use L1M1_CDNS_524688791851062  L1M1_CDNS_524688791851062_4
timestamp 1704896540
transform 1 0 8112 0 -1 10418
box 0 0 1 1
use L1M1_CDNS_524688791851062  L1M1_CDNS_524688791851062_5
timestamp 1704896540
transform 1 0 6023 0 -1 9514
box 0 0 1 1
use L1M1_CDNS_524688791851063  L1M1_CDNS_524688791851063_0
timestamp 1704896540
transform 1 0 8226 0 -1 10624
box -12 -6 46 1768
use L1M1_CDNS_524688791851064  L1M1_CDNS_524688791851064_0
timestamp 1704896540
transform 1 0 1646 0 -1 7083
box -12 -6 46 688
use L1M1_CDNS_524688791851065  L1M1_CDNS_524688791851065_0
timestamp 1704896540
transform 1 0 1646 0 1 2291
box -12 -6 46 3928
use L1M1_CDNS_524688791851066  L1M1_CDNS_524688791851066_0
timestamp 1704896540
transform 0 -1 1776 1 0 2363
box -12 -6 3862 40
use L1M1_CDNS_524688791851067  L1M1_CDNS_524688791851067_0
timestamp 1704896540
transform 1 0 8415 0 -1 10831
box -12 -6 46 2056
use L1M1_CDNS_524688791851068  L1M1_CDNS_524688791851068_0
timestamp 1704896540
transform 1 0 9 0 1 328
box -12 -6 46 10408
use L1M1_CDNS_524688791851069  L1M1_CDNS_524688791851069_0
timestamp 1704896540
transform 1 0 1457 0 -1 6243
box -12 -6 46 4144
use L1M1_CDNS_524688791851070  L1M1_CDNS_524688791851070_0
timestamp 1704896540
transform 0 1 3805 -1 0 7008
box -12 -6 3502 40
use L1M1_CDNS_524688791851071  L1M1_CDNS_524688791851071_0
timestamp 1704896540
transform 1 0 1457 0 1 7245
box -12 -6 46 1264
use L1M1_CDNS_524688791851072  L1M1_CDNS_524688791851072_0
timestamp 1704896540
transform -1 0 1807 0 1 8988
box 0 0 1 1
use L1M1_CDNS_524688791851073  L1M1_CDNS_524688791851073_0
timestamp 1704896540
transform -1 0 8376 0 -1 10906
box -12 -6 6886 40
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1704896540
transform 0 -1 2721 -1 0 5915
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_1
timestamp 1704896540
transform 0 -1 2721 -1 0 3531
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_2
timestamp 1704896540
transform 0 -1 1392 -1 0 2034
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_3
timestamp 1704896540
transform 0 -1 1204 -1 0 2034
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_4
timestamp 1704896540
transform -1 0 1677 0 1 7275
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_5
timestamp 1704896540
transform -1 0 1121 0 1 10681
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_6
timestamp 1704896540
transform -1 0 1121 0 1 423
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_7
timestamp 1704896540
transform -1 0 2856 0 -1 2304
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_8
timestamp 1704896540
transform 0 1 2669 1 0 7386
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_9
timestamp 1704896540
transform 0 1 2863 1 0 7386
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_10
timestamp 1704896540
transform 0 1 2971 1 0 4525
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_11
timestamp 1704896540
transform 0 1 2971 1 0 6909
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_12
timestamp 1704896540
transform 0 1 2863 1 0 5717
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_13
timestamp 1704896540
transform 0 1 2863 1 0 3333
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_14
timestamp 1704896540
transform 0 1 3517 1 0 7386
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_15
timestamp 1704896540
transform 0 1 2015 1 0 7386
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_16
timestamp 1704896540
transform 0 1 2669 1 0 5468
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_17
timestamp 1704896540
transform 0 1 2453 1 0 5468
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_18
timestamp 1704896540
transform 0 1 2669 1 0 3652
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_19
timestamp 1704896540
transform 0 1 2453 1 0 3652
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_20
timestamp 1704896540
transform 0 -1 1204 1 0 10699
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_21
timestamp 1704896540
transform 0 -1 3569 1 0 2297
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_22
timestamp 1704896540
transform 0 -1 3569 1 0 1808
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_23
timestamp 1704896540
transform 0 -1 2067 1 0 2297
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_24
timestamp 1704896540
transform 0 -1 2067 1 0 1808
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_25
timestamp 1704896540
transform 0 -1 2613 1 0 6909
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_26
timestamp 1704896540
transform 0 -1 2613 1 0 4525
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_27
timestamp 1704896540
transform 0 -1 2915 1 0 5468
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_28
timestamp 1704896540
transform 0 -1 3131 1 0 5468
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_29
timestamp 1704896540
transform 0 -1 3131 1 0 3652
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_30
timestamp 1704896540
transform 0 -1 2915 1 0 3652
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_31
timestamp 1704896540
transform 1 0 1549 0 -1 10911
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_32
timestamp 1704896540
transform 1 0 3907 0 1 7275
box 0 0 1 1
use M1M2_CDNS_52468879185200  M1M2_CDNS_52468879185200_0
timestamp 1704896540
transform 0 1 3648 1 0 7386
box 0 0 1 1
use M1M2_CDNS_52468879185200  M1M2_CDNS_52468879185200_1
timestamp 1704896540
transform 0 1 1756 1 0 7386
box 0 0 1 1
use M1M2_CDNS_52468879185200  M1M2_CDNS_52468879185200_2
timestamp 1704896540
transform 0 1 3924 1 0 7386
box 0 0 1 1
use M1M2_CDNS_52468879185200  M1M2_CDNS_52468879185200_3
timestamp 1704896540
transform 1 0 7816 0 1 8740
box 0 0 1 1
use M1M2_CDNS_52468879185200  M1M2_CDNS_52468879185200_4
timestamp 1704896540
transform 1 0 7816 0 1 10546
box 0 0 1 1
use M1M2_CDNS_52468879185200  M1M2_CDNS_52468879185200_5
timestamp 1704896540
transform 1 0 7816 0 1 9643
box 0 0 1 1
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_0
timestamp 1704896540
transform 0 -1 1501 -1 0 10887
box 0 0 1 1
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_1
timestamp 1704896540
transform -1 0 8071 0 1 11020
box 0 0 1 1
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_2
timestamp 1704896540
transform 0 -1 1284 1 0 6430
box 0 0 1 1
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_3
timestamp 1704896540
transform 1 0 4790 0 1 11100
box 0 0 1 1
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_4
timestamp 1704896540
transform 1 0 4790 0 1 10940
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_0
timestamp 1704896540
transform 0 -1 1204 -1 0 8844
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_1
timestamp 1704896540
transform 0 -1 1204 -1 0 8624
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_2
timestamp 1704896540
transform 0 -1 1284 -1 0 6237
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_3
timestamp 1704896540
transform 0 -1 1284 -1 0 10610
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_4
timestamp 1704896540
transform 0 1 3517 -1 0 9829
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_5
timestamp 1704896540
transform 0 1 4651 -1 0 10732
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_6
timestamp 1704896540
transform 0 1 4651 -1 0 9829
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_7
timestamp 1704896540
transform 0 1 4651 -1 0 8926
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_8
timestamp 1704896540
transform 0 1 3517 -1 0 8926
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_9
timestamp 1704896540
transform 0 1 2015 -1 0 8926
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_10
timestamp 1704896540
transform 0 1 2015 -1 0 9829
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_11
timestamp 1704896540
transform 0 1 3517 -1 0 10732
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_12
timestamp 1704896540
transform 0 1 2015 -1 0 10732
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_13
timestamp 1704896540
transform 0 -1 1501 1 0 8734
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_14
timestamp 1704896540
transform 0 -1 1501 1 0 9637
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_15
timestamp 1704896540
transform 0 -1 1284 1 0 557
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_16
timestamp 1704896540
transform 0 -1 1284 1 0 6936
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_17
timestamp 1704896540
transform 1 0 2696 0 1 11100
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_18
timestamp 1704896540
transform 1 0 2696 0 1 10940
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_19
timestamp 1704896540
transform 1 0 5467 0 1 10786
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_20
timestamp 1704896540
transform 1 0 2971 0 1 10786
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_21
timestamp 1704896540
transform 1 0 4511 0 1 10786
box 0 0 1 1
use M1M2_CDNS_52468879185204  M1M2_CDNS_52468879185204_0
timestamp 1704896540
transform 0 1 1340 1 0 6824
box 0 0 1 1
use M1M2_CDNS_52468879185208  M1M2_CDNS_52468879185208_0
timestamp 1704896540
transform 0 1 5306 -1 0 10732
box 0 0 192 244
use M1M2_CDNS_52468879185208  M1M2_CDNS_52468879185208_1
timestamp 1704896540
transform 0 1 5306 -1 0 9829
box 0 0 192 244
use M1M2_CDNS_52468879185208  M1M2_CDNS_52468879185208_2
timestamp 1704896540
transform 0 1 2670 -1 0 9829
box 0 0 192 244
use M1M2_CDNS_52468879185208  M1M2_CDNS_52468879185208_3
timestamp 1704896540
transform 0 1 2670 -1 0 10732
box 0 0 192 244
use M1M2_CDNS_52468879185297  M1M2_CDNS_52468879185297_0
timestamp 1704896540
transform 0 -1 1121 -1 0 6718
box 0 0 1 1
use M1M2_CDNS_52468879185297  M1M2_CDNS_52468879185297_1
timestamp 1704896540
transform 1 0 8132 0 -1 10911
box 0 0 1 1
use M1M2_CDNS_52468879185297  M1M2_CDNS_52468879185297_2
timestamp 1704896540
transform 1 0 7161 0 1 11100
box 0 0 1 1
use M1M2_CDNS_52468879185297  M1M2_CDNS_52468879185297_3
timestamp 1704896540
transform 1 0 7161 0 1 10940
box 0 0 1 1
use M1M2_CDNS_52468879185299  M1M2_CDNS_52468879185299_0
timestamp 1704896540
transform 0 -1 1500 -1 0 7107
box 0 0 704 52
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_0
timestamp 1704896540
transform 0 -1 2641 1 0 7144
box 0 0 1 1
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_0
timestamp 1704896540
transform 0 1 4392 -1 0 10732
box 0 0 192 180
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_1
timestamp 1704896540
transform 0 1 3648 -1 0 9829
box 0 0 192 180
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_2
timestamp 1704896540
transform 0 1 1756 -1 0 9829
box 0 0 192 180
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_3
timestamp 1704896540
transform 0 1 4392 -1 0 9829
box 0 0 192 180
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_4
timestamp 1704896540
transform 0 1 3648 -1 0 10732
box 0 0 192 180
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_5
timestamp 1704896540
transform 0 1 1756 -1 0 10732
box 0 0 192 180
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_6
timestamp 1704896540
transform 1 0 5342 0 1 8740
box 0 0 192 180
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_7
timestamp 1704896540
transform 1 0 4386 0 1 8740
box 0 0 192 180
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_8
timestamp 1704896540
transform 1 0 6278 0 1 8740
box 0 0 192 180
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_9
timestamp 1704896540
transform 1 0 6562 0 1 8740
box 0 0 192 180
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_10
timestamp 1704896540
transform 1 0 6278 0 1 9643
box 0 0 192 180
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_11
timestamp 1704896540
transform 1 0 6562 0 1 9643
box 0 0 192 180
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_12
timestamp 1704896540
transform 1 0 4110 0 1 8740
box 0 0 192 180
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_13
timestamp 1704896540
transform 1 0 6562 0 1 10546
box 0 0 192 180
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_14
timestamp 1704896540
transform 1 0 1750 0 1 8740
box 0 0 192 180
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_15
timestamp 1704896540
transform 1 0 2696 0 1 8740
box 0 0 192 180
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_16
timestamp 1704896540
transform 1 0 3642 0 1 8740
box 0 0 192 180
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_17
timestamp 1704896540
transform 1 0 3918 0 1 8740
box 0 0 192 180
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_18
timestamp 1704896540
transform 1 0 6278 0 1 10546
box 0 0 192 180
use M1M2_CDNS_524688791851020  M1M2_CDNS_524688791851020_0
timestamp 1704896540
transform 0 -1 8272 1 0 8734
box 0 0 1984 52
use M1M2_CDNS_524688791851022  M1M2_CDNS_524688791851022_0
timestamp 1704896540
transform 0 1 1448 1 0 7239
box 0 0 1280 52
use M1M2_CDNS_524688791851031  M1M2_CDNS_524688791851031_0
timestamp 1704896540
transform 0 1 3084 1 0 7386
box 0 0 128 372
use M1M2_CDNS_524688791851031  M1M2_CDNS_524688791851031_1
timestamp 1704896540
transform 0 1 2128 1 0 7386
box 0 0 128 372
use M1M2_CDNS_524688791851032  M1M2_CDNS_524688791851032_0
timestamp 1704896540
transform 0 1 4764 -1 0 10732
box 0 0 192 372
use M1M2_CDNS_524688791851032  M1M2_CDNS_524688791851032_1
timestamp 1704896540
transform 0 1 5720 -1 0 10732
box 0 0 192 372
use M1M2_CDNS_524688791851032  M1M2_CDNS_524688791851032_2
timestamp 1704896540
transform 0 1 3924 -1 0 10732
box 0 0 192 372
use M1M2_CDNS_524688791851032  M1M2_CDNS_524688791851032_3
timestamp 1704896540
transform 0 1 3924 -1 0 9829
box 0 0 192 372
use M1M2_CDNS_524688791851032  M1M2_CDNS_524688791851032_4
timestamp 1704896540
transform 0 1 4764 -1 0 9829
box 0 0 192 372
use M1M2_CDNS_524688791851032  M1M2_CDNS_524688791851032_5
timestamp 1704896540
transform 0 1 2128 -1 0 9829
box 0 0 192 372
use M1M2_CDNS_524688791851032  M1M2_CDNS_524688791851032_6
timestamp 1704896540
transform 0 1 3084 -1 0 9829
box 0 0 192 372
use M1M2_CDNS_524688791851032  M1M2_CDNS_524688791851032_7
timestamp 1704896540
transform 0 1 5720 -1 0 9829
box 0 0 192 372
use M1M2_CDNS_524688791851032  M1M2_CDNS_524688791851032_8
timestamp 1704896540
transform 0 1 2128 -1 0 10732
box 0 0 192 372
use M1M2_CDNS_524688791851032  M1M2_CDNS_524688791851032_9
timestamp 1704896540
transform 0 1 3084 -1 0 10732
box 0 0 192 372
use M1M2_CDNS_524688791851033  M1M2_CDNS_524688791851033_0
timestamp 1704896540
transform 0 -1 3851 1 0 2348
box 0 0 4672 52
use M1M2_CDNS_524688791851035  M1M2_CDNS_524688791851035_0
timestamp 1704896540
transform 0 -1 4136 -1 0 7276
box 0 0 5056 52
use M1M2_CDNS_524688791851074  M1M2_CDNS_524688791851074_0
timestamp 1704896540
transform 0 1 189 -1 0 10640
box 0 0 10112 52
use M1M2_CDNS_524688791851075  M1M2_CDNS_524688791851075_0
timestamp 1704896540
transform 0 1 1069 -1 0 6198
box 0 0 5568 52
use M1M2_CDNS_524688791851076  M1M2_CDNS_524688791851076_0
timestamp 1704896540
transform 0 1 1069 1 0 7000
box 0 0 3520 52
use M1M2_CDNS_524688791851077  M1M2_CDNS_524688791851077_0
timestamp 1704896540
transform 1 0 5746 0 1 8740
box 0 0 320 180
use M1M2_CDNS_524688791851077  M1M2_CDNS_524688791851077_1
timestamp 1704896540
transform 1 0 4790 0 1 8740
box 0 0 320 180
use M1M2_CDNS_524688791851077  M1M2_CDNS_524688791851077_2
timestamp 1704896540
transform 1 0 2154 0 1 8740
box 0 0 320 180
use M1M2_CDNS_524688791851077  M1M2_CDNS_524688791851077_3
timestamp 1704896540
transform 1 0 3110 0 1 8740
box 0 0 320 180
use M1M2_CDNS_524688791851078  M1M2_CDNS_524688791851078_0
timestamp 1704896540
transform 0 -1 1785 -1 0 7020
box 0 0 576 52
use M1M2_CDNS_524688791851079  M1M2_CDNS_524688791851079_0
timestamp 1704896540
transform 0 -1 1785 1 0 2348
box 0 0 3840 52
use M1M2_CDNS_524688791851080  M1M2_CDNS_524688791851080_0
timestamp 1704896540
transform 0 1 8406 -1 0 10887
box 0 0 2112 116
use M1M2_CDNS_524688791851081  M1M2_CDNS_524688791851081_0
timestamp 1704896540
transform 1 0 6837 0 1 8740
box 0 0 256 180
use M1M2_CDNS_524688791851081  M1M2_CDNS_524688791851081_1
timestamp 1704896540
transform 1 0 7161 0 1 8740
box 0 0 256 180
use M1M2_CDNS_524688791851081  M1M2_CDNS_524688791851081_2
timestamp 1704896540
transform 1 0 6837 0 1 9643
box 0 0 256 180
use M1M2_CDNS_524688791851081  M1M2_CDNS_524688791851081_3
timestamp 1704896540
transform 1 0 7161 0 1 9643
box 0 0 256 180
use M1M2_CDNS_524688791851081  M1M2_CDNS_524688791851081_4
timestamp 1704896540
transform 1 0 7161 0 1 10546
box 0 0 256 180
use M1M2_CDNS_524688791851081  M1M2_CDNS_524688791851081_5
timestamp 1704896540
transform 1 0 6837 0 1 10546
box 0 0 256 180
use M1M2_CDNS_524688791851082  M1M2_CDNS_524688791851082_0
timestamp 1704896540
transform 0 -1 52 1 0 318
box 0 0 10368 52
use M1M2_CDNS_524688791851083  M1M2_CDNS_524688791851083_0
timestamp 1704896540
transform 0 1 1448 -1 0 6188
box 0 0 5760 52
use M1M2_CDNS_524688791851084  M1M2_CDNS_524688791851084_0
timestamp 1704896540
transform 1 0 399 0 1 503
box 0 0 512 52
use M1M2_CDNS_524688791851085  M1M2_CDNS_524688791851085_0
timestamp 1704896540
transform 0 1 1340 1 0 9012
box 0 0 1408 52
use nDFres_CDNS_524688791851094  nDFres_CDNS_524688791851094_0
timestamp 1704896540
transform 0 1 433 1 0 685
box -68 -26 1803 92
use nDFres_CDNS_524688791851094  nDFres_CDNS_524688791851094_1
timestamp 1704896540
transform 0 1 811 1 0 685
box -68 -26 1803 92
use nDFres_CDNS_524688791851094  nDFres_CDNS_524688791851094_2
timestamp 1704896540
transform 0 1 685 1 0 685
box -68 -26 1803 92
use nDFres_CDNS_524688791851094  nDFres_CDNS_524688791851094_3
timestamp 1704896540
transform 0 1 433 1 0 6730
box -68 -26 1803 92
use nDFres_CDNS_524688791851094  nDFres_CDNS_524688791851094_4
timestamp 1704896540
transform 0 1 559 1 0 6730
box -68 -26 1803 92
use nDFres_CDNS_524688791851094  nDFres_CDNS_524688791851094_5
timestamp 1704896540
transform 0 1 559 1 0 2700
box -68 -26 1803 92
use nDFres_CDNS_524688791851094  nDFres_CDNS_524688791851094_6
timestamp 1704896540
transform 0 1 433 1 0 2700
box -68 -26 1803 92
use nDFres_CDNS_524688791851094  nDFres_CDNS_524688791851094_7
timestamp 1704896540
transform 0 1 685 1 0 2700
box -68 -26 1803 92
use nDFres_CDNS_524688791851094  nDFres_CDNS_524688791851094_8
timestamp 1704896540
transform 0 1 811 1 0 6730
box -68 -26 1803 92
use nDFres_CDNS_524688791851094  nDFres_CDNS_524688791851094_9
timestamp 1704896540
transform 0 1 811 1 0 2700
box -68 -26 1803 92
use nDFres_CDNS_524688791851094  nDFres_CDNS_524688791851094_10
timestamp 1704896540
transform 0 1 811 1 0 8745
box -68 -26 1803 92
use nDFres_CDNS_524688791851094  nDFres_CDNS_524688791851094_11
timestamp 1704896540
transform 0 1 811 1 0 4715
box -68 -26 1803 92
use nDFres_CDNS_524688791851094  nDFres_CDNS_524688791851094_12
timestamp 1704896540
transform 0 1 685 1 0 4715
box -68 -26 1803 92
use nDFres_CDNS_524688791851094  nDFres_CDNS_524688791851094_13
timestamp 1704896540
transform 0 1 433 1 0 4715
box -68 -26 1803 92
use nDFres_CDNS_524688791851094  nDFres_CDNS_524688791851094_14
timestamp 1704896540
transform 0 1 559 1 0 4715
box -68 -26 1803 92
use nDFres_CDNS_524688791851094  nDFres_CDNS_524688791851094_15
timestamp 1704896540
transform 0 1 559 1 0 8745
box -68 -26 1803 92
use nDFres_CDNS_524688791851094  nDFres_CDNS_524688791851094_16
timestamp 1704896540
transform 0 1 433 1 0 8745
box -68 -26 1803 92
use nDFres_CDNS_524688791851094  nDFres_CDNS_524688791851094_17
timestamp 1704896540
transform 0 1 685 1 0 8745
box -68 -26 1803 92
use nDFres_CDNS_524688791851094  nDFres_CDNS_524688791851094_18
timestamp 1704896540
transform 0 1 685 1 0 6730
box -68 -26 1803 92
use nDFres_CDNS_524688791851094  nDFres_CDNS_524688791851094_19
timestamp 1704896540
transform 0 1 559 1 0 685
box -68 -26 1803 92
use nDFres_CDNS_524688791851094  nDFres_CDNS_524688791851094_20
timestamp 1704896540
transform 0 1 937 1 0 685
box -68 -26 1803 92
use nDFres_CDNS_524688791851094  nDFres_CDNS_524688791851094_21
timestamp 1704896540
transform 0 1 937 1 0 2700
box -68 -26 1803 92
use nDFres_CDNS_524688791851094  nDFres_CDNS_524688791851094_22
timestamp 1704896540
transform 0 1 937 1 0 4715
box -68 -26 1803 92
use nDFres_CDNS_524688791851094  nDFres_CDNS_524688791851094_23
timestamp 1704896540
transform 0 1 937 1 0 6730
box -68 -26 1803 92
use nDFres_CDNS_524688791851094  nDFres_CDNS_524688791851094_24
timestamp 1704896540
transform 0 1 937 1 0 8745
box -68 -26 1803 92
use nDFres_CDNS_524688791851094  nDFres_CDNS_524688791851094_25
timestamp 1704896540
transform 0 -1 373 1 0 685
box -68 -26 1803 92
use nDFres_CDNS_524688791851094  nDFres_CDNS_524688791851094_26
timestamp 1704896540
transform 0 -1 373 1 0 2700
box -68 -26 1803 92
use nDFres_CDNS_524688791851094  nDFres_CDNS_524688791851094_27
timestamp 1704896540
transform 0 -1 373 1 0 4715
box -68 -26 1803 92
use nDFres_CDNS_524688791851094  nDFres_CDNS_524688791851094_28
timestamp 1704896540
transform 0 -1 373 1 0 6730
box -68 -26 1803 92
use nDFres_CDNS_524688791851094  nDFres_CDNS_524688791851094_29
timestamp 1704896540
transform 0 -1 373 1 0 8745
box -68 -26 1803 92
use nfet_CDNS_524688791851024  nfet_CDNS_524688791851024_0
timestamp 1704896540
transform 1 0 2160 0 1 7610
box -79 -52 535 1052
use nfet_CDNS_524688791851024  nfet_CDNS_524688791851024_1
timestamp 1704896540
transform 1 0 2672 0 1 7610
box -79 -52 535 1052
use nfet_CDNS_524688791851024  nfet_CDNS_524688791851024_2
timestamp 1704896540
transform 1 0 3184 0 1 7610
box -79 -52 535 1052
use nfet_CDNS_524688791851024  nfet_CDNS_524688791851024_3
timestamp 1704896540
transform 1 0 3696 0 1 7610
box -79 -52 535 1052
use nfet_CDNS_524688791851046  nfet_CDNS_524688791851046_0
timestamp 1704896540
transform -1 0 2764 0 1 2367
box -79 -52 879 1052
use nfet_CDNS_524688791851046  nfet_CDNS_524688791851046_1
timestamp 1704896540
transform -1 0 3620 0 1 2367
box -79 -52 879 1052
use nfet_CDNS_524688791851046  nfet_CDNS_524688791851046_2
timestamp 1704896540
transform -1 0 3620 0 1 4751
box -79 -52 879 1052
use nfet_CDNS_524688791851046  nfet_CDNS_524688791851046_3
timestamp 1704896540
transform -1 0 2764 0 1 4751
box -79 -52 879 1052
use nfet_CDNS_524688791851046  nfet_CDNS_524688791851046_4
timestamp 1704896540
transform 1 0 1964 0 1 3559
box -79 -52 879 1052
use nfet_CDNS_524688791851046  nfet_CDNS_524688791851046_5
timestamp 1704896540
transform 1 0 1964 0 1 5943
box -79 -52 879 1052
use nfet_CDNS_524688791851046  nfet_CDNS_524688791851046_6
timestamp 1704896540
transform 1 0 2820 0 1 3559
box -79 -52 879 1052
use nfet_CDNS_524688791851046  nfet_CDNS_524688791851046_7
timestamp 1704896540
transform 1 0 2820 0 1 5943
box -79 -52 879 1052
use nfet_CDNS_524688791851047  nfet_CDNS_524688791851047_0
timestamp 1704896540
transform -1 0 3776 0 1 4751
box -79 -52 182 1052
use nfet_CDNS_524688791851047  nfet_CDNS_524688791851047_1
timestamp 1704896540
transform -1 0 3776 0 1 3559
box -79 -52 182 1052
use nfet_CDNS_524688791851047  nfet_CDNS_524688791851047_2
timestamp 1704896540
transform -1 0 3776 0 1 2367
box -79 -52 182 1052
use nfet_CDNS_524688791851047  nfet_CDNS_524688791851047_3
timestamp 1704896540
transform -1 0 3776 0 1 5943
box -79 -52 182 1052
use nfet_CDNS_524688791851047  nfet_CDNS_524688791851047_4
timestamp 1704896540
transform 1 0 1808 0 1 5943
box -79 -52 182 1052
use nfet_CDNS_524688791851047  nfet_CDNS_524688791851047_5
timestamp 1704896540
transform 1 0 1808 0 1 4751
box -79 -52 182 1052
use nfet_CDNS_524688791851047  nfet_CDNS_524688791851047_6
timestamp 1704896540
transform 1 0 1808 0 1 3559
box -79 -52 182 1052
use nfet_CDNS_524688791851047  nfet_CDNS_524688791851047_7
timestamp 1704896540
transform 1 0 1808 0 1 2367
box -79 -52 182 1052
use nfet_CDNS_524688791851090  nfet_CDNS_524688791851090_0
timestamp 1704896540
transform 0 -1 3845 1 0 8905
box -79 -26 879 2026
use nfet_CDNS_524688791851090  nfet_CDNS_524688791851090_1
timestamp 1704896540
transform 0 -1 8105 1 0 8905
box -79 -26 879 2026
use nfet_CDNS_524688791851090  nfet_CDNS_524688791851090_2
timestamp 1704896540
transform 0 -1 8105 1 0 9761
box -79 -26 879 2026
use nfet_CDNS_524688791851090  nfet_CDNS_524688791851090_3
timestamp 1704896540
transform 0 -1 5975 1 0 8905
box -79 -26 879 2026
use nfet_CDNS_524688791851090  nfet_CDNS_524688791851090_4
timestamp 1704896540
transform 0 -1 5975 1 0 9761
box -79 -26 879 2026
use nfet_CDNS_524688791851090  nfet_CDNS_524688791851090_5
timestamp 1704896540
transform 0 -1 3845 1 0 9761
box -79 -26 879 2026
use nfet_CDNS_524688791851091  nfet_CDNS_524688791851091_0
timestamp 1704896540
transform -1 0 1928 0 1 7610
box -79 -52 199 1052
use nfet_CDNS_524688791851091  nfet_CDNS_524688791851091_1
timestamp 1704896540
transform -1 0 4328 0 1 7610
box -79 -52 199 1052
use nfet_CDNS_524688791851091  nfet_CDNS_524688791851091_2
timestamp 1704896540
transform 1 0 1984 0 1 7610
box -79 -52 199 1052
use pfet_CDNS_524688791851092  pfet_CDNS_524688791851092_0
timestamp 1704896540
transform 1 0 2364 0 1 536
box -119 -66 519 1466
use pfet_CDNS_524688791851092  pfet_CDNS_524688791851092_1
timestamp 1704896540
transform 1 0 3276 0 1 536
box -119 -66 519 1466
use pfet_CDNS_524688791851092  pfet_CDNS_524688791851092_2
timestamp 1704896540
transform 1 0 1908 0 1 536
box -119 -66 519 1466
use pfet_CDNS_524688791851092  pfet_CDNS_524688791851092_3
timestamp 1704896540
transform 1 0 2820 0 1 536
box -119 -66 519 1466
use pfet_CDNS_524688791851093  pfet_CDNS_524688791851093_0
timestamp 1704896540
transform -1 0 1852 0 1 536
box -119 -66 319 1466
use pfet_CDNS_524688791851093  pfet_CDNS_524688791851093_1
timestamp 1704896540
transform 1 0 3732 0 1 536
box -119 -66 319 1466
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_0
timestamp 1704896540
transform 0 1 4235 -1 0 8708
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_0
timestamp 1704896540
transform -1 0 3932 0 -1 2034
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_1
timestamp 1704896540
transform 1 0 3676 0 -1 3465
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_2
timestamp 1704896540
transform 1 0 3676 0 -1 7041
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_3
timestamp 1704896540
transform 1 0 3676 0 -1 4657
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_4
timestamp 1704896540
transform 1 0 1774 0 -1 3465
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_5
timestamp 1704896540
transform 1 0 3676 0 -1 5849
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_6
timestamp 1704896540
transform 1 0 1774 0 -1 4657
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_7
timestamp 1704896540
transform 1 0 1774 0 -1 5849
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_8
timestamp 1704896540
transform 1 0 1774 0 -1 7041
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_9
timestamp 1704896540
transform 1 0 1652 0 -1 2034
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_0
timestamp 1704896540
transform 0 1 1808 1 0 8642
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_1
timestamp 1704896540
transform 0 -1 2327 1 0 8642
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_2
timestamp 1704896540
transform 0 -1 4119 1 0 8642
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_3
timestamp 1704896540
transform 0 -1 3863 1 0 8642
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_4
timestamp 1704896540
transform 0 -1 3607 1 0 8642
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_5
timestamp 1704896540
transform 0 -1 3351 1 0 8642
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_6
timestamp 1704896540
transform 0 -1 3095 1 0 8642
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_7
timestamp 1704896540
transform 0 -1 2839 1 0 8642
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_8
timestamp 1704896540
transform 0 -1 2583 1 0 8642
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_9
timestamp 1704896540
transform 0 -1 2104 1 0 8642
box 0 0 1 1
use PYL1_CDNS_52468879185317  PYL1_CDNS_52468879185317_0
timestamp 1704896540
transform -1 0 1823 0 1 9788
box 0 0 66 746
use PYL1_CDNS_52468879185317  PYL1_CDNS_52468879185317_1
timestamp 1704896540
transform -1 0 1823 0 1 8932
box 0 0 66 746
use PYL1_CDNS_52468879185317  PYL1_CDNS_52468879185317_2
timestamp 1704896540
transform -1 0 6073 0 1 8932
box 0 0 66 746
use PYL1_CDNS_52468879185317  PYL1_CDNS_52468879185317_3
timestamp 1704896540
transform -1 0 6073 0 1 9788
box 0 0 66 746
use PYL1_CDNS_52468879185317  PYL1_CDNS_52468879185317_4
timestamp 1704896540
transform -1 0 3943 0 1 9788
box 0 0 66 746
use PYL1_CDNS_52468879185317  PYL1_CDNS_52468879185317_5
timestamp 1704896540
transform 1 0 8127 0 1 8932
box 0 0 66 746
use PYL1_CDNS_52468879185317  PYL1_CDNS_52468879185317_6
timestamp 1704896540
transform 1 0 8127 0 1 9788
box 0 0 66 746
use PYL1_CDNS_52468879185447  PYL1_CDNS_52468879185447_0
timestamp 1704896540
transform 1 0 1939 0 -1 2034
box 0 0 1 1
use PYL1_CDNS_52468879185447  PYL1_CDNS_52468879185447_1
timestamp 1704896540
transform 1 0 2395 0 -1 2034
box 0 0 1 1
use PYL1_CDNS_52468879185447  PYL1_CDNS_52468879185447_2
timestamp 1704896540
transform 1 0 2851 0 -1 2034
box 0 0 1 1
use PYL1_CDNS_52468879185447  PYL1_CDNS_52468879185447_3
timestamp 1704896540
transform 1 0 3307 0 -1 2034
box 0 0 1 1
use PYL1_CDNS_524688791851028  PYL1_CDNS_524688791851028_0
timestamp 1704896540
transform 1 0 2847 0 -1 7041
box 0 0 746 66
use PYL1_CDNS_524688791851028  PYL1_CDNS_524688791851028_1
timestamp 1704896540
transform 1 0 1991 0 -1 7041
box 0 0 746 66
use PYL1_CDNS_524688791851028  PYL1_CDNS_524688791851028_2
timestamp 1704896540
transform 1 0 2847 0 -1 5849
box 0 0 746 66
use PYL1_CDNS_524688791851028  PYL1_CDNS_524688791851028_3
timestamp 1704896540
transform 1 0 1991 0 -1 5849
box 0 0 746 66
use PYL1_CDNS_524688791851028  PYL1_CDNS_524688791851028_4
timestamp 1704896540
transform 1 0 2847 0 -1 4657
box 0 0 746 66
use PYL1_CDNS_524688791851028  PYL1_CDNS_524688791851028_5
timestamp 1704896540
transform 1 0 1991 0 -1 4657
box 0 0 746 66
use PYL1_CDNS_524688791851028  PYL1_CDNS_524688791851028_6
timestamp 1704896540
transform 1 0 2847 0 -1 3465
box 0 0 746 66
use PYL1_CDNS_524688791851028  PYL1_CDNS_524688791851028_7
timestamp 1704896540
transform 1 0 1991 0 -1 3465
box 0 0 746 66
use sky130_fd_io__tk_em1o_CDNS_52468879185315  sky130_fd_io__tk_em1o_CDNS_52468879185315_0
timestamp 1704896540
transform 0 1 1563 -1 0 9041
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_0
timestamp 1704896540
transform 0 -1 2231 -1 0 2158
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_1
timestamp 1704896540
transform 0 -1 3143 -1 0 2158
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_2
timestamp 1704896540
transform 0 -1 2417 -1 0 7772
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_3
timestamp 1704896540
transform 0 -1 3441 -1 0 7772
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_4
timestamp 1704896540
transform 0 -1 3953 -1 0 7772
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_524688791851088  sky130_fd_io__tk_em1o_CDNS_524688791851088_0
timestamp 1704896540
transform 1 0 1363 0 -1 9551
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_524688791851089  sky130_fd_io__tk_em1o_CDNS_524688791851089_0
timestamp 1704896540
transform 1 0 1363 0 -1 10428
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185314  sky130_fd_io__tk_em1s_CDNS_52468879185314_0
timestamp 1704896540
transform 0 1 1563 -1 0 9944
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185314  sky130_fd_io__tk_em1s_CDNS_52468879185314_1
timestamp 1704896540
transform 0 1 1563 1 0 9522
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185978  sky130_fd_io__tk_em1s_CDNS_52468879185978_0
timestamp 1704896540
transform 0 -1 873 -1 0 6662
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185978  sky130_fd_io__tk_em1s_CDNS_52468879185978_1
timestamp 1704896540
transform 1 0 2045 0 -1 2030
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185978  sky130_fd_io__tk_em1s_CDNS_52468879185978_2
timestamp 1704896540
transform 1 0 2957 0 -1 2030
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_524688791851086  sky130_fd_io__tk_em1s_CDNS_524688791851086_0
timestamp 1704896540
transform 1 0 1363 0 -1 9182
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_524688791851087  sky130_fd_io__tk_em1s_CDNS_524688791851087_0
timestamp 1704896540
transform -1 0 2352 0 -1 8568
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_524688791851087  sky130_fd_io__tk_em1s_CDNS_524688791851087_1
timestamp 1704896540
transform 1 0 3963 0 -1 8568
box 0 0 1 1
<< labels >>
flabel comment s 1953 7140 1953 7140 0 FreeSans 1000 0 0 0 condiode
flabel comment s 8513 11047 8513 11047 3 FreeSans 200 180 0 0 voutref
flabel comment s 15 11048 15 11048 3 FreeSans 200 0 0 0 voutref
flabel comment s 8044 8792 8044 8792 3 FreeSans 200 90 0 0 voutref
flabel metal1 s 4128 2146 4154 2192 3 FreeSans 200 180 0 0 ibuf_sel_h_n
port 2 nsew
flabel metal1 s -3 10781 77 10827 3 FreeSans 200 0 0 0 ngate
port 4 nsew
flabel metal1 s 1396 7144 1417 7208 3 FreeSans 200 180 0 0 out
port 3 nsew
flabel metal1 s -3 10940 27 10992 3 FreeSans 200 0 0 0 vgnd
port 5 nsew
flabel metal1 s -3 11100 27 11152 3 FreeSans 200 0 0 0 vgnd
port 5 nsew
flabel metal1 s 8490 11100 8522 11152 3 FreeSans 200 180 0 0 vgnd
port 5 nsew
flabel metal1 s 8490 10940 8522 10992 3 FreeSans 200 180 0 0 vgnd
port 5 nsew
flabel metal2 s 189 226 317 247 3 FreeSans 200 90 0 0 vgnd
port 5 nsew
flabel metal2 s 3517 400 3851 421 3 FreeSans 200 90 0 0 vgnd
port 5 nsew
flabel metal2 s 3079 400 3461 421 3 FreeSans 200 90 0 0 vgnd
port 5 nsew
flabel metal2 s 2669 400 2915 421 3 FreeSans 200 90 0 0 vgnd
port 5 nsew
flabel metal2 s 373 226 937 247 3 FreeSans 200 90 0 0 vgnd
port 5 nsew
flabel metal2 s 8325 8734 8522 8756 3 FreeSans 200 90 0 0 vcc
port 6 nsew
flabel metal2 s 4015 400 4136 421 3 FreeSans 200 90 0 0 vcc
port 6 nsew
flabel metal2 s 1780 400 2009 421 3 FreeSans 200 90 0 0 vcc
port 6 nsew
flabel metal2 s 993 226 1121 247 3 FreeSans 200 90 0 0 vgnd
port 5 nsew
flabel metal2 s 0 226 133 247 3 FreeSans 200 90 0 0 vcc
port 6 nsew
flabel metal2 s 2971 400 3023 421 3 FreeSans 200 90 0 0 inp
port 7 nsew
flabel metal2 s 2561 400 2613 421 3 FreeSans 200 90 0 0 inn
port 8 nsew
flabel metal2 s 2997 411 2997 411 3 FreeSans 200 90 0 0 inp
flabel metal2 s 1340 226 1392 247 3 FreeSans 200 90 0 0 en_inpop_h
port 9 nsew
<< properties >>
string GDS_END 80239638
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 80073746
string path 0.650 7.350 0.650 9.475 
<< end >>
