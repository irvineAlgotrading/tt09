VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_hvl__a21o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__a21o_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.125000 ;
    PORT
      LAYER li1 ;
        RECT 2.805 1.505 3.715 1.835 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.125000 ;
    PORT
      LAYER li1 ;
        RECT 3.895 1.505 4.195 1.835 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.125000 ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.505 2.275 1.750 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 4.320 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.100 0.215 4.280 1.415 ;
        RECT -0.130 -0.215 4.450 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 4.320 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 4.650 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 4.320 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 4.320 3.815 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.611250 ;
    PORT
      LAYER li1 ;
        RECT 0.110 1.325 0.360 3.735 ;
        RECT 0.110 0.495 0.460 1.325 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 4.320 4.155 ;
        RECT 0.540 2.280 1.440 3.755 ;
        RECT 1.620 2.100 1.870 3.755 ;
        RECT 2.320 2.450 2.650 3.755 ;
        RECT 2.830 2.630 3.780 3.755 ;
        RECT 3.960 2.450 4.210 3.735 ;
        RECT 2.320 2.280 4.210 2.450 ;
        RECT 3.960 2.195 4.210 2.280 ;
        RECT 0.565 1.930 2.625 2.100 ;
        RECT 0.565 1.725 0.895 1.930 ;
        RECT 2.455 1.325 2.625 1.930 ;
        RECT 0.640 0.365 2.250 1.325 ;
        RECT 2.430 0.495 2.680 1.325 ;
        RECT 2.860 0.365 4.170 1.325 ;
        RECT 0.000 -0.085 4.320 0.085 ;
  END
END sky130_fd_sc_hvl__a21o_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__a21oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__a21oi_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.125000 ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.505 1.915 1.750 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.125000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.505 1.315 1.750 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.125000 ;
    PORT
      LAYER li1 ;
        RECT 2.470 1.805 2.800 3.260 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 3.360 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.440 0.215 3.340 1.415 ;
        RECT -0.130 -0.215 3.490 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 3.360 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 3.690 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 3.360 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 3.360 3.815 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.832500 ;
    PORT
      LAYER li1 ;
        RECT 2.980 1.625 3.235 3.755 ;
        RECT 2.220 1.455 3.235 1.625 ;
        RECT 2.220 0.495 2.470 1.455 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 3.360 4.155 ;
        RECT 0.260 2.100 0.510 3.755 ;
        RECT 0.690 2.280 1.940 3.755 ;
        RECT 2.120 2.100 2.290 3.755 ;
        RECT 0.260 1.930 2.290 2.100 ;
        RECT 0.330 0.365 2.040 1.325 ;
        RECT 2.675 0.365 3.265 1.275 ;
        RECT 0.000 -0.085 3.360 0.085 ;
  END
END sky130_fd_sc_hvl__a21oi_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__a22o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__a22o_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.280 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.125000 ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.505 4.645 1.750 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.125000 ;
    PORT
      LAYER li1 ;
        RECT 4.825 1.505 5.155 1.750 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.125000 ;
    PORT
      LAYER li1 ;
        RECT 3.035 0.810 3.205 1.750 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.125000 ;
    PORT
      LAYER li1 ;
        RECT 1.990 1.775 2.320 3.260 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 5.280 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.020 0.215 5.235 1.415 ;
        RECT -0.130 -0.215 5.410 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 5.280 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 5.610 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 5.280 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 5.280 3.815 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.626250 ;
    PORT
      LAYER li1 ;
        RECT 0.105 0.495 0.380 3.755 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 5.280 4.155 ;
        RECT 0.560 2.175 1.460 3.755 ;
        RECT 1.640 3.635 3.530 3.805 ;
        RECT 1.640 2.175 1.810 3.635 ;
        RECT 0.585 1.595 0.915 1.755 ;
        RECT 2.500 1.595 2.830 3.455 ;
        RECT 3.280 2.100 3.530 3.635 ;
        RECT 3.710 2.280 4.660 3.755 ;
        RECT 4.840 2.100 5.170 3.735 ;
        RECT 3.280 1.930 5.170 2.100 ;
        RECT 0.585 1.425 2.855 1.595 ;
        RECT 0.550 0.365 2.260 1.245 ;
        RECT 2.685 0.630 2.855 1.425 ;
        RECT 3.385 0.630 3.635 1.325 ;
        RECT 2.685 0.460 3.635 0.630 ;
        RECT 3.815 0.365 5.125 1.325 ;
        RECT 0.000 -0.085 5.280 0.085 ;
  END
END sky130_fd_sc_hvl__a22o_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__a22oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__a22oi_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.840 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.125000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.505 2.755 1.750 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.125000 ;
    PORT
      LAYER li1 ;
        RECT 2.940 1.505 3.715 1.750 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.125000 ;
    PORT
      LAYER li1 ;
        RECT 1.465 1.505 1.795 1.750 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.125000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.505 0.835 1.835 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 3.840 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.105 0.215 3.635 1.415 ;
        RECT -0.130 -0.215 3.970 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 3.840 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 4.170 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 3.840 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 3.840 3.815 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.630000 ;
    PORT
      LAYER li1 ;
        RECT 0.925 2.175 1.285 3.455 ;
        RECT 1.085 0.980 1.285 2.175 ;
        RECT 1.705 0.980 1.955 1.325 ;
        RECT 1.085 0.810 1.955 0.980 ;
        RECT 1.705 0.495 1.955 0.810 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 3.840 4.155 ;
        RECT 0.145 3.635 1.955 3.805 ;
        RECT 0.145 2.175 0.475 3.635 ;
        RECT 1.705 2.100 1.955 3.635 ;
        RECT 2.135 2.280 3.085 3.755 ;
        RECT 3.265 2.100 3.595 3.755 ;
        RECT 1.705 1.930 3.595 2.100 ;
        RECT 0.090 0.365 0.680 1.325 ;
        RECT 2.135 0.365 3.750 1.325 ;
        RECT 0.000 -0.085 3.840 0.085 ;
  END
END sky130_fd_sc_hvl__a22oi_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__and2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__and2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.175 0.535 1.845 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER li1 ;
        RECT 1.065 0.810 1.455 1.725 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 3.360 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.030 1.085 3.340 1.415 ;
        RECT 0.020 0.215 3.340 1.085 ;
        RECT -0.130 -0.215 3.490 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 3.360 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 3.690 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 3.360 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 3.360 3.815 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.626250 ;
    PORT
      LAYER li1 ;
        RECT 2.980 0.495 3.255 3.755 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 3.360 4.155 ;
        RECT 0.090 2.255 1.020 3.705 ;
        RECT 1.200 2.075 1.370 2.675 ;
        RECT 1.550 2.255 2.800 3.755 ;
        RECT 0.715 1.905 2.775 2.075 ;
        RECT 0.715 0.995 0.885 1.905 ;
        RECT 2.445 1.725 2.775 1.905 ;
        RECT 0.130 0.825 0.885 0.995 ;
        RECT 0.130 0.495 0.380 0.825 ;
        RECT 1.635 0.365 2.625 1.325 ;
        RECT 0.000 -0.085 3.360 0.085 ;
  END
END sky130_fd_sc_hvl__and2_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__and3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__and3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.840 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER li1 ;
        RECT 0.605 0.810 0.935 1.645 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER li1 ;
        RECT 0.605 2.175 1.565 2.490 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER li1 ;
        RECT 1.115 0.810 2.255 1.645 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 3.840 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.065 0.215 3.820 1.415 ;
        RECT -0.130 -0.215 3.970 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 3.840 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 4.170 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 3.840 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 3.840 3.815 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.626250 ;
    PORT
      LAYER li1 ;
        RECT 3.365 2.175 3.715 3.755 ;
        RECT 3.410 0.495 3.715 2.175 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 3.840 4.155 ;
        RECT 0.130 1.995 0.380 3.045 ;
        RECT 0.560 2.670 1.510 3.705 ;
        RECT 1.770 1.995 2.020 3.045 ;
        RECT 2.200 2.175 3.150 3.755 ;
        RECT 0.130 1.825 3.240 1.995 ;
        RECT 0.130 0.825 0.425 1.825 ;
        RECT 2.910 1.665 3.240 1.825 ;
        RECT 2.435 0.365 3.240 1.325 ;
        RECT 0.000 -0.085 3.840 0.085 ;
  END
END sky130_fd_sc_hvl__and3_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__buf_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__buf_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.400 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.585000 ;
    PORT
      LAYER li1 ;
        RECT 1.465 1.465 1.795 3.260 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 2.400 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.025 1.085 1.335 1.415 ;
        RECT 0.025 0.215 2.335 1.085 ;
        RECT -0.130 -0.215 2.530 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 2.400 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 2.730 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 2.400 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 2.400 3.815 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.626250 ;
    PORT
      LAYER li1 ;
        RECT 0.115 2.175 0.550 3.755 ;
        RECT 0.115 0.495 0.365 2.175 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 2.400 4.155 ;
        RECT 0.730 2.175 1.285 3.755 ;
        RECT 0.675 1.285 1.005 1.745 ;
        RECT 1.975 1.285 2.225 3.005 ;
        RECT 0.675 1.115 2.225 1.285 ;
        RECT 0.545 0.365 1.795 0.935 ;
        RECT 1.975 0.495 2.225 1.115 ;
        RECT 0.000 -0.085 2.400 0.085 ;
  END
END sky130_fd_sc_hvl__buf_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__buf_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__buf_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.585000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.775 2.775 2.120 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 3.360 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.250 0.215 3.340 1.415 ;
        RECT -0.130 -0.215 3.490 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 3.360 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 3.690 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 3.360 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 3.360 3.815 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.630000 ;
    PORT
      LAYER li1 ;
        RECT 1.200 1.780 1.370 3.755 ;
        RECT 0.125 1.720 1.370 1.780 ;
        RECT 0.125 1.550 1.390 1.720 ;
        RECT 1.220 0.495 1.390 1.550 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 3.360 4.155 ;
        RECT 0.090 2.175 1.020 3.755 ;
        RECT 1.550 2.300 2.800 3.755 ;
        RECT 1.570 1.595 1.865 1.755 ;
        RECT 2.980 1.595 3.250 3.005 ;
        RECT 1.570 1.425 3.250 1.595 ;
        RECT 0.090 0.365 1.040 1.325 ;
        RECT 1.570 0.365 2.820 1.245 ;
        RECT 3.000 0.825 3.250 1.425 ;
        RECT 0.000 -0.085 3.360 0.085 ;
  END
END sky130_fd_sc_hvl__buf_2

#--------EOF---------

MACRO sky130_fd_sc_hvl__buf_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__buf_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.800 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.125000 ;
    PORT
      LAYER li1 ;
        RECT 3.885 1.775 4.215 2.120 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 4.800 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.330 0.215 4.780 1.415 ;
        RECT -0.130 -0.215 4.930 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 4.800 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 5.130 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 4.800 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 4.800 3.815 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.260000 ;
    PORT
      LAYER li1 ;
        RECT 1.220 2.075 1.470 3.755 ;
        RECT 2.780 2.075 3.110 3.755 ;
        RECT 1.220 1.905 3.110 2.075 ;
        RECT 1.220 1.780 1.390 1.905 ;
        RECT 0.125 1.550 1.390 1.780 ;
        RECT 1.220 1.375 1.390 1.550 ;
        RECT 1.220 1.205 3.030 1.375 ;
        RECT 1.220 0.495 1.470 1.205 ;
        RECT 2.780 0.495 3.030 1.205 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 4.800 4.155 ;
        RECT 0.090 2.175 1.040 3.755 ;
        RECT 1.650 2.255 2.600 3.755 ;
        RECT 3.290 2.300 4.240 3.755 ;
        RECT 1.570 1.595 3.600 1.725 ;
        RECT 4.420 1.595 4.670 3.755 ;
        RECT 1.570 1.555 4.670 1.595 ;
        RECT 3.430 1.425 4.670 1.555 ;
        RECT 0.090 0.365 1.040 1.325 ;
        RECT 1.650 0.365 2.600 1.025 ;
        RECT 3.210 0.365 4.160 1.245 ;
        RECT 4.340 0.495 4.670 1.425 ;
        RECT 0.000 -0.085 4.800 0.085 ;
  END
END sky130_fd_sc_hvl__buf_4

#--------EOF---------

MACRO sky130_fd_sc_hvl__buf_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__buf_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.600 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.375000 ;
    PORT
      LAYER li1 ;
        RECT 0.635 1.580 2.245 1.815 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 9.600 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.115 0.215 9.505 1.585 ;
        RECT -0.130 -0.215 9.730 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 9.600 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 9.930 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 9.600 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 9.600 3.815 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.520000 ;
    PORT
      LAYER li1 ;
        RECT 3.605 2.205 3.935 3.445 ;
        RECT 5.165 2.205 5.495 3.445 ;
        RECT 6.725 2.205 7.055 3.445 ;
        RECT 8.285 3.230 8.735 3.445 ;
        RECT 8.285 2.205 8.965 3.230 ;
        RECT 3.605 2.035 8.965 2.205 ;
        RECT 3.665 1.625 8.555 1.795 ;
        RECT 3.665 0.805 3.875 1.625 ;
        RECT 5.225 0.805 5.435 1.625 ;
        RECT 6.785 0.805 6.995 1.625 ;
        RECT 8.345 0.975 8.555 1.625 ;
        RECT 8.735 0.975 8.965 2.035 ;
        RECT 8.345 0.805 8.965 0.975 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 9.600 4.155 ;
        RECT 0.615 3.625 9.505 3.795 ;
        RECT 0.245 2.265 0.435 3.545 ;
        RECT 0.615 2.445 1.865 3.625 ;
        RECT 2.045 2.265 2.595 3.445 ;
        RECT 2.765 2.385 3.435 3.625 ;
        RECT 4.105 2.385 4.995 3.625 ;
        RECT 5.665 2.385 6.555 3.625 ;
        RECT 7.225 2.385 8.115 3.625 ;
        RECT 8.905 3.475 9.505 3.625 ;
        RECT 9.135 2.385 9.505 3.475 ;
        RECT 0.245 2.095 2.595 2.265 ;
        RECT 0.245 1.475 0.435 2.095 ;
        RECT 2.425 1.955 2.595 2.095 ;
        RECT 2.425 1.625 3.380 1.955 ;
        RECT 0.245 0.805 0.455 1.475 ;
        RECT 2.425 1.400 2.595 1.625 ;
        RECT 0.675 0.550 1.925 1.385 ;
        RECT 2.105 1.230 2.595 1.400 ;
        RECT 2.105 0.730 2.315 1.230 ;
        RECT 2.765 0.760 3.495 1.445 ;
        RECT 2.605 0.550 3.495 0.760 ;
        RECT 4.045 0.550 5.055 1.445 ;
        RECT 5.605 0.550 6.615 1.445 ;
        RECT 7.165 0.550 8.175 1.445 ;
        RECT 9.135 0.600 9.505 1.445 ;
        RECT 8.975 0.550 9.505 0.600 ;
        RECT 0.675 0.380 9.505 0.550 ;
        RECT 0.000 -0.085 9.600 0.085 ;
  END
END sky130_fd_sc_hvl__buf_8

#--------EOF---------

MACRO sky130_fd_sc_hvl__buf_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__buf_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.760 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.750000 ;
    PORT
      LAYER li1 ;
        RECT 0.220 1.580 4.630 1.815 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 17.760 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.020 0.215 17.690 1.585 ;
        RECT -0.130 -0.215 17.890 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 17.760 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 18.090 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 17.760 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 17.760 3.815 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.040000 ;
    PORT
      LAYER met1 ;
        RECT 5.590 2.490 5.880 2.520 ;
        RECT 7.150 2.490 7.440 2.520 ;
        RECT 8.710 2.490 9.000 2.520 ;
        RECT 10.270 2.490 10.560 2.520 ;
        RECT 11.830 2.490 12.120 2.520 ;
        RECT 13.390 2.490 13.680 2.520 ;
        RECT 14.950 2.490 15.240 2.520 ;
        RECT 16.510 2.490 16.800 2.520 ;
        RECT 5.590 2.320 16.800 2.490 ;
        RECT 5.590 2.290 5.880 2.320 ;
        RECT 7.150 2.290 7.440 2.320 ;
        RECT 8.710 2.290 9.000 2.320 ;
        RECT 10.270 2.290 10.560 2.320 ;
        RECT 11.830 2.290 12.120 2.320 ;
        RECT 13.390 2.290 13.680 2.320 ;
        RECT 14.950 2.290 15.240 2.320 ;
        RECT 16.510 2.290 16.800 2.320 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 17.760 4.155 ;
        RECT 0.110 2.175 0.680 3.755 ;
        RECT 0.850 2.265 1.160 3.755 ;
        RECT 1.340 2.445 2.230 3.675 ;
        RECT 2.400 2.265 2.710 3.755 ;
        RECT 2.880 2.445 3.770 3.675 ;
        RECT 3.940 2.265 4.290 3.755 ;
        RECT 4.460 2.445 5.350 3.675 ;
        RECT 0.850 1.985 5.350 2.265 ;
        RECT 4.800 1.410 5.350 1.985 ;
        RECT 0.110 0.425 0.645 1.410 ;
        RECT 0.815 1.195 5.350 1.410 ;
        RECT 0.815 0.755 1.170 1.195 ;
        RECT 1.340 0.415 2.230 1.025 ;
        RECT 2.400 0.730 2.790 1.195 ;
        RECT 2.960 0.425 3.855 1.025 ;
        RECT 4.025 0.730 4.270 1.195 ;
        RECT 4.440 0.425 5.330 1.025 ;
        RECT 5.570 0.790 5.900 3.755 ;
        RECT 6.070 2.175 6.960 3.755 ;
        RECT 6.160 1.565 6.830 1.895 ;
        RECT 6.070 0.425 6.960 1.395 ;
        RECT 7.130 0.790 7.460 3.755 ;
        RECT 7.630 2.175 8.520 3.755 ;
        RECT 7.720 1.565 8.390 1.895 ;
        RECT 7.630 0.425 8.520 1.395 ;
        RECT 8.690 0.790 9.020 3.755 ;
        RECT 9.190 2.175 10.080 3.755 ;
        RECT 9.280 1.565 9.950 1.895 ;
        RECT 9.190 0.425 10.080 1.395 ;
        RECT 10.250 0.790 10.580 3.755 ;
        RECT 10.750 2.175 11.640 3.755 ;
        RECT 10.840 1.565 11.510 1.895 ;
        RECT 10.750 0.425 11.640 1.395 ;
        RECT 11.810 0.790 12.140 3.755 ;
        RECT 12.310 2.175 13.200 3.755 ;
        RECT 12.400 1.565 13.070 1.895 ;
        RECT 12.310 0.425 13.200 1.395 ;
        RECT 13.370 0.790 13.700 3.755 ;
        RECT 13.870 2.175 14.760 3.755 ;
        RECT 13.960 1.565 14.630 1.895 ;
        RECT 13.870 0.425 14.760 1.395 ;
        RECT 14.930 0.790 15.260 3.755 ;
        RECT 15.430 2.175 16.320 3.755 ;
        RECT 15.520 1.565 16.190 1.895 ;
        RECT 15.430 0.425 16.320 1.395 ;
        RECT 16.490 0.790 16.900 3.755 ;
        RECT 17.070 2.175 17.600 3.755 ;
        RECT 17.070 0.425 17.600 1.495 ;
        RECT 0.000 -0.085 17.760 0.085 ;
      LAYER met1 ;
        RECT 4.740 1.750 5.360 1.780 ;
        RECT 6.170 1.750 6.820 1.780 ;
        RECT 7.730 1.750 8.380 1.780 ;
        RECT 9.290 1.750 9.940 1.780 ;
        RECT 10.850 1.750 11.500 1.780 ;
        RECT 12.410 1.750 13.060 1.780 ;
        RECT 13.970 1.750 14.620 1.780 ;
        RECT 15.530 1.750 16.180 1.780 ;
        RECT 4.740 1.580 16.250 1.750 ;
        RECT 4.740 1.550 5.360 1.580 ;
        RECT 6.170 1.550 6.820 1.580 ;
        RECT 7.730 1.550 8.380 1.580 ;
        RECT 9.290 1.550 9.940 1.580 ;
        RECT 10.850 1.550 11.500 1.580 ;
        RECT 12.410 1.550 13.060 1.580 ;
        RECT 13.970 1.550 14.620 1.580 ;
        RECT 15.530 1.550 16.180 1.580 ;
  END
END sky130_fd_sc_hvl__buf_16

#--------EOF---------

MACRO sky130_fd_sc_hvl__buf_32
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__buf_32 ;
  ORIGIN 0.000 0.000 ;
  SIZE 33.600 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 11.250000 ;
    PORT
      LAYER li1 ;
        RECT 0.220 1.580 4.630 1.815 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 33.600 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.020 0.215 33.530 1.585 ;
        RECT -0.130 -0.215 33.730 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 33.600 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 33.930 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 33.600 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 33.600 3.815 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 10.080000 ;
    PORT
      LAYER met1 ;
        RECT 8.950 2.290 32.640 2.520 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 33.600 4.155 ;
        RECT 0.110 2.175 0.680 3.755 ;
        RECT 0.850 2.265 1.160 3.755 ;
        RECT 1.340 2.445 2.230 3.675 ;
        RECT 2.400 2.265 2.710 3.755 ;
        RECT 2.880 2.445 3.770 3.675 ;
        RECT 3.940 2.265 4.290 3.755 ;
        RECT 4.460 2.445 5.350 3.675 ;
        RECT 5.520 2.265 5.830 3.755 ;
        RECT 6.000 2.445 6.890 3.675 ;
        RECT 7.060 2.265 7.410 3.755 ;
        RECT 0.850 1.985 7.410 2.265 ;
        RECT 7.580 2.235 8.480 3.675 ;
        RECT 4.800 1.410 7.410 1.985 ;
        RECT 0.110 0.425 0.645 1.410 ;
        RECT 0.815 1.195 7.410 1.410 ;
        RECT 0.815 0.755 1.170 1.195 ;
        RECT 1.340 0.415 2.230 1.025 ;
        RECT 2.400 0.730 2.790 1.195 ;
        RECT 2.960 0.425 3.855 1.025 ;
        RECT 4.025 0.730 4.270 1.195 ;
        RECT 4.440 0.425 5.330 1.025 ;
        RECT 5.520 0.730 5.910 1.195 ;
        RECT 6.080 0.425 6.975 1.025 ;
        RECT 7.145 0.730 7.390 1.195 ;
        RECT 7.580 1.025 8.480 1.395 ;
        RECT 7.560 0.425 8.480 1.025 ;
        RECT 8.930 0.790 9.260 3.755 ;
        RECT 9.430 2.175 10.320 3.755 ;
        RECT 9.520 1.565 10.190 1.895 ;
        RECT 9.430 0.425 10.320 1.395 ;
        RECT 10.490 0.790 10.820 3.755 ;
        RECT 10.990 2.175 11.880 3.755 ;
        RECT 11.080 1.565 11.750 1.895 ;
        RECT 10.990 0.425 11.880 1.395 ;
        RECT 12.050 0.790 12.380 3.755 ;
        RECT 12.550 2.175 13.440 3.755 ;
        RECT 12.640 1.565 13.310 1.895 ;
        RECT 12.550 0.425 13.440 1.395 ;
        RECT 13.610 0.790 13.940 3.755 ;
        RECT 14.110 2.175 15.000 3.755 ;
        RECT 14.200 1.565 14.870 1.895 ;
        RECT 14.110 0.425 15.000 1.395 ;
        RECT 15.170 0.790 15.500 3.755 ;
        RECT 15.670 2.175 16.560 3.755 ;
        RECT 15.760 1.565 16.430 1.895 ;
        RECT 15.670 0.425 16.560 1.395 ;
        RECT 16.730 0.790 17.060 3.755 ;
        RECT 17.230 2.175 18.120 3.755 ;
        RECT 17.320 1.565 17.990 1.895 ;
        RECT 17.230 0.425 18.120 1.395 ;
        RECT 18.290 0.790 18.620 3.755 ;
        RECT 18.790 2.175 19.680 3.755 ;
        RECT 18.880 1.565 19.550 1.895 ;
        RECT 18.790 0.425 19.680 1.395 ;
        RECT 19.850 0.790 20.260 3.755 ;
        RECT 20.430 2.175 20.960 3.755 ;
        RECT 20.430 1.565 21.100 1.895 ;
        RECT 20.430 0.425 20.960 1.395 ;
        RECT 21.410 0.790 21.740 3.755 ;
        RECT 21.910 2.175 22.800 3.755 ;
        RECT 22.000 1.565 22.670 1.895 ;
        RECT 21.910 0.425 22.800 1.395 ;
        RECT 22.970 0.790 23.300 3.755 ;
        RECT 23.470 2.175 24.360 3.755 ;
        RECT 23.560 1.565 24.230 1.895 ;
        RECT 23.470 0.425 24.360 1.395 ;
        RECT 24.530 0.790 24.860 3.755 ;
        RECT 25.030 2.175 25.920 3.755 ;
        RECT 25.120 1.565 25.790 1.895 ;
        RECT 25.030 0.425 25.920 1.395 ;
        RECT 26.090 0.790 26.420 3.755 ;
        RECT 26.590 2.175 27.480 3.755 ;
        RECT 26.680 1.565 27.350 1.895 ;
        RECT 26.590 0.425 27.480 1.395 ;
        RECT 27.650 0.790 27.980 3.755 ;
        RECT 28.150 2.175 29.040 3.755 ;
        RECT 28.240 1.565 28.910 1.895 ;
        RECT 28.150 0.425 29.040 1.395 ;
        RECT 29.210 0.790 29.540 3.755 ;
        RECT 29.710 2.175 30.600 3.755 ;
        RECT 29.800 1.565 30.470 1.895 ;
        RECT 29.710 0.425 30.600 1.395 ;
        RECT 30.770 0.790 31.100 3.755 ;
        RECT 31.270 2.175 32.160 3.755 ;
        RECT 31.360 1.565 32.030 1.895 ;
        RECT 31.270 0.425 32.160 1.395 ;
        RECT 32.330 0.790 32.740 3.755 ;
        RECT 32.910 2.175 33.440 3.755 ;
        RECT 32.910 0.425 33.440 1.495 ;
        RECT 0.000 -0.085 33.600 0.085 ;
      LAYER met1 ;
        RECT 4.960 1.550 32.090 1.780 ;
  END
END sky130_fd_sc_hvl__buf_32

#--------EOF---------

MACRO sky130_fd_sc_hvl__conb_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__conb_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.400 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 2.400 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.130 -0.215 2.530 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 2.400 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 2.730 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 2.400 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 2.400 3.815 ;
    END
  END VPWR
  PIN HI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.075 2.185 1.325 3.530 ;
        RECT 0.615 1.935 1.325 2.185 ;
        RECT 0.615 1.070 0.865 1.935 ;
        RECT 0.290 0.430 0.865 1.070 ;
    END
  END HI
  PIN LO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.530 3.175 2.110 3.815 ;
        RECT 1.530 1.765 1.795 3.175 ;
        RECT 1.035 1.500 1.795 1.765 ;
        RECT 1.035 0.500 1.365 1.500 ;
    END
  END LO
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 2.400 4.155 ;
        RECT 0.215 3.445 0.865 3.785 ;
        RECT 0.215 3.175 0.620 3.445 ;
        RECT 1.780 0.625 2.185 1.070 ;
        RECT 1.535 0.285 2.185 0.625 ;
        RECT 0.000 -0.085 2.400 0.085 ;
  END
END sky130_fd_sc_hvl__conb_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__decap_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__decap_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.920 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 1.920 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.080 0.215 1.890 1.475 ;
        RECT -0.130 -0.215 2.050 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 1.920 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 2.250 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 1.920 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 1.920 3.815 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 1.920 4.155 ;
        RECT 0.250 2.685 1.700 3.755 ;
        RECT 0.475 1.250 0.805 2.030 ;
        RECT 1.015 1.700 1.345 2.685 ;
        RECT 0.475 0.845 1.780 1.250 ;
        RECT 0.170 0.365 1.780 0.845 ;
        RECT 0.000 -0.085 1.920 0.085 ;
  END
END sky130_fd_sc_hvl__decap_4

#--------EOF---------

MACRO sky130_fd_sc_hvl__decap_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__decap_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.840 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 3.840 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.405 0.215 3.495 1.470 ;
        RECT -0.130 -0.215 3.970 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 3.840 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 4.170 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 3.840 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 3.840 3.815 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 3.840 4.155 ;
        RECT 0.500 2.680 3.240 3.750 ;
        RECT 0.735 1.360 1.065 2.025 ;
        RECT 1.470 1.695 1.800 2.680 ;
        RECT 2.015 1.360 2.345 2.025 ;
        RECT 2.750 1.695 3.080 2.680 ;
        RECT 0.575 0.360 3.305 1.360 ;
        RECT 0.000 -0.085 3.840 0.085 ;
  END
END sky130_fd_sc_hvl__decap_8

#--------EOF---------

MACRO sky130_fd_sc_hvl__dfrbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__dfrbp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.800 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.585000 ;
    PORT
      LAYER li1 ;
        RECT 0.595 1.175 0.925 1.720 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER li1 ;
        RECT 3.850 0.810 4.165 2.105 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.260000 ;
    PORT
      LAYER li1 ;
        RECT 2.980 1.505 3.665 2.120 ;
        RECT 7.165 1.825 8.515 1.995 ;
        RECT 3.495 0.630 3.665 1.505 ;
        RECT 8.345 1.295 8.515 1.825 ;
        RECT 6.455 1.125 8.515 1.295 ;
        RECT 11.510 1.130 11.840 1.350 ;
        RECT 6.455 0.630 6.625 1.125 ;
        RECT 3.495 0.460 6.625 0.630 ;
        RECT 8.345 0.435 8.515 1.125 ;
        RECT 10.905 0.960 11.840 1.130 ;
        RECT 10.905 0.435 11.075 0.960 ;
        RECT 8.345 0.265 11.075 0.435 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 16.800 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 13.205 1.415 14.535 1.585 ;
        RECT 2.725 1.085 9.880 1.415 ;
        RECT 13.205 1.085 16.780 1.415 ;
        RECT 0.055 0.215 16.780 1.085 ;
        RECT -0.130 -0.215 16.930 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 16.800 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 17.130 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 16.800 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 16.800 3.815 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.626250 ;
    PORT
      LAYER li1 ;
        RECT 16.340 0.515 16.690 3.755 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.641250 ;
    PORT
      LAYER li1 ;
        RECT 14.130 1.780 14.380 3.755 ;
        RECT 14.045 1.495 14.380 1.780 ;
        RECT 14.045 0.665 14.425 1.495 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 16.800 4.155 ;
        RECT 0.165 2.445 0.415 3.455 ;
        RECT 0.595 2.625 1.485 3.705 ;
        RECT 1.665 3.635 3.205 3.805 ;
        RECT 1.665 2.445 1.835 3.635 ;
        RECT 0.165 2.275 1.835 2.445 ;
        RECT 0.165 0.995 0.415 2.275 ;
        RECT 1.505 1.900 1.835 2.275 ;
        RECT 2.015 1.550 2.275 3.455 ;
        RECT 2.525 2.470 2.855 3.420 ;
        RECT 3.035 2.820 3.205 3.635 ;
        RECT 3.385 3.000 3.555 3.705 ;
        RECT 3.735 3.600 5.565 3.770 ;
        RECT 3.735 2.820 3.905 3.600 ;
        RECT 4.085 3.000 4.515 3.420 ;
        RECT 4.865 3.000 5.215 3.420 ;
        RECT 3.035 2.650 3.905 2.820 ;
        RECT 4.345 2.470 4.515 3.000 ;
        RECT 2.525 2.300 4.515 2.470 ;
        RECT 2.015 0.995 2.185 1.550 ;
        RECT 4.345 1.325 4.515 2.300 ;
        RECT 4.695 1.780 4.865 2.820 ;
        RECT 5.045 2.370 5.215 3.000 ;
        RECT 5.395 3.045 5.565 3.600 ;
        RECT 5.745 3.225 6.685 3.705 ;
        RECT 6.865 3.635 7.735 3.805 ;
        RECT 6.865 3.045 7.035 3.635 ;
        RECT 5.395 2.875 7.035 3.045 ;
        RECT 5.395 2.550 5.650 2.875 ;
        RECT 7.215 2.695 7.385 3.455 ;
        RECT 7.565 2.870 7.735 3.635 ;
        RECT 7.915 3.050 8.865 3.705 ;
        RECT 7.565 2.700 9.375 2.870 ;
        RECT 6.105 2.525 7.385 2.695 ;
        RECT 6.105 2.370 6.275 2.525 ;
        RECT 5.045 2.200 6.275 2.370 ;
        RECT 8.695 2.345 9.025 2.520 ;
        RECT 5.595 1.780 5.925 2.020 ;
        RECT 4.695 1.505 5.925 1.780 ;
        RECT 6.105 1.645 6.275 2.200 ;
        RECT 6.455 2.175 9.025 2.345 ;
        RECT 6.455 1.825 6.785 2.175 ;
        RECT 6.105 1.475 8.165 1.645 ;
        RECT 6.105 1.325 6.275 1.475 ;
        RECT 0.165 0.495 0.495 0.995 ;
        RECT 0.675 0.365 1.625 0.995 ;
        RECT 1.805 0.495 2.185 0.995 ;
        RECT 2.365 0.365 3.315 1.325 ;
        RECT 4.345 0.825 4.655 1.325 ;
        RECT 5.270 1.155 6.275 1.325 ;
        RECT 5.270 0.825 5.600 1.155 ;
        RECT 7.215 0.365 8.165 0.945 ;
        RECT 8.695 0.615 9.025 2.175 ;
        RECT 9.205 1.400 9.375 2.700 ;
        RECT 9.555 2.440 9.805 3.350 ;
        RECT 9.555 2.270 10.410 2.440 ;
        RECT 10.590 2.350 11.540 3.705 ;
        RECT 11.965 2.520 12.295 2.770 ;
        RECT 11.965 2.350 12.880 2.520 ;
        RECT 10.240 2.170 10.410 2.270 ;
        RECT 9.725 1.580 10.060 2.090 ;
        RECT 10.240 2.000 12.530 2.170 ;
        RECT 9.205 1.230 10.375 1.400 ;
        RECT 10.090 1.070 10.375 1.230 ;
        RECT 9.580 0.785 9.910 0.995 ;
        RECT 10.555 0.785 10.725 2.000 ;
        RECT 12.200 1.880 12.530 2.000 ;
        RECT 10.930 1.700 11.260 1.820 ;
        RECT 12.710 1.700 12.880 2.350 ;
        RECT 13.060 2.175 13.950 3.755 ;
        RECT 10.930 1.530 12.880 1.700 ;
        RECT 10.930 1.310 11.260 1.530 ;
        RECT 9.580 0.615 10.725 0.785 ;
        RECT 12.710 0.975 12.880 1.530 ;
        RECT 14.665 1.835 14.995 3.005 ;
        RECT 15.175 2.175 16.125 3.755 ;
        RECT 14.665 1.505 16.160 1.835 ;
        RECT 11.255 0.365 12.205 0.780 ;
        RECT 12.710 0.515 13.075 0.975 ;
        RECT 13.255 0.365 13.845 1.495 ;
        RECT 14.665 0.825 15.015 1.505 ;
        RECT 15.195 0.365 16.145 1.325 ;
        RECT 0.000 -0.085 16.800 0.085 ;
      LAYER met1 ;
        RECT 2.015 1.735 2.305 1.780 ;
        RECT 4.895 1.735 5.185 1.780 ;
        RECT 9.695 1.735 9.985 1.780 ;
        RECT 2.015 1.595 9.985 1.735 ;
        RECT 2.015 1.550 2.305 1.595 ;
        RECT 4.895 1.550 5.185 1.595 ;
        RECT 9.695 1.550 9.985 1.595 ;
  END
END sky130_fd_sc_hvl__dfrbp_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__dfrtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__dfrtp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.360 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.585000 ;
    PORT
      LAYER li1 ;
        RECT 0.560 1.175 0.890 2.150 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER li1 ;
        RECT 3.415 0.810 3.745 2.105 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.260000 ;
    PORT
      LAYER li1 ;
        RECT 2.695 1.620 3.235 2.490 ;
        RECT 6.605 1.825 8.460 1.995 ;
        RECT 3.065 0.630 3.235 1.620 ;
        RECT 8.290 1.295 8.460 1.825 ;
        RECT 5.840 1.125 8.460 1.295 ;
        RECT 11.455 1.265 11.785 1.655 ;
        RECT 5.840 0.630 6.010 1.125 ;
        RECT 3.065 0.460 6.010 0.630 ;
        RECT 8.290 0.435 8.460 1.125 ;
        RECT 10.780 1.095 11.785 1.265 ;
        RECT 10.780 0.435 10.950 1.095 ;
        RECT 8.290 0.265 10.950 0.435 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 15.360 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.270 1.085 9.870 1.415 ;
        RECT 13.115 1.085 15.340 1.585 ;
        RECT 0.020 0.215 15.340 1.085 ;
        RECT -0.130 -0.215 15.490 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 15.360 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 15.690 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 15.360 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 15.360 3.815 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.611250 ;
    PORT
      LAYER li1 ;
        RECT 14.900 0.665 15.235 3.735 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 15.360 4.155 ;
        RECT 0.110 2.525 0.440 3.455 ;
        RECT 0.630 2.725 1.220 3.705 ;
        RECT 1.400 3.635 2.840 3.805 ;
        RECT 1.400 2.525 1.570 3.635 ;
        RECT 0.110 2.355 1.570 2.525 ;
        RECT 0.110 0.495 0.380 2.355 ;
        RECT 1.240 1.855 1.570 2.355 ;
        RECT 1.750 2.150 2.000 3.455 ;
        RECT 2.240 2.840 2.490 3.455 ;
        RECT 2.670 3.190 2.840 3.635 ;
        RECT 3.020 3.370 3.350 3.705 ;
        RECT 3.530 3.635 5.270 3.805 ;
        RECT 3.530 3.190 3.700 3.635 ;
        RECT 2.670 3.020 3.700 3.190 ;
        RECT 3.880 2.840 4.050 3.455 ;
        RECT 4.580 3.200 4.910 3.455 ;
        RECT 2.240 2.670 4.050 2.840 ;
        RECT 4.230 2.670 4.450 3.000 ;
        RECT 3.880 2.490 4.050 2.670 ;
        RECT 3.880 2.320 4.100 2.490 ;
        RECT 1.750 1.920 2.275 2.150 ;
        RECT 1.750 0.995 2.020 1.920 ;
        RECT 3.930 1.325 4.100 2.320 ;
        RECT 4.280 2.150 4.450 2.670 ;
        RECT 4.630 2.500 4.800 3.200 ;
        RECT 5.100 3.045 5.270 3.635 ;
        RECT 5.450 3.225 6.400 3.705 ;
        RECT 6.580 3.635 7.610 3.805 ;
        RECT 6.580 3.045 6.750 3.635 ;
        RECT 5.100 3.000 6.750 3.045 ;
        RECT 4.980 2.875 6.750 3.000 ;
        RECT 4.980 2.680 5.310 2.875 ;
        RECT 6.930 2.695 7.260 3.455 ;
        RECT 7.440 3.275 7.610 3.635 ;
        RECT 7.790 3.455 8.740 3.755 ;
        RECT 7.440 3.105 9.250 3.275 ;
        RECT 5.490 2.525 7.260 2.695 ;
        RECT 5.490 2.500 5.660 2.525 ;
        RECT 4.630 2.330 5.660 2.500 ;
        RECT 8.570 2.345 8.900 2.925 ;
        RECT 4.280 1.920 5.305 2.150 ;
        RECT 4.975 1.425 5.305 1.920 ;
        RECT 5.490 1.645 5.660 2.330 ;
        RECT 5.840 2.175 8.900 2.345 ;
        RECT 5.840 1.825 6.170 2.175 ;
        RECT 5.490 1.475 8.110 1.645 ;
        RECT 0.560 0.365 1.510 0.995 ;
        RECT 1.690 0.495 2.020 0.995 ;
        RECT 2.200 0.365 2.790 1.245 ;
        RECT 3.930 0.825 4.200 1.325 ;
        RECT 5.490 1.245 5.660 1.475 ;
        RECT 4.650 1.075 5.660 1.245 ;
        RECT 8.640 1.325 8.900 2.175 ;
        RECT 9.080 1.755 9.250 3.105 ;
        RECT 9.430 2.845 9.680 3.755 ;
        RECT 9.430 2.675 10.305 2.845 ;
        RECT 10.485 2.675 11.435 3.705 ;
        RECT 11.840 2.705 12.090 3.175 ;
        RECT 12.270 2.885 13.165 3.705 ;
        RECT 9.625 1.935 9.955 2.435 ;
        RECT 10.135 2.355 10.305 2.675 ;
        RECT 11.840 2.535 12.845 2.705 ;
        RECT 10.135 2.185 12.495 2.355 ;
        RECT 9.080 1.585 10.250 1.755 ;
        RECT 4.650 0.825 4.980 1.075 ;
        RECT 7.160 0.365 8.110 0.945 ;
        RECT 8.640 0.615 8.970 1.325 ;
        RECT 9.430 0.785 9.760 1.325 ;
        RECT 9.965 1.085 10.250 1.585 ;
        RECT 10.430 0.785 10.600 2.185 ;
        RECT 12.675 2.005 12.845 2.535 ;
        RECT 10.805 1.835 12.845 2.005 ;
        RECT 10.805 1.445 11.135 1.835 ;
        RECT 12.620 0.995 12.845 1.835 ;
        RECT 13.345 2.005 13.595 3.005 ;
        RECT 13.775 2.195 14.720 3.735 ;
        RECT 13.345 1.675 14.720 2.005 ;
        RECT 13.345 1.495 13.555 1.675 ;
        RECT 13.225 0.995 13.555 1.495 ;
        RECT 9.430 0.615 10.600 0.785 ;
        RECT 11.130 0.365 12.080 0.915 ;
        RECT 12.620 0.495 12.950 0.995 ;
        RECT 13.735 0.365 14.685 1.495 ;
        RECT 0.000 -0.085 15.360 0.085 ;
      LAYER met1 ;
        RECT 2.015 2.105 2.305 2.150 ;
        RECT 4.415 2.105 4.705 2.150 ;
        RECT 9.695 2.105 9.985 2.150 ;
        RECT 2.015 1.965 9.985 2.105 ;
        RECT 2.015 1.920 2.305 1.965 ;
        RECT 4.415 1.920 4.705 1.965 ;
        RECT 9.695 1.920 9.985 1.965 ;
  END
END sky130_fd_sc_hvl__dfrtp_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__dfsbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__dfsbp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 17.760 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.585000 ;
    PORT
      LAYER li1 ;
        RECT 0.560 1.550 0.890 2.520 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.515 2.875 2.145 ;
    END
  END D
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.840000 ;
    PORT
      LAYER li1 ;
        RECT 10.715 1.975 12.830 2.145 ;
        RECT 10.715 1.775 10.885 1.975 ;
        RECT 10.160 1.605 10.885 1.775 ;
        RECT 10.160 1.325 10.330 1.605 ;
        RECT 12.150 1.555 12.830 1.975 ;
        RECT 6.985 1.155 10.330 1.325 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 17.760 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 9.540 1.645 10.090 1.845 ;
        RECT 7.315 1.315 8.605 1.415 ;
        RECT 9.540 1.315 11.200 1.645 ;
        RECT 0.020 1.095 2.090 1.110 ;
        RECT 0.020 1.085 5.690 1.095 ;
        RECT 7.315 1.085 11.200 1.315 ;
        RECT 13.280 1.085 17.740 1.415 ;
        RECT 0.020 0.215 17.740 1.085 ;
        RECT -0.130 -0.215 17.890 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 17.760 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 2.385 18.090 4.485 ;
        RECT -0.330 1.885 5.990 2.385 ;
        RECT 11.500 1.885 18.090 2.385 ;
      LAYER met1 ;
        RECT 0.000 3.955 17.760 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 17.760 3.815 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.498750 ;
    PORT
      LAYER li1 ;
        RECT 17.300 2.355 17.635 3.435 ;
        RECT 17.405 1.325 17.635 2.355 ;
        RECT 17.300 0.495 17.635 1.325 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.641250 ;
    PORT
      LAYER li1 ;
        RECT 15.015 0.495 15.375 3.755 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 17.760 4.155 ;
        RECT 0.110 1.370 0.380 3.450 ;
        RECT 0.650 2.700 1.240 3.705 ;
        RECT 1.420 3.630 2.290 3.800 ;
        RECT 1.420 1.870 1.590 3.630 ;
        RECT 1.260 1.370 1.590 1.870 ;
        RECT 0.110 1.200 1.590 1.370 ;
        RECT 1.770 1.335 1.940 3.450 ;
        RECT 2.120 2.495 2.290 3.630 ;
        RECT 2.470 2.675 2.675 3.705 ;
        RECT 2.855 3.355 5.500 3.525 ;
        RECT 2.855 2.495 3.025 3.355 ;
        RECT 2.120 2.325 3.025 2.495 ;
        RECT 3.205 2.675 3.545 3.175 ;
        RECT 0.110 0.540 0.360 1.200 ;
        RECT 1.770 1.165 2.820 1.335 ;
        RECT 0.540 0.365 1.490 1.020 ;
        RECT 1.770 1.000 2.000 1.165 ;
        RECT 1.670 0.540 2.000 1.000 ;
        RECT 2.220 0.365 2.470 0.985 ;
        RECT 2.650 0.435 2.820 1.165 ;
        RECT 3.205 1.005 3.375 2.675 ;
        RECT 3.725 2.395 3.895 3.355 ;
        RECT 4.075 3.005 5.150 3.175 ;
        RECT 4.075 2.675 4.405 3.005 ;
        RECT 4.585 2.395 4.800 2.555 ;
        RECT 3.555 2.225 4.800 2.395 ;
        RECT 3.555 1.105 3.725 2.225 ;
        RECT 4.980 2.025 5.150 3.005 ;
        RECT 5.330 2.725 5.500 3.355 ;
        RECT 5.680 2.905 6.245 3.705 ;
        RECT 6.425 3.355 7.675 3.525 ;
        RECT 6.425 2.725 6.595 3.355 ;
        RECT 5.330 2.555 6.595 2.725 ;
        RECT 6.775 2.375 7.025 3.175 ;
        RECT 7.505 2.715 7.675 3.355 ;
        RECT 7.855 2.895 8.805 3.705 ;
        RECT 9.345 3.585 10.535 3.755 ;
        RECT 7.505 2.545 9.120 2.715 ;
        RECT 9.345 2.675 9.675 3.585 ;
        RECT 5.330 2.205 7.025 2.375 ;
        RECT 7.730 2.025 8.060 2.365 ;
        RECT 3.905 1.855 8.060 2.025 ;
        RECT 8.870 1.885 9.120 2.545 ;
        RECT 9.855 2.475 10.185 2.555 ;
        RECT 9.300 2.305 10.185 2.475 ;
        RECT 10.365 2.495 10.535 3.585 ;
        RECT 10.715 2.675 11.665 3.705 ;
        RECT 12.035 2.495 13.180 3.175 ;
        RECT 10.365 2.325 13.180 2.495 ;
        RECT 3.000 0.615 3.375 1.005 ;
        RECT 3.905 0.925 4.075 1.855 ;
        RECT 9.300 1.675 9.470 2.305 ;
        RECT 10.365 2.125 10.535 2.325 ;
        RECT 4.255 1.505 9.470 1.675 ;
        RECT 9.650 1.955 10.535 2.125 ;
        RECT 9.650 1.505 9.980 1.955 ;
        RECT 4.255 1.105 4.585 1.505 ;
        RECT 3.780 0.615 4.110 0.925 ;
        RECT 4.290 0.435 4.460 1.105 ;
        RECT 4.945 1.085 6.150 1.325 ;
        RECT 2.650 0.265 4.460 0.435 ;
        RECT 4.650 0.365 5.600 0.905 ;
        RECT 5.820 0.515 6.150 1.085 ;
        RECT 10.510 1.255 11.460 1.425 ;
        RECT 10.510 0.975 10.680 1.255 ;
        RECT 6.785 0.365 7.735 0.975 ;
        RECT 8.185 0.545 8.515 0.975 ;
        RECT 8.755 0.725 10.680 0.975 ;
        RECT 10.860 0.545 11.110 1.075 ;
        RECT 8.185 0.375 11.110 0.545 ;
        RECT 11.290 0.975 11.460 1.255 ;
        RECT 11.640 1.375 11.970 1.795 ;
        RECT 13.010 1.725 13.180 2.325 ;
        RECT 13.360 2.075 13.690 2.675 ;
        RECT 13.870 2.255 14.820 3.755 ;
        RECT 13.360 1.905 14.395 2.075 ;
        RECT 13.010 1.555 14.045 1.725 ;
        RECT 14.225 1.375 14.395 1.905 ;
        RECT 11.640 1.205 14.395 1.375 ;
        RECT 15.625 1.675 15.955 3.185 ;
        RECT 16.135 2.355 17.085 3.705 ;
        RECT 16.845 1.675 17.175 2.175 ;
        RECT 15.625 1.505 17.175 1.675 ;
        RECT 11.640 1.155 11.970 1.205 ;
        RECT 11.290 0.515 11.660 0.975 ;
        RECT 12.200 0.365 13.150 0.975 ;
        RECT 13.390 0.825 13.720 1.205 ;
        RECT 13.900 0.365 14.835 1.025 ;
        RECT 15.625 0.825 15.975 1.505 ;
        RECT 16.155 0.365 17.105 1.305 ;
        RECT 0.000 -0.085 17.760 0.085 ;
  END
END sky130_fd_sc_hvl__dfsbp_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__dfstp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__dfstp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.880 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.585000 ;
    PORT
      LAYER li1 ;
        RECT 0.545 2.075 0.875 2.745 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER li1 ;
        RECT 2.505 1.525 2.835 2.095 ;
    END
  END D
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.840000 ;
    PORT
      LAYER li1 ;
        RECT 7.165 1.555 8.100 1.795 ;
        RECT 7.930 1.010 8.100 1.555 ;
        RECT 10.885 1.010 11.160 1.040 ;
        RECT 7.930 0.840 11.160 1.010 ;
        RECT 8.285 0.555 11.160 0.840 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 14.880 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 5.445 1.565 6.870 1.805 ;
        RECT 0.020 1.085 2.130 1.205 ;
        RECT 5.445 1.085 14.860 1.565 ;
        RECT 0.020 0.215 14.860 1.085 ;
        RECT -0.130 -0.215 15.010 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 14.880 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 2.245 15.210 4.485 ;
        RECT -0.330 1.885 5.145 2.245 ;
        RECT 7.170 1.885 15.210 2.245 ;
      LAYER met1 ;
        RECT 0.000 3.955 14.880 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 14.880 3.815 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.478750 ;
    PORT
      LAYER li1 ;
        RECT 14.420 0.645 14.770 3.615 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 14.880 4.155 ;
        RECT 0.115 1.465 0.365 3.735 ;
        RECT 0.545 2.925 1.495 3.755 ;
        RECT 1.675 2.945 2.005 3.735 ;
        RECT 1.690 2.445 2.005 2.945 ;
        RECT 2.235 2.625 2.485 3.705 ;
        RECT 2.665 2.445 2.835 3.755 ;
        RECT 1.690 2.275 2.835 2.445 ;
        RECT 3.015 3.285 5.005 3.615 ;
        RECT 1.180 1.465 1.510 1.895 ;
        RECT 0.115 1.295 1.510 1.465 ;
        RECT 0.115 0.615 0.380 1.295 ;
        RECT 0.570 0.365 1.160 1.115 ;
        RECT 1.340 0.435 1.510 1.295 ;
        RECT 1.690 0.615 1.940 2.275 ;
        RECT 3.015 1.345 3.185 3.285 ;
        RECT 2.120 1.175 3.185 1.345 ;
        RECT 2.120 0.435 2.290 1.175 ;
        RECT 3.365 0.995 3.535 3.105 ;
        RECT 3.715 1.085 3.885 3.285 ;
        RECT 4.065 2.605 4.395 3.105 ;
        RECT 4.065 1.135 4.235 2.605 ;
        RECT 4.835 2.325 5.005 3.285 ;
        RECT 5.185 2.675 5.425 3.555 ;
        RECT 5.605 2.855 5.935 3.705 ;
        RECT 6.565 2.845 6.895 3.105 ;
        RECT 6.115 2.675 6.895 2.845 ;
        RECT 7.075 2.675 8.025 3.705 ;
        RECT 8.695 3.595 9.825 3.805 ;
        RECT 8.695 2.845 8.865 3.595 ;
        RECT 9.045 3.025 9.660 3.415 ;
        RECT 8.695 2.675 9.310 2.845 ;
        RECT 5.185 2.505 6.285 2.675 ;
        RECT 6.465 2.325 8.960 2.495 ;
        RECT 4.415 1.975 4.655 2.165 ;
        RECT 4.835 2.155 6.635 2.325 ;
        RECT 6.815 1.975 8.450 2.145 ;
        RECT 8.630 2.085 8.960 2.325 ;
        RECT 4.415 1.805 6.985 1.975 ;
        RECT 8.280 1.875 8.450 1.975 ;
        RECT 9.140 1.875 9.310 2.675 ;
        RECT 4.415 1.495 4.655 1.805 ;
        RECT 8.280 1.705 9.310 1.875 ;
        RECT 9.490 2.485 9.660 3.025 ;
        RECT 10.010 2.665 10.960 3.705 ;
        RECT 11.300 3.255 11.550 3.755 ;
        RECT 11.730 3.355 12.680 3.735 ;
        RECT 11.380 3.175 11.550 3.255 ;
        RECT 11.380 3.005 12.560 3.175 ;
        RECT 11.410 2.675 11.740 2.825 ;
        RECT 11.410 2.485 12.210 2.675 ;
        RECT 9.490 2.315 12.210 2.485 ;
        RECT 5.135 1.315 5.865 1.625 ;
        RECT 8.280 1.545 8.785 1.705 ;
        RECT 9.490 1.475 9.660 2.315 ;
        RECT 10.305 1.825 10.635 2.135 ;
        RECT 11.880 2.005 12.210 2.315 ;
        RECT 12.390 1.825 12.560 3.005 ;
        RECT 10.305 1.655 12.560 1.825 ;
        RECT 12.865 2.395 13.115 3.365 ;
        RECT 13.295 2.575 14.240 3.705 ;
        RECT 12.865 2.225 14.240 2.395 ;
        RECT 10.305 1.545 10.635 1.655 ;
        RECT 1.340 0.265 2.290 0.435 ;
        RECT 2.470 0.365 3.005 0.995 ;
        RECT 3.185 0.495 3.535 0.995 ;
        RECT 4.065 0.965 6.315 1.135 ;
        RECT 4.065 0.495 4.315 0.965 ;
        RECT 4.855 0.365 5.805 0.785 ;
        RECT 5.985 0.265 6.315 0.965 ;
        RECT 6.800 0.365 7.750 1.375 ;
        RECT 9.025 1.190 9.660 1.475 ;
        RECT 11.340 0.365 11.930 1.475 ;
        RECT 12.120 0.975 12.450 1.655 ;
        RECT 12.865 1.475 13.075 2.225 ;
        RECT 13.910 1.725 14.240 2.225 ;
        RECT 12.745 0.975 13.075 1.475 ;
        RECT 13.255 0.365 14.205 1.475 ;
        RECT 0.000 -0.085 14.880 0.085 ;
  END
END sky130_fd_sc_hvl__dfstp_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__dfxbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__dfxbp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.920 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.585000 ;
    PORT
      LAYER li1 ;
        RECT 0.560 1.550 0.890 2.220 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.545 3.350 2.125 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 13.920 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 10.365 1.435 13.900 1.575 ;
        RECT 0.020 1.105 2.110 1.110 ;
        RECT 5.795 1.105 7.085 1.435 ;
        RECT 9.035 1.105 13.900 1.435 ;
        RECT 0.020 0.215 13.900 1.105 ;
        RECT -0.130 -0.215 14.050 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 13.920 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 14.250 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 13.920 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 13.920 3.815 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.596250 ;
    PORT
      LAYER li1 ;
        RECT 10.455 2.195 10.890 3.735 ;
        RECT 10.685 1.465 10.890 2.195 ;
        RECT 10.455 0.675 10.890 1.465 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.626250 ;
    PORT
      LAYER li1 ;
        RECT 13.460 2.175 13.810 3.755 ;
        RECT 13.480 0.675 13.810 2.175 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 13.920 4.155 ;
        RECT 0.110 1.370 0.380 3.230 ;
        RECT 0.570 2.400 1.160 3.705 ;
        RECT 1.340 3.410 2.290 3.580 ;
        RECT 1.340 1.870 1.510 3.410 ;
        RECT 1.690 2.400 1.940 3.230 ;
        RECT 1.215 1.370 1.545 1.870 ;
        RECT 0.110 1.200 1.545 1.370 ;
        RECT 1.750 1.365 1.940 2.400 ;
        RECT 2.120 2.475 2.290 3.410 ;
        RECT 2.470 2.655 3.000 3.705 ;
        RECT 3.180 3.335 5.085 3.505 ;
        RECT 3.180 2.475 3.350 3.335 ;
        RECT 2.120 2.305 3.350 2.475 ;
        RECT 3.530 2.655 3.770 3.155 ;
        RECT 0.110 0.540 0.440 1.200 ;
        RECT 1.750 1.195 3.340 1.365 ;
        RECT 0.620 0.365 1.570 1.020 ;
        RECT 1.750 0.520 1.920 1.195 ;
        RECT 2.100 0.365 2.990 1.015 ;
        RECT 3.170 0.435 3.340 1.195 ;
        RECT 3.530 0.935 3.700 2.655 ;
        RECT 3.950 1.785 4.120 3.335 ;
        RECT 3.880 1.115 4.120 1.785 ;
        RECT 4.300 2.075 4.550 3.155 ;
        RECT 4.755 2.805 5.085 3.335 ;
        RECT 5.265 2.985 6.215 3.715 ;
        RECT 6.395 3.635 8.245 3.805 ;
        RECT 6.395 2.805 6.565 3.635 ;
        RECT 4.755 2.635 6.565 2.805 ;
        RECT 4.755 2.255 5.085 2.635 ;
        RECT 6.745 2.455 6.915 3.455 ;
        RECT 5.435 2.285 6.915 2.455 ;
        RECT 5.435 2.255 5.765 2.285 ;
        RECT 6.210 2.075 6.540 2.105 ;
        RECT 4.300 1.905 6.540 2.075 ;
        RECT 4.300 1.015 4.470 1.905 ;
        RECT 4.650 1.415 4.980 1.725 ;
        RECT 6.210 1.595 6.540 1.905 ;
        RECT 4.650 1.245 6.485 1.415 ;
        RECT 6.745 1.325 6.915 2.285 ;
        RECT 7.095 2.495 7.265 3.635 ;
        RECT 7.445 2.675 7.795 3.455 ;
        RECT 7.095 2.205 7.425 2.495 ;
        RECT 4.650 1.195 4.980 1.245 ;
        RECT 3.520 0.615 3.850 0.935 ;
        RECT 4.300 0.615 4.630 1.015 ;
        RECT 4.810 0.435 4.980 1.195 ;
        RECT 3.170 0.265 4.980 0.435 ;
        RECT 5.185 0.365 6.135 1.065 ;
        RECT 6.315 0.435 6.485 1.245 ;
        RECT 6.665 0.615 6.995 1.325 ;
        RECT 7.175 1.195 7.445 1.865 ;
        RECT 7.175 0.435 7.345 1.195 ;
        RECT 7.625 1.015 7.795 2.675 ;
        RECT 7.975 1.105 8.245 3.635 ;
        RECT 8.505 2.675 9.455 3.715 ;
        RECT 8.425 2.325 9.725 2.495 ;
        RECT 7.540 0.685 7.795 1.015 ;
        RECT 8.425 0.685 8.595 2.325 ;
        RECT 8.775 1.675 9.105 2.145 ;
        RECT 9.395 1.855 9.725 2.325 ;
        RECT 9.905 1.975 10.235 3.715 ;
        RECT 11.070 2.195 11.605 3.735 ;
        RECT 11.785 2.195 12.115 2.985 ;
        RECT 11.805 1.995 12.115 2.195 ;
        RECT 12.295 2.175 13.245 3.755 ;
        RECT 9.905 1.675 10.505 1.975 ;
        RECT 8.775 1.645 10.505 1.675 ;
        RECT 11.805 1.665 13.300 1.995 ;
        RECT 8.775 1.505 10.235 1.645 ;
        RECT 7.540 0.515 8.595 0.685 ;
        RECT 6.315 0.265 7.345 0.435 ;
        RECT 8.775 0.365 9.725 1.325 ;
        RECT 9.905 0.535 10.235 1.505 ;
        RECT 11.070 0.365 11.625 1.485 ;
        RECT 11.805 1.005 12.135 1.665 ;
        RECT 12.315 0.365 13.265 1.485 ;
        RECT 0.000 -0.085 13.920 0.085 ;
  END
END sky130_fd_sc_hvl__dfxbp_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__dfxtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__dfxtp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.000 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.585000 ;
    PORT
      LAYER li1 ;
        RECT 0.540 1.905 0.870 2.575 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER li1 ;
        RECT 1.595 1.555 2.470 1.750 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 12.000 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 10.670 1.445 11.980 1.585 ;
        RECT 0.020 1.115 2.130 1.185 ;
        RECT 5.765 1.115 7.175 1.445 ;
        RECT 9.310 1.115 11.980 1.445 ;
        RECT 0.020 0.215 11.980 1.115 ;
        RECT -0.130 -0.215 12.130 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 12.000 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 12.330 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 12.000 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 12.000 3.815 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.596250 ;
    PORT
      LAYER li1 ;
        RECT 11.560 2.185 11.890 3.735 ;
        RECT 11.640 0.685 11.890 2.185 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 12.000 4.155 ;
        RECT 0.110 1.725 0.360 3.565 ;
        RECT 0.540 2.755 1.490 3.705 ;
        RECT 1.670 2.615 2.000 3.565 ;
        RECT 2.220 2.795 2.470 3.705 ;
        RECT 5.070 3.485 6.020 3.735 ;
        RECT 2.650 3.305 3.680 3.475 ;
        RECT 2.650 2.615 2.820 3.305 ;
        RECT 3.510 3.135 7.655 3.305 ;
        RECT 1.670 2.445 2.820 2.615 ;
        RECT 3.000 2.280 3.330 3.125 ;
        RECT 3.510 2.460 3.840 3.135 ;
        RECT 4.055 2.675 4.385 2.955 ;
        RECT 6.470 2.755 7.305 2.955 ;
        RECT 1.165 1.930 2.820 2.225 ;
        RECT 3.000 2.110 4.035 2.280 ;
        RECT 1.165 1.725 1.415 1.930 ;
        RECT 2.650 1.760 3.685 1.930 ;
        RECT 0.110 1.555 1.415 1.725 ;
        RECT 0.110 0.595 0.380 1.555 ;
        RECT 1.690 1.205 3.115 1.375 ;
        RECT 3.430 1.205 3.685 1.760 ;
        RECT 0.560 0.365 1.510 1.095 ;
        RECT 1.690 0.595 2.020 1.205 ;
        RECT 2.200 0.365 2.765 1.025 ;
        RECT 2.945 0.435 3.115 1.205 ;
        RECT 3.865 1.025 4.035 2.110 ;
        RECT 3.295 0.615 4.035 1.025 ;
        RECT 4.215 1.695 4.385 2.675 ;
        RECT 4.565 2.385 6.955 2.555 ;
        RECT 4.565 1.885 4.890 2.385 ;
        RECT 6.705 2.225 6.955 2.385 ;
        RECT 5.435 2.045 5.765 2.205 ;
        RECT 7.135 2.045 7.305 2.755 ;
        RECT 5.435 1.875 7.305 2.045 ;
        RECT 7.485 2.515 7.655 3.135 ;
        RECT 7.835 2.865 8.085 3.735 ;
        RECT 7.835 2.695 8.600 2.865 ;
        RECT 8.815 2.695 9.765 3.735 ;
        RECT 7.485 2.225 8.250 2.515 ;
        RECT 8.430 2.445 8.600 2.695 ;
        RECT 8.430 2.275 10.035 2.445 ;
        RECT 4.215 1.525 6.345 1.695 ;
        RECT 4.215 0.615 4.545 1.525 ;
        RECT 4.725 1.175 6.555 1.345 ;
        RECT 4.725 0.435 5.055 1.175 ;
        RECT 2.945 0.265 5.055 0.435 ;
        RECT 5.255 0.365 6.205 0.995 ;
        RECT 6.385 0.435 6.555 1.175 ;
        RECT 6.735 0.615 7.065 1.875 ;
        RECT 7.485 1.445 7.655 2.225 ;
        RECT 7.280 1.125 7.655 1.445 ;
        RECT 7.280 0.435 7.450 1.125 ;
        RECT 8.430 1.025 8.600 2.275 ;
        RECT 9.000 1.595 9.330 2.015 ;
        RECT 9.705 1.775 10.035 2.275 ;
        RECT 10.215 2.005 10.545 3.735 ;
        RECT 10.725 2.195 11.315 3.735 ;
        RECT 10.215 1.675 11.460 2.005 ;
        RECT 10.215 1.595 10.510 1.675 ;
        RECT 9.000 1.425 10.510 1.595 ;
        RECT 7.835 0.945 8.600 1.025 ;
        RECT 7.630 0.855 8.600 0.945 ;
        RECT 7.630 0.525 8.005 0.855 ;
        RECT 6.385 0.265 7.450 0.435 ;
        RECT 8.780 0.365 9.730 1.245 ;
        RECT 10.180 0.525 10.510 1.425 ;
        RECT 10.690 0.365 11.280 1.495 ;
        RECT 0.000 -0.085 12.000 0.085 ;
  END
END sky130_fd_sc_hvl__dfxtp_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__diode_2
  CLASS CORE ANTENNACELL ;
  FOREIGN sky130_fd_sc_hvl__diode_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.960 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN DIODE
    DIRECTION INPUT ;
    ANTENNADIFFAREA 0.607200 ;
    PORT
      LAYER li1 ;
        RECT 0.105 0.515 0.855 3.280 ;
    END
  END DIODE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 0.960 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.020 0.215 0.940 1.585 ;
        RECT -0.130 -0.215 1.090 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 0.960 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 1.290 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 0.960 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 0.960 3.815 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 0.960 4.155 ;
        RECT 0.000 -0.085 0.960 0.085 ;
  END
END sky130_fd_sc_hvl__diode_2

#--------EOF---------

MACRO sky130_fd_sc_hvl__dlclkp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__dlclkp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.080 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.170000 ;
    PORT
      LAYER li1 ;
        RECT 8.235 3.125 8.600 3.445 ;
        RECT 8.350 2.025 8.600 3.125 ;
        RECT 3.360 1.465 3.690 1.975 ;
        RECT 8.350 1.725 8.680 2.025 ;
    END
  END CLK
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.585000 ;
    PORT
      LAYER li1 ;
        RECT 0.610 1.385 0.940 2.200 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 10.080 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 8.680 1.405 9.970 1.415 ;
        RECT 7.060 1.345 9.970 1.405 ;
        RECT 0.020 1.210 2.090 1.345 ;
        RECT 4.240 1.210 9.970 1.345 ;
        RECT 0.020 0.215 9.970 1.210 ;
        RECT -0.130 -0.215 10.210 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 10.080 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 10.410 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 10.080 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 10.080 3.815 ;
    END
  END VPWR
  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.596250 ;
    PORT
      LAYER li1 ;
        RECT 9.630 1.895 9.995 3.735 ;
        RECT 9.725 1.215 9.995 1.895 ;
        RECT 9.630 0.515 9.995 1.215 ;
    END
  END GCLK
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 10.080 4.155 ;
        RECT 0.110 3.555 3.330 3.815 ;
        RECT 5.685 3.615 9.460 3.815 ;
        RECT 0.110 3.445 1.025 3.555 ;
        RECT 2.665 3.445 3.330 3.555 ;
        RECT 0.110 2.200 0.440 3.445 ;
        RECT 1.195 3.165 2.495 3.385 ;
        RECT 1.670 1.885 2.000 2.995 ;
        RECT 2.275 2.315 2.495 3.165 ;
        RECT 3.000 2.485 3.330 3.445 ;
        RECT 3.520 3.385 5.515 3.555 ;
        RECT 5.685 3.445 8.065 3.615 ;
        RECT 8.770 3.445 9.460 3.615 ;
        RECT 3.520 2.315 3.690 3.385 ;
        RECT 2.275 2.145 3.690 2.315 ;
        RECT 3.860 3.005 5.175 3.215 ;
        RECT 1.595 1.555 2.105 1.885 ;
        RECT 0.140 0.625 0.470 1.170 ;
        RECT 1.670 0.840 2.000 1.555 ;
        RECT 2.275 1.080 2.470 2.145 ;
        RECT 2.220 0.705 2.470 1.080 ;
        RECT 2.640 1.295 2.970 1.965 ;
        RECT 3.860 1.295 4.070 3.005 ;
        RECT 2.640 1.125 4.070 1.295 ;
        RECT 0.140 0.365 0.765 0.625 ;
        RECT 1.155 0.535 1.865 0.670 ;
        RECT 2.640 0.535 2.810 1.125 ;
        RECT 1.155 0.365 2.810 0.535 ;
        RECT 2.980 0.625 3.330 0.955 ;
        RECT 3.820 0.705 4.070 1.125 ;
        RECT 4.375 2.330 4.660 2.660 ;
        RECT 5.345 2.595 5.515 3.385 ;
        RECT 5.135 2.425 5.515 2.595 ;
        RECT 4.375 1.365 4.545 2.330 ;
        RECT 5.135 1.945 5.305 2.425 ;
        RECT 5.820 2.330 6.150 3.445 ;
        RECT 6.660 2.085 6.930 2.660 ;
        RECT 7.150 2.225 7.480 3.445 ;
        RECT 4.715 1.615 5.305 1.945 ;
        RECT 5.515 1.875 6.930 2.085 ;
        RECT 5.515 1.535 5.845 1.875 ;
        RECT 6.660 1.825 6.930 1.875 ;
        RECT 7.455 1.825 7.785 2.055 ;
        RECT 6.125 1.365 6.490 1.655 ;
        RECT 4.375 1.195 6.490 1.365 ;
        RECT 2.980 0.535 3.650 0.625 ;
        RECT 4.375 0.535 4.660 1.195 ;
        RECT 5.820 0.625 6.150 1.025 ;
        RECT 2.980 0.255 3.925 0.535 ;
        RECT 4.095 0.255 4.660 0.535 ;
        RECT 4.830 0.255 6.150 0.625 ;
        RECT 6.320 0.670 6.490 1.195 ;
        RECT 6.660 1.615 7.785 1.825 ;
        RECT 6.660 0.840 6.930 1.615 ;
        RECT 7.455 1.385 7.785 1.615 ;
        RECT 7.955 1.555 8.180 2.955 ;
        RECT 8.770 2.195 9.100 3.445 ;
        RECT 8.945 1.555 9.555 1.725 ;
        RECT 7.955 1.385 9.555 1.555 ;
        RECT 7.955 1.215 8.180 1.385 ;
        RECT 7.150 0.885 8.180 1.215 ;
        RECT 6.320 0.355 6.910 0.670 ;
        RECT 8.770 0.625 9.100 1.215 ;
        RECT 7.080 0.255 9.460 0.625 ;
        RECT 0.000 -0.085 10.080 0.085 ;
  END
END sky130_fd_sc_hvl__dlclkp_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__dlrtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__dlrtp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.600 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.585000 ;
    PORT
      LAYER li1 ;
        RECT 0.570 1.930 0.900 2.600 ;
    END
  END D
  PIN GATE
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.585000 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.175 1.795 1.400 ;
    END
  END GATE
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.585000 ;
    PORT
      LAYER li1 ;
        RECT 7.515 1.780 7.845 1.855 ;
        RECT 7.515 0.810 8.120 1.780 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 9.600 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 8.250 1.085 9.580 1.415 ;
        RECT 0.030 0.215 9.580 1.085 ;
        RECT -0.130 -0.215 9.730 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 9.600 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 9.930 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 9.600 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 9.600 3.815 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.641250 ;
    PORT
      LAYER li1 ;
        RECT 8.735 2.175 9.475 3.755 ;
        RECT 9.140 0.495 9.475 2.175 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 9.600 4.155 ;
        RECT 0.140 1.750 0.390 3.610 ;
        RECT 0.570 2.780 1.520 3.705 ;
        RECT 1.700 2.195 2.030 3.610 ;
        RECT 2.290 2.545 2.620 3.245 ;
        RECT 2.800 2.725 3.750 3.705 ;
        RECT 4.560 2.895 4.890 3.245 ;
        RECT 4.560 2.725 5.525 2.895 ;
        RECT 2.290 2.375 4.785 2.545 ;
        RECT 4.615 2.295 4.785 2.375 ;
        RECT 1.700 2.025 4.435 2.195 ;
        RECT 1.625 1.750 3.655 1.845 ;
        RECT 0.140 1.675 3.655 1.750 ;
        RECT 0.140 1.580 1.795 1.675 ;
        RECT 3.835 1.605 4.435 2.025 ;
        RECT 4.615 1.965 5.175 2.295 ;
        RECT 0.140 0.495 0.390 1.580 ;
        RECT 3.835 1.495 4.005 1.605 ;
        RECT 1.975 1.325 4.005 1.495 ;
        RECT 4.615 1.395 4.785 1.965 ;
        RECT 1.975 0.995 2.145 1.325 ;
        RECT 4.185 1.225 4.785 1.395 ;
        RECT 5.355 1.345 5.525 2.725 ;
        RECT 5.705 2.255 6.655 3.705 ;
        RECT 6.960 2.205 7.390 3.005 ;
        RECT 7.570 2.385 8.520 3.755 ;
        RECT 6.960 2.075 8.470 2.205 ;
        RECT 5.810 2.035 8.470 2.075 ;
        RECT 5.810 1.905 7.130 2.035 ;
        RECT 5.810 1.525 6.140 1.905 ;
        RECT 6.450 1.345 6.780 1.725 ;
        RECT 4.185 1.145 4.495 1.225 ;
        RECT 0.570 0.365 1.520 0.995 ;
        RECT 1.700 0.495 2.145 0.995 ;
        RECT 2.370 0.975 4.495 1.145 ;
        RECT 4.965 1.175 6.780 1.345 ;
        RECT 4.965 0.995 5.135 1.175 ;
        RECT 6.960 0.995 7.130 1.905 ;
        RECT 8.300 1.995 8.470 2.035 ;
        RECT 8.300 1.665 8.630 1.995 ;
        RECT 2.370 0.495 2.620 0.975 ;
        RECT 2.800 0.365 3.750 0.795 ;
        RECT 4.675 0.495 5.135 0.995 ;
        RECT 5.545 0.365 6.495 0.995 ;
        RECT 6.755 0.495 7.130 0.995 ;
        RECT 8.300 0.365 8.890 1.325 ;
        RECT 0.000 -0.085 9.600 0.085 ;
  END
END sky130_fd_sc_hvl__dlrtp_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__dlxtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__dlxtp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.160 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.585000 ;
    PORT
      LAYER li1 ;
        RECT 2.525 1.795 3.100 2.465 ;
    END
  END D
  PIN GATE
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.585000 ;
    PORT
      LAYER li1 ;
        RECT 0.540 1.175 0.870 1.725 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 8.160 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 5.955 1.085 8.140 1.415 ;
        RECT 0.225 0.215 8.140 1.085 ;
        RECT -0.130 -0.215 8.290 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 8.160 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 8.490 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 8.160 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 8.160 3.815 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.626250 ;
    PORT
      LAYER li1 ;
        RECT 7.700 0.515 8.050 3.755 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 8.160 4.155 ;
        RECT 0.110 2.075 0.360 2.985 ;
        RECT 0.540 2.255 1.430 3.705 ;
        RECT 1.890 2.995 2.840 3.705 ;
        RECT 3.020 3.635 4.050 3.805 ;
        RECT 3.020 2.815 3.190 3.635 ;
        RECT 1.610 2.645 3.190 2.815 ;
        RECT 3.370 2.895 3.700 3.455 ;
        RECT 1.610 2.075 1.780 2.645 ;
        RECT 1.960 2.195 2.290 2.465 ;
        RECT 0.110 2.015 1.780 2.075 ;
        RECT 0.110 1.905 1.795 2.015 ;
        RECT 0.110 0.995 0.360 1.905 ;
        RECT 1.540 1.345 1.795 1.905 ;
        RECT 1.975 1.615 2.290 2.195 ;
        RECT 3.370 2.335 3.540 2.895 ;
        RECT 3.880 2.715 4.050 3.635 ;
        RECT 4.230 3.065 4.480 3.725 ;
        RECT 4.230 2.895 5.090 3.065 ;
        RECT 5.270 2.895 6.220 3.705 ;
        RECT 3.720 2.515 4.740 2.715 ;
        RECT 3.370 2.165 4.230 2.335 ;
        RECT 3.550 1.615 3.880 1.985 ;
        RECT 1.975 1.445 3.880 1.615 ;
        RECT 0.110 0.495 0.665 0.995 ;
        RECT 0.845 0.365 1.795 0.995 ;
        RECT 1.975 0.515 2.225 1.445 ;
        RECT 4.060 1.265 4.230 2.165 ;
        RECT 3.385 1.095 4.230 1.265 ;
        RECT 4.410 1.095 4.740 2.515 ;
        RECT 4.920 2.005 5.090 2.895 ;
        RECT 6.025 2.355 6.355 2.675 ;
        RECT 6.535 2.535 7.485 3.755 ;
        RECT 6.025 2.185 7.030 2.355 ;
        RECT 4.920 1.835 6.680 2.005 ;
        RECT 3.385 0.995 3.555 1.095 ;
        RECT 2.405 0.365 2.995 0.975 ;
        RECT 3.225 0.495 3.555 0.995 ;
        RECT 4.920 0.915 5.090 1.835 ;
        RECT 6.350 1.775 6.680 1.835 ;
        RECT 5.430 1.595 5.760 1.655 ;
        RECT 6.860 1.595 7.030 2.185 ;
        RECT 5.430 1.425 7.030 1.595 ;
        RECT 5.430 1.075 5.760 1.425 ;
        RECT 4.005 0.745 5.090 0.915 ;
        RECT 4.005 0.495 4.335 0.745 ;
        RECT 5.270 0.365 5.860 0.895 ;
        RECT 6.045 0.845 6.375 1.425 ;
        RECT 6.555 0.365 7.505 1.245 ;
        RECT 0.000 -0.085 8.160 0.085 ;
  END
END sky130_fd_sc_hvl__dlxtp_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__einvn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__einvn_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.125000 ;
    PORT
      LAYER li1 ;
        RECT 2.275 1.725 2.780 2.540 ;
        RECT 2.505 1.160 2.780 1.725 ;
    END
  END A
  PIN TE_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.335000 ;
    PORT
      LAYER li1 ;
        RECT 0.635 2.025 1.795 2.120 ;
        RECT 0.515 1.825 1.795 2.025 ;
    END
  END TE_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 3.360 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.020 0.215 3.310 1.415 ;
        RECT -0.130 -0.215 3.490 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 3.360 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 3.690 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 3.360 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 3.360 3.815 ;
    END
  END VPWR
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.641250 ;
    PORT
      LAYER li1 ;
        RECT 2.950 0.495 3.235 3.755 ;
    END
  END Z
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 3.360 4.155 ;
        RECT 0.090 2.300 0.535 3.025 ;
        RECT 0.740 2.710 2.770 3.755 ;
        RECT 0.740 2.300 2.105 2.710 ;
        RECT 0.090 2.195 0.455 2.300 ;
        RECT 0.090 1.645 0.345 2.195 ;
        RECT 0.090 1.425 2.065 1.645 ;
        RECT 0.090 0.910 0.440 1.425 ;
        RECT 0.610 0.900 2.335 1.245 ;
        RECT 0.610 0.740 2.770 0.900 ;
        RECT 0.440 0.365 2.770 0.740 ;
        RECT 0.000 -0.085 3.360 0.085 ;
  END
END sky130_fd_sc_hvl__einvn_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__einvp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__einvp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.125000 ;
    PORT
      LAYER li1 ;
        RECT 2.445 1.955 2.810 2.540 ;
        RECT 2.275 1.625 2.865 1.955 ;
        RECT 2.445 1.160 2.810 1.625 ;
    END
  END A
  PIN TE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.960000 ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.505 1.305 1.750 ;
    END
  END TE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 3.360 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.020 0.215 3.340 1.495 ;
        RECT -0.130 -0.215 3.490 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 3.360 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 3.690 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 3.360 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 3.360 3.815 ;
    END
  END VPWR
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.641250 ;
    PORT
      LAYER li1 ;
        RECT 2.980 2.125 3.235 3.755 ;
        RECT 3.035 1.455 3.235 2.125 ;
        RECT 2.980 0.575 3.235 1.455 ;
    END
  END Z
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 3.360 4.155 ;
        RECT 0.175 2.100 0.650 3.005 ;
        RECT 0.830 2.710 2.800 3.755 ;
        RECT 0.830 2.280 2.275 2.710 ;
        RECT 0.175 1.930 2.065 2.100 ;
        RECT 0.175 1.335 0.345 1.930 ;
        RECT 1.475 1.725 2.065 1.930 ;
        RECT 0.175 0.905 0.380 1.335 ;
        RECT 0.550 0.990 2.275 1.335 ;
        RECT 0.550 0.735 2.800 0.990 ;
        RECT 0.470 0.365 2.800 0.735 ;
        RECT 0.000 -0.085 3.360 0.085 ;
  END
END sky130_fd_sc_hvl__einvp_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__fill_1
  CLASS CORE SPACER ;
  FOREIGN sky130_fd_sc_hvl__fill_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.480 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 0.480 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.130 -0.215 0.610 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 0.480 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 0.810 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 0.480 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 0.480 3.815 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 0.480 4.155 ;
        RECT 0.000 -0.085 0.480 0.085 ;
  END
END sky130_fd_sc_hvl__fill_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__fill_2
  CLASS CORE SPACER ;
  FOREIGN sky130_fd_sc_hvl__fill_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.960 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 0.960 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.130 -0.215 1.090 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 0.960 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 1.290 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 0.960 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 0.960 3.815 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 0.960 4.155 ;
        RECT 0.000 -0.085 0.960 0.085 ;
  END
END sky130_fd_sc_hvl__fill_2

#--------EOF---------

MACRO sky130_fd_sc_hvl__fill_4
  CLASS CORE SPACER ;
  FOREIGN sky130_fd_sc_hvl__fill_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.920 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 1.920 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.130 -0.215 2.050 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 1.920 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 2.250 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 1.920 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 1.920 3.815 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 1.920 4.155 ;
        RECT 0.000 -0.085 1.920 0.085 ;
  END
END sky130_fd_sc_hvl__fill_4

#--------EOF---------

MACRO sky130_fd_sc_hvl__fill_8
  CLASS CORE SPACER ;
  FOREIGN sky130_fd_sc_hvl__fill_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.840 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 3.840 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.130 -0.215 3.970 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 3.840 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 4.170 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 3.840 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 3.840 3.815 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 3.840 4.155 ;
        RECT 0.000 -0.085 3.840 0.085 ;
  END
END sky130_fd_sc_hvl__fill_8

#--------EOF---------

MACRO sky130_fd_sc_hvl__inv_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__inv_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.440 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.125000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.550 0.835 1.935 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 1.440 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.090 0.215 1.420 1.415 ;
        RECT -0.130 -0.215 1.570 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 1.440 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 1.770 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 1.440 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 1.440 3.815 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.641250 ;
    PORT
      LAYER li1 ;
        RECT 0.960 2.175 1.345 3.755 ;
        RECT 1.015 0.495 1.345 2.175 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 1.440 4.155 ;
        RECT 0.090 2.175 0.680 3.755 ;
        RECT 0.090 0.365 0.680 1.325 ;
        RECT 0.000 -0.085 1.440 0.085 ;
  END
END sky130_fd_sc_hvl__inv_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__inv_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__inv_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.400 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.250000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.550 1.070 1.880 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 2.400 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.270 0.215 2.380 1.460 ;
        RECT -0.130 -0.215 2.530 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 2.400 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 2.730 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 2.400 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 2.400 3.815 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.630000 ;
    PORT
      LAYER li1 ;
        RECT 1.240 1.780 1.490 3.755 ;
        RECT 1.240 1.610 1.795 1.780 ;
        RECT 1.565 1.370 1.795 1.610 ;
        RECT 1.200 0.540 1.795 1.370 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 2.400 4.155 ;
        RECT 0.110 2.175 1.060 3.755 ;
        RECT 1.680 2.175 2.270 3.755 ;
        RECT 0.090 0.365 1.020 1.370 ;
        RECT 1.980 0.365 2.310 1.370 ;
        RECT 0.000 -0.085 2.400 0.085 ;
  END
END sky130_fd_sc_hvl__inv_2

#--------EOF---------

MACRO sky130_fd_sc_hvl__inv_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__inv_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.840 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.500000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.580 2.835 1.750 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 3.840 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150 0.215 3.820 1.415 ;
        RECT -0.130 -0.215 3.970 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 3.840 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 4.170 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 3.840 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 3.840 3.815 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.260000 ;
    PORT
      LAYER li1 ;
        RECT 1.040 2.100 1.370 3.755 ;
        RECT 2.680 2.100 2.930 3.755 ;
        RECT 1.040 1.930 3.715 2.100 ;
        RECT 3.015 1.550 3.715 1.930 ;
        RECT 3.015 1.400 3.185 1.550 ;
        RECT 1.040 1.230 3.185 1.400 ;
        RECT 1.040 0.495 1.290 1.230 ;
        RECT 2.600 0.495 3.185 1.230 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 3.840 4.155 ;
        RECT 0.090 2.175 0.680 3.755 ;
        RECT 1.550 2.280 2.500 3.755 ;
        RECT 3.120 2.280 3.710 3.755 ;
        RECT 0.090 0.365 0.680 1.325 ;
        RECT 1.470 0.365 2.420 1.050 ;
        RECT 3.380 0.365 3.710 1.325 ;
        RECT 0.000 -0.085 3.840 0.085 ;
  END
END sky130_fd_sc_hvl__inv_4

#--------EOF---------

MACRO sky130_fd_sc_hvl__inv_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__inv_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.200 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 9.000000 ;
    PORT
      LAYER li1 ;
        RECT 0.310 1.580 6.760 1.815 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 7.200 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.265 0.215 7.165 1.585 ;
        RECT -0.130 -0.215 7.330 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 7.200 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 7.530 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 7.200 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 7.200 3.815 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.520000 ;
    PORT
      LAYER li1 ;
        RECT 1.275 2.205 1.605 3.445 ;
        RECT 2.835 2.205 3.165 3.445 ;
        RECT 4.395 2.205 4.725 3.445 ;
        RECT 5.955 2.205 6.285 3.445 ;
        RECT 1.275 2.035 7.110 2.205 ;
        RECT 1.195 1.395 6.225 1.400 ;
        RECT 6.940 1.395 7.110 2.035 ;
        RECT 1.195 1.230 7.110 1.395 ;
        RECT 1.195 0.730 1.405 1.230 ;
        RECT 2.755 0.730 2.965 1.230 ;
        RECT 4.315 0.730 4.525 1.230 ;
        RECT 5.915 1.225 7.110 1.230 ;
        RECT 5.915 0.730 6.565 1.225 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 7.200 4.155 ;
        RECT 0.095 3.625 7.025 3.795 ;
        RECT 0.095 2.445 0.985 3.625 ;
        RECT 1.775 2.385 2.665 3.625 ;
        RECT 3.335 2.385 4.225 3.625 ;
        RECT 4.895 2.385 5.785 3.625 ;
        RECT 6.455 2.385 7.025 3.625 ;
        RECT 0.095 0.550 0.985 1.385 ;
        RECT 1.575 0.550 2.585 1.045 ;
        RECT 3.135 0.550 4.145 1.045 ;
        RECT 4.695 0.550 5.745 1.045 ;
        RECT 6.735 0.550 7.105 1.045 ;
        RECT 0.095 0.380 7.105 0.550 ;
        RECT 0.000 -0.085 7.200 0.085 ;
  END
END sky130_fd_sc_hvl__inv_8

#--------EOF---------

MACRO sky130_fd_sc_hvl__inv_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__inv_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.440 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 18.000000 ;
    PORT
      LAYER met1 ;
        RECT 1.535 1.750 2.185 1.780 ;
        RECT 3.085 1.750 3.735 1.780 ;
        RECT 4.645 1.750 5.295 1.780 ;
        RECT 6.205 1.750 6.855 1.780 ;
        RECT 7.765 1.750 8.415 1.780 ;
        RECT 9.325 1.750 9.975 1.780 ;
        RECT 10.885 1.750 11.535 1.780 ;
        RECT 1.535 1.580 11.535 1.750 ;
        RECT 1.535 1.550 2.185 1.580 ;
        RECT 3.085 1.550 3.735 1.580 ;
        RECT 4.645 1.550 5.295 1.580 ;
        RECT 6.205 1.550 6.855 1.580 ;
        RECT 7.765 1.550 8.415 1.580 ;
        RECT 9.325 1.550 9.975 1.580 ;
        RECT 10.885 1.550 11.535 1.580 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 13.440 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.030 0.215 13.025 1.585 ;
        RECT -0.130 -0.215 13.570 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 13.440 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 13.770 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 13.440 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 13.440 3.815 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 5.040000 ;
    PORT
      LAYER met1 ;
        RECT 0.925 2.490 1.215 2.520 ;
        RECT 2.485 2.490 2.775 2.520 ;
        RECT 4.045 2.490 4.335 2.520 ;
        RECT 5.605 2.490 5.895 2.520 ;
        RECT 7.165 2.490 7.455 2.520 ;
        RECT 8.725 2.490 9.015 2.520 ;
        RECT 10.285 2.490 10.575 2.520 ;
        RECT 11.845 2.490 12.135 2.520 ;
        RECT 0.925 2.320 12.135 2.490 ;
        RECT 0.925 2.290 1.215 2.320 ;
        RECT 2.485 2.290 2.775 2.320 ;
        RECT 4.045 2.290 4.335 2.320 ;
        RECT 5.605 2.290 5.895 2.320 ;
        RECT 7.165 2.290 7.455 2.320 ;
        RECT 8.725 2.290 9.015 2.320 ;
        RECT 10.285 2.290 10.575 2.320 ;
        RECT 11.845 2.290 12.135 2.320 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 13.440 4.155 ;
        RECT 0.125 2.175 0.655 3.755 ;
        RECT 0.095 0.375 0.630 1.475 ;
        RECT 0.900 0.795 1.230 3.755 ;
        RECT 1.400 2.175 2.290 3.755 ;
        RECT 1.400 1.565 2.290 1.895 ;
        RECT 1.400 0.375 2.290 1.395 ;
        RECT 2.460 0.795 2.790 3.755 ;
        RECT 2.960 2.175 3.850 3.755 ;
        RECT 2.960 1.565 3.850 1.895 ;
        RECT 2.960 0.375 3.850 1.395 ;
        RECT 4.020 0.795 4.350 3.755 ;
        RECT 4.520 2.175 5.410 3.755 ;
        RECT 4.520 1.565 5.410 1.895 ;
        RECT 4.520 0.375 5.410 1.395 ;
        RECT 5.580 0.795 5.910 3.755 ;
        RECT 6.080 2.175 6.970 3.755 ;
        RECT 6.080 1.565 6.970 1.895 ;
        RECT 6.080 0.375 6.970 1.395 ;
        RECT 7.140 0.795 7.470 3.755 ;
        RECT 7.640 2.175 8.530 3.755 ;
        RECT 7.640 1.565 8.530 1.895 ;
        RECT 7.640 0.375 8.530 1.395 ;
        RECT 8.700 0.795 9.030 3.755 ;
        RECT 9.200 2.175 10.090 3.755 ;
        RECT 9.200 1.565 10.090 1.895 ;
        RECT 9.200 0.375 10.090 1.395 ;
        RECT 10.260 0.795 10.590 3.755 ;
        RECT 10.760 2.175 11.650 3.755 ;
        RECT 10.760 1.565 11.650 1.895 ;
        RECT 10.760 0.375 11.650 1.395 ;
        RECT 11.820 0.795 12.150 3.755 ;
        RECT 12.320 2.175 12.935 3.675 ;
        RECT 12.320 0.375 12.935 1.395 ;
        RECT 0.000 -0.085 13.440 0.085 ;
  END
END sky130_fd_sc_hvl__inv_16

#--------EOF---------

MACRO sky130_fd_sc_hvl__lsbufhv2hv_hl_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__lsbufhv2hv_hl_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.640 BY 8.140 ;
  SYMMETRY X Y ;
  SITE unithvdbl ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.585000 ;
    PORT
      LAYER li1 ;
        RECT 4.355 1.775 4.685 2.900 ;
    END
  END A
  PIN LOWHVPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 2.800 1.885 5.425 5.135 ;
      LAYER met1 ;
        RECT 0.070 3.020 8.570 3.305 ;
    END
  END LOWHVPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 7.515 8.640 7.885 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 8.640 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.915 1.085 4.225 1.415 ;
        RECT 2.915 0.215 5.225 1.085 ;
        RECT -0.130 -0.215 8.770 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 8.640 0.115 ;
    END
    PORT
      LAYER pwell ;
        RECT -0.130 7.925 8.770 8.355 ;
      LAYER met1 ;
        RECT 0.000 8.025 8.640 8.255 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.000 8.055 8.640 8.225 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.000 -0.085 8.640 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 0.800 6.255 ;
        RECT 7.425 1.885 8.970 6.255 ;
      LAYER met1 ;
        RECT 0.000 3.955 8.640 4.185 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.425 3.985 8.640 4.155 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.000 3.985 0.800 4.155 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 8.640 3.815 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 4.325 8.640 4.695 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.626250 ;
    PORT
      LAYER li1 ;
        RECT 2.995 0.495 3.395 4.065 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 3.130 4.265 5.095 4.835 ;
        RECT 3.565 2.485 4.185 4.265 ;
        RECT 3.565 1.605 3.895 2.065 ;
        RECT 4.865 1.605 5.115 3.315 ;
        RECT 3.565 1.435 5.115 1.605 ;
        RECT 3.565 0.365 4.515 1.265 ;
        RECT 4.865 0.495 5.115 1.435 ;
  END
END sky130_fd_sc_hvl__lsbufhv2hv_hl_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__lsbufhv2hv_lh_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__lsbufhv2hv_lh_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.560 BY 8.140 ;
  SYMMETRY X Y ;
  SITE unithvdbl ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.750000 ;
    PORT
      LAYER li1 ;
        RECT 2.495 1.530 2.805 2.200 ;
    END
  END A
  PIN LOWHVPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 2.800 2.015 5.270 4.315 ;
      LAYER met1 ;
        RECT 0.070 3.020 10.490 3.305 ;
    END
  END LOWHVPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 7.515 10.560 7.885 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 10.560 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 5.870 1.585 9.500 2.165 ;
        RECT 3.000 0.215 9.500 1.585 ;
        RECT -0.130 -0.215 10.690 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 10.560 0.115 ;
    END
    PORT
      LAYER pwell ;
        RECT -0.130 7.925 10.690 8.355 ;
        RECT 3.340 5.975 6.970 7.925 ;
        RECT 9.250 6.725 10.540 7.925 ;
      LAYER met1 ;
        RECT 0.000 8.025 10.560 8.255 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.000 8.055 10.560 8.225 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.000 -0.085 10.560 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 0.800 6.255 ;
        RECT 7.270 2.465 10.890 6.255 ;
        RECT 9.800 1.885 10.890 2.465 ;
      LAYER met1 ;
        RECT 0.000 3.955 10.560 4.185 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.715 3.985 10.560 4.155 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.000 3.985 0.800 4.155 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 4.325 10.560 4.695 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 10.560 3.815 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.596250 ;
    PORT
      LAYER li1 ;
        RECT 10.120 4.405 10.450 7.625 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 3.300 7.715 7.010 7.885 ;
        RECT 3.300 6.085 3.890 7.715 ;
        RECT 4.210 5.995 4.540 7.545 ;
        RECT 4.860 6.165 5.450 7.715 ;
        RECT 5.770 5.995 6.100 7.545 ;
        RECT 6.420 6.165 7.010 7.715 ;
        RECT 9.210 6.835 9.800 7.745 ;
        RECT 4.210 5.665 7.930 5.995 ;
        RECT 3.090 5.165 5.660 5.495 ;
        RECT 3.090 1.995 3.420 5.165 ;
        RECT 3.590 3.355 4.780 4.025 ;
        RECT 7.600 3.935 7.930 5.665 ;
        RECT 8.635 5.535 8.965 6.555 ;
        RECT 8.215 5.205 8.965 5.535 ;
        RECT 7.375 3.605 8.045 3.935 ;
        RECT 3.740 2.325 4.330 3.355 ;
        RECT 7.600 3.125 7.930 3.435 ;
        RECT 8.215 3.125 8.545 5.205 ;
        RECT 9.210 4.800 9.800 5.945 ;
        RECT 8.790 4.405 9.800 4.800 ;
        RECT 4.650 2.475 4.980 3.115 ;
        RECT 7.600 2.795 8.545 3.125 ;
        RECT 8.940 2.795 9.530 3.705 ;
        RECT 8.215 2.475 8.545 2.795 ;
        RECT 4.650 2.165 6.570 2.475 ;
        RECT 5.330 2.145 6.570 2.165 ;
        RECT 6.740 2.145 8.630 2.475 ;
        RECT 3.090 1.745 4.845 1.995 ;
        RECT 3.090 0.685 3.420 1.745 ;
        RECT 5.330 1.475 5.660 2.145 ;
        RECT 3.740 0.425 4.330 1.475 ;
        RECT 4.650 1.145 5.660 1.475 ;
        RECT 4.650 0.685 4.980 1.145 ;
        RECT 5.830 0.425 6.420 1.975 ;
        RECT 6.740 0.595 7.070 2.145 ;
        RECT 7.390 0.425 7.980 1.975 ;
        RECT 8.300 0.595 8.630 2.145 ;
        RECT 8.950 0.425 9.540 1.975 ;
        RECT 3.740 0.255 9.540 0.425 ;
  END
END sky130_fd_sc_hvl__lsbufhv2hv_lh_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__lsbufhv2lv_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__lsbufhv2lv_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.160 BY 8.140 ;
  SYMMETRY X Y ;
  SITE unithvdbl ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER li1 ;
        RECT 0.630 4.870 1.300 5.200 ;
    END
  END A
  PIN LVPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 3.530 1.925 5.000 5.575 ;
      LAYER met1 ;
        RECT 0.070 3.020 8.090 3.305 ;
    END
  END LVPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 7.515 8.160 7.885 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 8.160 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.830 1.625 3.120 4.055 ;
        RECT 1.830 1.585 4.520 1.625 ;
        RECT 0.020 0.215 4.520 1.585 ;
        RECT -0.130 -0.215 8.290 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 8.160 0.115 ;
    END
    PORT
      LAYER pwell ;
        RECT -0.130 7.925 8.290 8.355 ;
        RECT 0.020 6.555 3.900 7.925 ;
        RECT 1.830 5.505 3.120 6.555 ;
      LAYER met1 ;
        RECT 0.000 8.025 8.160 8.255 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.000 8.055 8.160 8.225 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.000 -0.085 8.160 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 1.530 6.255 ;
        RECT 7.000 1.885 8.490 6.255 ;
      LAYER met1 ;
        RECT 0.000 3.955 8.160 4.185 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.275 3.985 8.160 4.155 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.000 3.985 0.885 4.155 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 8.160 3.815 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 4.325 8.160 4.695 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.492900 ;
    PORT
      LAYER li1 ;
        RECT 3.485 0.735 3.960 3.245 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.170 6.575 0.420 7.060 ;
        RECT 0.895 6.745 1.485 7.745 ;
        RECT 0.170 6.220 1.750 6.575 ;
        RECT 0.130 4.695 0.460 5.880 ;
        RECT 0.950 5.550 1.750 6.220 ;
        RECT 0.130 4.465 0.720 4.695 ;
        RECT 0.130 3.445 0.720 3.675 ;
        RECT 0.130 2.260 0.460 3.445 ;
        RECT 1.470 3.085 1.750 5.550 ;
        RECT 1.920 5.445 2.250 7.455 ;
        RECT 2.530 5.615 3.120 7.745 ;
        RECT 3.480 5.845 3.810 7.455 ;
        RECT 3.290 5.595 5.170 5.845 ;
        RECT 3.290 5.445 3.540 5.595 ;
        RECT 1.920 5.195 3.540 5.445 ;
        RECT 3.710 4.595 3.960 5.415 ;
        RECT 0.630 2.835 1.750 3.085 ;
        RECT 1.920 4.255 3.960 4.595 ;
        RECT 0.950 1.895 1.200 2.590 ;
        RECT 1.445 1.895 1.750 2.235 ;
        RECT 0.170 1.565 1.750 1.895 ;
        RECT 0.170 1.080 0.420 1.565 ;
        RECT 0.895 0.395 1.485 1.395 ;
        RECT 1.920 0.685 2.250 4.255 ;
        RECT 4.130 4.085 4.400 5.415 ;
        RECT 2.570 0.395 3.160 3.910 ;
        RECT 3.780 3.415 4.750 4.085 ;
        RECT 4.130 3.075 4.750 3.415 ;
        RECT 4.130 2.085 4.400 3.075 ;
        RECT 4.920 2.905 5.170 5.595 ;
        RECT 4.570 2.655 5.170 2.905 ;
        RECT 4.570 2.085 4.820 2.655 ;
        RECT 4.130 0.395 4.720 1.515 ;
  END
END sky130_fd_sc_hvl__lsbufhv2lv_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__lsbufhv2lv_simple_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__lsbufhv2lv_simple_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.640 BY 8.140 ;
  SYMMETRY X Y ;
  SITE unithvdbl ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.585000 ;
    PORT
      LAYER li1 ;
        RECT 4.355 1.465 4.685 3.260 ;
    END
  END A
  PIN LVPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 2.800 1.885 5.425 4.825 ;
      LAYER met1 ;
        RECT 0.070 3.020 8.570 3.305 ;
    END
  END LVPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 7.515 8.640 7.885 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 8.640 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.915 1.085 4.225 1.415 ;
        RECT 2.915 0.215 5.225 1.085 ;
        RECT -0.130 -0.215 8.770 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 8.640 0.115 ;
    END
    PORT
      LAYER pwell ;
        RECT -0.130 7.925 8.770 8.355 ;
      LAYER met1 ;
        RECT 0.000 8.025 8.640 8.255 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.000 8.055 8.640 8.225 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.000 -0.085 8.640 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 0.800 6.255 ;
        RECT 7.425 1.885 8.970 6.255 ;
      LAYER met1 ;
        RECT 0.000 3.955 8.640 4.185 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.425 3.985 8.640 4.155 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.000 3.985 0.800 4.155 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 8.640 3.815 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 4.325 8.640 4.695 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.626250 ;
    PORT
      LAYER li1 ;
        RECT 2.995 2.175 3.440 3.755 ;
        RECT 2.995 0.495 3.255 2.175 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 3.130 3.955 5.095 4.525 ;
        RECT 3.620 2.175 4.175 3.955 ;
        RECT 3.565 1.285 3.895 1.745 ;
        RECT 4.865 1.285 5.115 3.005 ;
        RECT 3.565 1.115 5.115 1.285 ;
        RECT 3.435 0.365 4.685 0.935 ;
        RECT 4.865 0.495 5.115 1.115 ;
  END
END sky130_fd_sc_hvl__lsbufhv2lv_simple_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__lsbuflv2hv_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__lsbuflv2hv_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.560 BY 8.140 ;
  SYMMETRY X Y ;
  SITE unithvdbl ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER li1 ;
        RECT 2.495 1.530 2.805 2.200 ;
    END
  END A
  PIN LVPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 2.800 2.015 4.335 4.325 ;
      LAYER met1 ;
        RECT 0.070 3.020 10.490 3.305 ;
    END
  END LVPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 7.515 10.560 7.885 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 10.560 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 5.090 1.725 9.500 2.165 ;
        RECT 2.855 0.215 9.500 1.725 ;
        RECT -0.130 -0.215 10.690 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 10.560 0.115 ;
    END
    PORT
      LAYER pwell ;
        RECT -0.130 7.925 10.690 8.355 ;
        RECT 1.625 5.975 6.035 7.925 ;
        RECT 8.425 6.725 10.540 7.925 ;
      LAYER met1 ;
        RECT 0.000 8.025 10.560 8.255 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.000 8.055 10.560 8.225 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.000 -0.085 10.560 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 0.800 6.255 ;
        RECT 6.335 2.465 10.890 6.255 ;
        RECT 9.800 1.885 10.890 2.465 ;
      LAYER met1 ;
        RECT 0.000 3.955 10.560 4.185 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.755 3.985 10.560 4.155 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.000 3.985 0.800 4.155 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 4.325 10.560 4.695 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 10.560 3.815 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.596250 ;
    PORT
      LAYER li1 ;
        RECT 10.120 6.725 10.450 7.625 ;
        RECT 10.210 6.055 10.450 6.725 ;
        RECT 10.120 4.405 10.450 6.055 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 1.585 7.715 5.295 7.885 ;
        RECT 1.585 6.085 2.175 7.715 ;
        RECT 2.495 5.995 2.825 7.545 ;
        RECT 3.145 6.165 3.735 7.715 ;
        RECT 4.055 5.995 4.385 7.545 ;
        RECT 4.705 6.165 5.295 7.715 ;
        RECT 5.615 5.995 5.945 7.625 ;
        RECT 8.515 6.555 8.845 7.625 ;
        RECT 9.210 6.835 9.800 7.745 ;
        RECT 7.660 5.995 7.990 6.555 ;
        RECT 2.495 5.665 7.990 5.995 ;
        RECT 2.885 3.055 3.175 5.495 ;
        RECT 3.345 3.225 4.115 4.200 ;
        RECT 3.435 3.075 4.115 3.225 ;
        RECT 6.185 3.465 6.515 5.665 ;
        RECT 7.660 5.205 7.990 5.665 ;
        RECT 8.515 6.225 10.040 6.555 ;
        RECT 6.685 4.470 7.495 4.800 ;
        RECT 7.165 3.805 7.495 4.470 ;
        RECT 7.755 4.405 8.345 4.800 ;
        RECT 8.515 4.405 8.845 6.225 ;
        RECT 9.210 4.405 9.800 5.945 ;
        RECT 6.185 3.135 6.995 3.465 ;
        RECT 2.885 2.765 3.265 3.055 ;
        RECT 2.975 1.995 3.265 2.765 ;
        RECT 3.435 2.165 3.705 3.075 ;
        RECT 3.875 2.475 4.185 2.905 ;
        RECT 6.665 2.795 6.995 3.135 ;
        RECT 7.165 3.395 7.835 3.805 ;
        RECT 7.165 2.475 7.495 3.395 ;
        RECT 8.005 2.795 8.595 3.705 ;
        RECT 3.875 2.165 5.790 2.475 ;
        RECT 4.480 2.145 5.790 2.165 ;
        RECT 5.960 2.145 9.410 2.475 ;
        RECT 2.975 1.745 4.310 1.995 ;
        RECT 2.975 0.735 3.265 1.745 ;
        RECT 4.480 1.575 4.810 2.145 ;
        RECT 3.435 0.565 3.705 1.575 ;
        RECT 3.875 1.245 4.810 1.575 ;
        RECT 3.875 0.735 4.185 1.245 ;
        RECT 3.095 0.335 4.045 0.565 ;
        RECT 5.050 0.425 5.640 1.975 ;
        RECT 5.960 0.595 6.290 2.145 ;
        RECT 6.610 0.425 7.200 1.975 ;
        RECT 7.520 0.595 7.850 2.145 ;
        RECT 8.170 0.425 8.760 1.975 ;
        RECT 9.080 0.515 9.410 2.145 ;
        RECT 5.050 0.255 8.760 0.425 ;
  END
END sky130_fd_sc_hvl__lsbuflv2hv_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__lsbuflv2hv_clkiso_hlkg_3
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__lsbuflv2hv_clkiso_hlkg_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 24.960 BY 8.140 ;
  SYMMETRY X Y ;
  SITE unithvdbl ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.558000 ;
    PORT
      LAYER li1 ;
        RECT 21.070 5.975 21.400 6.455 ;
    END
  END A
  PIN SLEEP_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.750000 ;
    PORT
      LAYER li1 ;
        RECT 14.315 5.545 14.985 5.875 ;
    END
  END SLEEP_B
  PIN LVPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 17.395 2.045 21.695 6.095 ;
      LAYER met1 ;
        RECT 0.070 3.020 24.890 3.305 ;
    END
  END LVPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 24.960 0.625 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 7.515 24.960 7.885 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.130 7.925 25.090 8.355 ;
        RECT 2.245 6.765 12.195 7.925 ;
        RECT 13.740 6.765 15.030 7.925 ;
        RECT 0.915 6.085 15.030 6.765 ;
        RECT 17.670 6.515 21.485 7.925 ;
      LAYER met1 ;
        RECT 0.000 8.025 24.960 8.255 ;
    END
    PORT
      LAYER pwell ;
        RECT 0.915 0.215 5.875 1.795 ;
        RECT 17.670 0.215 20.060 1.625 ;
        RECT -0.130 -0.215 25.090 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 24.960 0.115 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.000 8.055 24.960 8.225 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.000 -0.085 24.960 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 5.755 0.510 6.255 ;
        RECT -0.330 2.095 15.395 5.755 ;
        RECT -0.330 1.885 0.510 2.095 ;
        RECT 9.415 1.705 15.395 2.095 ;
      LAYER met1 ;
        RECT 0.000 3.955 24.960 4.185 ;
    END
    PORT
      LAYER li1 ;
        RECT 9.135 3.985 9.925 4.155 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.360 4.155 0.530 5.180 ;
        RECT 0.000 3.985 0.685 4.155 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 4.325 24.960 4.695 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 24.960 3.815 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.180000 ;
    PORT
      LAYER li1 ;
        RECT 1.060 2.140 1.280 5.115 ;
        RECT 2.620 2.140 2.840 5.115 ;
        RECT 1.060 1.920 2.840 2.140 ;
        RECT 1.060 0.645 1.280 1.920 ;
        RECT 2.620 0.645 2.840 1.920 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 1.060 7.570 14.885 7.800 ;
        RECT 1.060 7.180 1.280 7.570 ;
        RECT 2.360 7.205 2.580 7.570 ;
        RECT 1.060 6.850 1.810 7.180 ;
        RECT 1.060 6.195 1.280 6.850 ;
        RECT 1.840 5.975 2.060 6.525 ;
        RECT 2.360 6.195 2.585 7.205 ;
        RECT 3.570 5.975 3.790 7.205 ;
        RECT 4.750 6.195 4.970 7.570 ;
        RECT 5.930 5.975 6.150 7.205 ;
        RECT 7.110 6.195 7.330 7.570 ;
        RECT 8.290 5.975 8.510 7.205 ;
        RECT 9.470 6.195 9.690 7.570 ;
        RECT 10.650 5.975 10.870 7.205 ;
        RECT 11.830 6.195 12.050 7.570 ;
        RECT 12.555 5.975 12.775 6.525 ;
        RECT 13.335 6.195 13.555 7.570 ;
        RECT 1.840 5.755 6.520 5.975 ;
        RECT 1.835 4.625 2.065 5.115 ;
        RECT 3.395 4.625 3.625 5.115 ;
        RECT 1.655 4.395 2.245 4.625 ;
        RECT 3.215 4.395 3.805 4.625 ;
        RECT 1.835 2.405 2.065 4.395 ;
        RECT 3.395 2.405 3.625 4.395 ;
        RECT 3.950 2.195 4.170 3.755 ;
        RECT 4.725 3.515 5.310 3.755 ;
        RECT 4.725 2.405 4.955 3.515 ;
        RECT 3.010 2.140 4.170 2.195 ;
        RECT 5.510 2.140 5.730 3.755 ;
        RECT 6.300 2.515 6.520 5.755 ;
        RECT 7.860 5.755 12.775 5.975 ;
        RECT 13.885 5.755 14.105 6.865 ;
        RECT 14.665 6.195 14.885 7.570 ;
        RECT 17.780 7.515 21.375 7.745 ;
        RECT 17.780 6.915 18.110 7.515 ;
        RECT 18.290 6.745 18.460 7.345 ;
        RECT 18.690 6.915 19.020 7.515 ;
        RECT 19.200 6.745 19.450 7.345 ;
        RECT 17.790 6.575 19.450 6.745 ;
        RECT 19.620 6.625 19.950 7.515 ;
        RECT 20.185 6.625 20.435 7.515 ;
        RECT 20.615 6.625 20.945 7.345 ;
        RECT 21.125 6.625 21.375 7.515 ;
        RECT 17.790 5.855 18.020 6.575 ;
        RECT 20.615 6.405 20.900 6.625 ;
        RECT 18.265 6.185 20.900 6.405 ;
        RECT 18.265 5.975 19.940 6.185 ;
        RECT 7.860 5.235 8.080 5.755 ;
        RECT 13.090 5.425 14.105 5.755 ;
        RECT 7.345 4.905 8.080 5.235 ;
        RECT 7.075 3.065 7.305 4.345 ;
        RECT 7.075 2.835 7.435 3.065 ;
        RECT 7.860 2.835 8.080 4.905 ;
        RECT 10.210 5.035 13.550 5.255 ;
        RECT 10.210 3.745 10.430 5.035 ;
        RECT 10.025 3.515 10.615 3.745 ;
        RECT 7.205 2.655 7.435 2.835 ;
        RECT 6.300 2.185 6.995 2.515 ;
        RECT 7.205 2.425 7.805 2.655 ;
        RECT 3.010 1.920 5.730 2.140 ;
        RECT 3.010 1.865 4.170 1.920 ;
        RECT 1.835 0.485 2.065 1.655 ;
        RECT 3.395 0.485 3.625 1.655 ;
        RECT 3.950 0.645 4.170 1.865 ;
        RECT 4.725 0.485 4.955 1.655 ;
        RECT 5.510 0.645 5.730 1.920 ;
        RECT 7.575 1.805 7.805 2.425 ;
        RECT 10.210 2.015 10.430 3.515 ;
        RECT 10.990 1.805 11.210 4.725 ;
        RECT 11.770 3.745 11.990 5.035 ;
        RECT 11.585 3.515 12.175 3.745 ;
        RECT 11.770 2.015 11.990 3.515 ;
        RECT 12.550 1.805 12.770 4.725 ;
        RECT 13.330 3.745 13.550 5.035 ;
        RECT 13.885 4.265 14.105 5.425 ;
        RECT 17.160 5.805 18.020 5.855 ;
        RECT 20.170 5.805 20.420 5.935 ;
        RECT 17.160 5.635 19.465 5.805 ;
        RECT 14.655 4.625 14.885 5.055 ;
        RECT 14.295 4.395 14.885 4.625 ;
        RECT 14.655 4.265 14.885 4.395 ;
        RECT 13.145 3.515 13.735 3.745 ;
        RECT 13.330 2.015 13.550 3.515 ;
        RECT 7.575 1.585 12.770 1.805 ;
        RECT 13.965 1.565 14.295 2.285 ;
        RECT 17.160 2.165 17.380 5.635 ;
        RECT 17.785 4.605 18.035 5.465 ;
        RECT 18.235 4.775 18.565 5.635 ;
        RECT 18.765 4.605 18.935 5.465 ;
        RECT 19.135 4.775 19.465 5.635 ;
        RECT 19.665 4.605 20.420 5.805 ;
        RECT 20.615 4.775 20.900 6.185 ;
        RECT 21.070 4.605 21.400 5.805 ;
        RECT 17.785 4.435 21.400 4.605 ;
        RECT 19.665 4.235 20.420 4.435 ;
        RECT 17.795 3.905 20.420 4.235 ;
        RECT 19.665 3.705 20.420 3.905 ;
        RECT 17.815 3.535 20.420 3.705 ;
        RECT 17.815 2.335 18.065 3.535 ;
        RECT 18.265 2.505 18.595 3.365 ;
        RECT 18.795 2.675 18.965 3.535 ;
        RECT 19.165 2.505 19.495 3.365 ;
        RECT 19.695 3.020 20.420 3.535 ;
        RECT 19.695 2.675 19.945 3.020 ;
        RECT 18.265 2.335 19.940 2.505 ;
        RECT 17.160 1.735 19.465 2.165 ;
        RECT 19.710 1.565 19.940 2.335 ;
        RECT 13.965 1.395 19.940 1.565 ;
        RECT 13.965 1.345 18.530 1.395 ;
        RECT 17.780 0.625 18.110 1.175 ;
        RECT 18.280 0.795 18.530 1.345 ;
        RECT 18.710 0.625 19.040 1.225 ;
        RECT 19.270 0.795 19.440 1.395 ;
        RECT 19.620 0.625 19.950 1.225 ;
        RECT 1.835 0.255 2.425 0.485 ;
        RECT 3.035 0.255 3.625 0.485 ;
        RECT 4.545 0.255 5.135 0.485 ;
        RECT 17.780 0.395 19.950 0.625 ;
  END
END sky130_fd_sc_hvl__lsbuflv2hv_clkiso_hlkg_3

#--------EOF---------

MACRO sky130_fd_sc_hvl__lsbuflv2hv_isosrchvaon_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__lsbuflv2hv_isosrchvaon_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.920 BY 8.140 ;
  SYMMETRY X Y ;
  SITE unithvdbl ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER li1 ;
        RECT 9.205 1.685 9.895 2.015 ;
    END
  END A
  PIN SLEEP_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 7.125000 ;
    PORT
      LAYER li1 ;
        RECT 4.730 1.830 5.400 2.160 ;
    END
  END SLEEP_B
  PIN LVPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 8.890 2.045 10.710 6.095 ;
      LAYER met1 ;
        RECT 0.070 3.020 13.850 3.305 ;
    END
  END LVPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 13.920 0.625 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 7.515 13.920 7.885 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.130 7.925 14.050 8.355 ;
        RECT 0.810 6.335 4.440 7.925 ;
        RECT 9.095 6.515 10.145 7.925 ;
      LAYER met1 ;
        RECT 0.000 8.025 13.920 8.255 ;
    END
    PORT
      LAYER pwell ;
        RECT 0.810 1.545 3.730 1.795 ;
        RECT 0.810 0.215 4.570 1.545 ;
        RECT 9.455 0.215 10.505 1.625 ;
        RECT -0.130 -0.215 14.050 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 13.920 0.115 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.000 8.055 13.920 8.225 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.000 -0.085 13.920 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 6.005 0.510 6.255 ;
        RECT -0.330 2.095 6.020 6.005 ;
        RECT -0.330 1.885 0.510 2.095 ;
      LAYER met1 ;
        RECT 0.000 3.955 13.920 4.185 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.360 4.155 0.530 5.280 ;
        RECT 0.000 3.985 0.685 4.155 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 4.325 13.920 4.695 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 13.920 3.815 ;
    END
    PORT
      LAYER li1 ;
        RECT 3.175 4.630 3.395 5.405 ;
        RECT 3.175 4.410 3.645 4.630 ;
        RECT 3.425 3.735 3.645 4.410 ;
        RECT 3.060 3.445 3.645 3.735 ;
        RECT 3.425 2.405 3.645 3.445 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.397500 ;
    PORT
      LAYER li1 ;
        RECT 0.955 2.695 1.175 3.075 ;
        RECT 0.755 2.405 1.175 2.695 ;
        RECT 0.755 1.605 0.975 2.405 ;
        RECT 0.755 1.315 1.175 1.605 ;
        RECT 0.955 0.895 1.175 1.315 ;
    END
  END X
  OBS
      LAYER pwell ;
        RECT 6.320 1.195 8.590 6.455 ;
      LAYER li1 ;
        RECT 0.955 7.625 4.900 7.845 ;
        RECT 0.955 6.445 1.175 7.625 ;
        RECT 1.735 6.275 1.955 7.455 ;
        RECT 2.515 6.445 2.735 7.625 ;
        RECT 0.895 6.055 1.955 6.275 ;
        RECT 0.895 4.795 1.115 6.055 ;
        RECT 3.295 5.885 3.515 7.455 ;
        RECT 4.075 6.445 4.295 7.625 ;
        RECT 4.680 6.515 4.900 7.625 ;
        RECT 9.705 7.520 10.295 7.750 ;
        RECT 7.750 7.075 9.535 7.405 ;
        RECT 4.680 6.295 8.445 6.515 ;
        RECT 1.365 5.665 5.675 5.885 ;
        RECT 1.365 5.555 2.035 5.665 ;
        RECT 5.455 4.945 5.675 5.665 ;
        RECT 0.895 4.575 2.780 4.795 ;
        RECT 2.110 4.295 2.780 4.575 ;
        RECT 1.760 3.445 2.350 3.735 ;
        RECT 1.760 2.405 1.930 3.445 ;
        RECT 2.560 3.085 2.780 4.295 ;
        RECT 2.260 2.860 2.780 3.085 ;
        RECT 1.760 0.625 1.990 1.565 ;
        RECT 2.260 0.645 2.480 2.860 ;
        RECT 4.205 2.160 4.425 3.755 ;
        RECT 2.650 1.940 4.425 2.160 ;
        RECT 2.650 1.830 3.320 1.940 ;
        RECT 3.360 0.625 3.590 1.655 ;
        RECT 4.205 0.645 4.425 1.940 ;
        RECT 6.465 1.305 6.685 6.295 ;
        RECT 7.340 0.625 7.570 6.055 ;
        RECT 8.225 1.305 8.445 6.295 ;
        RECT 9.205 4.775 9.535 7.075 ;
        RECT 9.705 6.625 10.035 7.520 ;
        RECT 9.705 6.125 10.535 6.455 ;
        RECT 9.705 4.235 10.035 5.805 ;
        RECT 9.100 3.905 10.035 4.235 ;
        RECT 9.565 3.365 9.895 3.905 ;
        RECT 10.205 3.365 10.535 6.125 ;
        RECT 9.305 3.020 9.895 3.365 ;
        RECT 9.565 2.335 9.895 3.020 ;
        RECT 10.065 3.035 10.535 3.365 ;
        RECT 9.565 0.625 9.895 1.515 ;
        RECT 10.065 0.735 10.395 3.035 ;
        RECT 1.400 0.395 1.990 0.625 ;
        RECT 3.175 0.395 3.765 0.625 ;
        RECT 7.155 0.395 7.745 0.625 ;
        RECT 9.305 0.395 9.895 0.625 ;
  END
END sky130_fd_sc_hvl__lsbuflv2hv_isosrchvaon_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__lsbuflv2hv_symmetric_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__lsbuflv2hv_symmetric_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.040 BY 8.140 ;
  SYMMETRY X Y ;
  SITE unithvdbl ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER li1 ;
        RECT 2.495 1.530 2.805 2.200 ;
    END
  END A
  PIN LVPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 2.800 2.015 4.335 4.325 ;
      LAYER met1 ;
        RECT 0.070 3.020 10.970 3.305 ;
    END
  END LVPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 7.515 11.040 7.885 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 11.040 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT -0.130 7.925 11.170 8.355 ;
        RECT 3.185 5.975 5.255 7.925 ;
        RECT 8.905 6.725 11.020 7.925 ;
      LAYER met1 ;
        RECT 0.000 8.025 11.040 8.255 ;
    END
    PORT
      LAYER pwell ;
        RECT 5.090 1.725 9.500 2.165 ;
        RECT 2.855 0.215 9.500 1.725 ;
        RECT -0.130 -0.215 11.170 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 11.040 0.115 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.000 8.055 11.040 8.225 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.000 -0.085 11.040 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 0.800 6.255 ;
        RECT 6.335 2.465 11.370 6.255 ;
        RECT 9.800 1.885 11.370 2.465 ;
      LAYER met1 ;
        RECT 0.000 3.955 11.040 4.185 ;
    END
    PORT
      LAYER li1 ;
        RECT 8.235 3.985 11.040 4.155 ;
    END
    PORT
      LAYER li1 ;
        RECT 0.000 3.985 0.800 4.155 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 11.040 3.815 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 4.325 11.040 4.695 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.596250 ;
    PORT
      LAYER li1 ;
        RECT 10.600 6.725 10.930 7.625 ;
        RECT 10.690 6.055 10.930 6.725 ;
        RECT 10.600 4.405 10.930 6.055 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 3.145 7.715 5.295 7.885 ;
        RECT 3.145 6.165 3.735 7.715 ;
        RECT 4.055 5.995 4.385 7.545 ;
        RECT 4.705 6.165 5.295 7.715 ;
        RECT 8.535 6.615 8.815 6.955 ;
        RECT 6.695 6.285 8.815 6.615 ;
        RECT 8.995 6.555 9.325 7.625 ;
        RECT 9.690 6.835 10.280 7.745 ;
        RECT 6.695 5.995 7.025 6.285 ;
        RECT 4.055 5.665 7.025 5.995 ;
        RECT 2.885 3.055 3.175 5.495 ;
        RECT 6.695 4.735 7.025 5.665 ;
        RECT 6.565 4.405 7.025 4.735 ;
        RECT 7.390 4.405 7.980 5.945 ;
        RECT 8.300 4.405 8.630 6.285 ;
        RECT 8.995 6.225 10.520 6.555 ;
        RECT 8.995 4.405 9.325 6.225 ;
        RECT 9.690 4.405 10.280 5.945 ;
        RECT 3.345 3.225 4.115 4.200 ;
        RECT 3.435 3.075 4.115 3.225 ;
        RECT 2.885 2.765 3.265 3.055 ;
        RECT 2.975 1.995 3.265 2.765 ;
        RECT 3.435 2.165 3.705 3.075 ;
        RECT 3.875 2.475 4.185 2.905 ;
        RECT 6.565 2.795 6.895 4.405 ;
        RECT 7.095 2.705 7.765 4.215 ;
        RECT 7.955 2.875 8.545 3.705 ;
        RECT 8.915 2.705 9.835 3.465 ;
        RECT 10.125 2.795 10.715 3.705 ;
        RECT 7.095 2.495 9.835 2.705 ;
        RECT 3.875 2.165 5.790 2.475 ;
        RECT 4.480 2.145 5.790 2.165 ;
        RECT 5.960 2.145 7.850 2.325 ;
        RECT 2.975 1.745 4.310 1.995 ;
        RECT 2.975 0.735 3.265 1.745 ;
        RECT 4.480 1.575 4.810 2.145 ;
        RECT 3.435 0.565 3.705 1.575 ;
        RECT 3.875 1.245 4.810 1.575 ;
        RECT 3.875 0.735 4.185 1.245 ;
        RECT 3.095 0.335 4.045 0.565 ;
        RECT 5.050 0.425 5.640 1.975 ;
        RECT 5.960 0.595 6.290 2.145 ;
        RECT 6.610 0.425 7.200 1.975 ;
        RECT 5.050 0.255 7.200 0.425 ;
        RECT 7.520 0.425 7.850 2.145 ;
        RECT 8.170 0.595 8.760 2.495 ;
        RECT 9.080 0.425 9.410 2.055 ;
        RECT 7.520 0.255 9.410 0.425 ;
  END
END sky130_fd_sc_hvl__lsbuflv2hv_symmetric_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__mux2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__mux2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.280 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER li1 ;
        RECT 2.295 1.955 2.625 2.235 ;
        RECT 2.295 1.785 2.905 1.955 ;
        RECT 2.735 1.390 2.905 1.785 ;
        RECT 2.735 1.095 3.685 1.390 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER li1 ;
        RECT 3.085 1.570 3.685 1.955 ;
    END
  END A1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.840000 ;
    PORT
      LAYER li1 ;
        RECT 1.435 3.095 3.230 3.265 ;
        RECT 1.435 1.705 1.765 3.095 ;
        RECT 3.060 2.305 3.230 3.095 ;
        RECT 3.060 2.135 4.675 2.305 ;
        RECT 4.365 1.550 4.675 2.135 ;
    END
  END S
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 5.280 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.055 1.085 1.385 1.415 ;
        RECT 0.055 0.215 5.260 1.085 ;
        RECT -0.130 -0.215 5.410 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 5.280 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 5.610 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 5.280 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 5.280 3.815 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.641250 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.925 0.495 3.755 ;
        RECT 0.125 0.495 0.415 1.925 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 5.280 4.155 ;
        RECT 0.675 2.175 1.255 3.755 ;
        RECT 2.550 2.585 2.880 2.915 ;
        RECT 1.945 2.415 2.880 2.585 ;
        RECT 3.410 2.495 4.720 3.705 ;
        RECT 0.620 1.525 0.950 1.745 ;
        RECT 1.945 1.525 2.115 2.415 ;
        RECT 0.620 1.355 2.555 1.525 ;
        RECT 0.595 0.365 2.205 1.175 ;
        RECT 2.385 0.915 2.555 1.355 ;
        RECT 3.865 1.275 4.115 1.775 ;
        RECT 4.900 1.275 5.150 2.915 ;
        RECT 3.865 1.105 5.150 1.275 ;
        RECT 2.385 0.495 2.880 0.915 ;
        RECT 3.060 0.365 4.720 0.915 ;
        RECT 4.900 0.495 5.150 1.105 ;
        RECT 0.000 -0.085 5.280 0.085 ;
  END
END sky130_fd_sc_hvl__mux2_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__mux4_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__mux4_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.480 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER li1 ;
        RECT 6.770 1.550 7.100 2.520 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER li1 ;
        RECT 4.400 2.300 4.730 3.260 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.525 1.515 2.150 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER li1 ;
        RECT 3.485 2.300 3.845 2.915 ;
    END
  END A3
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.260000 ;
    PORT
      LAYER li1 ;
        RECT 1.905 3.635 3.060 3.805 ;
        RECT 0.565 2.500 0.895 2.915 ;
        RECT 1.905 2.500 2.155 3.635 ;
        RECT 2.890 2.970 3.060 3.635 ;
        RECT 0.565 2.330 2.155 2.500 ;
        RECT 1.905 2.305 2.155 2.330 ;
        RECT 2.685 2.800 3.060 2.970 ;
        RECT 2.685 1.770 2.855 2.800 ;
        RECT 2.685 1.445 5.420 1.770 ;
        RECT 4.925 0.810 5.420 1.445 ;
    END
  END S0
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.840000 ;
    PORT
      LAYER li1 ;
        RECT 8.050 2.915 9.290 3.055 ;
        RECT 7.810 2.885 9.290 2.915 ;
        RECT 7.810 1.920 8.220 2.885 ;
        RECT 9.120 1.985 9.290 2.885 ;
        RECT 9.120 1.315 9.370 1.985 ;
    END
  END S1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 12.480 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 10.160 1.125 12.460 1.505 ;
        RECT 7.990 1.085 12.460 1.125 ;
        RECT 0.020 0.215 12.460 1.085 ;
        RECT -0.130 -0.215 12.610 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 12.480 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 12.810 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 12.480 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 12.480 3.815 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.596250 ;
    PORT
      LAYER li1 ;
        RECT 12.120 0.605 12.370 3.735 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 12.480 4.155 ;
        RECT 0.110 3.115 0.440 3.575 ;
        RECT 0.110 1.345 0.280 3.115 ;
        RECT 0.620 3.095 1.570 3.705 ;
        RECT 2.335 3.175 2.710 3.455 ;
        RECT 1.905 1.345 2.155 2.035 ;
        RECT 0.110 1.175 2.155 1.345 ;
        RECT 2.335 1.265 2.505 3.175 ;
        RECT 3.270 3.095 4.220 3.705 ;
        RECT 5.460 3.095 5.790 3.595 ;
        RECT 6.330 3.095 7.280 3.705 ;
        RECT 8.320 3.635 10.870 3.805 ;
        RECT 7.460 3.115 7.870 3.535 ;
        RECT 8.320 3.235 8.650 3.635 ;
        RECT 9.470 3.115 9.800 3.455 ;
        RECT 5.620 2.915 5.790 3.095 ;
        RECT 7.460 2.915 7.630 3.115 ;
        RECT 3.035 2.120 3.285 2.620 ;
        RECT 5.005 2.120 5.335 2.915 ;
        RECT 5.620 2.745 7.630 2.915 ;
        RECT 3.035 1.950 6.240 2.120 ;
        RECT 0.110 0.515 0.440 1.175 ;
        RECT 2.335 1.095 4.550 1.265 ;
        RECT 5.910 1.095 6.240 1.950 ;
        RECT 0.620 0.365 1.570 0.995 ;
        RECT 2.335 0.495 2.710 1.095 ;
        RECT 3.250 0.365 4.200 0.915 ;
        RECT 4.380 0.435 4.550 1.095 ;
        RECT 6.420 0.915 6.590 2.745 ;
        RECT 7.460 1.740 7.630 2.745 ;
        RECT 7.460 1.570 8.350 1.740 ;
        RECT 5.600 0.615 6.590 0.915 ;
        RECT 6.770 1.175 8.000 1.345 ;
        RECT 6.770 0.435 6.940 1.175 ;
        RECT 4.380 0.265 6.940 0.435 ;
        RECT 7.120 0.365 7.650 0.995 ;
        RECT 7.830 0.435 8.000 1.175 ;
        RECT 8.180 0.615 8.350 1.570 ;
        RECT 9.550 1.135 9.720 3.115 ;
        RECT 9.900 2.655 10.150 2.915 ;
        RECT 9.900 2.115 10.520 2.655 ;
        RECT 8.530 1.035 9.720 1.135 ;
        RECT 8.530 0.965 9.990 1.035 ;
        RECT 8.530 0.435 8.700 0.965 ;
        RECT 7.830 0.265 8.700 0.435 ;
        RECT 8.880 0.435 9.210 0.785 ;
        RECT 9.550 0.615 9.990 0.965 ;
        RECT 10.270 0.915 10.520 2.115 ;
        RECT 10.700 1.925 10.870 3.635 ;
        RECT 11.050 2.175 11.940 3.755 ;
        RECT 10.700 1.595 11.915 1.925 ;
        RECT 10.700 0.435 10.870 1.595 ;
        RECT 8.880 0.265 10.870 0.435 ;
        RECT 11.050 0.365 11.940 1.415 ;
        RECT 0.000 -0.085 12.480 0.085 ;
  END
END sky130_fd_sc_hvl__mux4_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__nand2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__nand2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.400 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.125000 ;
    PORT
      LAYER li1 ;
        RECT 1.975 1.525 2.275 1.855 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.125000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.550 1.015 1.935 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 2.400 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.250 0.215 2.290 1.435 ;
        RECT -0.130 -0.215 2.530 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 2.400 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 2.730 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 2.400 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 2.400 3.815 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.633750 ;
    PORT
      LAYER li1 ;
        RECT 1.220 1.695 1.470 3.755 ;
        RECT 1.220 1.525 1.795 1.695 ;
        RECT 1.580 1.345 1.795 1.525 ;
        RECT 1.580 1.175 2.180 1.345 ;
        RECT 1.850 0.515 2.180 1.175 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 2.400 4.155 ;
        RECT 0.090 2.175 1.040 3.755 ;
        RECT 1.660 2.175 2.250 3.755 ;
        RECT 0.090 0.365 1.400 1.345 ;
        RECT 0.000 -0.085 2.400 0.085 ;
  END
END sky130_fd_sc_hvl__nand2_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__nand3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__nand3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.125000 ;
    PORT
      LAYER li1 ;
        RECT 2.455 0.810 2.725 1.725 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.125000 ;
    PORT
      LAYER li1 ;
        RECT 1.885 0.810 2.275 1.725 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.125000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.505 0.995 1.835 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 3.360 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.300 0.215 3.265 1.415 ;
        RECT -0.130 -0.215 3.490 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 3.360 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 3.690 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 3.360 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 3.360 3.815 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.065000 ;
    PORT
      LAYER li1 ;
        RECT 1.200 2.075 1.370 3.755 ;
        RECT 2.980 2.075 3.235 3.755 ;
        RECT 1.200 1.905 3.235 2.075 ;
        RECT 2.980 1.325 3.235 1.905 ;
        RECT 2.905 0.495 3.235 1.325 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 3.360 4.155 ;
        RECT 0.090 2.175 1.020 3.755 ;
        RECT 1.550 2.255 2.800 3.755 ;
        RECT 0.090 0.365 1.705 1.325 ;
        RECT 0.000 -0.085 3.360 0.085 ;
  END
END sky130_fd_sc_hvl__nand3_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__nor2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__nor2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.400 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.125000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.775 1.315 2.120 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.125000 ;
    PORT
      LAYER li1 ;
        RECT 1.495 1.775 1.825 2.120 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 2.400 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.270 0.215 2.380 1.415 ;
        RECT -0.130 -0.215 2.530 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 2.400 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 2.730 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 2.400 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 2.400 3.815 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.637500 ;
    PORT
      LAYER li1 ;
        RECT 2.020 1.595 2.275 3.755 ;
        RECT 1.200 1.425 2.275 1.595 ;
        RECT 1.200 0.495 1.530 1.425 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 2.400 4.155 ;
        RECT 0.090 2.300 1.760 3.755 ;
        RECT 0.090 0.365 1.020 1.325 ;
        RECT 1.720 0.365 2.310 1.245 ;
        RECT 0.000 -0.085 2.400 0.085 ;
  END
END sky130_fd_sc_hvl__nor2_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__nor3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__nor3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.125000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.525 0.425 2.120 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.125000 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.775 1.795 2.120 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.125000 ;
    PORT
      LAYER li1 ;
        RECT 1.975 1.775 2.305 3.260 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 3.360 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.060 0.215 2.910 1.415 ;
        RECT -0.130 -0.215 3.490 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 3.360 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 3.690 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 3.360 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 3.360 3.815 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.836250 ;
    PORT
      LAYER li1 ;
        RECT 2.490 1.595 2.755 3.755 ;
        RECT 0.930 1.425 2.755 1.595 ;
        RECT 0.930 0.495 1.180 1.425 ;
        RECT 2.490 0.495 2.755 1.425 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 3.360 4.155 ;
        RECT 0.090 2.300 1.760 3.755 ;
        RECT 0.090 0.365 0.680 1.325 ;
        RECT 1.360 0.365 2.310 1.245 ;
        RECT 0.000 -0.085 3.360 0.085 ;
  END
END sky130_fd_sc_hvl__nor3_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__o21a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__o21a_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.320 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.125000 ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.505 4.195 1.835 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.125000 ;
    PORT
      LAYER li1 ;
        RECT 2.555 1.550 2.785 3.260 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.125000 ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.805 2.000 2.120 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 4.320 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.020 1.415 1.330 1.445 ;
        RECT 0.020 0.215 4.295 1.415 ;
        RECT -0.130 -0.215 4.450 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 4.320 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 4.650 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 4.320 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 4.320 3.815 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.626250 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.975 0.595 3.755 ;
        RECT 0.125 0.525 0.380 1.975 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 4.320 4.155 ;
        RECT 0.775 2.300 2.025 3.755 ;
        RECT 0.550 1.625 0.835 1.795 ;
        RECT 2.205 1.625 2.375 3.755 ;
        RECT 2.965 2.175 4.230 3.755 ;
        RECT 0.550 1.455 2.375 1.625 ;
        RECT 0.550 0.365 1.315 1.275 ;
        RECT 1.495 0.495 1.825 1.455 ;
        RECT 3.855 1.275 4.185 1.325 ;
        RECT 2.275 1.105 4.185 1.275 ;
        RECT 2.275 0.495 2.605 1.105 ;
        RECT 2.785 0.365 3.675 0.925 ;
        RECT 3.855 0.495 4.185 1.105 ;
        RECT 0.000 -0.085 4.320 0.085 ;
  END
END sky130_fd_sc_hvl__o21a_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__o21ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__o21ai_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.125000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.505 0.855 1.835 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.125000 ;
    PORT
      LAYER li1 ;
        RECT 1.065 1.505 1.795 1.760 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.125000 ;
    PORT
      LAYER li1 ;
        RECT 2.325 1.805 3.235 2.120 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 3.360 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.020 0.215 2.930 1.415 ;
        RECT -0.130 -0.215 3.490 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 3.360 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 3.690 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 3.360 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 3.360 3.815 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.633750 ;
    PORT
      LAYER li1 ;
        RECT 1.565 2.110 2.040 3.755 ;
        RECT 1.565 1.940 2.145 2.110 ;
        RECT 1.975 1.625 2.145 1.940 ;
        RECT 1.975 1.455 2.820 1.625 ;
        RECT 2.490 0.495 2.820 1.455 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 3.360 4.155 ;
        RECT 0.090 2.175 1.040 3.755 ;
        RECT 2.220 2.300 3.170 3.755 ;
        RECT 0.130 1.275 0.460 1.325 ;
        RECT 0.130 1.105 2.040 1.275 ;
        RECT 0.130 0.495 0.460 1.105 ;
        RECT 0.640 0.365 1.530 0.925 ;
        RECT 1.710 0.495 2.040 1.105 ;
        RECT 0.000 -0.085 3.360 0.085 ;
  END
END sky130_fd_sc_hvl__o21ai_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__o22a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__o22a_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.280 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.125000 ;
    PORT
      LAYER li1 ;
        RECT 1.420 1.775 2.150 2.055 ;
        RECT 1.980 1.570 2.150 1.775 ;
        RECT 1.980 1.400 2.775 1.570 ;
        RECT 4.550 1.400 4.880 2.015 ;
        RECT 2.605 1.230 4.880 1.400 ;
        RECT 3.035 1.210 3.710 1.230 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.125000 ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.580 4.195 1.910 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.125000 ;
    PORT
      LAYER li1 ;
        RECT 2.330 1.750 2.755 2.120 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.125000 ;
    PORT
      LAYER li1 ;
        RECT 2.955 1.580 3.250 2.120 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 5.280 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.020 0.215 4.570 1.415 ;
        RECT -0.130 -0.215 5.410 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 5.280 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 5.610 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 5.280 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 5.280 3.815 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.641250 ;
    PORT
      LAYER li1 ;
        RECT 0.125 0.495 0.380 3.755 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 5.280 4.155 ;
        RECT 0.560 2.650 3.250 3.755 ;
        RECT 3.430 2.470 3.680 3.755 ;
        RECT 0.585 2.300 3.680 2.470 ;
        RECT 0.585 1.595 0.915 2.300 ;
        RECT 3.430 2.175 3.680 2.300 ;
        RECT 3.860 2.195 5.170 3.735 ;
        RECT 0.585 1.425 1.800 1.595 ;
        RECT 0.560 0.365 1.450 1.245 ;
        RECT 1.630 1.220 1.800 1.425 ;
        RECT 1.630 1.050 2.425 1.220 ;
        RECT 2.255 0.880 2.855 1.050 ;
        RECT 1.745 0.435 2.075 0.870 ;
        RECT 2.525 0.615 2.855 0.880 ;
        RECT 3.350 0.435 3.680 1.030 ;
        RECT 1.745 0.265 3.680 0.435 ;
        RECT 3.890 0.365 5.190 1.050 ;
        RECT 0.000 -0.085 5.280 0.085 ;
  END
END sky130_fd_sc_hvl__o22a_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__o22ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__o22ai_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.840 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.125000 ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.805 3.715 2.120 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.125000 ;
    PORT
      LAYER li1 ;
        RECT 2.250 1.805 2.755 2.120 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.125000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.535 0.550 1.865 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.125000 ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.535 1.595 1.750 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 3.840 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.050 0.215 3.820 1.445 ;
        RECT -0.130 -0.215 3.970 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 3.840 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 4.170 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 3.840 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 3.840 3.815 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.742500 ;
    PORT
      LAYER li1 ;
        RECT 1.875 3.260 2.045 3.755 ;
        RECT 1.525 2.175 2.045 3.260 ;
        RECT 1.525 2.100 1.795 2.175 ;
        RECT 0.735 1.930 1.795 2.100 ;
        RECT 0.735 1.355 0.905 1.930 ;
        RECT 0.735 0.615 1.270 1.355 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 3.840 4.155 ;
        RECT 0.090 2.280 1.345 3.755 ;
        RECT 2.305 2.300 3.615 3.755 ;
        RECT 1.800 1.455 3.670 1.625 ;
        RECT 0.160 0.435 0.490 1.355 ;
        RECT 1.800 0.435 1.970 1.455 ;
        RECT 0.160 0.265 1.970 0.435 ;
        RECT 2.150 0.365 3.250 1.275 ;
        RECT 3.420 0.525 3.670 1.455 ;
        RECT 0.000 -0.085 3.840 0.085 ;
  END
END sky130_fd_sc_hvl__o22ai_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__or2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__or2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.360 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER li1 ;
        RECT 1.530 1.175 1.860 1.725 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.175 0.935 1.725 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 3.360 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.010 1.085 3.340 1.415 ;
        RECT 0.290 0.215 3.340 1.085 ;
        RECT -0.130 -0.215 3.490 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 3.360 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 3.690 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 3.360 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 3.360 3.815 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.641250 ;
    PORT
      LAYER li1 ;
        RECT 2.980 0.495 3.235 3.755 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 3.360 4.155 ;
        RECT 0.400 2.075 0.650 2.675 ;
        RECT 0.830 2.255 2.800 3.755 ;
        RECT 0.400 1.905 2.775 2.075 ;
        RECT 1.180 0.995 1.350 1.905 ;
        RECT 2.445 1.725 2.775 1.905 ;
        RECT 0.090 0.365 1.000 0.995 ;
        RECT 1.180 0.495 1.510 0.995 ;
        RECT 2.040 0.365 2.630 1.325 ;
        RECT 0.000 -0.085 3.360 0.085 ;
  END
END sky130_fd_sc_hvl__or2_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__or3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__or3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.840 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER li1 ;
        RECT 1.915 1.080 2.450 1.390 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.910 1.535 3.260 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER li1 ;
        RECT 0.530 1.080 1.315 1.390 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 3.840 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.510 1.085 3.820 1.415 ;
        RECT 0.020 0.215 3.820 1.085 ;
        RECT -0.130 -0.215 3.970 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 3.840 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 4.170 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 3.840 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 3.840 3.815 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.626250 ;
    PORT
      LAYER li1 ;
        RECT 3.460 0.495 3.715 3.755 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 3.840 4.155 ;
        RECT 1.620 3.430 3.280 3.755 ;
        RECT 0.145 1.730 0.395 2.780 ;
        RECT 1.705 2.175 3.280 3.430 ;
        RECT 2.925 1.730 3.255 1.935 ;
        RECT 0.145 1.560 3.255 1.730 ;
        RECT 0.145 0.495 0.360 1.560 ;
        RECT 1.565 0.910 1.735 1.560 ;
        RECT 0.530 0.365 1.385 0.910 ;
        RECT 1.565 0.495 1.965 0.910 ;
        RECT 2.620 0.365 3.290 1.325 ;
        RECT 0.000 -0.085 3.840 0.085 ;
  END
END sky130_fd_sc_hvl__or3_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__probe_p_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__probe_p_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.600 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.375000 ;
    PORT
      LAYER li1 ;
        RECT 0.635 1.580 2.245 1.815 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 9.600 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.115 0.215 9.505 1.585 ;
        RECT -0.130 -0.215 9.730 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 9.600 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 9.930 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 9.600 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 9.600 3.815 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3.290 2.625 6.310 2.835 ;
    END
    PORT
      LAYER met5 ;
        RECT 3.290 1.235 6.310 2.620 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 9.600 4.155 ;
        RECT 0.615 3.625 9.505 3.795 ;
        RECT 0.245 2.265 0.435 3.545 ;
        RECT 0.615 2.445 1.865 3.625 ;
        RECT 2.045 2.265 2.595 3.445 ;
        RECT 2.765 2.385 3.435 3.625 ;
        RECT 0.245 2.095 2.595 2.265 ;
        RECT 0.245 1.475 0.435 2.095 ;
        RECT 2.425 1.955 2.595 2.095 ;
        RECT 3.605 2.205 3.935 3.445 ;
        RECT 4.105 2.385 4.995 3.625 ;
        RECT 5.165 2.205 5.495 3.445 ;
        RECT 5.665 2.385 6.555 3.625 ;
        RECT 6.725 2.205 7.055 3.445 ;
        RECT 7.225 2.385 8.115 3.625 ;
        RECT 8.905 3.475 9.505 3.625 ;
        RECT 8.285 3.230 8.735 3.445 ;
        RECT 8.285 2.205 8.965 3.230 ;
        RECT 9.135 2.385 9.505 3.475 ;
        RECT 3.605 2.035 8.965 2.205 ;
        RECT 2.425 1.625 3.380 1.955 ;
        RECT 3.665 1.625 8.555 1.795 ;
        RECT 0.245 0.805 0.455 1.475 ;
        RECT 2.425 1.400 2.595 1.625 ;
        RECT 0.675 0.550 1.925 1.385 ;
        RECT 2.105 1.230 2.595 1.400 ;
        RECT 2.105 0.730 2.315 1.230 ;
        RECT 2.765 0.760 3.495 1.445 ;
        RECT 3.665 0.805 3.875 1.625 ;
        RECT 2.605 0.550 3.495 0.760 ;
        RECT 4.045 0.550 5.055 1.445 ;
        RECT 5.225 0.805 5.435 1.625 ;
        RECT 5.605 0.550 6.615 1.445 ;
        RECT 6.785 0.805 6.995 1.625 ;
        RECT 7.165 0.550 8.175 1.445 ;
        RECT 8.345 0.975 8.555 1.625 ;
        RECT 8.735 0.975 8.965 2.035 ;
        RECT 8.345 0.805 8.965 0.975 ;
        RECT 9.135 0.600 9.505 1.445 ;
        RECT 8.975 0.550 9.505 0.600 ;
        RECT 0.675 0.380 9.505 0.550 ;
        RECT 0.000 -0.085 9.600 0.085 ;
      LAYER met1 ;
        RECT 5.505 2.005 7.315 2.235 ;
        RECT 5.505 1.975 6.145 2.005 ;
      LAYER met2 ;
        RECT 5.485 1.865 6.165 2.235 ;
      LAYER met3 ;
        RECT 5.435 1.885 6.215 2.215 ;
      LAYER met4 ;
        RECT 3.410 1.355 6.190 2.535 ;
  END
END sky130_fd_sc_hvl__probe_p_8

#--------EOF---------

MACRO sky130_fd_sc_hvl__probec_p_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__probec_p_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.600 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.375000 ;
    PORT
      LAYER li1 ;
        RECT 0.635 1.580 2.245 1.815 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 7.910 -0.365 10.410 1.235 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.115 0.215 9.505 1.585 ;
        RECT -0.130 -0.215 9.730 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 9.600 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 9.930 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 9.600 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 7.910 2.835 10.410 4.435 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 2.290 1.235 4.160 2.835 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.710 2.835 6.310 4.435 ;
        RECT 4.260 1.235 6.310 2.835 ;
        RECT 4.710 -0.365 6.310 1.235 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 9.600 4.155 ;
        RECT 0.615 3.625 9.505 3.795 ;
        RECT 0.245 2.265 0.435 3.545 ;
        RECT 0.615 2.445 1.865 3.625 ;
        RECT 2.045 2.265 2.595 3.445 ;
        RECT 2.765 2.385 3.435 3.625 ;
        RECT 0.245 2.095 2.595 2.265 ;
        RECT 0.245 1.475 0.435 2.095 ;
        RECT 2.425 1.955 2.595 2.095 ;
        RECT 3.605 2.205 3.935 3.445 ;
        RECT 4.105 2.385 4.995 3.625 ;
        RECT 5.165 2.205 5.495 3.445 ;
        RECT 5.665 2.385 6.555 3.625 ;
        RECT 6.725 2.205 7.055 3.445 ;
        RECT 7.225 2.385 8.115 3.625 ;
        RECT 8.905 3.475 9.505 3.625 ;
        RECT 8.285 3.230 8.735 3.445 ;
        RECT 8.285 2.205 8.965 3.230 ;
        RECT 9.135 2.385 9.505 3.475 ;
        RECT 3.605 1.955 8.965 2.205 ;
        RECT 2.425 1.625 3.380 1.955 ;
        RECT 3.665 1.625 8.965 1.955 ;
        RECT 0.245 0.805 0.455 1.475 ;
        RECT 2.425 1.400 2.595 1.625 ;
        RECT 0.675 0.550 1.925 1.385 ;
        RECT 2.105 1.230 2.595 1.400 ;
        RECT 2.105 0.730 2.315 1.230 ;
        RECT 2.765 0.760 3.495 1.445 ;
        RECT 3.665 0.805 3.875 1.625 ;
        RECT 2.605 0.550 3.495 0.760 ;
        RECT 4.045 0.550 5.055 1.445 ;
        RECT 5.225 0.805 5.435 1.625 ;
        RECT 5.605 0.550 6.615 1.445 ;
        RECT 6.785 0.805 6.995 1.625 ;
        RECT 7.165 0.550 8.175 1.445 ;
        RECT 8.345 0.805 8.965 1.625 ;
        RECT 9.135 0.600 9.505 1.445 ;
        RECT 8.975 0.550 9.505 0.600 ;
        RECT 0.675 0.380 9.505 0.550 ;
        RECT 0.000 -0.085 9.600 0.085 ;
      LAYER met1 ;
        RECT 0.000 3.765 9.600 3.815 ;
        RECT 0.000 3.505 9.920 3.765 ;
        RECT 0.000 3.445 9.600 3.505 ;
        RECT 5.560 1.905 6.210 2.165 ;
        RECT 0.000 0.565 9.600 0.625 ;
        RECT 0.000 0.305 9.920 0.565 ;
        RECT 0.000 0.255 9.600 0.305 ;
      LAYER met2 ;
        RECT 9.215 3.505 9.985 3.785 ;
        RECT 5.440 1.895 6.210 2.175 ;
        RECT 9.215 0.285 9.985 0.565 ;
      LAYER met3 ;
        RECT 9.210 3.480 9.990 3.810 ;
        RECT 2.835 1.875 3.615 2.195 ;
        RECT 5.435 1.870 6.215 2.200 ;
        RECT 9.210 0.260 9.990 0.590 ;
      LAYER met4 ;
        RECT 9.010 3.045 10.190 4.225 ;
        RECT 2.410 1.445 3.590 2.625 ;
        RECT 5.010 1.445 6.190 2.625 ;
        RECT 9.010 -0.155 10.190 1.025 ;
  END
END sky130_fd_sc_hvl__probec_p_8

#--------EOF---------

MACRO sky130_fd_sc_hvl__schmittbuf_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__schmittbuf_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.280 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.170000 ;
    PORT
      LAYER li1 ;
        RECT 2.015 1.855 3.305 2.150 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 5.280 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.520 1.585 3.575 1.675 ;
        RECT 0.190 1.575 3.575 1.585 ;
        RECT 0.190 1.415 3.940 1.575 ;
        RECT 0.190 0.215 5.260 1.415 ;
        RECT -0.130 -0.215 5.410 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 5.280 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.975 5.610 4.485 ;
        RECT -0.330 1.885 1.340 1.975 ;
        RECT 3.885 1.885 5.610 1.975 ;
      LAYER met1 ;
        RECT 0.000 3.955 5.280 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 5.280 3.815 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.596250 ;
    PORT
      LAYER li1 ;
        RECT 4.860 0.515 5.195 3.715 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 5.280 4.155 ;
        RECT 0.740 3.655 1.030 3.735 ;
        RECT 0.085 3.485 1.030 3.655 ;
        RECT 0.085 1.975 0.255 3.485 ;
        RECT 0.740 3.405 1.030 3.485 ;
        RECT 3.130 3.405 4.570 3.735 ;
        RECT 1.200 3.235 2.790 3.405 ;
        RECT 0.430 2.335 0.680 3.085 ;
        RECT 0.430 2.165 0.875 2.335 ;
        RECT 1.200 2.295 1.460 3.235 ;
        RECT 1.655 2.330 2.010 3.065 ;
        RECT 0.085 1.805 0.530 1.975 ;
        RECT 0.280 1.090 0.530 1.805 ;
        RECT 0.705 0.795 0.875 2.165 ;
        RECT 1.655 1.985 1.835 2.330 ;
        RECT 2.460 2.320 2.790 3.235 ;
        RECT 3.235 2.320 4.570 3.405 ;
        RECT 1.045 1.685 1.835 1.985 ;
        RECT 3.855 1.685 4.690 2.055 ;
        RECT 1.045 1.655 4.690 1.685 ;
        RECT 1.600 1.645 4.690 1.655 ;
        RECT 1.600 1.505 4.210 1.645 ;
        RECT 1.060 1.145 1.390 1.410 ;
        RECT 1.600 1.315 1.940 1.505 ;
        RECT 2.390 1.145 2.720 1.335 ;
        RECT 1.060 0.975 2.720 1.145 ;
        RECT 0.705 0.570 2.010 0.795 ;
        RECT 3.120 0.375 4.630 1.285 ;
        RECT 0.000 -0.085 5.280 0.085 ;
  END
END sky130_fd_sc_hvl__schmittbuf_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__sdfrbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__sdfrbp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.160 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.585000 ;
    PORT
      LAYER li1 ;
        RECT 5.870 1.850 6.200 2.520 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.625 2.330 2.135 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.260000 ;
    PORT
      LAYER met1 ;
        RECT 5.375 2.105 5.665 2.150 ;
        RECT 10.655 2.105 10.945 2.150 ;
        RECT 14.975 2.105 15.265 2.150 ;
        RECT 5.375 1.965 15.265 2.105 ;
        RECT 5.375 1.920 5.665 1.965 ;
        RECT 10.655 1.920 10.945 1.965 ;
        RECT 14.975 1.920 15.265 1.965 ;
    END
  END RESET_B
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER li1 ;
        RECT 3.710 2.155 4.040 2.480 ;
        RECT 3.710 1.975 4.705 2.155 ;
        RECT 4.375 1.295 4.705 1.975 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.840000 ;
    PORT
      LAYER li1 ;
        RECT 1.515 2.835 1.765 2.995 ;
        RECT 1.515 2.665 3.040 2.835 ;
        RECT 0.655 1.295 0.985 1.965 ;
        RECT 3.485 1.445 4.195 1.795 ;
        RECT 0.815 0.435 0.985 1.295 ;
        RECT 1.515 1.275 4.195 1.445 ;
        RECT 1.515 0.435 1.685 1.275 ;
        RECT 0.815 0.265 1.685 0.435 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 20.160 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.195 1.085 1.525 1.205 ;
        RECT 11.460 1.180 13.515 1.415 ;
        RECT 4.735 1.085 13.515 1.180 ;
        RECT 16.635 1.255 17.925 1.415 ;
        RECT 18.840 1.255 20.130 1.585 ;
        RECT 16.635 1.085 20.130 1.255 ;
        RECT 0.195 0.215 20.130 1.085 ;
        RECT -0.130 -0.215 20.290 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 20.160 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 20.490 4.485 ;
        RECT 16.405 1.720 18.095 1.885 ;
      LAYER met1 ;
        RECT 0.000 3.955 20.160 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 20.160 3.815 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.626250 ;
    PORT
      LAYER li1 ;
        RECT 19.700 0.685 20.040 3.755 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.596250 ;
    PORT
      LAYER li1 ;
        RECT 17.435 0.515 17.835 3.570 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 20.160 4.155 ;
        RECT 0.090 3.205 0.985 3.705 ;
        RECT 1.165 3.205 1.415 3.705 ;
        RECT 1.675 3.235 2.115 3.735 ;
        RECT 2.545 3.365 3.495 3.735 ;
        RECT 1.165 2.485 1.335 3.205 ;
        RECT 1.945 3.185 2.115 3.235 ;
        RECT 4.655 3.185 4.905 3.735 ;
        RECT 5.085 3.365 5.975 3.755 ;
        RECT 6.155 3.635 7.025 3.805 ;
        RECT 6.155 3.185 6.325 3.635 ;
        RECT 1.945 3.015 6.325 3.185 ;
        RECT 3.270 2.665 4.680 2.835 ;
        RECT 3.270 2.485 3.440 2.665 ;
        RECT 1.165 2.315 3.440 2.485 ;
        RECT 4.350 2.325 4.680 2.665 ;
        RECT 0.090 0.365 0.635 1.115 ;
        RECT 1.165 0.615 1.335 2.315 ;
        RECT 2.730 1.625 3.060 2.315 ;
        RECT 4.885 1.095 5.055 3.015 ;
        RECT 5.235 1.295 5.635 2.150 ;
        RECT 6.505 1.675 6.675 3.455 ;
        RECT 6.855 2.025 7.025 3.635 ;
        RECT 7.205 2.205 7.375 3.705 ;
        RECT 8.275 3.425 8.605 3.755 ;
        RECT 7.555 3.255 8.955 3.425 ;
        RECT 7.555 2.025 7.725 3.255 ;
        RECT 8.355 3.015 8.605 3.075 ;
        RECT 6.855 1.855 7.725 2.025 ;
        RECT 7.905 2.225 8.605 3.015 ;
        RECT 6.505 1.505 7.695 1.675 ;
        RECT 1.865 0.435 2.115 0.995 ;
        RECT 3.275 0.925 5.055 1.095 ;
        RECT 3.275 0.615 3.605 0.925 ;
        RECT 4.765 0.435 5.095 0.755 ;
        RECT 1.865 0.265 5.095 0.435 ;
        RECT 5.275 0.365 6.225 0.995 ;
        RECT 6.505 0.495 6.675 1.505 ;
        RECT 7.365 1.345 7.695 1.505 ;
        RECT 7.905 0.995 8.150 2.225 ;
        RECT 8.785 0.995 8.955 3.255 ;
        RECT 6.870 0.365 7.720 0.915 ;
        RECT 7.900 0.435 8.150 0.995 ;
        RECT 8.410 0.615 8.955 0.995 ;
        RECT 9.135 3.075 9.385 3.755 ;
        RECT 9.925 3.255 10.875 3.755 ;
        RECT 11.325 3.075 11.775 3.735 ;
        RECT 9.135 2.905 11.775 3.075 ;
        RECT 11.955 3.015 12.545 3.735 ;
        RECT 9.135 0.995 9.305 2.905 ;
        RECT 11.325 2.835 11.775 2.905 ;
        RECT 9.510 2.485 9.840 2.675 ;
        RECT 11.325 2.665 11.945 2.835 ;
        RECT 9.510 2.315 11.595 2.485 ;
        RECT 9.510 2.005 9.840 2.315 ;
        RECT 9.700 1.095 9.975 1.755 ;
        RECT 10.225 1.445 10.505 1.945 ;
        RECT 10.685 1.625 11.245 2.135 ;
        RECT 11.425 2.045 11.595 2.315 ;
        RECT 11.775 2.225 11.945 2.665 ;
        RECT 12.735 2.695 12.985 3.755 ;
        RECT 13.435 3.045 13.765 3.755 ;
        RECT 13.435 2.875 14.620 3.045 ;
        RECT 12.735 2.525 13.570 2.695 ;
        RECT 12.125 2.175 13.220 2.345 ;
        RECT 12.125 2.045 12.295 2.175 ;
        RECT 11.425 1.875 12.295 2.045 ;
        RECT 13.400 1.995 13.570 2.525 ;
        RECT 12.475 1.825 13.570 1.995 ;
        RECT 12.475 1.445 12.645 1.825 ;
        RECT 10.225 1.275 12.645 1.445 ;
        RECT 9.135 0.615 9.520 0.995 ;
        RECT 9.700 0.925 12.145 1.095 ;
        RECT 9.700 0.435 9.975 0.925 ;
        RECT 7.900 0.265 9.975 0.435 ;
        RECT 10.770 0.365 11.805 0.745 ;
        RECT 11.975 0.435 12.145 0.925 ;
        RECT 12.315 0.615 12.645 1.275 ;
        RECT 12.825 1.475 13.155 1.645 ;
        RECT 12.825 0.435 12.995 1.475 ;
        RECT 13.750 1.295 13.920 2.875 ;
        RECT 13.175 1.125 13.920 1.295 ;
        RECT 13.175 0.615 13.425 1.125 ;
        RECT 14.100 0.435 14.270 2.555 ;
        RECT 14.450 1.245 14.620 2.875 ;
        RECT 14.800 2.675 15.720 3.705 ;
        RECT 15.900 2.495 16.150 3.175 ;
        RECT 14.800 2.300 16.150 2.495 ;
        RECT 15.005 1.425 15.685 2.120 ;
        RECT 15.980 2.005 16.150 2.300 ;
        RECT 16.330 2.185 17.255 3.705 ;
        RECT 15.980 1.835 16.545 2.005 ;
        RECT 15.865 1.245 16.195 1.655 ;
        RECT 14.450 1.075 16.195 1.245 ;
        RECT 16.375 0.895 16.545 1.835 ;
        RECT 18.025 1.985 18.355 2.985 ;
        RECT 18.535 2.175 19.485 3.755 ;
        RECT 18.025 1.655 19.520 1.985 ;
        RECT 11.975 0.265 14.270 0.435 ;
        RECT 14.450 0.365 15.400 0.895 ;
        RECT 16.175 0.515 16.545 0.895 ;
        RECT 16.725 0.365 17.255 1.305 ;
        RECT 18.025 0.685 18.385 1.655 ;
        RECT 18.565 0.365 19.515 1.475 ;
        RECT 0.000 -0.085 20.160 0.085 ;
  END
END sky130_fd_sc_hvl__sdfrbp_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__sdfrtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__sdfrtp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 19.200 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.585000 ;
    PORT
      LAYER li1 ;
        RECT 15.485 1.955 16.140 2.495 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER li1 ;
        RECT 2.910 2.660 3.205 3.260 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.260000 ;
    PORT
      LAYER met1 ;
        RECT 4.415 2.475 4.705 2.520 ;
        RECT 8.255 2.475 8.545 2.520 ;
        RECT 14.015 2.475 14.305 2.520 ;
        RECT 4.415 2.335 14.305 2.475 ;
        RECT 4.415 2.290 4.705 2.335 ;
        RECT 8.255 2.290 8.545 2.335 ;
        RECT 14.015 2.290 14.305 2.335 ;
    END
  END RESET_B
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.180 1.115 1.510 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.840000 ;
    PORT
      LAYER li1 ;
        RECT 1.995 2.005 2.380 2.575 ;
        RECT 1.995 1.835 3.175 2.005 ;
        RECT 4.880 1.835 5.635 2.525 ;
        RECT 1.995 1.445 2.245 1.835 ;
        RECT 3.005 1.550 5.635 1.835 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 19.200 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 9.215 1.180 15.625 1.455 ;
        RECT 0.555 1.105 15.625 1.180 ;
        RECT 16.995 1.105 19.180 1.415 ;
        RECT 0.555 0.215 19.180 1.105 ;
        RECT -0.130 -0.215 19.330 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 19.200 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 19.530 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 19.200 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 19.200 3.815 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.626250 ;
    PORT
      LAYER li1 ;
        RECT 18.820 0.515 19.075 3.755 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 19.200 4.155 ;
        RECT 0.305 3.275 0.635 3.705 ;
        RECT 1.420 3.455 2.370 3.705 ;
        RECT 2.560 3.535 3.555 3.705 ;
        RECT 2.560 3.275 2.730 3.535 ;
        RECT 0.305 3.105 2.730 3.275 ;
        RECT 3.385 3.225 3.555 3.535 ;
        RECT 3.735 3.405 4.625 3.705 ;
        RECT 4.805 3.635 6.005 3.805 ;
        RECT 4.805 3.225 4.975 3.635 ;
        RECT 0.305 1.860 0.475 3.105 ;
        RECT 3.385 3.055 4.975 3.225 ;
        RECT 0.730 2.755 2.730 2.925 ;
        RECT 5.155 2.875 5.485 3.455 ;
        RECT 5.755 3.165 6.005 3.635 ;
        RECT 0.730 2.255 1.060 2.755 ;
        RECT 0.305 1.690 1.465 1.860 ;
        RECT 0.665 0.435 0.995 0.995 ;
        RECT 1.295 0.915 1.465 1.690 ;
        RECT 1.645 1.265 1.815 2.755 ;
        RECT 2.560 2.480 2.730 2.755 ;
        RECT 3.385 2.705 5.485 2.875 ;
        RECT 3.385 2.480 3.555 2.705 ;
        RECT 2.560 2.310 3.555 2.480 ;
        RECT 3.965 2.290 4.675 2.525 ;
        RECT 3.965 2.015 4.300 2.290 ;
        RECT 2.480 1.345 2.810 1.655 ;
        RECT 2.480 1.265 5.535 1.345 ;
        RECT 1.645 1.175 5.535 1.265 ;
        RECT 1.645 1.095 2.810 1.175 ;
        RECT 1.295 0.615 2.485 0.915 ;
        RECT 3.645 0.435 3.975 0.995 ;
        RECT 0.665 0.265 3.975 0.435 ;
        RECT 4.155 0.365 5.105 0.995 ;
        RECT 5.285 0.515 5.535 1.175 ;
        RECT 5.835 1.005 6.005 3.165 ;
        RECT 5.755 0.515 6.005 1.005 ;
        RECT 6.185 3.635 7.215 3.805 ;
        RECT 6.185 0.435 6.355 3.635 ;
        RECT 6.535 2.885 6.865 3.455 ;
        RECT 7.045 3.235 7.215 3.635 ;
        RECT 7.405 3.415 8.355 3.705 ;
        RECT 8.535 3.635 9.785 3.805 ;
        RECT 8.535 3.235 8.705 3.635 ;
        RECT 7.045 3.065 8.705 3.235 ;
        RECT 8.885 2.885 9.215 3.455 ;
        RECT 6.535 2.715 9.215 2.885 ;
        RECT 6.535 0.995 6.705 2.715 ;
        RECT 6.950 2.085 7.280 2.535 ;
        RECT 6.950 1.915 7.605 2.085 ;
        RECT 7.045 1.345 7.255 1.735 ;
        RECT 7.435 1.695 7.605 1.915 ;
        RECT 7.785 2.045 8.115 2.535 ;
        RECT 8.295 2.225 8.760 2.535 ;
        RECT 9.045 2.395 9.215 2.715 ;
        RECT 9.455 3.305 9.785 3.635 ;
        RECT 9.965 3.485 10.915 3.735 ;
        RECT 13.015 3.370 13.965 3.705 ;
        RECT 14.145 3.355 15.095 3.525 ;
        RECT 9.455 3.135 12.810 3.305 ;
        RECT 14.145 3.190 14.315 3.355 ;
        RECT 9.455 2.695 9.785 3.135 ;
        RECT 10.960 2.675 11.440 2.955 ;
        RECT 10.490 2.395 10.780 2.555 ;
        RECT 9.045 2.225 10.780 2.395 ;
        RECT 10.960 2.045 11.130 2.675 ;
        RECT 11.620 2.455 11.790 3.135 ;
        RECT 7.785 1.875 11.130 2.045 ;
        RECT 7.435 1.525 10.780 1.695 ;
        RECT 7.045 1.175 9.635 1.345 ;
        RECT 6.535 0.615 6.865 0.995 ;
        RECT 7.045 0.435 7.255 1.175 ;
        RECT 6.185 0.265 7.255 0.435 ;
        RECT 8.115 0.365 9.065 0.995 ;
        RECT 9.305 0.885 9.635 1.175 ;
        RECT 9.840 0.365 10.430 1.345 ;
        RECT 10.610 0.435 10.780 1.525 ;
        RECT 10.960 1.285 11.130 1.875 ;
        RECT 11.310 2.285 11.790 2.455 ;
        RECT 11.310 1.465 11.480 2.285 ;
        RECT 11.970 2.105 12.300 2.955 ;
        RECT 12.480 2.285 12.810 3.135 ;
        RECT 13.030 3.020 14.315 3.190 ;
        RECT 13.030 2.105 13.200 3.020 ;
        RECT 14.495 2.840 14.745 3.175 ;
        RECT 11.660 1.935 13.200 2.105 ;
        RECT 13.380 2.670 14.745 2.840 ;
        RECT 11.660 1.365 11.830 1.935 ;
        RECT 13.380 1.895 13.710 2.670 ;
        RECT 14.040 1.895 14.370 2.490 ;
        RECT 12.010 1.715 13.020 1.755 ;
        RECT 12.010 1.545 14.395 1.715 ;
        RECT 10.960 0.615 11.325 1.285 ;
        RECT 11.660 0.615 12.105 1.365 ;
        RECT 12.285 0.435 12.455 1.545 ;
        RECT 10.610 0.265 12.455 0.435 ;
        RECT 13.085 0.365 14.035 1.365 ;
        RECT 14.225 0.705 14.395 1.545 ;
        RECT 14.575 1.345 14.745 2.670 ;
        RECT 14.925 2.275 15.095 3.355 ;
        RECT 15.275 2.675 16.165 3.705 ;
        RECT 14.925 1.775 15.255 2.275 ;
        RECT 16.345 2.125 16.595 3.505 ;
        RECT 17.065 2.305 17.550 3.005 ;
        RECT 16.345 1.955 17.200 2.125 ;
        RECT 14.925 1.605 16.850 1.775 ;
        RECT 17.030 1.425 17.200 1.955 ;
        RECT 14.575 1.175 15.535 1.345 ;
        RECT 15.205 0.885 15.535 1.175 ;
        RECT 15.755 1.255 17.200 1.425 ;
        RECT 17.380 1.815 17.550 2.305 ;
        RECT 17.730 2.175 18.640 3.755 ;
        RECT 17.380 1.485 18.615 1.815 ;
        RECT 15.755 0.705 16.085 1.255 ;
        RECT 17.380 1.075 17.550 1.485 ;
        RECT 14.225 0.535 16.085 0.705 ;
        RECT 16.275 0.365 16.865 0.995 ;
        RECT 17.105 0.825 17.550 1.075 ;
        RECT 17.730 0.365 18.640 1.305 ;
        RECT 0.000 -0.085 19.200 0.085 ;
  END
END sky130_fd_sc_hvl__sdfrtp_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__sdfsbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__sdfsbp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.160 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.585000 ;
    PORT
      LAYER li1 ;
        RECT 4.380 1.180 4.710 2.150 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER li1 ;
        RECT 1.975 1.845 2.305 2.355 ;
    END
  END D
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER li1 ;
        RECT 3.485 0.810 3.690 2.150 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.840000 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.665 1.795 2.165 ;
        RECT 2.680 1.665 2.955 1.765 ;
        RECT 0.605 1.495 2.955 1.665 ;
        RECT 2.680 1.095 2.955 1.495 ;
    END
  END SCE
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.840000 ;
    PORT
      LAYER li1 ;
        RECT 14.000 1.425 14.845 1.645 ;
        RECT 10.205 1.210 12.355 1.380 ;
        RECT 12.185 0.435 12.355 1.210 ;
        RECT 14.000 0.435 14.170 1.425 ;
        RECT 12.185 0.265 14.170 0.435 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 20.160 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 6.650 1.130 9.450 1.150 ;
        RECT 5.320 1.085 9.450 1.130 ;
        RECT 11.075 1.085 20.140 1.415 ;
        RECT 0.045 0.215 20.140 1.085 ;
        RECT -0.130 -0.215 20.290 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 20.160 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 20.490 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 20.160 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 20.160 3.815 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.498750 ;
    PORT
      LAYER li1 ;
        RECT 19.700 2.355 20.035 3.435 ;
        RECT 19.805 1.325 20.035 2.355 ;
        RECT 19.700 0.495 20.035 1.325 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.611250 ;
    PORT
      LAYER li1 ;
        RECT 17.405 0.495 17.785 3.735 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 20.160 4.155 ;
        RECT 0.130 2.705 0.460 3.305 ;
        RECT 0.640 2.885 1.590 3.705 ;
        RECT 2.400 3.055 2.730 3.305 ;
        RECT 2.400 2.885 3.235 3.055 ;
        RECT 0.130 2.535 2.885 2.705 ;
        RECT 0.130 1.315 0.300 2.535 ;
        RECT 2.635 2.015 2.885 2.535 ;
        RECT 3.065 2.625 3.235 2.885 ;
        RECT 3.415 2.805 4.305 3.705 ;
        RECT 4.485 3.635 5.515 3.805 ;
        RECT 4.485 2.625 4.655 3.635 ;
        RECT 4.835 2.805 5.165 3.455 ;
        RECT 3.065 2.455 4.655 2.625 ;
        RECT 0.130 1.095 2.300 1.315 ;
        RECT 0.130 0.495 0.485 1.095 ;
        RECT 3.135 0.915 3.305 2.455 ;
        RECT 4.940 1.870 5.165 2.805 ;
        RECT 5.345 2.220 5.515 3.635 ;
        RECT 5.695 2.400 5.865 3.705 ;
        RECT 6.045 3.390 7.295 3.560 ;
        RECT 6.045 2.220 6.215 3.390 ;
        RECT 5.345 2.050 6.215 2.220 ;
        RECT 6.395 2.290 6.645 3.210 ;
        RECT 6.840 2.740 7.295 3.390 ;
        RECT 4.940 1.700 6.065 1.870 ;
        RECT 0.665 0.365 1.615 0.915 ;
        RECT 2.425 0.745 3.305 0.915 ;
        RECT 2.425 0.495 2.755 0.745 ;
        RECT 3.870 0.365 4.760 0.995 ;
        RECT 4.940 0.515 5.190 1.700 ;
        RECT 5.735 1.200 6.065 1.700 ;
        RECT 6.395 1.020 6.565 2.290 ;
        RECT 6.840 1.060 7.010 2.740 ;
        RECT 5.370 0.365 5.960 1.020 ;
        RECT 6.190 0.435 6.565 1.020 ;
        RECT 6.760 0.615 7.010 1.060 ;
        RECT 7.190 2.290 7.520 2.560 ;
        RECT 7.190 0.435 7.360 2.290 ;
        RECT 7.700 2.080 7.995 3.240 ;
        RECT 8.615 2.960 9.565 3.705 ;
        RECT 10.955 3.350 11.905 3.755 ;
        RECT 9.745 3.170 10.775 3.340 ;
        RECT 9.745 2.780 9.915 3.170 ;
        RECT 10.605 3.000 12.335 3.170 ;
        RECT 8.200 2.610 9.915 2.780 ;
        RECT 8.200 2.290 8.530 2.610 ;
        RECT 10.095 2.430 10.425 2.990 ;
        RECT 8.910 2.260 10.425 2.430 ;
        RECT 11.315 2.080 11.645 2.555 ;
        RECT 12.025 2.295 12.335 3.000 ;
        RECT 12.515 2.695 12.845 3.755 ;
        RECT 13.500 2.875 14.450 3.705 ;
        RECT 14.970 2.695 15.300 3.175 ;
        RECT 12.515 2.525 15.300 2.695 ;
        RECT 12.025 2.125 13.405 2.295 ;
        RECT 7.700 1.910 11.645 2.080 ;
        RECT 7.700 1.060 7.870 1.910 ;
        RECT 12.200 1.730 12.530 1.875 ;
        RECT 7.540 0.640 7.870 1.060 ;
        RECT 8.050 1.560 12.530 1.730 ;
        RECT 8.050 1.150 8.325 1.560 ;
        RECT 13.165 1.415 13.405 2.125 ;
        RECT 13.585 1.995 13.755 2.525 ;
        RECT 15.685 2.345 16.060 2.675 ;
        RECT 13.935 2.175 16.060 2.345 ;
        RECT 16.240 2.195 17.190 3.735 ;
        RECT 13.585 1.825 15.545 1.995 ;
        RECT 8.050 0.435 8.220 1.150 ;
        RECT 8.910 1.140 9.910 1.380 ;
        RECT 6.190 0.265 8.220 0.435 ;
        RECT 8.410 0.365 9.360 0.960 ;
        RECT 9.580 0.515 9.910 1.140 ;
        RECT 10.545 0.365 11.495 1.030 ;
        RECT 12.655 0.785 12.985 1.325 ;
        RECT 13.585 0.785 13.755 1.825 ;
        RECT 15.215 1.425 15.545 1.825 ;
        RECT 12.655 0.615 13.755 0.785 ;
        RECT 14.350 0.365 15.300 1.245 ;
        RECT 15.730 0.825 16.060 2.175 ;
        RECT 18.025 1.675 18.355 3.185 ;
        RECT 18.535 2.355 19.485 3.705 ;
        RECT 19.245 1.675 19.575 2.175 ;
        RECT 18.025 1.505 19.575 1.675 ;
        RECT 16.240 0.365 17.190 1.325 ;
        RECT 18.025 0.825 18.355 1.505 ;
        RECT 18.535 0.365 19.485 1.325 ;
        RECT 0.000 -0.085 20.160 0.085 ;
  END
END sky130_fd_sc_hvl__sdfsbp_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__sdfstp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__sdfstp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.720 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.585000 ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.175 4.525 2.150 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER li1 ;
        RECT 1.945 1.845 2.275 2.355 ;
    END
  END D
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER li1 ;
        RECT 3.420 1.175 3.750 2.150 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.840000 ;
    PORT
      LAYER li1 ;
        RECT 0.565 1.665 0.895 2.165 ;
        RECT 2.525 1.665 2.890 1.780 ;
        RECT 0.565 1.495 2.890 1.665 ;
        RECT 2.525 1.095 2.890 1.495 ;
    END
  END SCE
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.840000 ;
    PORT
      LAYER li1 ;
        RECT 10.535 1.175 11.635 1.345 ;
        RECT 11.465 0.435 11.635 1.175 ;
        RECT 14.045 0.810 14.520 1.760 ;
        RECT 14.045 0.435 14.215 0.810 ;
        RECT 11.465 0.265 14.215 0.435 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 18.720 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 5.110 1.115 6.400 1.165 ;
        RECT 5.110 1.085 9.240 1.115 ;
        RECT 10.865 1.085 18.700 1.415 ;
        RECT 0.020 0.215 18.700 1.085 ;
        RECT -0.130 -0.215 18.850 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 18.720 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 19.050 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 18.720 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 18.720 3.815 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.478750 ;
    PORT
      LAYER li1 ;
        RECT 18.260 0.495 18.610 3.395 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 18.720 4.155 ;
        RECT 0.110 2.705 0.440 3.285 ;
        RECT 0.620 2.885 1.570 3.705 ;
        RECT 2.380 3.055 2.710 3.305 ;
        RECT 2.380 2.885 3.240 3.055 ;
        RECT 0.110 2.535 2.890 2.705 ;
        RECT 0.110 1.315 0.280 2.535 ;
        RECT 2.635 2.015 2.890 2.535 ;
        RECT 3.070 2.625 3.240 2.885 ;
        RECT 3.420 2.805 4.315 3.705 ;
        RECT 4.495 3.635 5.365 3.805 ;
        RECT 4.495 2.625 4.665 3.635 ;
        RECT 3.070 2.455 4.665 2.625 ;
        RECT 0.110 1.095 2.255 1.315 ;
        RECT 0.110 0.515 0.440 1.095 ;
        RECT 3.070 0.915 3.240 2.455 ;
        RECT 4.845 1.905 5.015 3.455 ;
        RECT 5.195 2.445 5.365 3.635 ;
        RECT 5.545 2.625 5.725 3.705 ;
        RECT 5.905 3.635 7.095 3.805 ;
        RECT 5.905 2.445 6.075 3.635 ;
        RECT 5.195 2.275 6.075 2.445 ;
        RECT 6.255 2.095 6.530 3.455 ;
        RECT 4.845 1.735 5.835 1.905 ;
        RECT 0.620 0.365 1.570 0.915 ;
        RECT 2.380 0.745 3.240 0.915 ;
        RECT 2.380 0.495 2.710 0.745 ;
        RECT 3.420 0.365 4.370 0.995 ;
        RECT 4.845 0.975 5.015 1.735 ;
        RECT 5.505 1.235 5.835 1.735 ;
        RECT 6.140 1.425 6.530 2.095 ;
        RECT 6.710 2.675 7.095 3.635 ;
        RECT 7.275 3.355 8.305 3.525 ;
        RECT 4.650 0.515 5.015 0.975 ;
        RECT 5.200 0.365 5.450 1.055 ;
        RECT 5.630 0.435 5.800 1.235 ;
        RECT 6.140 1.055 6.310 1.425 ;
        RECT 5.980 0.675 6.310 1.055 ;
        RECT 6.710 1.025 6.880 2.675 ;
        RECT 7.275 1.775 7.445 3.355 ;
        RECT 6.550 0.615 6.880 1.025 ;
        RECT 7.060 1.605 7.445 1.775 ;
        RECT 7.625 2.675 7.955 3.175 ;
        RECT 8.135 2.745 8.305 3.355 ;
        RECT 8.495 2.925 9.445 3.705 ;
        RECT 10.835 3.285 11.785 3.755 ;
        RECT 9.625 3.105 10.655 3.275 ;
        RECT 9.625 2.745 9.795 3.105 ;
        RECT 10.485 2.935 12.180 3.105 ;
        RECT 7.060 0.435 7.230 1.605 ;
        RECT 7.625 1.525 7.795 2.675 ;
        RECT 8.135 2.575 9.795 2.745 ;
        RECT 8.135 2.225 8.410 2.575 ;
        RECT 9.975 2.395 10.305 2.925 ;
        RECT 8.790 2.225 10.305 2.395 ;
        RECT 11.905 2.395 12.180 2.935 ;
        RECT 12.360 2.845 12.690 3.755 ;
        RECT 12.360 2.675 12.920 2.845 ;
        RECT 13.265 2.675 14.215 3.705 ;
        RECT 14.395 3.335 15.625 3.505 ;
        RECT 11.905 2.225 12.570 2.395 ;
        RECT 7.975 1.875 12.220 2.045 ;
        RECT 7.975 1.705 8.305 1.875 ;
        RECT 8.485 1.525 11.525 1.695 ;
        RECT 11.970 1.685 12.220 1.875 ;
        RECT 7.625 1.355 8.655 1.525 ;
        RECT 9.520 1.455 9.850 1.525 ;
        RECT 12.400 1.505 12.570 2.225 ;
        RECT 7.625 1.025 7.795 1.355 ;
        RECT 8.835 1.275 9.165 1.345 ;
        RECT 12.095 1.335 12.570 1.505 ;
        RECT 12.750 2.110 12.920 2.675 ;
        RECT 14.395 2.495 14.565 3.335 ;
        RECT 13.710 2.290 14.565 2.495 ;
        RECT 14.745 2.175 15.075 3.155 ;
        RECT 15.295 2.865 15.625 3.335 ;
        RECT 15.815 3.045 16.405 3.705 ;
        RECT 15.295 2.695 16.020 2.865 ;
        RECT 14.745 2.110 15.585 2.175 ;
        RECT 12.750 1.940 15.585 2.110 ;
        RECT 8.835 1.105 9.700 1.275 ;
        RECT 7.410 0.525 7.795 1.025 ;
        RECT 5.630 0.265 7.230 0.435 ;
        RECT 8.200 0.365 9.150 0.925 ;
        RECT 9.370 0.515 9.700 1.105 ;
        RECT 10.335 0.365 11.285 0.995 ;
        RECT 12.095 0.785 12.265 1.335 ;
        RECT 12.750 1.155 12.920 1.940 ;
        RECT 12.445 0.965 12.920 1.155 ;
        RECT 13.100 0.785 13.350 1.745 ;
        RECT 15.255 1.505 15.585 1.940 ;
        RECT 12.095 0.615 13.350 0.785 ;
        RECT 14.700 0.365 15.590 1.325 ;
        RECT 15.770 0.825 16.020 2.695 ;
        RECT 16.585 2.355 16.955 3.145 ;
        RECT 17.135 2.355 18.080 3.705 ;
        RECT 16.585 1.675 16.915 2.355 ;
        RECT 17.750 1.675 18.080 2.175 ;
        RECT 16.585 1.505 18.080 1.675 ;
        RECT 16.585 0.825 16.915 1.505 ;
        RECT 17.095 0.365 18.045 1.325 ;
        RECT 0.000 -0.085 18.720 0.085 ;
  END
END sky130_fd_sc_hvl__sdfstp_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__sdfxbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__sdfxbp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 19.680 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.585000 ;
    PORT
      LAYER li1 ;
        RECT 10.685 1.895 11.395 2.120 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER li1 ;
        RECT 4.165 1.175 4.675 2.150 ;
    END
  END D
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER li1 ;
        RECT 1.565 1.930 1.975 2.440 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.840000 ;
    PORT
      LAYER li1 ;
        RECT 0.565 1.750 0.895 2.220 ;
        RECT 2.425 1.750 2.755 2.745 ;
        RECT 0.565 1.550 2.755 1.750 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 19.680 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 7.725 1.415 9.835 1.450 ;
        RECT 5.205 1.085 9.835 1.415 ;
        RECT 12.040 1.085 17.175 1.415 ;
        RECT 18.330 1.085 19.660 1.415 ;
        RECT 0.430 0.215 19.660 1.085 ;
        RECT -0.130 -0.215 19.810 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 19.680 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 20.010 4.485 ;
        RECT 15.925 1.715 18.490 1.885 ;
      LAYER met1 ;
        RECT 0.000 3.955 19.680 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 19.680 3.815 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.611250 ;
    PORT
      LAYER li1 ;
        RECT 16.215 2.515 16.545 3.455 ;
        RECT 15.955 2.025 16.545 2.515 ;
        RECT 15.955 0.495 16.285 2.025 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.641250 ;
    PORT
      LAYER li1 ;
        RECT 19.220 0.495 19.555 3.755 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 19.680 4.155 ;
        RECT 0.110 2.555 0.440 3.015 ;
        RECT 0.630 2.620 1.220 3.705 ;
        RECT 1.400 3.095 1.570 3.755 ;
        RECT 1.750 3.335 2.700 3.755 ;
        RECT 2.880 3.610 4.030 3.780 ;
        RECT 2.880 3.275 3.210 3.610 ;
        RECT 3.430 3.095 3.680 3.430 ;
        RECT 1.400 2.925 3.680 3.095 ;
        RECT 3.860 2.850 4.030 3.610 ;
        RECT 4.210 3.635 6.140 3.805 ;
        RECT 4.210 3.030 4.540 3.635 ;
        RECT 4.990 2.850 5.240 3.430 ;
        RECT 3.860 2.680 5.240 2.850 ;
        RECT 0.110 1.345 0.280 2.555 ;
        RECT 3.510 2.330 5.135 2.500 ;
        RECT 3.065 1.345 3.330 1.845 ;
        RECT 0.110 1.175 3.330 1.345 ;
        RECT 0.540 0.495 0.870 1.175 ;
        RECT 3.510 0.995 3.680 2.330 ;
        RECT 1.050 0.365 2.000 0.995 ;
        RECT 2.810 0.825 3.680 0.995 ;
        RECT 2.810 0.495 3.140 0.825 ;
        RECT 3.860 0.365 4.785 0.995 ;
        RECT 4.965 0.435 5.135 2.330 ;
        RECT 5.420 1.775 5.790 3.455 ;
        RECT 5.970 3.285 6.140 3.635 ;
        RECT 6.320 3.465 7.210 3.755 ;
        RECT 7.390 3.285 9.435 3.455 ;
        RECT 5.970 3.115 7.560 3.285 ;
        RECT 5.970 2.125 6.140 3.115 ;
        RECT 7.740 2.855 8.655 3.105 ;
        RECT 9.105 3.100 9.435 3.285 ;
        RECT 7.740 2.555 7.910 2.855 ;
        RECT 8.835 2.750 10.355 2.920 ;
        RECT 8.835 2.675 9.005 2.750 ;
        RECT 6.320 2.305 7.910 2.555 ;
        RECT 8.090 2.485 9.005 2.675 ;
        RECT 9.675 2.320 10.005 2.570 ;
        RECT 10.185 2.470 10.355 2.750 ;
        RECT 10.535 2.650 11.125 3.705 ;
        RECT 11.785 3.635 14.340 3.805 ;
        RECT 11.315 2.470 11.565 3.110 ;
        RECT 7.740 2.135 8.785 2.305 ;
        RECT 5.970 1.955 7.470 2.125 ;
        RECT 5.315 1.605 7.120 1.775 ;
        RECT 5.315 0.615 5.645 1.605 ;
        RECT 7.300 1.425 7.470 1.955 ;
        RECT 5.825 1.255 8.165 1.425 ;
        RECT 5.825 0.435 5.995 1.255 ;
        RECT 4.965 0.265 5.995 0.435 ;
        RECT 6.175 0.365 7.065 1.075 ;
        RECT 7.245 0.760 7.575 1.075 ;
        RECT 7.835 0.940 8.165 1.255 ;
        RECT 8.615 1.360 8.785 2.135 ;
        RECT 9.070 1.715 9.400 2.215 ;
        RECT 9.675 1.715 9.845 2.320 ;
        RECT 10.185 2.300 11.565 2.470 ;
        RECT 10.185 2.140 10.355 2.300 ;
        RECT 11.785 2.205 12.115 3.635 ;
        RECT 12.310 3.285 13.795 3.455 ;
        RECT 10.025 1.895 10.355 2.140 ;
        RECT 11.800 1.715 12.130 2.025 ;
        RECT 9.070 1.545 12.130 1.715 ;
        RECT 8.615 0.940 8.945 1.360 ;
        RECT 9.395 0.760 9.725 1.360 ;
        RECT 7.245 0.590 9.725 0.760 ;
        RECT 9.985 0.495 10.315 1.545 ;
        RECT 11.800 1.445 12.130 1.545 ;
        RECT 10.495 1.265 10.825 1.365 ;
        RECT 10.495 1.095 11.875 1.265 ;
        RECT 12.310 1.245 12.480 3.285 ;
        RECT 12.660 2.205 12.990 3.105 ;
        RECT 13.440 2.265 13.795 3.285 ;
        RECT 14.010 2.695 14.340 3.635 ;
        RECT 14.520 2.695 15.425 3.735 ;
        RECT 15.605 3.635 16.895 3.805 ;
        RECT 15.605 2.695 15.995 3.635 ;
        RECT 15.605 2.515 15.775 2.695 ;
        RECT 14.465 2.265 15.775 2.515 ;
        RECT 10.495 0.365 11.445 0.915 ;
        RECT 11.625 0.645 11.875 1.095 ;
        RECT 12.150 0.825 12.480 1.245 ;
        RECT 12.820 2.085 12.990 2.205 ;
        RECT 12.820 1.915 15.135 2.085 ;
        RECT 12.820 1.325 12.990 1.915 ;
        RECT 13.280 1.505 13.610 1.735 ;
        RECT 14.805 1.545 15.135 1.915 ;
        RECT 12.820 0.825 13.260 1.325 ;
        RECT 13.440 0.645 13.610 1.505 ;
        RECT 11.625 0.475 13.610 0.645 ;
        RECT 13.915 0.365 14.865 1.325 ;
        RECT 15.315 0.495 15.775 2.265 ;
        RECT 16.725 1.835 16.895 3.635 ;
        RECT 17.075 2.025 17.665 3.705 ;
        RECT 17.870 2.025 18.200 2.815 ;
        RECT 18.380 2.175 18.970 3.755 ;
        RECT 18.030 1.835 18.200 2.025 ;
        RECT 16.725 1.505 17.055 1.835 ;
        RECT 18.030 1.675 19.040 1.835 ;
        RECT 17.630 1.505 19.040 1.675 ;
        RECT 16.465 0.365 17.415 1.325 ;
        RECT 17.630 0.495 17.960 1.505 ;
        RECT 18.140 0.365 19.040 1.325 ;
        RECT 0.000 -0.085 19.680 0.085 ;
      LAYER met1 ;
        RECT 5.375 3.215 5.665 3.260 ;
        RECT 13.535 3.215 13.825 3.260 ;
        RECT 5.375 3.075 13.825 3.215 ;
        RECT 5.375 3.030 5.665 3.075 ;
        RECT 13.535 3.030 13.825 3.075 ;
  END
END sky130_fd_sc_hvl__sdfxbp_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__sdfxtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__sdfxtp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.880 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.585000 ;
    PORT
      LAYER li1 ;
        RECT 4.345 1.175 4.675 1.685 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER li1 ;
        RECT 0.605 2.205 2.755 2.520 ;
    END
  END D
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER li1 ;
        RECT 3.600 2.215 4.195 2.765 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.840000 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.855 3.050 2.025 ;
        RECT 0.605 1.445 1.795 1.855 ;
        RECT 2.720 1.095 3.050 1.855 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 14.880 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 13.570 1.415 14.860 1.515 ;
        RECT 8.920 1.085 10.250 1.415 ;
        RECT 12.240 1.085 14.860 1.415 ;
        RECT 0.035 0.215 14.860 1.085 ;
        RECT -0.130 -0.215 15.010 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 14.880 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 15.210 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 14.880 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 14.880 3.815 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.596250 ;
    PORT
      LAYER li1 ;
        RECT 13.660 2.195 14.020 3.735 ;
        RECT 13.850 1.780 14.020 2.195 ;
        RECT 13.850 1.505 14.755 1.780 ;
        RECT 13.660 0.615 14.020 1.505 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 14.880 4.155 ;
        RECT 0.125 1.265 0.380 3.425 ;
        RECT 0.910 2.925 1.860 3.705 ;
        RECT 2.400 3.095 2.730 3.425 ;
        RECT 2.400 2.925 3.400 3.095 ;
        RECT 3.635 2.945 4.585 3.735 ;
        RECT 3.230 2.035 3.400 2.925 ;
        RECT 4.765 2.765 5.095 3.735 ;
        RECT 5.315 2.945 5.905 3.735 ;
        RECT 6.095 3.505 6.425 3.735 ;
        RECT 9.030 3.505 9.980 3.755 ;
        RECT 6.095 3.335 7.325 3.505 ;
        RECT 6.095 2.945 6.425 3.335 ;
        RECT 4.765 2.595 5.605 2.765 ;
        RECT 5.275 2.215 5.605 2.595 ;
        RECT 6.610 2.695 6.975 3.155 ;
        RECT 6.610 2.035 6.780 2.695 ;
        RECT 7.155 2.515 7.325 3.335 ;
        RECT 10.320 3.325 11.450 3.495 ;
        RECT 6.960 2.225 7.325 2.515 ;
        RECT 7.505 2.675 7.755 3.175 ;
        RECT 8.040 3.155 10.490 3.325 ;
        RECT 3.230 1.865 6.780 2.035 ;
        RECT 1.975 1.265 2.305 1.675 ;
        RECT 0.125 1.095 2.305 1.265 ;
        RECT 0.125 0.515 0.455 1.095 ;
        RECT 3.230 0.915 3.400 1.865 ;
        RECT 5.540 1.325 5.870 1.685 ;
        RECT 4.855 1.155 5.870 1.325 ;
        RECT 0.905 0.365 1.855 0.915 ;
        RECT 2.395 0.745 3.400 0.915 ;
        RECT 2.395 0.495 2.725 0.745 ;
        RECT 3.580 0.365 4.485 0.995 ;
        RECT 4.855 0.975 5.025 1.155 ;
        RECT 6.565 0.995 6.780 1.865 ;
        RECT 4.665 0.515 5.025 0.975 ;
        RECT 5.215 0.365 5.805 0.975 ;
        RECT 5.995 0.435 6.325 0.975 ;
        RECT 6.565 0.615 6.895 0.995 ;
        RECT 7.075 0.435 7.245 2.225 ;
        RECT 7.505 1.775 7.675 2.675 ;
        RECT 8.040 2.495 8.210 3.155 ;
        RECT 9.810 2.675 10.140 2.975 ;
        RECT 7.880 1.955 8.210 2.495 ;
        RECT 8.620 2.125 8.950 2.555 ;
        RECT 9.810 2.125 9.980 2.675 ;
        RECT 10.320 2.495 10.490 3.155 ;
        RECT 10.670 2.675 11.075 3.145 ;
        RECT 10.160 2.305 10.490 2.495 ;
        RECT 8.620 1.955 10.645 2.125 ;
        RECT 7.505 1.605 9.685 1.775 ;
        RECT 7.505 0.995 7.755 1.605 ;
        RECT 10.045 1.425 10.295 1.775 ;
        RECT 7.425 0.615 7.755 0.995 ;
        RECT 7.935 1.255 10.295 1.425 ;
        RECT 7.935 0.435 8.210 1.255 ;
        RECT 10.475 1.075 10.645 1.955 ;
        RECT 5.995 0.265 8.210 0.435 ;
        RECT 8.680 0.365 9.630 1.075 ;
        RECT 9.810 0.905 10.645 1.075 ;
        RECT 9.810 0.495 10.140 0.905 ;
        RECT 10.825 0.665 11.075 2.675 ;
        RECT 11.255 1.085 11.450 3.325 ;
        RECT 11.980 2.695 12.930 3.735 ;
        RECT 11.630 2.345 12.930 2.515 ;
        RECT 11.630 0.665 11.800 2.345 ;
        RECT 11.980 1.655 12.310 2.155 ;
        RECT 12.600 1.845 12.930 2.345 ;
        RECT 13.110 2.015 13.440 3.735 ;
        RECT 14.200 2.195 14.790 3.735 ;
        RECT 13.110 1.685 13.670 2.015 ;
        RECT 13.110 1.655 13.440 1.685 ;
        RECT 11.980 1.485 13.440 1.655 ;
        RECT 10.825 0.495 11.800 0.665 ;
        RECT 11.980 0.365 12.930 1.305 ;
        RECT 13.110 0.515 13.440 1.485 ;
        RECT 14.200 0.365 14.790 1.325 ;
        RECT 0.000 -0.085 14.880 0.085 ;
  END
END sky130_fd_sc_hvl__sdfxtp_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__sdlclkp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__sdlclkp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.040 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 1.170000 ;
    PORT
      LAYER li1 ;
        RECT 9.195 3.125 9.560 3.445 ;
        RECT 9.310 2.025 9.560 3.125 ;
        RECT 4.320 1.465 4.650 1.975 ;
        RECT 9.310 1.725 9.640 2.025 ;
    END
  END CLK
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.585000 ;
    PORT
      LAYER li1 ;
        RECT 1.475 1.535 1.805 2.125 ;
    END
  END GATE
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.585000 ;
    PORT
      LAYER li1 ;
        RECT 0.595 1.535 0.925 2.125 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 11.040 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 9.640 1.405 10.930 1.415 ;
        RECT 8.020 1.345 10.930 1.405 ;
        RECT 0.160 1.210 3.050 1.345 ;
        RECT 5.200 1.210 10.930 1.345 ;
        RECT 0.160 0.215 10.930 1.210 ;
        RECT -0.130 -0.215 11.170 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 11.040 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 11.370 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 11.040 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 11.040 3.815 ;
    END
  END VPWR
  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.596250 ;
    PORT
      LAYER li1 ;
        RECT 10.590 1.895 10.955 3.735 ;
        RECT 10.685 1.215 10.955 1.895 ;
        RECT 10.590 0.515 10.955 1.215 ;
    END
  END GCLK
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 11.040 4.155 ;
        RECT 0.290 3.615 4.290 3.815 ;
        RECT 0.290 3.445 1.985 3.615 ;
        RECT 3.625 3.445 4.290 3.615 ;
        RECT 6.645 3.615 10.420 3.815 ;
        RECT 0.290 2.295 0.620 3.445 ;
        RECT 2.155 3.225 3.455 3.445 ;
        RECT 1.850 2.295 2.145 3.055 ;
        RECT 1.975 1.365 2.145 2.295 ;
        RECT 2.630 1.885 2.960 3.055 ;
        RECT 3.235 2.315 3.455 3.225 ;
        RECT 3.960 2.485 4.290 3.445 ;
        RECT 4.480 3.385 6.475 3.555 ;
        RECT 6.645 3.445 9.025 3.615 ;
        RECT 9.730 3.445 10.420 3.615 ;
        RECT 4.480 2.315 4.650 3.385 ;
        RECT 3.235 2.145 4.650 2.315 ;
        RECT 4.820 3.005 6.135 3.215 ;
        RECT 2.555 1.555 3.065 1.885 ;
        RECT 0.290 1.195 2.145 1.365 ;
        RECT 0.290 0.840 0.620 1.195 ;
        RECT 1.070 0.625 1.400 1.025 ;
        RECT 1.850 0.840 2.145 1.195 ;
        RECT 2.630 0.840 2.960 1.555 ;
        RECT 3.235 1.080 3.430 2.145 ;
        RECT 3.180 0.705 3.430 1.080 ;
        RECT 3.600 1.295 3.930 1.965 ;
        RECT 4.820 1.295 5.030 3.005 ;
        RECT 3.600 1.125 5.030 1.295 ;
        RECT 0.730 0.365 1.740 0.625 ;
        RECT 2.115 0.535 2.825 0.670 ;
        RECT 3.600 0.535 3.770 1.125 ;
        RECT 2.115 0.365 3.770 0.535 ;
        RECT 3.940 0.625 4.290 0.955 ;
        RECT 4.780 0.705 5.030 1.125 ;
        RECT 5.335 2.330 5.620 2.660 ;
        RECT 6.305 2.595 6.475 3.385 ;
        RECT 6.095 2.425 6.475 2.595 ;
        RECT 5.335 1.365 5.505 2.330 ;
        RECT 6.095 1.945 6.265 2.425 ;
        RECT 6.780 2.330 7.110 3.445 ;
        RECT 7.620 2.085 7.890 2.660 ;
        RECT 8.110 2.225 8.440 3.445 ;
        RECT 5.675 1.615 6.265 1.945 ;
        RECT 6.475 1.875 7.890 2.085 ;
        RECT 6.475 1.535 6.805 1.875 ;
        RECT 7.620 1.825 7.890 1.875 ;
        RECT 8.415 1.825 8.745 2.055 ;
        RECT 7.085 1.365 7.450 1.655 ;
        RECT 5.335 1.195 7.450 1.365 ;
        RECT 3.940 0.535 4.610 0.625 ;
        RECT 5.335 0.535 5.620 1.195 ;
        RECT 6.780 0.625 7.110 1.025 ;
        RECT 3.940 0.255 4.885 0.535 ;
        RECT 5.055 0.255 5.620 0.535 ;
        RECT 5.790 0.255 7.110 0.625 ;
        RECT 7.280 0.670 7.450 1.195 ;
        RECT 7.620 1.615 8.745 1.825 ;
        RECT 7.620 0.840 7.890 1.615 ;
        RECT 8.415 1.385 8.745 1.615 ;
        RECT 8.915 1.555 9.140 2.955 ;
        RECT 9.730 2.195 10.060 3.445 ;
        RECT 9.905 1.555 10.515 1.725 ;
        RECT 8.915 1.385 10.515 1.555 ;
        RECT 8.915 1.215 9.140 1.385 ;
        RECT 8.110 0.885 9.140 1.215 ;
        RECT 7.280 0.355 7.870 0.670 ;
        RECT 9.730 0.625 10.060 1.215 ;
        RECT 8.040 0.255 10.420 0.625 ;
        RECT 0.000 -0.085 11.040 0.085 ;
  END
END sky130_fd_sc_hvl__sdlclkp_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__sdlxtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__sdlxtp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.520 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.585000 ;
    PORT
      LAYER li1 ;
        RECT 2.040 2.185 2.370 3.260 ;
    END
  END D
  PIN GATE
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.585000 ;
    PORT
      LAYER li1 ;
        RECT 4.370 1.145 4.665 2.495 ;
    END
  END GATE
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.585000 ;
    PORT
      LAYER li1 ;
        RECT 3.515 1.525 3.860 2.495 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.005000 ;
    PORT
      LAYER li1 ;
        RECT 0.585 2.005 1.795 2.775 ;
        RECT 0.585 1.835 2.770 2.005 ;
        RECT 2.600 1.695 2.770 1.835 ;
        RECT 2.600 1.445 2.985 1.695 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 11.520 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 9.325 1.085 11.490 1.415 ;
        RECT 0.040 0.215 11.490 1.085 ;
        RECT -0.130 -0.215 11.650 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 11.520 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 11.850 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 11.520 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 11.520 3.815 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.626250 ;
    PORT
      LAYER li1 ;
        RECT 11.060 0.515 11.400 3.755 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 11.520 4.155 ;
        RECT 0.130 1.345 0.380 3.395 ;
        RECT 0.560 2.995 1.510 3.705 ;
        RECT 2.575 2.845 2.825 3.725 ;
        RECT 3.365 3.025 4.315 3.725 ;
        RECT 4.495 3.635 5.365 3.805 ;
        RECT 4.495 2.845 4.665 3.635 ;
        RECT 2.575 2.675 4.665 2.845 ;
        RECT 2.950 1.905 3.335 2.495 ;
        RECT 1.965 1.345 2.295 1.655 ;
        RECT 0.130 1.265 2.295 1.345 ;
        RECT 3.165 1.265 3.335 1.905 ;
        RECT 4.030 1.345 4.200 2.675 ;
        RECT 0.130 1.175 3.335 1.265 ;
        RECT 0.130 0.495 0.480 1.175 ;
        RECT 1.965 1.095 3.335 1.175 ;
        RECT 3.515 1.175 4.200 1.345 ;
        RECT 4.845 1.345 5.015 3.455 ;
        RECT 5.195 2.405 5.365 3.635 ;
        RECT 5.545 2.585 5.715 3.705 ;
        RECT 5.895 3.595 7.250 3.765 ;
        RECT 5.895 2.405 6.065 3.595 ;
        RECT 5.195 2.235 6.065 2.405 ;
        RECT 6.245 2.585 6.575 3.415 ;
        RECT 6.755 2.925 7.250 3.595 ;
        RECT 7.700 2.925 8.030 3.755 ;
        RECT 8.685 3.005 9.635 3.705 ;
        RECT 5.590 1.345 5.920 1.845 ;
        RECT 4.845 1.175 5.920 1.345 ;
        RECT 0.660 0.365 1.610 0.995 ;
        RECT 3.515 0.915 3.685 1.175 ;
        RECT 4.845 0.975 5.015 1.175 ;
        RECT 2.420 0.745 3.685 0.915 ;
        RECT 2.420 0.495 2.750 0.745 ;
        RECT 3.865 0.365 4.455 0.975 ;
        RECT 4.695 0.515 5.025 0.975 ;
        RECT 5.205 0.365 5.795 0.995 ;
        RECT 6.245 0.975 6.415 2.585 ;
        RECT 6.755 0.975 6.925 2.925 ;
        RECT 7.860 2.825 8.030 2.925 ;
        RECT 7.860 2.655 8.920 2.825 ;
        RECT 7.840 2.215 8.570 2.475 ;
        RECT 7.840 1.755 8.010 2.215 ;
        RECT 8.750 2.005 8.920 2.655 ;
        RECT 9.385 2.355 9.715 2.675 ;
        RECT 9.895 2.535 10.845 3.755 ;
        RECT 9.385 2.185 10.550 2.355 ;
        RECT 6.045 0.435 6.415 0.975 ;
        RECT 6.595 0.615 6.925 0.975 ;
        RECT 7.105 1.585 8.010 1.755 ;
        RECT 8.190 1.835 10.200 2.005 ;
        RECT 7.105 0.435 7.275 1.585 ;
        RECT 8.190 1.245 8.360 1.835 ;
        RECT 9.870 1.755 10.200 1.835 ;
        RECT 7.455 1.075 8.360 1.245 ;
        RECT 8.540 1.575 8.870 1.655 ;
        RECT 10.380 1.575 10.550 2.185 ;
        RECT 8.540 1.405 10.550 1.575 ;
        RECT 8.540 1.075 8.870 1.405 ;
        RECT 7.455 0.495 7.705 1.075 ;
        RECT 6.045 0.265 7.275 0.435 ;
        RECT 8.245 0.365 9.195 0.895 ;
        RECT 9.415 0.845 9.745 1.405 ;
        RECT 9.925 0.365 10.875 1.225 ;
        RECT 0.000 -0.085 11.520 0.085 ;
  END
END sky130_fd_sc_hvl__sdlxtp_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__xnor2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__xnor2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.280 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.250000 ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.580 2.060 1.750 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.250000 ;
    PORT
      LAYER li1 ;
        RECT 1.565 2.100 3.255 2.120 ;
        RECT 0.575 1.930 3.255 2.100 ;
        RECT 0.575 1.725 0.905 1.930 ;
        RECT 2.925 1.805 3.255 1.930 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 5.280 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 3.860 1.415 5.190 1.455 ;
        RECT 0.020 0.215 5.190 1.415 ;
        RECT -0.130 -0.215 5.410 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 5.280 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 5.610 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 5.280 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 5.280 3.815 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.481250 ;
    PORT
      LAYER li1 ;
        RECT 4.025 2.075 4.275 3.755 ;
        RECT 4.025 1.905 5.155 2.075 ;
        RECT 4.445 1.545 5.155 1.905 ;
        RECT 4.750 0.535 5.155 1.545 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 5.280 4.155 ;
        RECT 0.090 2.630 0.985 3.755 ;
        RECT 1.165 2.450 1.335 3.755 ;
        RECT 0.110 2.280 1.335 2.450 ;
        RECT 1.515 2.300 3.845 3.755 ;
        RECT 0.110 1.400 0.360 2.280 ;
        RECT 4.465 2.255 5.055 3.755 ;
        RECT 3.650 1.625 3.980 1.725 ;
        RECT 2.240 1.455 3.980 1.625 ;
        RECT 2.240 1.400 2.410 1.455 ;
        RECT 0.110 1.230 2.410 1.400 ;
        RECT 0.110 0.495 0.440 1.230 ;
        RECT 2.590 1.105 4.300 1.285 ;
        RECT 0.610 0.365 2.410 1.050 ;
        RECT 2.590 0.495 2.920 1.105 ;
        RECT 3.100 0.365 3.630 0.925 ;
        RECT 3.970 0.535 4.300 1.105 ;
        RECT 0.000 -0.085 5.280 0.085 ;
  END
END sky130_fd_sc_hvl__xnor2_1

#--------EOF---------

MACRO sky130_fd_sc_hvl__xor2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__xor2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.280 BY 4.070 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.250000 ;
    PORT
      LAYER li1 ;
        RECT 2.045 1.775 3.235 2.150 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.250000 ;
    PORT
      LAYER li1 ;
        RECT 0.560 1.775 1.510 2.055 ;
        RECT 1.340 1.595 1.510 1.775 ;
        RECT 3.415 1.595 3.715 1.835 ;
        RECT 1.340 1.505 3.715 1.595 ;
        RECT 1.340 1.425 3.585 1.505 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000 0.255 5.280 0.625 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.020 0.215 4.990 1.415 ;
        RECT -0.130 -0.215 5.410 0.215 ;
      LAYER met1 ;
        RECT 0.000 -0.115 5.280 0.115 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.330 1.885 5.610 4.485 ;
      LAYER met1 ;
        RECT 0.000 3.955 5.280 4.185 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000 3.445 5.280 3.815 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.637500 ;
    PORT
      LAYER li1 ;
        RECT 3.965 1.325 4.370 2.425 ;
        RECT 3.850 0.495 4.370 1.325 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 3.985 5.280 4.155 ;
        RECT 0.130 2.605 0.380 3.755 ;
        RECT 0.560 2.785 2.530 3.755 ;
        RECT 2.710 3.125 2.880 3.755 ;
        RECT 3.060 3.305 4.720 3.755 ;
        RECT 4.900 3.125 5.150 3.755 ;
        RECT 2.710 2.955 5.150 3.125 ;
        RECT 2.710 2.785 2.880 2.955 ;
        RECT 3.060 2.605 4.720 2.775 ;
        RECT 0.130 2.435 3.230 2.605 ;
        RECT 0.130 1.595 0.380 2.435 ;
        RECT 4.550 1.995 4.720 2.605 ;
        RECT 4.900 2.175 5.150 2.955 ;
        RECT 4.550 1.665 4.880 1.995 ;
        RECT 0.130 1.425 1.160 1.595 ;
        RECT 0.090 0.365 0.680 1.245 ;
        RECT 0.910 0.495 1.160 1.425 ;
        RECT 1.340 0.365 3.670 1.245 ;
        RECT 4.550 0.365 5.140 1.325 ;
        RECT 0.000 -0.085 5.280 0.085 ;
  END
END sky130_fd_sc_hvl__xor2_1

#--------EOF---------


END LIBRARY
