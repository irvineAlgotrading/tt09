magic
tech sky130B
timestamp 1704896540
<< metal1 >>
rect 0 0 3 3418
rect 285 0 288 3418
<< via1 >>
rect 3 0 285 3418
<< metal2 >>
rect 0 0 3 3418
rect 285 0 288 3418
<< properties >>
string GDS_END 93836708
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 93774944
<< end >>
