magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< pwell >>
rect 896 -5162 1566 5162
<< mvpsubdiff >>
rect 922 5124 1540 5136
rect 922 5090 1113 5124
rect 1147 5090 1181 5124
rect 1215 5090 1249 5124
rect 1283 5090 1317 5124
rect 1351 5090 1540 5124
rect 922 5078 1540 5090
rect 922 5015 1054 5078
rect 922 4981 938 5015
rect 972 4981 1008 5015
rect 1042 4981 1054 5015
rect 1410 5015 1540 5078
rect 922 4947 1054 4981
rect 922 4913 938 4947
rect 972 4913 1008 4947
rect 1042 4913 1054 4947
rect 922 4879 1054 4913
rect 922 4845 938 4879
rect 972 4845 1008 4879
rect 1042 4845 1054 4879
rect 922 4811 1054 4845
rect 922 4777 938 4811
rect 972 4777 1008 4811
rect 1042 4777 1054 4811
rect 922 4743 1054 4777
rect 922 4709 938 4743
rect 972 4709 1008 4743
rect 1042 4709 1054 4743
rect 922 4675 1054 4709
rect 922 4641 938 4675
rect 972 4641 1008 4675
rect 1042 4641 1054 4675
rect 922 4607 1054 4641
rect 922 4573 938 4607
rect 972 4573 1008 4607
rect 1042 4573 1054 4607
rect 922 4539 1054 4573
rect 922 4505 938 4539
rect 972 4505 1008 4539
rect 1042 4505 1054 4539
rect 922 4471 1054 4505
rect 922 4437 938 4471
rect 972 4437 1008 4471
rect 1042 4437 1054 4471
rect 922 4403 1054 4437
rect 922 4369 938 4403
rect 972 4369 1008 4403
rect 1042 4369 1054 4403
rect 922 4335 1054 4369
rect 922 4301 938 4335
rect 972 4301 1008 4335
rect 1042 4301 1054 4335
rect 922 4267 1054 4301
rect 922 4233 938 4267
rect 972 4233 1008 4267
rect 1042 4233 1054 4267
rect 922 4199 1054 4233
rect 922 4165 938 4199
rect 972 4165 1008 4199
rect 1042 4165 1054 4199
rect 922 4131 1054 4165
rect 922 4097 938 4131
rect 972 4097 1008 4131
rect 1042 4097 1054 4131
rect 922 4063 1054 4097
rect 922 4029 938 4063
rect 972 4029 1008 4063
rect 1042 4029 1054 4063
rect 922 3995 1054 4029
rect 922 3961 938 3995
rect 972 3961 1008 3995
rect 1042 3961 1054 3995
rect 922 3927 1054 3961
rect 922 3893 938 3927
rect 972 3893 1008 3927
rect 1042 3893 1054 3927
rect 922 3859 1054 3893
rect 922 3825 938 3859
rect 972 3825 1008 3859
rect 1042 3825 1054 3859
rect 922 3791 1054 3825
rect 922 3757 938 3791
rect 972 3757 1008 3791
rect 1042 3757 1054 3791
rect 922 3723 1054 3757
rect 922 3689 938 3723
rect 972 3689 1008 3723
rect 1042 3689 1054 3723
rect 922 3655 1054 3689
rect 922 3621 938 3655
rect 972 3621 1008 3655
rect 1042 3621 1054 3655
rect 922 3587 1054 3621
rect 922 3553 938 3587
rect 972 3553 1008 3587
rect 1042 3553 1054 3587
rect 922 3519 1054 3553
rect 922 3485 938 3519
rect 972 3485 1008 3519
rect 1042 3485 1054 3519
rect 922 3451 1054 3485
rect 922 3417 938 3451
rect 972 3417 1008 3451
rect 1042 3417 1054 3451
rect 922 3383 1054 3417
rect 922 3349 938 3383
rect 972 3349 1008 3383
rect 1042 3349 1054 3383
rect 922 3315 1054 3349
rect 922 3281 938 3315
rect 972 3281 1008 3315
rect 1042 3281 1054 3315
rect 922 3247 1054 3281
rect 922 3213 938 3247
rect 972 3213 1008 3247
rect 1042 3213 1054 3247
rect 922 3179 1054 3213
rect 922 3145 938 3179
rect 972 3145 1008 3179
rect 1042 3145 1054 3179
rect 922 3111 1054 3145
rect 922 3077 938 3111
rect 972 3077 1008 3111
rect 1042 3077 1054 3111
rect 922 3043 1054 3077
rect 922 3009 938 3043
rect 972 3009 1008 3043
rect 1042 3009 1054 3043
rect 922 2975 1054 3009
rect 922 2941 938 2975
rect 972 2941 1008 2975
rect 1042 2941 1054 2975
rect 922 2907 1054 2941
rect 922 2873 938 2907
rect 972 2873 1008 2907
rect 1042 2873 1054 2907
rect 922 2839 1054 2873
rect 922 2805 938 2839
rect 972 2805 1008 2839
rect 1042 2805 1054 2839
rect 922 2771 1054 2805
rect 922 2737 938 2771
rect 972 2737 1008 2771
rect 1042 2737 1054 2771
rect 922 2703 1054 2737
rect 922 2669 938 2703
rect 972 2669 1008 2703
rect 1042 2669 1054 2703
rect 922 2635 1054 2669
rect 922 2601 938 2635
rect 972 2601 1008 2635
rect 1042 2601 1054 2635
rect 922 2567 1054 2601
rect 922 2533 938 2567
rect 972 2533 1008 2567
rect 1042 2533 1054 2567
rect 922 2499 1054 2533
rect 922 2465 938 2499
rect 972 2465 1008 2499
rect 1042 2465 1054 2499
rect 922 2431 1054 2465
rect 922 2397 938 2431
rect 972 2397 1008 2431
rect 1042 2397 1054 2431
rect 922 2363 1054 2397
rect 922 2329 938 2363
rect 972 2329 1008 2363
rect 1042 2329 1054 2363
rect 922 2295 1054 2329
rect 922 2261 938 2295
rect 972 2261 1008 2295
rect 1042 2261 1054 2295
rect 922 2227 1054 2261
rect 922 2193 938 2227
rect 972 2193 1008 2227
rect 1042 2193 1054 2227
rect 922 2159 1054 2193
rect 922 2125 938 2159
rect 972 2125 1008 2159
rect 1042 2125 1054 2159
rect 922 2091 1054 2125
rect 922 2057 938 2091
rect 972 2057 1008 2091
rect 1042 2057 1054 2091
rect 922 2023 1054 2057
rect 922 1989 938 2023
rect 972 1989 1008 2023
rect 1042 1989 1054 2023
rect 922 1955 1054 1989
rect 922 1921 938 1955
rect 972 1921 1008 1955
rect 1042 1921 1054 1955
rect 922 1887 1054 1921
rect 922 1853 938 1887
rect 972 1853 1008 1887
rect 1042 1853 1054 1887
rect 922 1819 1054 1853
rect 922 1785 938 1819
rect 972 1785 1008 1819
rect 1042 1785 1054 1819
rect 922 1751 1054 1785
rect 922 1717 938 1751
rect 972 1717 1008 1751
rect 1042 1717 1054 1751
rect 922 1683 1054 1717
rect 922 1649 938 1683
rect 972 1649 1008 1683
rect 1042 1649 1054 1683
rect 922 1615 1054 1649
rect 922 1581 938 1615
rect 972 1581 1008 1615
rect 1042 1581 1054 1615
rect 922 1547 1054 1581
rect 922 1513 938 1547
rect 972 1513 1008 1547
rect 1042 1513 1054 1547
rect 922 1479 1054 1513
rect 922 1445 938 1479
rect 972 1445 1008 1479
rect 1042 1445 1054 1479
rect 922 1411 1054 1445
rect 922 1377 938 1411
rect 972 1377 1008 1411
rect 1042 1377 1054 1411
rect 922 1343 1054 1377
rect 922 1309 938 1343
rect 972 1309 1008 1343
rect 1042 1309 1054 1343
rect 922 1275 1054 1309
rect 922 1241 938 1275
rect 972 1241 1008 1275
rect 1042 1241 1054 1275
rect 922 1207 1054 1241
rect 922 1173 938 1207
rect 972 1173 1008 1207
rect 1042 1173 1054 1207
rect 922 1139 1054 1173
rect 922 1105 938 1139
rect 972 1105 1008 1139
rect 1042 1105 1054 1139
rect 922 1071 1054 1105
rect 922 1037 938 1071
rect 972 1037 1008 1071
rect 1042 1037 1054 1071
rect 922 1003 1054 1037
rect 922 969 938 1003
rect 972 969 1008 1003
rect 1042 969 1054 1003
rect 922 935 1054 969
rect 922 901 938 935
rect 972 901 1008 935
rect 1042 901 1054 935
rect 922 867 1054 901
rect 922 833 938 867
rect 972 833 1008 867
rect 1042 833 1054 867
rect 922 799 1054 833
rect 922 765 938 799
rect 972 765 1008 799
rect 1042 765 1054 799
rect 922 731 1054 765
rect 922 697 938 731
rect 972 697 1008 731
rect 1042 697 1054 731
rect 922 663 1054 697
rect 922 629 938 663
rect 972 629 1008 663
rect 1042 629 1054 663
rect 922 595 1054 629
rect 922 561 938 595
rect 972 561 1008 595
rect 1042 561 1054 595
rect 922 527 1054 561
rect 922 493 938 527
rect 972 493 1008 527
rect 1042 493 1054 527
rect 922 459 1054 493
rect 922 425 938 459
rect 972 425 1008 459
rect 1042 425 1054 459
rect 922 391 1054 425
rect 922 357 938 391
rect 972 357 1008 391
rect 1042 357 1054 391
rect 922 323 1054 357
rect 922 289 938 323
rect 972 289 1008 323
rect 1042 289 1054 323
rect 922 255 1054 289
rect 922 221 938 255
rect 972 221 1008 255
rect 1042 221 1054 255
rect 922 187 1054 221
rect 922 153 938 187
rect 972 153 1008 187
rect 1042 153 1054 187
rect 922 119 1054 153
rect 922 85 938 119
rect 972 85 1008 119
rect 1042 85 1054 119
rect 922 51 1054 85
rect 922 17 938 51
rect 972 17 1008 51
rect 1042 17 1054 51
rect 922 -17 1054 17
rect 922 -51 938 -17
rect 972 -51 1008 -17
rect 1042 -51 1054 -17
rect 922 -85 1054 -51
rect 922 -119 938 -85
rect 972 -119 1008 -85
rect 1042 -119 1054 -85
rect 922 -153 1054 -119
rect 922 -187 938 -153
rect 972 -187 1008 -153
rect 1042 -187 1054 -153
rect 922 -221 1054 -187
rect 922 -255 938 -221
rect 972 -255 1008 -221
rect 1042 -255 1054 -221
rect 922 -289 1054 -255
rect 922 -323 938 -289
rect 972 -323 1008 -289
rect 1042 -323 1054 -289
rect 922 -357 1054 -323
rect 922 -391 938 -357
rect 972 -391 1008 -357
rect 1042 -391 1054 -357
rect 922 -425 1054 -391
rect 922 -459 938 -425
rect 972 -459 1008 -425
rect 1042 -459 1054 -425
rect 922 -493 1054 -459
rect 922 -527 938 -493
rect 972 -527 1008 -493
rect 1042 -527 1054 -493
rect 922 -561 1054 -527
rect 922 -595 938 -561
rect 972 -595 1008 -561
rect 1042 -595 1054 -561
rect 922 -629 1054 -595
rect 922 -663 938 -629
rect 972 -663 1008 -629
rect 1042 -663 1054 -629
rect 922 -697 1054 -663
rect 922 -731 938 -697
rect 972 -731 1008 -697
rect 1042 -731 1054 -697
rect 922 -765 1054 -731
rect 922 -799 938 -765
rect 972 -799 1008 -765
rect 1042 -799 1054 -765
rect 922 -833 1054 -799
rect 922 -867 938 -833
rect 972 -867 1008 -833
rect 1042 -867 1054 -833
rect 922 -901 1054 -867
rect 922 -935 938 -901
rect 972 -935 1008 -901
rect 1042 -935 1054 -901
rect 922 -969 1054 -935
rect 922 -1003 938 -969
rect 972 -1003 1008 -969
rect 1042 -1003 1054 -969
rect 922 -1037 1054 -1003
rect 922 -1071 938 -1037
rect 972 -1071 1008 -1037
rect 1042 -1071 1054 -1037
rect 922 -1105 1054 -1071
rect 922 -1139 938 -1105
rect 972 -1139 1008 -1105
rect 1042 -1139 1054 -1105
rect 922 -1173 1054 -1139
rect 922 -1207 938 -1173
rect 972 -1207 1008 -1173
rect 1042 -1207 1054 -1173
rect 922 -1241 1054 -1207
rect 922 -1275 938 -1241
rect 972 -1275 1008 -1241
rect 1042 -1275 1054 -1241
rect 922 -1309 1054 -1275
rect 922 -1343 938 -1309
rect 972 -1343 1008 -1309
rect 1042 -1343 1054 -1309
rect 922 -1377 1054 -1343
rect 922 -1411 938 -1377
rect 972 -1411 1008 -1377
rect 1042 -1411 1054 -1377
rect 922 -1445 1054 -1411
rect 922 -1479 938 -1445
rect 972 -1479 1008 -1445
rect 1042 -1479 1054 -1445
rect 922 -1513 1054 -1479
rect 922 -1547 938 -1513
rect 972 -1547 1008 -1513
rect 1042 -1547 1054 -1513
rect 922 -1581 1054 -1547
rect 922 -1615 938 -1581
rect 972 -1615 1008 -1581
rect 1042 -1615 1054 -1581
rect 922 -1649 1054 -1615
rect 922 -1683 938 -1649
rect 972 -1683 1008 -1649
rect 1042 -1683 1054 -1649
rect 922 -1717 1054 -1683
rect 922 -1751 938 -1717
rect 972 -1751 1008 -1717
rect 1042 -1751 1054 -1717
rect 922 -1785 1054 -1751
rect 922 -1819 938 -1785
rect 972 -1819 1008 -1785
rect 1042 -1819 1054 -1785
rect 922 -1853 1054 -1819
rect 922 -1887 938 -1853
rect 972 -1887 1008 -1853
rect 1042 -1887 1054 -1853
rect 922 -1921 1054 -1887
rect 922 -1955 938 -1921
rect 972 -1955 1008 -1921
rect 1042 -1955 1054 -1921
rect 922 -1989 1054 -1955
rect 922 -2023 938 -1989
rect 972 -2023 1008 -1989
rect 1042 -2023 1054 -1989
rect 922 -2057 1054 -2023
rect 922 -2091 938 -2057
rect 972 -2091 1008 -2057
rect 1042 -2091 1054 -2057
rect 922 -2125 1054 -2091
rect 922 -2159 938 -2125
rect 972 -2159 1008 -2125
rect 1042 -2159 1054 -2125
rect 922 -2193 1054 -2159
rect 922 -2227 938 -2193
rect 972 -2227 1008 -2193
rect 1042 -2227 1054 -2193
rect 922 -2261 1054 -2227
rect 922 -2295 938 -2261
rect 972 -2295 1008 -2261
rect 1042 -2295 1054 -2261
rect 922 -2329 1054 -2295
rect 922 -2363 938 -2329
rect 972 -2363 1008 -2329
rect 1042 -2363 1054 -2329
rect 922 -2397 1054 -2363
rect 922 -2431 938 -2397
rect 972 -2431 1008 -2397
rect 1042 -2431 1054 -2397
rect 922 -2465 1054 -2431
rect 922 -2499 938 -2465
rect 972 -2499 1008 -2465
rect 1042 -2499 1054 -2465
rect 922 -2533 1054 -2499
rect 922 -2567 938 -2533
rect 972 -2567 1008 -2533
rect 1042 -2567 1054 -2533
rect 922 -2601 1054 -2567
rect 922 -2635 938 -2601
rect 972 -2635 1008 -2601
rect 1042 -2635 1054 -2601
rect 922 -2669 1054 -2635
rect 922 -2703 938 -2669
rect 972 -2703 1008 -2669
rect 1042 -2703 1054 -2669
rect 922 -2737 1054 -2703
rect 922 -2771 938 -2737
rect 972 -2771 1008 -2737
rect 1042 -2771 1054 -2737
rect 922 -2805 1054 -2771
rect 922 -2839 938 -2805
rect 972 -2839 1008 -2805
rect 1042 -2839 1054 -2805
rect 922 -2873 1054 -2839
rect 922 -2907 938 -2873
rect 972 -2907 1008 -2873
rect 1042 -2907 1054 -2873
rect 922 -2941 1054 -2907
rect 922 -2975 938 -2941
rect 972 -2975 1008 -2941
rect 1042 -2975 1054 -2941
rect 922 -3009 1054 -2975
rect 922 -3043 938 -3009
rect 972 -3043 1008 -3009
rect 1042 -3043 1054 -3009
rect 922 -3077 1054 -3043
rect 922 -3111 938 -3077
rect 972 -3111 1008 -3077
rect 1042 -3111 1054 -3077
rect 922 -3145 1054 -3111
rect 922 -3179 938 -3145
rect 972 -3179 1008 -3145
rect 1042 -3179 1054 -3145
rect 922 -3213 1054 -3179
rect 922 -3247 938 -3213
rect 972 -3247 1008 -3213
rect 1042 -3247 1054 -3213
rect 922 -3281 1054 -3247
rect 922 -3315 938 -3281
rect 972 -3315 1008 -3281
rect 1042 -3315 1054 -3281
rect 922 -3349 1054 -3315
rect 922 -3383 938 -3349
rect 972 -3383 1008 -3349
rect 1042 -3383 1054 -3349
rect 922 -3417 1054 -3383
rect 922 -3451 938 -3417
rect 972 -3451 1008 -3417
rect 1042 -3451 1054 -3417
rect 922 -3485 1054 -3451
rect 922 -3519 938 -3485
rect 972 -3519 1008 -3485
rect 1042 -3519 1054 -3485
rect 922 -3553 1054 -3519
rect 922 -3587 938 -3553
rect 972 -3587 1008 -3553
rect 1042 -3587 1054 -3553
rect 922 -3621 1054 -3587
rect 922 -3655 938 -3621
rect 972 -3655 1008 -3621
rect 1042 -3655 1054 -3621
rect 922 -3689 1054 -3655
rect 922 -3723 938 -3689
rect 972 -3723 1008 -3689
rect 1042 -3723 1054 -3689
rect 922 -3757 1054 -3723
rect 922 -3791 938 -3757
rect 972 -3791 1008 -3757
rect 1042 -3791 1054 -3757
rect 922 -3825 1054 -3791
rect 922 -3859 938 -3825
rect 972 -3859 1008 -3825
rect 1042 -3859 1054 -3825
rect 922 -3893 1054 -3859
rect 922 -3927 938 -3893
rect 972 -3927 1008 -3893
rect 1042 -3927 1054 -3893
rect 922 -3961 1054 -3927
rect 922 -3995 938 -3961
rect 972 -3995 1008 -3961
rect 1042 -3995 1054 -3961
rect 922 -4029 1054 -3995
rect 922 -4063 938 -4029
rect 972 -4063 1008 -4029
rect 1042 -4063 1054 -4029
rect 922 -4097 1054 -4063
rect 922 -4131 938 -4097
rect 972 -4131 1008 -4097
rect 1042 -4131 1054 -4097
rect 922 -4165 1054 -4131
rect 922 -4199 938 -4165
rect 972 -4199 1008 -4165
rect 1042 -4199 1054 -4165
rect 922 -4233 1054 -4199
rect 922 -4267 938 -4233
rect 972 -4267 1008 -4233
rect 1042 -4267 1054 -4233
rect 922 -4301 1054 -4267
rect 922 -4335 938 -4301
rect 972 -4335 1008 -4301
rect 1042 -4335 1054 -4301
rect 922 -4369 1054 -4335
rect 922 -4403 938 -4369
rect 972 -4403 1008 -4369
rect 1042 -4403 1054 -4369
rect 922 -4437 1054 -4403
rect 922 -4471 938 -4437
rect 972 -4471 1008 -4437
rect 1042 -4471 1054 -4437
rect 922 -4505 1054 -4471
rect 922 -4539 938 -4505
rect 972 -4539 1008 -4505
rect 1042 -4539 1054 -4505
rect 922 -4573 1054 -4539
rect 922 -4607 938 -4573
rect 972 -4607 1008 -4573
rect 1042 -4607 1054 -4573
rect 922 -4641 1054 -4607
rect 922 -4675 938 -4641
rect 972 -4675 1008 -4641
rect 1042 -4675 1054 -4641
rect 922 -4709 1054 -4675
rect 922 -4743 938 -4709
rect 972 -4743 1008 -4709
rect 1042 -4743 1054 -4709
rect 922 -4777 1054 -4743
rect 922 -4811 938 -4777
rect 972 -4811 1008 -4777
rect 1042 -4811 1054 -4777
rect 922 -4845 1054 -4811
rect 922 -4879 938 -4845
rect 972 -4879 1008 -4845
rect 1042 -4879 1054 -4845
rect 922 -4913 1054 -4879
rect 922 -4947 938 -4913
rect 972 -4947 1008 -4913
rect 1042 -4947 1054 -4913
rect 922 -4981 1054 -4947
rect 922 -5015 938 -4981
rect 972 -5015 1008 -4981
rect 1042 -5015 1054 -4981
rect 922 -5078 1054 -5015
rect 1410 -5015 1422 5015
rect 1524 -5015 1540 5015
rect 1410 -5078 1540 -5015
rect 922 -5090 1540 -5078
rect 922 -5124 1113 -5090
rect 1147 -5124 1181 -5090
rect 1215 -5124 1249 -5090
rect 1283 -5124 1317 -5090
rect 1351 -5124 1540 -5090
rect 922 -5136 1540 -5124
<< mvpsubdiffcont >>
rect 1113 5090 1147 5124
rect 1181 5090 1215 5124
rect 1249 5090 1283 5124
rect 1317 5090 1351 5124
rect 938 4981 972 5015
rect 1008 4981 1042 5015
rect 938 4913 972 4947
rect 1008 4913 1042 4947
rect 938 4845 972 4879
rect 1008 4845 1042 4879
rect 938 4777 972 4811
rect 1008 4777 1042 4811
rect 938 4709 972 4743
rect 1008 4709 1042 4743
rect 938 4641 972 4675
rect 1008 4641 1042 4675
rect 938 4573 972 4607
rect 1008 4573 1042 4607
rect 938 4505 972 4539
rect 1008 4505 1042 4539
rect 938 4437 972 4471
rect 1008 4437 1042 4471
rect 938 4369 972 4403
rect 1008 4369 1042 4403
rect 938 4301 972 4335
rect 1008 4301 1042 4335
rect 938 4233 972 4267
rect 1008 4233 1042 4267
rect 938 4165 972 4199
rect 1008 4165 1042 4199
rect 938 4097 972 4131
rect 1008 4097 1042 4131
rect 938 4029 972 4063
rect 1008 4029 1042 4063
rect 938 3961 972 3995
rect 1008 3961 1042 3995
rect 938 3893 972 3927
rect 1008 3893 1042 3927
rect 938 3825 972 3859
rect 1008 3825 1042 3859
rect 938 3757 972 3791
rect 1008 3757 1042 3791
rect 938 3689 972 3723
rect 1008 3689 1042 3723
rect 938 3621 972 3655
rect 1008 3621 1042 3655
rect 938 3553 972 3587
rect 1008 3553 1042 3587
rect 938 3485 972 3519
rect 1008 3485 1042 3519
rect 938 3417 972 3451
rect 1008 3417 1042 3451
rect 938 3349 972 3383
rect 1008 3349 1042 3383
rect 938 3281 972 3315
rect 1008 3281 1042 3315
rect 938 3213 972 3247
rect 1008 3213 1042 3247
rect 938 3145 972 3179
rect 1008 3145 1042 3179
rect 938 3077 972 3111
rect 1008 3077 1042 3111
rect 938 3009 972 3043
rect 1008 3009 1042 3043
rect 938 2941 972 2975
rect 1008 2941 1042 2975
rect 938 2873 972 2907
rect 1008 2873 1042 2907
rect 938 2805 972 2839
rect 1008 2805 1042 2839
rect 938 2737 972 2771
rect 1008 2737 1042 2771
rect 938 2669 972 2703
rect 1008 2669 1042 2703
rect 938 2601 972 2635
rect 1008 2601 1042 2635
rect 938 2533 972 2567
rect 1008 2533 1042 2567
rect 938 2465 972 2499
rect 1008 2465 1042 2499
rect 938 2397 972 2431
rect 1008 2397 1042 2431
rect 938 2329 972 2363
rect 1008 2329 1042 2363
rect 938 2261 972 2295
rect 1008 2261 1042 2295
rect 938 2193 972 2227
rect 1008 2193 1042 2227
rect 938 2125 972 2159
rect 1008 2125 1042 2159
rect 938 2057 972 2091
rect 1008 2057 1042 2091
rect 938 1989 972 2023
rect 1008 1989 1042 2023
rect 938 1921 972 1955
rect 1008 1921 1042 1955
rect 938 1853 972 1887
rect 1008 1853 1042 1887
rect 938 1785 972 1819
rect 1008 1785 1042 1819
rect 938 1717 972 1751
rect 1008 1717 1042 1751
rect 938 1649 972 1683
rect 1008 1649 1042 1683
rect 938 1581 972 1615
rect 1008 1581 1042 1615
rect 938 1513 972 1547
rect 1008 1513 1042 1547
rect 938 1445 972 1479
rect 1008 1445 1042 1479
rect 938 1377 972 1411
rect 1008 1377 1042 1411
rect 938 1309 972 1343
rect 1008 1309 1042 1343
rect 938 1241 972 1275
rect 1008 1241 1042 1275
rect 938 1173 972 1207
rect 1008 1173 1042 1207
rect 938 1105 972 1139
rect 1008 1105 1042 1139
rect 938 1037 972 1071
rect 1008 1037 1042 1071
rect 938 969 972 1003
rect 1008 969 1042 1003
rect 938 901 972 935
rect 1008 901 1042 935
rect 938 833 972 867
rect 1008 833 1042 867
rect 938 765 972 799
rect 1008 765 1042 799
rect 938 697 972 731
rect 1008 697 1042 731
rect 938 629 972 663
rect 1008 629 1042 663
rect 938 561 972 595
rect 1008 561 1042 595
rect 938 493 972 527
rect 1008 493 1042 527
rect 938 425 972 459
rect 1008 425 1042 459
rect 938 357 972 391
rect 1008 357 1042 391
rect 938 289 972 323
rect 1008 289 1042 323
rect 938 221 972 255
rect 1008 221 1042 255
rect 938 153 972 187
rect 1008 153 1042 187
rect 938 85 972 119
rect 1008 85 1042 119
rect 938 17 972 51
rect 1008 17 1042 51
rect 938 -51 972 -17
rect 1008 -51 1042 -17
rect 938 -119 972 -85
rect 1008 -119 1042 -85
rect 938 -187 972 -153
rect 1008 -187 1042 -153
rect 938 -255 972 -221
rect 1008 -255 1042 -221
rect 938 -323 972 -289
rect 1008 -323 1042 -289
rect 938 -391 972 -357
rect 1008 -391 1042 -357
rect 938 -459 972 -425
rect 1008 -459 1042 -425
rect 938 -527 972 -493
rect 1008 -527 1042 -493
rect 938 -595 972 -561
rect 1008 -595 1042 -561
rect 938 -663 972 -629
rect 1008 -663 1042 -629
rect 938 -731 972 -697
rect 1008 -731 1042 -697
rect 938 -799 972 -765
rect 1008 -799 1042 -765
rect 938 -867 972 -833
rect 1008 -867 1042 -833
rect 938 -935 972 -901
rect 1008 -935 1042 -901
rect 938 -1003 972 -969
rect 1008 -1003 1042 -969
rect 938 -1071 972 -1037
rect 1008 -1071 1042 -1037
rect 938 -1139 972 -1105
rect 1008 -1139 1042 -1105
rect 938 -1207 972 -1173
rect 1008 -1207 1042 -1173
rect 938 -1275 972 -1241
rect 1008 -1275 1042 -1241
rect 938 -1343 972 -1309
rect 1008 -1343 1042 -1309
rect 938 -1411 972 -1377
rect 1008 -1411 1042 -1377
rect 938 -1479 972 -1445
rect 1008 -1479 1042 -1445
rect 938 -1547 972 -1513
rect 1008 -1547 1042 -1513
rect 938 -1615 972 -1581
rect 1008 -1615 1042 -1581
rect 938 -1683 972 -1649
rect 1008 -1683 1042 -1649
rect 938 -1751 972 -1717
rect 1008 -1751 1042 -1717
rect 938 -1819 972 -1785
rect 1008 -1819 1042 -1785
rect 938 -1887 972 -1853
rect 1008 -1887 1042 -1853
rect 938 -1955 972 -1921
rect 1008 -1955 1042 -1921
rect 938 -2023 972 -1989
rect 1008 -2023 1042 -1989
rect 938 -2091 972 -2057
rect 1008 -2091 1042 -2057
rect 938 -2159 972 -2125
rect 1008 -2159 1042 -2125
rect 938 -2227 972 -2193
rect 1008 -2227 1042 -2193
rect 938 -2295 972 -2261
rect 1008 -2295 1042 -2261
rect 938 -2363 972 -2329
rect 1008 -2363 1042 -2329
rect 938 -2431 972 -2397
rect 1008 -2431 1042 -2397
rect 938 -2499 972 -2465
rect 1008 -2499 1042 -2465
rect 938 -2567 972 -2533
rect 1008 -2567 1042 -2533
rect 938 -2635 972 -2601
rect 1008 -2635 1042 -2601
rect 938 -2703 972 -2669
rect 1008 -2703 1042 -2669
rect 938 -2771 972 -2737
rect 1008 -2771 1042 -2737
rect 938 -2839 972 -2805
rect 1008 -2839 1042 -2805
rect 938 -2907 972 -2873
rect 1008 -2907 1042 -2873
rect 938 -2975 972 -2941
rect 1008 -2975 1042 -2941
rect 938 -3043 972 -3009
rect 1008 -3043 1042 -3009
rect 938 -3111 972 -3077
rect 1008 -3111 1042 -3077
rect 938 -3179 972 -3145
rect 1008 -3179 1042 -3145
rect 938 -3247 972 -3213
rect 1008 -3247 1042 -3213
rect 938 -3315 972 -3281
rect 1008 -3315 1042 -3281
rect 938 -3383 972 -3349
rect 1008 -3383 1042 -3349
rect 938 -3451 972 -3417
rect 1008 -3451 1042 -3417
rect 938 -3519 972 -3485
rect 1008 -3519 1042 -3485
rect 938 -3587 972 -3553
rect 1008 -3587 1042 -3553
rect 938 -3655 972 -3621
rect 1008 -3655 1042 -3621
rect 938 -3723 972 -3689
rect 1008 -3723 1042 -3689
rect 938 -3791 972 -3757
rect 1008 -3791 1042 -3757
rect 938 -3859 972 -3825
rect 1008 -3859 1042 -3825
rect 938 -3927 972 -3893
rect 1008 -3927 1042 -3893
rect 938 -3995 972 -3961
rect 1008 -3995 1042 -3961
rect 938 -4063 972 -4029
rect 1008 -4063 1042 -4029
rect 938 -4131 972 -4097
rect 1008 -4131 1042 -4097
rect 938 -4199 972 -4165
rect 1008 -4199 1042 -4165
rect 938 -4267 972 -4233
rect 1008 -4267 1042 -4233
rect 938 -4335 972 -4301
rect 1008 -4335 1042 -4301
rect 938 -4403 972 -4369
rect 1008 -4403 1042 -4369
rect 938 -4471 972 -4437
rect 1008 -4471 1042 -4437
rect 938 -4539 972 -4505
rect 1008 -4539 1042 -4505
rect 938 -4607 972 -4573
rect 1008 -4607 1042 -4573
rect 938 -4675 972 -4641
rect 1008 -4675 1042 -4641
rect 938 -4743 972 -4709
rect 1008 -4743 1042 -4709
rect 938 -4811 972 -4777
rect 1008 -4811 1042 -4777
rect 938 -4879 972 -4845
rect 1008 -4879 1042 -4845
rect 938 -4947 972 -4913
rect 1008 -4947 1042 -4913
rect 938 -5015 972 -4981
rect 1008 -5015 1042 -4981
rect 1422 -5015 1524 5015
rect 1113 -5124 1147 -5090
rect 1181 -5124 1215 -5090
rect 1249 -5124 1283 -5090
rect 1317 -5124 1351 -5090
<< mvndiode >>
rect 1132 4981 1332 5000
rect 1132 -4981 1147 4981
rect 1317 -4981 1332 4981
rect 1132 -5000 1332 -4981
<< mvndiodec >>
rect 1147 -4981 1317 4981
<< locali >>
rect 922 5124 1540 5188
rect 922 5090 1107 5124
rect 1147 5090 1179 5124
rect 1215 5090 1249 5124
rect 1285 5090 1317 5124
rect 1357 5090 1540 5124
rect 922 5057 1042 5090
rect 922 5023 934 5057
rect 968 5023 1042 5057
rect 922 5021 1042 5023
rect 922 5015 1008 5021
rect 922 4985 938 5015
rect 922 4951 934 4985
rect 972 4981 1008 5015
rect 1422 5057 1540 5090
rect 1422 5023 1494 5057
rect 1528 5023 1540 5057
rect 1422 5021 1540 5023
rect 968 4951 1042 4981
rect 922 4949 1042 4951
rect 922 4947 1008 4949
rect 922 4913 938 4947
rect 972 4913 1008 4947
rect 922 4879 934 4913
rect 968 4879 1042 4913
rect 922 4845 938 4879
rect 972 4845 1008 4879
rect 922 4843 1008 4845
rect 922 4841 1042 4843
rect 922 4807 934 4841
rect 968 4811 1042 4841
rect 922 4777 938 4807
rect 972 4777 1008 4811
rect 922 4771 1008 4777
rect 922 4769 1042 4771
rect 922 4735 934 4769
rect 968 4743 1042 4769
rect 922 4709 938 4735
rect 972 4709 1008 4743
rect 922 4699 1008 4709
rect 922 4697 1042 4699
rect 922 4663 934 4697
rect 968 4675 1042 4697
rect 922 4641 938 4663
rect 972 4641 1008 4675
rect 922 4627 1008 4641
rect 922 4625 1042 4627
rect 922 4591 934 4625
rect 968 4607 1042 4625
rect 922 4573 938 4591
rect 972 4573 1008 4607
rect 922 4555 1008 4573
rect 922 4553 1042 4555
rect 922 4519 934 4553
rect 968 4539 1042 4553
rect 922 4505 938 4519
rect 972 4505 1008 4539
rect 922 4483 1008 4505
rect 922 4481 1042 4483
rect 922 4447 934 4481
rect 968 4471 1042 4481
rect 922 4437 938 4447
rect 972 4437 1008 4471
rect 922 4411 1008 4437
rect 922 4409 1042 4411
rect 922 4375 934 4409
rect 968 4403 1042 4409
rect 922 4369 938 4375
rect 972 4369 1008 4403
rect 922 4339 1008 4369
rect 922 4337 1042 4339
rect 922 4303 934 4337
rect 968 4335 1042 4337
rect 922 4301 938 4303
rect 972 4301 1008 4335
rect 922 4267 1008 4301
rect 922 4265 938 4267
rect 922 4231 934 4265
rect 972 4233 1008 4267
rect 968 4231 1042 4233
rect 922 4229 1042 4231
rect 922 4199 1008 4229
rect 922 4193 938 4199
rect 922 4159 934 4193
rect 972 4165 1008 4199
rect 968 4159 1042 4165
rect 922 4157 1042 4159
rect 922 4131 1008 4157
rect 922 4121 938 4131
rect 922 4087 934 4121
rect 972 4097 1008 4131
rect 968 4087 1042 4097
rect 922 4085 1042 4087
rect 922 4063 1008 4085
rect 922 4049 938 4063
rect 922 4015 934 4049
rect 972 4029 1008 4063
rect 968 4015 1042 4029
rect 922 4013 1042 4015
rect 922 3995 1008 4013
rect 922 3977 938 3995
rect 922 3943 934 3977
rect 972 3961 1008 3995
rect 968 3943 1042 3961
rect 922 3941 1042 3943
rect 922 3927 1008 3941
rect 922 3905 938 3927
rect 922 3871 934 3905
rect 972 3893 1008 3927
rect 968 3871 1042 3893
rect 922 3869 1042 3871
rect 922 3859 1008 3869
rect 922 3833 938 3859
rect 922 3799 934 3833
rect 972 3825 1008 3859
rect 968 3799 1042 3825
rect 922 3797 1042 3799
rect 922 3791 1008 3797
rect 922 3761 938 3791
rect 922 3727 934 3761
rect 972 3757 1008 3791
rect 968 3727 1042 3757
rect 922 3725 1042 3727
rect 922 3723 1008 3725
rect 922 3689 938 3723
rect 972 3689 1008 3723
rect 922 3655 934 3689
rect 968 3655 1042 3689
rect 922 3621 938 3655
rect 972 3621 1008 3655
rect 922 3619 1008 3621
rect 922 3617 1042 3619
rect 922 3583 934 3617
rect 968 3587 1042 3617
rect 922 3553 938 3583
rect 972 3553 1008 3587
rect 922 3547 1008 3553
rect 922 3545 1042 3547
rect 922 3511 934 3545
rect 968 3519 1042 3545
rect 922 3485 938 3511
rect 972 3485 1008 3519
rect 922 3475 1008 3485
rect 922 3473 1042 3475
rect 922 3439 934 3473
rect 968 3451 1042 3473
rect 922 3417 938 3439
rect 972 3417 1008 3451
rect 922 3403 1008 3417
rect 922 3401 1042 3403
rect 922 3367 934 3401
rect 968 3383 1042 3401
rect 922 3349 938 3367
rect 972 3349 1008 3383
rect 922 3331 1008 3349
rect 922 3329 1042 3331
rect 922 3295 934 3329
rect 968 3315 1042 3329
rect 922 3281 938 3295
rect 972 3281 1008 3315
rect 922 3259 1008 3281
rect 922 3257 1042 3259
rect 922 3223 934 3257
rect 968 3247 1042 3257
rect 922 3213 938 3223
rect 972 3213 1008 3247
rect 922 3187 1008 3213
rect 922 3185 1042 3187
rect 922 3151 934 3185
rect 968 3179 1042 3185
rect 922 3145 938 3151
rect 972 3145 1008 3179
rect 922 3115 1008 3145
rect 922 3113 1042 3115
rect 922 3079 934 3113
rect 968 3111 1042 3113
rect 922 3077 938 3079
rect 972 3077 1008 3111
rect 922 3043 1008 3077
rect 922 3041 938 3043
rect 922 3007 934 3041
rect 972 3009 1008 3043
rect 968 3007 1042 3009
rect 922 3005 1042 3007
rect 922 2975 1008 3005
rect 922 2969 938 2975
rect 922 2935 934 2969
rect 972 2941 1008 2975
rect 968 2935 1042 2941
rect 922 2933 1042 2935
rect 922 2907 1008 2933
rect 922 2897 938 2907
rect 922 2863 934 2897
rect 972 2873 1008 2907
rect 968 2863 1042 2873
rect 922 2861 1042 2863
rect 922 2839 1008 2861
rect 922 2825 938 2839
rect 922 2791 934 2825
rect 972 2805 1008 2839
rect 968 2791 1042 2805
rect 922 2789 1042 2791
rect 922 2771 1008 2789
rect 922 2753 938 2771
rect 922 2719 934 2753
rect 972 2737 1008 2771
rect 968 2719 1042 2737
rect 922 2717 1042 2719
rect 922 2703 1008 2717
rect 922 2681 938 2703
rect 922 2647 934 2681
rect 972 2669 1008 2703
rect 968 2647 1042 2669
rect 922 2645 1042 2647
rect 922 2635 1008 2645
rect 922 2609 938 2635
rect 922 2575 934 2609
rect 972 2601 1008 2635
rect 968 2575 1042 2601
rect 922 2573 1042 2575
rect 922 2567 1008 2573
rect 922 2537 938 2567
rect 922 2503 934 2537
rect 972 2533 1008 2567
rect 968 2503 1042 2533
rect 922 2501 1042 2503
rect 922 2499 1008 2501
rect 922 2465 938 2499
rect 972 2465 1008 2499
rect 922 2431 934 2465
rect 968 2431 1042 2465
rect 922 2397 938 2431
rect 972 2397 1008 2431
rect 922 2395 1008 2397
rect 922 2393 1042 2395
rect 922 2359 934 2393
rect 968 2363 1042 2393
rect 922 2329 938 2359
rect 972 2329 1008 2363
rect 922 2323 1008 2329
rect 922 2321 1042 2323
rect 922 2287 934 2321
rect 968 2295 1042 2321
rect 922 2261 938 2287
rect 972 2261 1008 2295
rect 922 2251 1008 2261
rect 922 2249 1042 2251
rect 922 2215 934 2249
rect 968 2227 1042 2249
rect 922 2193 938 2215
rect 972 2193 1008 2227
rect 922 2179 1008 2193
rect 922 2177 1042 2179
rect 922 2143 934 2177
rect 968 2159 1042 2177
rect 922 2125 938 2143
rect 972 2125 1008 2159
rect 922 2107 1008 2125
rect 922 2105 1042 2107
rect 922 2071 934 2105
rect 968 2091 1042 2105
rect 922 2057 938 2071
rect 972 2057 1008 2091
rect 922 2035 1008 2057
rect 922 2033 1042 2035
rect 922 1999 934 2033
rect 968 2023 1042 2033
rect 922 1989 938 1999
rect 972 1989 1008 2023
rect 922 1963 1008 1989
rect 922 1961 1042 1963
rect 922 1927 934 1961
rect 968 1955 1042 1961
rect 922 1921 938 1927
rect 972 1921 1008 1955
rect 922 1891 1008 1921
rect 922 1889 1042 1891
rect 922 1855 934 1889
rect 968 1887 1042 1889
rect 922 1853 938 1855
rect 972 1853 1008 1887
rect 922 1819 1008 1853
rect 922 1817 938 1819
rect 922 1783 934 1817
rect 972 1785 1008 1819
rect 968 1783 1042 1785
rect 922 1781 1042 1783
rect 922 1751 1008 1781
rect 922 1745 938 1751
rect 922 1711 934 1745
rect 972 1717 1008 1751
rect 968 1711 1042 1717
rect 922 1709 1042 1711
rect 922 1683 1008 1709
rect 922 1673 938 1683
rect 922 1639 934 1673
rect 972 1649 1008 1683
rect 968 1639 1042 1649
rect 922 1637 1042 1639
rect 922 1615 1008 1637
rect 922 1601 938 1615
rect 922 1567 934 1601
rect 972 1581 1008 1615
rect 968 1567 1042 1581
rect 922 1565 1042 1567
rect 922 1547 1008 1565
rect 922 1529 938 1547
rect 922 1495 934 1529
rect 972 1513 1008 1547
rect 968 1495 1042 1513
rect 922 1493 1042 1495
rect 922 1479 1008 1493
rect 922 1457 938 1479
rect 922 1423 934 1457
rect 972 1445 1008 1479
rect 968 1423 1042 1445
rect 922 1421 1042 1423
rect 922 1411 1008 1421
rect 922 1385 938 1411
rect 922 1351 934 1385
rect 972 1377 1008 1411
rect 968 1351 1042 1377
rect 922 1349 1042 1351
rect 922 1343 1008 1349
rect 922 1313 938 1343
rect 922 1279 934 1313
rect 972 1309 1008 1343
rect 968 1279 1042 1309
rect 922 1277 1042 1279
rect 922 1275 1008 1277
rect 922 1241 938 1275
rect 972 1241 1008 1275
rect 922 1207 934 1241
rect 968 1207 1042 1241
rect 922 1173 938 1207
rect 972 1173 1008 1207
rect 922 1171 1008 1173
rect 922 1169 1042 1171
rect 922 1135 934 1169
rect 968 1139 1042 1169
rect 922 1105 938 1135
rect 972 1105 1008 1139
rect 922 1099 1008 1105
rect 922 1097 1042 1099
rect 922 1063 934 1097
rect 968 1071 1042 1097
rect 922 1037 938 1063
rect 972 1037 1008 1071
rect 922 1027 1008 1037
rect 922 1025 1042 1027
rect 922 991 934 1025
rect 968 1003 1042 1025
rect 922 969 938 991
rect 972 969 1008 1003
rect 922 955 1008 969
rect 922 953 1042 955
rect 922 919 934 953
rect 968 935 1042 953
rect 922 901 938 919
rect 972 901 1008 935
rect 922 883 1008 901
rect 922 881 1042 883
rect 922 847 934 881
rect 968 867 1042 881
rect 922 833 938 847
rect 972 833 1008 867
rect 922 811 1008 833
rect 922 809 1042 811
rect 922 775 934 809
rect 968 799 1042 809
rect 922 765 938 775
rect 972 765 1008 799
rect 922 739 1008 765
rect 922 737 1042 739
rect 922 703 934 737
rect 968 731 1042 737
rect 922 697 938 703
rect 972 697 1008 731
rect 922 667 1008 697
rect 922 665 1042 667
rect 922 631 934 665
rect 968 663 1042 665
rect 922 629 938 631
rect 972 629 1008 663
rect 922 595 1008 629
rect 922 593 938 595
rect 922 559 934 593
rect 972 561 1008 595
rect 968 559 1042 561
rect 922 557 1042 559
rect 922 527 1008 557
rect 922 521 938 527
rect 922 487 934 521
rect 972 493 1008 527
rect 968 487 1042 493
rect 922 485 1042 487
rect 922 459 1008 485
rect 922 449 938 459
rect 922 415 934 449
rect 972 425 1008 459
rect 968 415 1042 425
rect 922 413 1042 415
rect 922 391 1008 413
rect 922 377 938 391
rect 922 343 934 377
rect 972 357 1008 391
rect 968 343 1042 357
rect 922 341 1042 343
rect 922 323 1008 341
rect 922 305 938 323
rect 922 271 934 305
rect 972 289 1008 323
rect 968 271 1042 289
rect 922 269 1042 271
rect 922 255 1008 269
rect 922 233 938 255
rect 922 199 934 233
rect 972 221 1008 255
rect 968 199 1042 221
rect 922 197 1042 199
rect 922 187 1008 197
rect 922 161 938 187
rect 922 127 934 161
rect 972 153 1008 187
rect 968 127 1042 153
rect 922 125 1042 127
rect 922 119 1008 125
rect 922 89 938 119
rect 922 55 934 89
rect 972 85 1008 119
rect 968 55 1042 85
rect 922 53 1042 55
rect 922 51 1008 53
rect 922 17 938 51
rect 972 17 1008 51
rect 922 -17 934 17
rect 968 -17 1042 17
rect 922 -51 938 -17
rect 972 -51 1008 -17
rect 922 -53 1008 -51
rect 922 -55 1042 -53
rect 922 -89 934 -55
rect 968 -85 1042 -55
rect 922 -119 938 -89
rect 972 -119 1008 -85
rect 922 -125 1008 -119
rect 922 -127 1042 -125
rect 922 -161 934 -127
rect 968 -153 1042 -127
rect 922 -187 938 -161
rect 972 -187 1008 -153
rect 922 -197 1008 -187
rect 922 -199 1042 -197
rect 922 -233 934 -199
rect 968 -221 1042 -199
rect 922 -255 938 -233
rect 972 -255 1008 -221
rect 922 -269 1008 -255
rect 922 -271 1042 -269
rect 922 -305 934 -271
rect 968 -289 1042 -271
rect 922 -323 938 -305
rect 972 -323 1008 -289
rect 922 -341 1008 -323
rect 922 -343 1042 -341
rect 922 -377 934 -343
rect 968 -357 1042 -343
rect 922 -391 938 -377
rect 972 -391 1008 -357
rect 922 -413 1008 -391
rect 922 -415 1042 -413
rect 922 -449 934 -415
rect 968 -425 1042 -415
rect 922 -459 938 -449
rect 972 -459 1008 -425
rect 922 -485 1008 -459
rect 922 -487 1042 -485
rect 922 -521 934 -487
rect 968 -493 1042 -487
rect 922 -527 938 -521
rect 972 -527 1008 -493
rect 922 -557 1008 -527
rect 922 -559 1042 -557
rect 922 -593 934 -559
rect 968 -561 1042 -559
rect 922 -595 938 -593
rect 972 -595 1008 -561
rect 922 -629 1008 -595
rect 922 -631 938 -629
rect 922 -665 934 -631
rect 972 -663 1008 -629
rect 968 -665 1042 -663
rect 922 -667 1042 -665
rect 922 -697 1008 -667
rect 922 -703 938 -697
rect 922 -737 934 -703
rect 972 -731 1008 -697
rect 968 -737 1042 -731
rect 922 -739 1042 -737
rect 922 -765 1008 -739
rect 922 -775 938 -765
rect 922 -809 934 -775
rect 972 -799 1008 -765
rect 968 -809 1042 -799
rect 922 -811 1042 -809
rect 922 -833 1008 -811
rect 922 -847 938 -833
rect 922 -881 934 -847
rect 972 -867 1008 -833
rect 968 -881 1042 -867
rect 922 -883 1042 -881
rect 922 -901 1008 -883
rect 922 -919 938 -901
rect 922 -953 934 -919
rect 972 -935 1008 -901
rect 968 -953 1042 -935
rect 922 -955 1042 -953
rect 922 -969 1008 -955
rect 922 -991 938 -969
rect 922 -1025 934 -991
rect 972 -1003 1008 -969
rect 968 -1025 1042 -1003
rect 922 -1027 1042 -1025
rect 922 -1037 1008 -1027
rect 922 -1063 938 -1037
rect 922 -1097 934 -1063
rect 972 -1071 1008 -1037
rect 968 -1097 1042 -1071
rect 922 -1099 1042 -1097
rect 922 -1105 1008 -1099
rect 922 -1135 938 -1105
rect 922 -1169 934 -1135
rect 972 -1139 1008 -1105
rect 968 -1169 1042 -1139
rect 922 -1171 1042 -1169
rect 922 -1173 1008 -1171
rect 922 -1207 938 -1173
rect 972 -1207 1008 -1173
rect 922 -1241 934 -1207
rect 968 -1241 1042 -1207
rect 922 -1275 938 -1241
rect 972 -1275 1008 -1241
rect 922 -1277 1008 -1275
rect 922 -1279 1042 -1277
rect 922 -1313 934 -1279
rect 968 -1309 1042 -1279
rect 922 -1343 938 -1313
rect 972 -1343 1008 -1309
rect 922 -1349 1008 -1343
rect 922 -1351 1042 -1349
rect 922 -1385 934 -1351
rect 968 -1377 1042 -1351
rect 922 -1411 938 -1385
rect 972 -1411 1008 -1377
rect 922 -1421 1008 -1411
rect 922 -1423 1042 -1421
rect 922 -1457 934 -1423
rect 968 -1445 1042 -1423
rect 922 -1479 938 -1457
rect 972 -1479 1008 -1445
rect 922 -1493 1008 -1479
rect 922 -1495 1042 -1493
rect 922 -1529 934 -1495
rect 968 -1513 1042 -1495
rect 922 -1547 938 -1529
rect 972 -1547 1008 -1513
rect 922 -1565 1008 -1547
rect 922 -1567 1042 -1565
rect 922 -1601 934 -1567
rect 968 -1581 1042 -1567
rect 922 -1615 938 -1601
rect 972 -1615 1008 -1581
rect 922 -1637 1008 -1615
rect 922 -1639 1042 -1637
rect 922 -1673 934 -1639
rect 968 -1649 1042 -1639
rect 922 -1683 938 -1673
rect 972 -1683 1008 -1649
rect 922 -1709 1008 -1683
rect 922 -1711 1042 -1709
rect 922 -1745 934 -1711
rect 968 -1717 1042 -1711
rect 922 -1751 938 -1745
rect 972 -1751 1008 -1717
rect 922 -1781 1008 -1751
rect 922 -1783 1042 -1781
rect 922 -1817 934 -1783
rect 968 -1785 1042 -1783
rect 922 -1819 938 -1817
rect 972 -1819 1008 -1785
rect 922 -1853 1008 -1819
rect 922 -1855 938 -1853
rect 922 -1889 934 -1855
rect 972 -1887 1008 -1853
rect 968 -1889 1042 -1887
rect 922 -1891 1042 -1889
rect 922 -1921 1008 -1891
rect 922 -1927 938 -1921
rect 922 -1961 934 -1927
rect 972 -1955 1008 -1921
rect 968 -1961 1042 -1955
rect 922 -1963 1042 -1961
rect 922 -1989 1008 -1963
rect 922 -1999 938 -1989
rect 922 -2033 934 -1999
rect 972 -2023 1008 -1989
rect 968 -2033 1042 -2023
rect 922 -2035 1042 -2033
rect 922 -2057 1008 -2035
rect 922 -2071 938 -2057
rect 922 -2105 934 -2071
rect 972 -2091 1008 -2057
rect 968 -2105 1042 -2091
rect 922 -2107 1042 -2105
rect 922 -2125 1008 -2107
rect 922 -2143 938 -2125
rect 922 -2177 934 -2143
rect 972 -2159 1008 -2125
rect 968 -2177 1042 -2159
rect 922 -2179 1042 -2177
rect 922 -2193 1008 -2179
rect 922 -2215 938 -2193
rect 922 -2249 934 -2215
rect 972 -2227 1008 -2193
rect 968 -2249 1042 -2227
rect 922 -2251 1042 -2249
rect 922 -2261 1008 -2251
rect 922 -2287 938 -2261
rect 922 -2321 934 -2287
rect 972 -2295 1008 -2261
rect 968 -2321 1042 -2295
rect 922 -2323 1042 -2321
rect 922 -2329 1008 -2323
rect 922 -2359 938 -2329
rect 922 -2393 934 -2359
rect 972 -2363 1008 -2329
rect 968 -2393 1042 -2363
rect 922 -2395 1042 -2393
rect 922 -2397 1008 -2395
rect 922 -2431 938 -2397
rect 972 -2431 1008 -2397
rect 922 -2465 934 -2431
rect 968 -2465 1042 -2431
rect 922 -2499 938 -2465
rect 972 -2499 1008 -2465
rect 922 -2501 1008 -2499
rect 922 -2503 1042 -2501
rect 922 -2537 934 -2503
rect 968 -2533 1042 -2503
rect 922 -2567 938 -2537
rect 972 -2567 1008 -2533
rect 922 -2573 1008 -2567
rect 922 -2575 1042 -2573
rect 922 -2609 934 -2575
rect 968 -2601 1042 -2575
rect 922 -2635 938 -2609
rect 972 -2635 1008 -2601
rect 922 -2645 1008 -2635
rect 922 -2647 1042 -2645
rect 922 -2681 934 -2647
rect 968 -2669 1042 -2647
rect 922 -2703 938 -2681
rect 972 -2703 1008 -2669
rect 922 -2717 1008 -2703
rect 922 -2719 1042 -2717
rect 922 -2753 934 -2719
rect 968 -2737 1042 -2719
rect 922 -2771 938 -2753
rect 972 -2771 1008 -2737
rect 922 -2789 1008 -2771
rect 922 -2791 1042 -2789
rect 922 -2825 934 -2791
rect 968 -2805 1042 -2791
rect 922 -2839 938 -2825
rect 972 -2839 1008 -2805
rect 922 -2861 1008 -2839
rect 922 -2863 1042 -2861
rect 922 -2897 934 -2863
rect 968 -2873 1042 -2863
rect 922 -2907 938 -2897
rect 972 -2907 1008 -2873
rect 922 -2933 1008 -2907
rect 922 -2935 1042 -2933
rect 922 -2969 934 -2935
rect 968 -2941 1042 -2935
rect 922 -2975 938 -2969
rect 972 -2975 1008 -2941
rect 922 -3005 1008 -2975
rect 922 -3007 1042 -3005
rect 922 -3041 934 -3007
rect 968 -3009 1042 -3007
rect 922 -3043 938 -3041
rect 972 -3043 1008 -3009
rect 922 -3077 1008 -3043
rect 922 -3079 938 -3077
rect 922 -3113 934 -3079
rect 972 -3111 1008 -3077
rect 968 -3113 1042 -3111
rect 922 -3115 1042 -3113
rect 922 -3145 1008 -3115
rect 922 -3151 938 -3145
rect 922 -3185 934 -3151
rect 972 -3179 1008 -3145
rect 968 -3185 1042 -3179
rect 922 -3187 1042 -3185
rect 922 -3213 1008 -3187
rect 922 -3223 938 -3213
rect 922 -3257 934 -3223
rect 972 -3247 1008 -3213
rect 968 -3257 1042 -3247
rect 922 -3259 1042 -3257
rect 922 -3281 1008 -3259
rect 922 -3295 938 -3281
rect 922 -3329 934 -3295
rect 972 -3315 1008 -3281
rect 968 -3329 1042 -3315
rect 922 -3331 1042 -3329
rect 922 -3349 1008 -3331
rect 922 -3367 938 -3349
rect 922 -3401 934 -3367
rect 972 -3383 1008 -3349
rect 968 -3401 1042 -3383
rect 922 -3403 1042 -3401
rect 922 -3417 1008 -3403
rect 922 -3439 938 -3417
rect 922 -3473 934 -3439
rect 972 -3451 1008 -3417
rect 968 -3473 1042 -3451
rect 922 -3475 1042 -3473
rect 922 -3485 1008 -3475
rect 922 -3511 938 -3485
rect 922 -3545 934 -3511
rect 972 -3519 1008 -3485
rect 968 -3545 1042 -3519
rect 922 -3547 1042 -3545
rect 922 -3553 1008 -3547
rect 922 -3583 938 -3553
rect 922 -3617 934 -3583
rect 972 -3587 1008 -3553
rect 968 -3617 1042 -3587
rect 922 -3619 1042 -3617
rect 922 -3621 1008 -3619
rect 922 -3655 938 -3621
rect 972 -3655 1008 -3621
rect 922 -3689 934 -3655
rect 968 -3689 1042 -3655
rect 922 -3723 938 -3689
rect 972 -3723 1008 -3689
rect 922 -3725 1008 -3723
rect 922 -3727 1042 -3725
rect 922 -3761 934 -3727
rect 968 -3757 1042 -3727
rect 922 -3791 938 -3761
rect 972 -3791 1008 -3757
rect 922 -3797 1008 -3791
rect 922 -3799 1042 -3797
rect 922 -3833 934 -3799
rect 968 -3825 1042 -3799
rect 922 -3859 938 -3833
rect 972 -3859 1008 -3825
rect 922 -3869 1008 -3859
rect 922 -3871 1042 -3869
rect 922 -3905 934 -3871
rect 968 -3893 1042 -3871
rect 922 -3927 938 -3905
rect 972 -3927 1008 -3893
rect 922 -3941 1008 -3927
rect 922 -3943 1042 -3941
rect 922 -3977 934 -3943
rect 968 -3961 1042 -3943
rect 922 -3995 938 -3977
rect 972 -3995 1008 -3961
rect 922 -4013 1008 -3995
rect 922 -4015 1042 -4013
rect 922 -4049 934 -4015
rect 968 -4029 1042 -4015
rect 922 -4063 938 -4049
rect 972 -4063 1008 -4029
rect 922 -4085 1008 -4063
rect 922 -4087 1042 -4085
rect 922 -4121 934 -4087
rect 968 -4097 1042 -4087
rect 922 -4131 938 -4121
rect 972 -4131 1008 -4097
rect 922 -4157 1008 -4131
rect 922 -4159 1042 -4157
rect 922 -4193 934 -4159
rect 968 -4165 1042 -4159
rect 922 -4199 938 -4193
rect 972 -4199 1008 -4165
rect 922 -4229 1008 -4199
rect 922 -4231 1042 -4229
rect 922 -4265 934 -4231
rect 968 -4233 1042 -4231
rect 922 -4267 938 -4265
rect 972 -4267 1008 -4233
rect 922 -4301 1008 -4267
rect 922 -4303 938 -4301
rect 922 -4337 934 -4303
rect 972 -4335 1008 -4301
rect 968 -4337 1042 -4335
rect 922 -4339 1042 -4337
rect 922 -4369 1008 -4339
rect 922 -4375 938 -4369
rect 922 -4409 934 -4375
rect 972 -4403 1008 -4369
rect 968 -4409 1042 -4403
rect 922 -4411 1042 -4409
rect 922 -4437 1008 -4411
rect 922 -4447 938 -4437
rect 922 -4481 934 -4447
rect 972 -4471 1008 -4437
rect 968 -4481 1042 -4471
rect 922 -4483 1042 -4481
rect 922 -4505 1008 -4483
rect 922 -4519 938 -4505
rect 922 -4553 934 -4519
rect 972 -4539 1008 -4505
rect 968 -4553 1042 -4539
rect 922 -4555 1042 -4553
rect 922 -4573 1008 -4555
rect 922 -4591 938 -4573
rect 922 -4625 934 -4591
rect 972 -4607 1008 -4573
rect 968 -4625 1042 -4607
rect 922 -4627 1042 -4625
rect 922 -4641 1008 -4627
rect 922 -4663 938 -4641
rect 922 -4697 934 -4663
rect 972 -4675 1008 -4641
rect 968 -4697 1042 -4675
rect 922 -4699 1042 -4697
rect 922 -4709 1008 -4699
rect 922 -4735 938 -4709
rect 922 -4769 934 -4735
rect 972 -4743 1008 -4709
rect 968 -4769 1042 -4743
rect 922 -4771 1042 -4769
rect 922 -4777 1008 -4771
rect 922 -4807 938 -4777
rect 922 -4841 934 -4807
rect 972 -4811 1008 -4777
rect 968 -4841 1042 -4811
rect 922 -4843 1042 -4841
rect 922 -4845 1008 -4843
rect 922 -4879 938 -4845
rect 972 -4879 1008 -4845
rect 922 -4913 934 -4879
rect 968 -4913 1042 -4879
rect 922 -4947 938 -4913
rect 972 -4947 1008 -4913
rect 922 -4949 1008 -4947
rect 922 -4951 1042 -4949
rect 922 -4985 934 -4951
rect 968 -4981 1042 -4951
rect 922 -5015 938 -4985
rect 972 -5015 1008 -4981
rect 1144 4985 1320 5004
rect 1144 4981 1179 4985
rect 1285 4981 1320 4985
rect 1144 -4981 1147 4981
rect 1317 -4981 1320 4981
rect 1144 -4985 1179 -4981
rect 1285 -4985 1320 -4981
rect 1144 -5004 1320 -4985
rect 922 -5021 1008 -5015
rect 922 -5023 1042 -5021
rect 922 -5057 934 -5023
rect 968 -5057 1042 -5023
rect 922 -5090 1042 -5057
rect 1528 -5021 1540 5021
rect 1422 -5023 1540 -5021
rect 1422 -5057 1494 -5023
rect 1528 -5057 1540 -5023
rect 1422 -5090 1540 -5057
rect 922 -5124 1107 -5090
rect 1147 -5124 1179 -5090
rect 1215 -5124 1249 -5090
rect 1285 -5124 1317 -5090
rect 1357 -5124 1540 -5090
rect 922 -5188 1540 -5124
<< viali >>
rect 1107 5090 1113 5124
rect 1113 5090 1141 5124
rect 1179 5090 1181 5124
rect 1181 5090 1213 5124
rect 1251 5090 1283 5124
rect 1283 5090 1285 5124
rect 1323 5090 1351 5124
rect 1351 5090 1357 5124
rect 934 5023 968 5057
rect 1008 5015 1042 5021
rect 934 4981 938 4985
rect 938 4981 968 4985
rect 1008 4987 1042 5015
rect 1494 5023 1528 5057
rect 1422 5015 1528 5021
rect 934 4951 968 4981
rect 1008 4947 1042 4949
rect 1008 4915 1042 4947
rect 934 4879 968 4913
rect 1008 4845 1042 4877
rect 1008 4843 1042 4845
rect 934 4811 968 4841
rect 934 4807 938 4811
rect 938 4807 968 4811
rect 1008 4777 1042 4805
rect 1008 4771 1042 4777
rect 934 4743 968 4769
rect 934 4735 938 4743
rect 938 4735 968 4743
rect 1008 4709 1042 4733
rect 1008 4699 1042 4709
rect 934 4675 968 4697
rect 934 4663 938 4675
rect 938 4663 968 4675
rect 1008 4641 1042 4661
rect 1008 4627 1042 4641
rect 934 4607 968 4625
rect 934 4591 938 4607
rect 938 4591 968 4607
rect 1008 4573 1042 4589
rect 1008 4555 1042 4573
rect 934 4539 968 4553
rect 934 4519 938 4539
rect 938 4519 968 4539
rect 1008 4505 1042 4517
rect 1008 4483 1042 4505
rect 934 4471 968 4481
rect 934 4447 938 4471
rect 938 4447 968 4471
rect 1008 4437 1042 4445
rect 1008 4411 1042 4437
rect 934 4403 968 4409
rect 934 4375 938 4403
rect 938 4375 968 4403
rect 1008 4369 1042 4373
rect 1008 4339 1042 4369
rect 934 4335 968 4337
rect 934 4303 938 4335
rect 938 4303 968 4335
rect 1008 4267 1042 4301
rect 934 4233 938 4265
rect 938 4233 968 4265
rect 934 4231 968 4233
rect 1008 4199 1042 4229
rect 934 4165 938 4193
rect 938 4165 968 4193
rect 1008 4195 1042 4199
rect 934 4159 968 4165
rect 1008 4131 1042 4157
rect 934 4097 938 4121
rect 938 4097 968 4121
rect 1008 4123 1042 4131
rect 934 4087 968 4097
rect 1008 4063 1042 4085
rect 934 4029 938 4049
rect 938 4029 968 4049
rect 1008 4051 1042 4063
rect 934 4015 968 4029
rect 1008 3995 1042 4013
rect 934 3961 938 3977
rect 938 3961 968 3977
rect 1008 3979 1042 3995
rect 934 3943 968 3961
rect 1008 3927 1042 3941
rect 934 3893 938 3905
rect 938 3893 968 3905
rect 1008 3907 1042 3927
rect 934 3871 968 3893
rect 1008 3859 1042 3869
rect 934 3825 938 3833
rect 938 3825 968 3833
rect 1008 3835 1042 3859
rect 934 3799 968 3825
rect 1008 3791 1042 3797
rect 934 3757 938 3761
rect 938 3757 968 3761
rect 1008 3763 1042 3791
rect 934 3727 968 3757
rect 1008 3723 1042 3725
rect 1008 3691 1042 3723
rect 934 3655 968 3689
rect 1008 3621 1042 3653
rect 1008 3619 1042 3621
rect 934 3587 968 3617
rect 934 3583 938 3587
rect 938 3583 968 3587
rect 1008 3553 1042 3581
rect 1008 3547 1042 3553
rect 934 3519 968 3545
rect 934 3511 938 3519
rect 938 3511 968 3519
rect 1008 3485 1042 3509
rect 1008 3475 1042 3485
rect 934 3451 968 3473
rect 934 3439 938 3451
rect 938 3439 968 3451
rect 1008 3417 1042 3437
rect 1008 3403 1042 3417
rect 934 3383 968 3401
rect 934 3367 938 3383
rect 938 3367 968 3383
rect 1008 3349 1042 3365
rect 1008 3331 1042 3349
rect 934 3315 968 3329
rect 934 3295 938 3315
rect 938 3295 968 3315
rect 1008 3281 1042 3293
rect 1008 3259 1042 3281
rect 934 3247 968 3257
rect 934 3223 938 3247
rect 938 3223 968 3247
rect 1008 3213 1042 3221
rect 1008 3187 1042 3213
rect 934 3179 968 3185
rect 934 3151 938 3179
rect 938 3151 968 3179
rect 1008 3145 1042 3149
rect 1008 3115 1042 3145
rect 934 3111 968 3113
rect 934 3079 938 3111
rect 938 3079 968 3111
rect 1008 3043 1042 3077
rect 934 3009 938 3041
rect 938 3009 968 3041
rect 934 3007 968 3009
rect 1008 2975 1042 3005
rect 934 2941 938 2969
rect 938 2941 968 2969
rect 1008 2971 1042 2975
rect 934 2935 968 2941
rect 1008 2907 1042 2933
rect 934 2873 938 2897
rect 938 2873 968 2897
rect 1008 2899 1042 2907
rect 934 2863 968 2873
rect 1008 2839 1042 2861
rect 934 2805 938 2825
rect 938 2805 968 2825
rect 1008 2827 1042 2839
rect 934 2791 968 2805
rect 1008 2771 1042 2789
rect 934 2737 938 2753
rect 938 2737 968 2753
rect 1008 2755 1042 2771
rect 934 2719 968 2737
rect 1008 2703 1042 2717
rect 934 2669 938 2681
rect 938 2669 968 2681
rect 1008 2683 1042 2703
rect 934 2647 968 2669
rect 1008 2635 1042 2645
rect 934 2601 938 2609
rect 938 2601 968 2609
rect 1008 2611 1042 2635
rect 934 2575 968 2601
rect 1008 2567 1042 2573
rect 934 2533 938 2537
rect 938 2533 968 2537
rect 1008 2539 1042 2567
rect 934 2503 968 2533
rect 1008 2499 1042 2501
rect 1008 2467 1042 2499
rect 934 2431 968 2465
rect 1008 2397 1042 2429
rect 1008 2395 1042 2397
rect 934 2363 968 2393
rect 934 2359 938 2363
rect 938 2359 968 2363
rect 1008 2329 1042 2357
rect 1008 2323 1042 2329
rect 934 2295 968 2321
rect 934 2287 938 2295
rect 938 2287 968 2295
rect 1008 2261 1042 2285
rect 1008 2251 1042 2261
rect 934 2227 968 2249
rect 934 2215 938 2227
rect 938 2215 968 2227
rect 1008 2193 1042 2213
rect 1008 2179 1042 2193
rect 934 2159 968 2177
rect 934 2143 938 2159
rect 938 2143 968 2159
rect 1008 2125 1042 2141
rect 1008 2107 1042 2125
rect 934 2091 968 2105
rect 934 2071 938 2091
rect 938 2071 968 2091
rect 1008 2057 1042 2069
rect 1008 2035 1042 2057
rect 934 2023 968 2033
rect 934 1999 938 2023
rect 938 1999 968 2023
rect 1008 1989 1042 1997
rect 1008 1963 1042 1989
rect 934 1955 968 1961
rect 934 1927 938 1955
rect 938 1927 968 1955
rect 1008 1921 1042 1925
rect 1008 1891 1042 1921
rect 934 1887 968 1889
rect 934 1855 938 1887
rect 938 1855 968 1887
rect 1008 1819 1042 1853
rect 934 1785 938 1817
rect 938 1785 968 1817
rect 934 1783 968 1785
rect 1008 1751 1042 1781
rect 934 1717 938 1745
rect 938 1717 968 1745
rect 1008 1747 1042 1751
rect 934 1711 968 1717
rect 1008 1683 1042 1709
rect 934 1649 938 1673
rect 938 1649 968 1673
rect 1008 1675 1042 1683
rect 934 1639 968 1649
rect 1008 1615 1042 1637
rect 934 1581 938 1601
rect 938 1581 968 1601
rect 1008 1603 1042 1615
rect 934 1567 968 1581
rect 1008 1547 1042 1565
rect 934 1513 938 1529
rect 938 1513 968 1529
rect 1008 1531 1042 1547
rect 934 1495 968 1513
rect 1008 1479 1042 1493
rect 934 1445 938 1457
rect 938 1445 968 1457
rect 1008 1459 1042 1479
rect 934 1423 968 1445
rect 1008 1411 1042 1421
rect 934 1377 938 1385
rect 938 1377 968 1385
rect 1008 1387 1042 1411
rect 934 1351 968 1377
rect 1008 1343 1042 1349
rect 934 1309 938 1313
rect 938 1309 968 1313
rect 1008 1315 1042 1343
rect 934 1279 968 1309
rect 1008 1275 1042 1277
rect 1008 1243 1042 1275
rect 934 1207 968 1241
rect 1008 1173 1042 1205
rect 1008 1171 1042 1173
rect 934 1139 968 1169
rect 934 1135 938 1139
rect 938 1135 968 1139
rect 1008 1105 1042 1133
rect 1008 1099 1042 1105
rect 934 1071 968 1097
rect 934 1063 938 1071
rect 938 1063 968 1071
rect 1008 1037 1042 1061
rect 1008 1027 1042 1037
rect 934 1003 968 1025
rect 934 991 938 1003
rect 938 991 968 1003
rect 1008 969 1042 989
rect 1008 955 1042 969
rect 934 935 968 953
rect 934 919 938 935
rect 938 919 968 935
rect 1008 901 1042 917
rect 1008 883 1042 901
rect 934 867 968 881
rect 934 847 938 867
rect 938 847 968 867
rect 1008 833 1042 845
rect 1008 811 1042 833
rect 934 799 968 809
rect 934 775 938 799
rect 938 775 968 799
rect 1008 765 1042 773
rect 1008 739 1042 765
rect 934 731 968 737
rect 934 703 938 731
rect 938 703 968 731
rect 1008 697 1042 701
rect 1008 667 1042 697
rect 934 663 968 665
rect 934 631 938 663
rect 938 631 968 663
rect 1008 595 1042 629
rect 934 561 938 593
rect 938 561 968 593
rect 934 559 968 561
rect 1008 527 1042 557
rect 934 493 938 521
rect 938 493 968 521
rect 1008 523 1042 527
rect 934 487 968 493
rect 1008 459 1042 485
rect 934 425 938 449
rect 938 425 968 449
rect 1008 451 1042 459
rect 934 415 968 425
rect 1008 391 1042 413
rect 934 357 938 377
rect 938 357 968 377
rect 1008 379 1042 391
rect 934 343 968 357
rect 1008 323 1042 341
rect 934 289 938 305
rect 938 289 968 305
rect 1008 307 1042 323
rect 934 271 968 289
rect 1008 255 1042 269
rect 934 221 938 233
rect 938 221 968 233
rect 1008 235 1042 255
rect 934 199 968 221
rect 1008 187 1042 197
rect 934 153 938 161
rect 938 153 968 161
rect 1008 163 1042 187
rect 934 127 968 153
rect 1008 119 1042 125
rect 934 85 938 89
rect 938 85 968 89
rect 1008 91 1042 119
rect 934 55 968 85
rect 1008 51 1042 53
rect 1008 19 1042 51
rect 934 -17 968 17
rect 1008 -51 1042 -19
rect 1008 -53 1042 -51
rect 934 -85 968 -55
rect 934 -89 938 -85
rect 938 -89 968 -85
rect 1008 -119 1042 -91
rect 1008 -125 1042 -119
rect 934 -153 968 -127
rect 934 -161 938 -153
rect 938 -161 968 -153
rect 1008 -187 1042 -163
rect 1008 -197 1042 -187
rect 934 -221 968 -199
rect 934 -233 938 -221
rect 938 -233 968 -221
rect 1008 -255 1042 -235
rect 1008 -269 1042 -255
rect 934 -289 968 -271
rect 934 -305 938 -289
rect 938 -305 968 -289
rect 1008 -323 1042 -307
rect 1008 -341 1042 -323
rect 934 -357 968 -343
rect 934 -377 938 -357
rect 938 -377 968 -357
rect 1008 -391 1042 -379
rect 1008 -413 1042 -391
rect 934 -425 968 -415
rect 934 -449 938 -425
rect 938 -449 968 -425
rect 1008 -459 1042 -451
rect 1008 -485 1042 -459
rect 934 -493 968 -487
rect 934 -521 938 -493
rect 938 -521 968 -493
rect 1008 -527 1042 -523
rect 1008 -557 1042 -527
rect 934 -561 968 -559
rect 934 -593 938 -561
rect 938 -593 968 -561
rect 1008 -629 1042 -595
rect 934 -663 938 -631
rect 938 -663 968 -631
rect 934 -665 968 -663
rect 1008 -697 1042 -667
rect 934 -731 938 -703
rect 938 -731 968 -703
rect 1008 -701 1042 -697
rect 934 -737 968 -731
rect 1008 -765 1042 -739
rect 934 -799 938 -775
rect 938 -799 968 -775
rect 1008 -773 1042 -765
rect 934 -809 968 -799
rect 1008 -833 1042 -811
rect 934 -867 938 -847
rect 938 -867 968 -847
rect 1008 -845 1042 -833
rect 934 -881 968 -867
rect 1008 -901 1042 -883
rect 934 -935 938 -919
rect 938 -935 968 -919
rect 1008 -917 1042 -901
rect 934 -953 968 -935
rect 1008 -969 1042 -955
rect 934 -1003 938 -991
rect 938 -1003 968 -991
rect 1008 -989 1042 -969
rect 934 -1025 968 -1003
rect 1008 -1037 1042 -1027
rect 934 -1071 938 -1063
rect 938 -1071 968 -1063
rect 1008 -1061 1042 -1037
rect 934 -1097 968 -1071
rect 1008 -1105 1042 -1099
rect 934 -1139 938 -1135
rect 938 -1139 968 -1135
rect 1008 -1133 1042 -1105
rect 934 -1169 968 -1139
rect 1008 -1173 1042 -1171
rect 1008 -1205 1042 -1173
rect 934 -1241 968 -1207
rect 1008 -1275 1042 -1243
rect 1008 -1277 1042 -1275
rect 934 -1309 968 -1279
rect 934 -1313 938 -1309
rect 938 -1313 968 -1309
rect 1008 -1343 1042 -1315
rect 1008 -1349 1042 -1343
rect 934 -1377 968 -1351
rect 934 -1385 938 -1377
rect 938 -1385 968 -1377
rect 1008 -1411 1042 -1387
rect 1008 -1421 1042 -1411
rect 934 -1445 968 -1423
rect 934 -1457 938 -1445
rect 938 -1457 968 -1445
rect 1008 -1479 1042 -1459
rect 1008 -1493 1042 -1479
rect 934 -1513 968 -1495
rect 934 -1529 938 -1513
rect 938 -1529 968 -1513
rect 1008 -1547 1042 -1531
rect 1008 -1565 1042 -1547
rect 934 -1581 968 -1567
rect 934 -1601 938 -1581
rect 938 -1601 968 -1581
rect 1008 -1615 1042 -1603
rect 1008 -1637 1042 -1615
rect 934 -1649 968 -1639
rect 934 -1673 938 -1649
rect 938 -1673 968 -1649
rect 1008 -1683 1042 -1675
rect 1008 -1709 1042 -1683
rect 934 -1717 968 -1711
rect 934 -1745 938 -1717
rect 938 -1745 968 -1717
rect 1008 -1751 1042 -1747
rect 1008 -1781 1042 -1751
rect 934 -1785 968 -1783
rect 934 -1817 938 -1785
rect 938 -1817 968 -1785
rect 1008 -1853 1042 -1819
rect 934 -1887 938 -1855
rect 938 -1887 968 -1855
rect 934 -1889 968 -1887
rect 1008 -1921 1042 -1891
rect 934 -1955 938 -1927
rect 938 -1955 968 -1927
rect 1008 -1925 1042 -1921
rect 934 -1961 968 -1955
rect 1008 -1989 1042 -1963
rect 934 -2023 938 -1999
rect 938 -2023 968 -1999
rect 1008 -1997 1042 -1989
rect 934 -2033 968 -2023
rect 1008 -2057 1042 -2035
rect 934 -2091 938 -2071
rect 938 -2091 968 -2071
rect 1008 -2069 1042 -2057
rect 934 -2105 968 -2091
rect 1008 -2125 1042 -2107
rect 934 -2159 938 -2143
rect 938 -2159 968 -2143
rect 1008 -2141 1042 -2125
rect 934 -2177 968 -2159
rect 1008 -2193 1042 -2179
rect 934 -2227 938 -2215
rect 938 -2227 968 -2215
rect 1008 -2213 1042 -2193
rect 934 -2249 968 -2227
rect 1008 -2261 1042 -2251
rect 934 -2295 938 -2287
rect 938 -2295 968 -2287
rect 1008 -2285 1042 -2261
rect 934 -2321 968 -2295
rect 1008 -2329 1042 -2323
rect 934 -2363 938 -2359
rect 938 -2363 968 -2359
rect 1008 -2357 1042 -2329
rect 934 -2393 968 -2363
rect 1008 -2397 1042 -2395
rect 1008 -2429 1042 -2397
rect 934 -2465 968 -2431
rect 1008 -2499 1042 -2467
rect 1008 -2501 1042 -2499
rect 934 -2533 968 -2503
rect 934 -2537 938 -2533
rect 938 -2537 968 -2533
rect 1008 -2567 1042 -2539
rect 1008 -2573 1042 -2567
rect 934 -2601 968 -2575
rect 934 -2609 938 -2601
rect 938 -2609 968 -2601
rect 1008 -2635 1042 -2611
rect 1008 -2645 1042 -2635
rect 934 -2669 968 -2647
rect 934 -2681 938 -2669
rect 938 -2681 968 -2669
rect 1008 -2703 1042 -2683
rect 1008 -2717 1042 -2703
rect 934 -2737 968 -2719
rect 934 -2753 938 -2737
rect 938 -2753 968 -2737
rect 1008 -2771 1042 -2755
rect 1008 -2789 1042 -2771
rect 934 -2805 968 -2791
rect 934 -2825 938 -2805
rect 938 -2825 968 -2805
rect 1008 -2839 1042 -2827
rect 1008 -2861 1042 -2839
rect 934 -2873 968 -2863
rect 934 -2897 938 -2873
rect 938 -2897 968 -2873
rect 1008 -2907 1042 -2899
rect 1008 -2933 1042 -2907
rect 934 -2941 968 -2935
rect 934 -2969 938 -2941
rect 938 -2969 968 -2941
rect 1008 -2975 1042 -2971
rect 1008 -3005 1042 -2975
rect 934 -3009 968 -3007
rect 934 -3041 938 -3009
rect 938 -3041 968 -3009
rect 1008 -3077 1042 -3043
rect 934 -3111 938 -3079
rect 938 -3111 968 -3079
rect 934 -3113 968 -3111
rect 1008 -3145 1042 -3115
rect 934 -3179 938 -3151
rect 938 -3179 968 -3151
rect 1008 -3149 1042 -3145
rect 934 -3185 968 -3179
rect 1008 -3213 1042 -3187
rect 934 -3247 938 -3223
rect 938 -3247 968 -3223
rect 1008 -3221 1042 -3213
rect 934 -3257 968 -3247
rect 1008 -3281 1042 -3259
rect 934 -3315 938 -3295
rect 938 -3315 968 -3295
rect 1008 -3293 1042 -3281
rect 934 -3329 968 -3315
rect 1008 -3349 1042 -3331
rect 934 -3383 938 -3367
rect 938 -3383 968 -3367
rect 1008 -3365 1042 -3349
rect 934 -3401 968 -3383
rect 1008 -3417 1042 -3403
rect 934 -3451 938 -3439
rect 938 -3451 968 -3439
rect 1008 -3437 1042 -3417
rect 934 -3473 968 -3451
rect 1008 -3485 1042 -3475
rect 934 -3519 938 -3511
rect 938 -3519 968 -3511
rect 1008 -3509 1042 -3485
rect 934 -3545 968 -3519
rect 1008 -3553 1042 -3547
rect 934 -3587 938 -3583
rect 938 -3587 968 -3583
rect 1008 -3581 1042 -3553
rect 934 -3617 968 -3587
rect 1008 -3621 1042 -3619
rect 1008 -3653 1042 -3621
rect 934 -3689 968 -3655
rect 1008 -3723 1042 -3691
rect 1008 -3725 1042 -3723
rect 934 -3757 968 -3727
rect 934 -3761 938 -3757
rect 938 -3761 968 -3757
rect 1008 -3791 1042 -3763
rect 1008 -3797 1042 -3791
rect 934 -3825 968 -3799
rect 934 -3833 938 -3825
rect 938 -3833 968 -3825
rect 1008 -3859 1042 -3835
rect 1008 -3869 1042 -3859
rect 934 -3893 968 -3871
rect 934 -3905 938 -3893
rect 938 -3905 968 -3893
rect 1008 -3927 1042 -3907
rect 1008 -3941 1042 -3927
rect 934 -3961 968 -3943
rect 934 -3977 938 -3961
rect 938 -3977 968 -3961
rect 1008 -3995 1042 -3979
rect 1008 -4013 1042 -3995
rect 934 -4029 968 -4015
rect 934 -4049 938 -4029
rect 938 -4049 968 -4029
rect 1008 -4063 1042 -4051
rect 1008 -4085 1042 -4063
rect 934 -4097 968 -4087
rect 934 -4121 938 -4097
rect 938 -4121 968 -4097
rect 1008 -4131 1042 -4123
rect 1008 -4157 1042 -4131
rect 934 -4165 968 -4159
rect 934 -4193 938 -4165
rect 938 -4193 968 -4165
rect 1008 -4199 1042 -4195
rect 1008 -4229 1042 -4199
rect 934 -4233 968 -4231
rect 934 -4265 938 -4233
rect 938 -4265 968 -4233
rect 1008 -4301 1042 -4267
rect 934 -4335 938 -4303
rect 938 -4335 968 -4303
rect 934 -4337 968 -4335
rect 1008 -4369 1042 -4339
rect 934 -4403 938 -4375
rect 938 -4403 968 -4375
rect 1008 -4373 1042 -4369
rect 934 -4409 968 -4403
rect 1008 -4437 1042 -4411
rect 934 -4471 938 -4447
rect 938 -4471 968 -4447
rect 1008 -4445 1042 -4437
rect 934 -4481 968 -4471
rect 1008 -4505 1042 -4483
rect 934 -4539 938 -4519
rect 938 -4539 968 -4519
rect 1008 -4517 1042 -4505
rect 934 -4553 968 -4539
rect 1008 -4573 1042 -4555
rect 934 -4607 938 -4591
rect 938 -4607 968 -4591
rect 1008 -4589 1042 -4573
rect 934 -4625 968 -4607
rect 1008 -4641 1042 -4627
rect 934 -4675 938 -4663
rect 938 -4675 968 -4663
rect 1008 -4661 1042 -4641
rect 934 -4697 968 -4675
rect 1008 -4709 1042 -4699
rect 934 -4743 938 -4735
rect 938 -4743 968 -4735
rect 1008 -4733 1042 -4709
rect 934 -4769 968 -4743
rect 1008 -4777 1042 -4771
rect 934 -4811 938 -4807
rect 938 -4811 968 -4807
rect 1008 -4805 1042 -4777
rect 934 -4841 968 -4811
rect 1008 -4845 1042 -4843
rect 1008 -4877 1042 -4845
rect 934 -4913 968 -4879
rect 1008 -4947 1042 -4915
rect 1008 -4949 1042 -4947
rect 934 -4981 968 -4951
rect 934 -4985 938 -4981
rect 938 -4985 968 -4981
rect 1008 -5015 1042 -4987
rect 1179 4981 1285 4985
rect 1179 -4981 1285 4981
rect 1179 -4985 1285 -4981
rect 1008 -5021 1042 -5015
rect 934 -5057 968 -5023
rect 1422 -5015 1524 5015
rect 1524 -5015 1528 5015
rect 1422 -5021 1528 -5015
rect 1494 -5057 1528 -5023
rect 1107 -5124 1113 -5090
rect 1113 -5124 1141 -5090
rect 1179 -5124 1181 -5090
rect 1181 -5124 1213 -5090
rect 1251 -5124 1283 -5090
rect 1283 -5124 1285 -5090
rect 1323 -5124 1351 -5090
rect 1351 -5124 1357 -5090
<< metal1 >>
rect 922 5124 1540 5188
rect 922 5090 1107 5124
rect 1141 5090 1179 5124
rect 1213 5090 1251 5124
rect 1285 5090 1323 5124
rect 1357 5090 1540 5124
rect 922 5084 1540 5090
rect 922 5057 1061 5084
tri 1061 5057 1088 5084 nw
tri 1376 5057 1403 5084 ne
rect 1403 5057 1540 5084
rect 922 5023 934 5057
rect 968 5023 1048 5057
tri 1048 5044 1061 5057 nw
tri 1403 5044 1416 5057 ne
rect 922 5021 1048 5023
rect 922 4987 1008 5021
rect 1042 4987 1048 5021
rect 1416 5023 1494 5057
rect 1528 5023 1540 5057
rect 1416 5021 1540 5023
rect 922 4985 1048 4987
rect 922 4951 934 4985
rect 968 4951 1048 4985
rect 922 4949 1048 4951
rect 922 4915 1008 4949
rect 1042 4915 1048 4949
rect 922 4913 1048 4915
rect 922 4879 934 4913
rect 968 4879 1048 4913
rect 922 4877 1048 4879
rect 922 4843 1008 4877
rect 1042 4843 1048 4877
rect 922 4841 1048 4843
rect 922 4807 934 4841
rect 968 4807 1048 4841
rect 922 4805 1048 4807
rect 922 4771 1008 4805
rect 1042 4771 1048 4805
rect 922 4769 1048 4771
rect 922 4735 934 4769
rect 968 4735 1048 4769
rect 922 4733 1048 4735
rect 922 4699 1008 4733
rect 1042 4699 1048 4733
rect 922 4697 1048 4699
rect 922 4663 934 4697
rect 968 4663 1048 4697
rect 922 4661 1048 4663
rect 922 4627 1008 4661
rect 1042 4627 1048 4661
rect 922 4625 1048 4627
rect 922 4591 934 4625
rect 968 4591 1048 4625
rect 922 4589 1048 4591
rect 922 4555 1008 4589
rect 1042 4555 1048 4589
rect 922 4553 1048 4555
rect 922 4519 934 4553
rect 968 4519 1048 4553
rect 922 4517 1048 4519
rect 922 4483 1008 4517
rect 1042 4483 1048 4517
rect 922 4481 1048 4483
rect 922 4447 934 4481
rect 968 4447 1048 4481
rect 922 4445 1048 4447
rect 922 4411 1008 4445
rect 1042 4411 1048 4445
rect 922 4409 1048 4411
rect 922 4375 934 4409
rect 968 4375 1048 4409
rect 922 4373 1048 4375
rect 922 4339 1008 4373
rect 1042 4339 1048 4373
rect 922 4337 1048 4339
rect 922 4303 934 4337
rect 968 4303 1048 4337
rect 922 4301 1048 4303
rect 922 4267 1008 4301
rect 1042 4267 1048 4301
rect 922 4265 1048 4267
rect 922 4231 934 4265
rect 968 4231 1048 4265
rect 922 4229 1048 4231
rect 922 4195 1008 4229
rect 1042 4195 1048 4229
rect 922 4193 1048 4195
rect 922 4159 934 4193
rect 968 4159 1048 4193
rect 922 4157 1048 4159
rect 922 4123 1008 4157
rect 1042 4123 1048 4157
rect 922 4121 1048 4123
rect 922 4087 934 4121
rect 968 4087 1048 4121
rect 922 4085 1048 4087
rect 922 4051 1008 4085
rect 1042 4051 1048 4085
rect 922 4049 1048 4051
rect 922 4015 934 4049
rect 968 4015 1048 4049
rect 922 4013 1048 4015
rect 922 3979 1008 4013
rect 1042 3979 1048 4013
rect 922 3977 1048 3979
rect 922 3943 934 3977
rect 968 3943 1048 3977
rect 922 3941 1048 3943
rect 922 3907 1008 3941
rect 1042 3907 1048 3941
rect 922 3905 1048 3907
rect 922 3871 934 3905
rect 968 3871 1048 3905
rect 922 3869 1048 3871
rect 922 3835 1008 3869
rect 1042 3835 1048 3869
rect 922 3833 1048 3835
rect 922 3799 934 3833
rect 968 3799 1048 3833
rect 922 3797 1048 3799
rect 922 3763 1008 3797
rect 1042 3763 1048 3797
rect 922 3761 1048 3763
rect 922 3727 934 3761
rect 968 3727 1048 3761
rect 922 3725 1048 3727
rect 922 3691 1008 3725
rect 1042 3691 1048 3725
rect 922 3689 1048 3691
rect 922 3655 934 3689
rect 968 3655 1048 3689
rect 922 3653 1048 3655
rect 922 3619 1008 3653
rect 1042 3619 1048 3653
rect 922 3617 1048 3619
rect 922 3583 934 3617
rect 968 3583 1048 3617
rect 922 3581 1048 3583
rect 922 3547 1008 3581
rect 1042 3547 1048 3581
rect 922 3545 1048 3547
rect 922 3511 934 3545
rect 968 3511 1048 3545
rect 922 3509 1048 3511
rect 922 3475 1008 3509
rect 1042 3475 1048 3509
rect 922 3473 1048 3475
rect 922 3439 934 3473
rect 968 3439 1048 3473
rect 922 3437 1048 3439
rect 922 3403 1008 3437
rect 1042 3403 1048 3437
rect 922 3401 1048 3403
rect 922 3367 934 3401
rect 968 3367 1048 3401
rect 922 3365 1048 3367
rect 922 3331 1008 3365
rect 1042 3331 1048 3365
rect 922 3329 1048 3331
rect 922 3295 934 3329
rect 968 3295 1048 3329
rect 922 3293 1048 3295
rect 922 3259 1008 3293
rect 1042 3259 1048 3293
rect 922 3257 1048 3259
rect 922 3223 934 3257
rect 968 3223 1048 3257
rect 922 3221 1048 3223
rect 922 3187 1008 3221
rect 1042 3187 1048 3221
rect 922 3185 1048 3187
rect 922 3151 934 3185
rect 968 3151 1048 3185
rect 922 3149 1048 3151
rect 922 3115 1008 3149
rect 1042 3115 1048 3149
rect 922 3113 1048 3115
rect 922 3079 934 3113
rect 968 3079 1048 3113
rect 922 3077 1048 3079
rect 922 3043 1008 3077
rect 1042 3043 1048 3077
rect 922 3041 1048 3043
rect 922 3007 934 3041
rect 968 3007 1048 3041
rect 922 3005 1048 3007
rect 922 2971 1008 3005
rect 1042 2971 1048 3005
rect 922 2969 1048 2971
rect 922 2935 934 2969
rect 968 2935 1048 2969
rect 922 2933 1048 2935
rect 922 2899 1008 2933
rect 1042 2899 1048 2933
rect 922 2897 1048 2899
rect 922 2863 934 2897
rect 968 2863 1048 2897
rect 922 2861 1048 2863
rect 922 2827 1008 2861
rect 1042 2827 1048 2861
rect 922 2825 1048 2827
rect 922 2791 934 2825
rect 968 2791 1048 2825
rect 922 2789 1048 2791
rect 922 2755 1008 2789
rect 1042 2755 1048 2789
rect 922 2753 1048 2755
rect 922 2719 934 2753
rect 968 2719 1048 2753
rect 922 2717 1048 2719
rect 922 2683 1008 2717
rect 1042 2683 1048 2717
rect 922 2681 1048 2683
rect 922 2647 934 2681
rect 968 2647 1048 2681
rect 922 2645 1048 2647
rect 922 2611 1008 2645
rect 1042 2611 1048 2645
rect 922 2609 1048 2611
rect 922 2575 934 2609
rect 968 2575 1048 2609
rect 922 2573 1048 2575
rect 922 2539 1008 2573
rect 1042 2539 1048 2573
rect 922 2537 1048 2539
rect 922 2503 934 2537
rect 968 2503 1048 2537
rect 922 2501 1048 2503
rect 922 2467 1008 2501
rect 1042 2467 1048 2501
rect 922 2465 1048 2467
rect 922 2431 934 2465
rect 968 2431 1048 2465
rect 922 2429 1048 2431
rect 922 2395 1008 2429
rect 1042 2395 1048 2429
rect 922 2393 1048 2395
rect 922 2359 934 2393
rect 968 2359 1048 2393
rect 922 2357 1048 2359
rect 922 2323 1008 2357
rect 1042 2323 1048 2357
rect 922 2321 1048 2323
rect 922 2287 934 2321
rect 968 2287 1048 2321
rect 922 2285 1048 2287
rect 922 2251 1008 2285
rect 1042 2251 1048 2285
rect 922 2249 1048 2251
rect 922 2215 934 2249
rect 968 2215 1048 2249
rect 922 2213 1048 2215
rect 922 2179 1008 2213
rect 1042 2179 1048 2213
rect 922 2177 1048 2179
rect 922 2143 934 2177
rect 968 2143 1048 2177
rect 922 2141 1048 2143
rect 922 2107 1008 2141
rect 1042 2107 1048 2141
rect 922 2105 1048 2107
rect 922 2071 934 2105
rect 968 2071 1048 2105
rect 922 2069 1048 2071
rect 922 2035 1008 2069
rect 1042 2035 1048 2069
rect 922 2033 1048 2035
rect 922 1999 934 2033
rect 968 1999 1048 2033
rect 922 1997 1048 1999
rect 922 1963 1008 1997
rect 1042 1963 1048 1997
rect 922 1961 1048 1963
rect 922 1927 934 1961
rect 968 1927 1048 1961
rect 922 1925 1048 1927
rect 922 1891 1008 1925
rect 1042 1891 1048 1925
rect 922 1889 1048 1891
rect 922 1855 934 1889
rect 968 1855 1048 1889
rect 922 1853 1048 1855
rect 922 1819 1008 1853
rect 1042 1819 1048 1853
rect 922 1817 1048 1819
rect 922 1783 934 1817
rect 968 1783 1048 1817
rect 922 1781 1048 1783
rect 922 1747 1008 1781
rect 1042 1747 1048 1781
rect 922 1745 1048 1747
rect 922 1711 934 1745
rect 968 1711 1048 1745
rect 922 1709 1048 1711
rect 922 1675 1008 1709
rect 1042 1675 1048 1709
rect 922 1673 1048 1675
rect 922 1639 934 1673
rect 968 1639 1048 1673
rect 922 1637 1048 1639
rect 922 1603 1008 1637
rect 1042 1603 1048 1637
rect 922 1601 1048 1603
rect 922 1567 934 1601
rect 968 1567 1048 1601
rect 922 1565 1048 1567
rect 922 1531 1008 1565
rect 1042 1531 1048 1565
rect 922 1529 1048 1531
rect 922 1495 934 1529
rect 968 1495 1048 1529
rect 922 1493 1048 1495
rect 922 1459 1008 1493
rect 1042 1459 1048 1493
rect 922 1457 1048 1459
rect 922 1423 934 1457
rect 968 1423 1048 1457
rect 922 1421 1048 1423
rect 922 1387 1008 1421
rect 1042 1387 1048 1421
rect 922 1385 1048 1387
rect 922 1351 934 1385
rect 968 1351 1048 1385
rect 922 1349 1048 1351
rect 922 1315 1008 1349
rect 1042 1315 1048 1349
rect 922 1313 1048 1315
rect 922 1279 934 1313
rect 968 1279 1048 1313
rect 922 1277 1048 1279
rect 922 1243 1008 1277
rect 1042 1243 1048 1277
rect 922 1241 1048 1243
rect 922 1207 934 1241
rect 968 1207 1048 1241
rect 922 1205 1048 1207
rect 922 1171 1008 1205
rect 1042 1171 1048 1205
rect 922 1169 1048 1171
rect 922 1135 934 1169
rect 968 1135 1048 1169
rect 922 1133 1048 1135
rect 922 1099 1008 1133
rect 1042 1099 1048 1133
rect 922 1097 1048 1099
rect 922 1063 934 1097
rect 968 1063 1048 1097
rect 922 1061 1048 1063
rect 922 1027 1008 1061
rect 1042 1027 1048 1061
rect 922 1025 1048 1027
rect 922 991 934 1025
rect 968 991 1048 1025
rect 922 989 1048 991
rect 922 955 1008 989
rect 1042 955 1048 989
rect 922 953 1048 955
rect 922 919 934 953
rect 968 919 1048 953
rect 922 917 1048 919
rect 922 883 1008 917
rect 1042 883 1048 917
rect 922 881 1048 883
rect 922 847 934 881
rect 968 847 1048 881
rect 922 845 1048 847
rect 922 811 1008 845
rect 1042 811 1048 845
rect 922 809 1048 811
rect 922 775 934 809
rect 968 775 1048 809
rect 922 773 1048 775
rect 922 739 1008 773
rect 1042 739 1048 773
rect 922 737 1048 739
rect 922 703 934 737
rect 968 703 1048 737
rect 922 701 1048 703
rect 922 667 1008 701
rect 1042 667 1048 701
rect 922 665 1048 667
rect 922 631 934 665
rect 968 631 1048 665
rect 922 629 1048 631
rect 922 595 1008 629
rect 1042 595 1048 629
rect 922 593 1048 595
rect 922 559 934 593
rect 968 559 1048 593
rect 922 557 1048 559
rect 922 523 1008 557
rect 1042 523 1048 557
rect 922 521 1048 523
rect 922 487 934 521
rect 968 487 1048 521
rect 922 485 1048 487
rect 922 451 1008 485
rect 1042 451 1048 485
rect 922 449 1048 451
rect 922 415 934 449
rect 968 415 1048 449
rect 922 413 1048 415
rect 922 379 1008 413
rect 1042 379 1048 413
rect 922 377 1048 379
rect 922 343 934 377
rect 968 343 1048 377
rect 922 341 1048 343
rect 922 307 1008 341
rect 1042 307 1048 341
rect 922 305 1048 307
rect 922 271 934 305
rect 968 271 1048 305
rect 922 269 1048 271
rect 922 235 1008 269
rect 1042 235 1048 269
rect 922 233 1048 235
rect 922 199 934 233
rect 968 199 1048 233
rect 922 197 1048 199
rect 922 163 1008 197
rect 1042 163 1048 197
rect 922 161 1048 163
rect 922 127 934 161
rect 968 127 1048 161
rect 922 125 1048 127
rect 922 91 1008 125
rect 1042 91 1048 125
rect 922 89 1048 91
rect 922 55 934 89
rect 968 55 1048 89
rect 922 53 1048 55
rect 922 19 1008 53
rect 1042 19 1048 53
rect 922 17 1048 19
rect 922 -17 934 17
rect 968 -17 1048 17
rect 922 -19 1048 -17
rect 922 -53 1008 -19
rect 1042 -53 1048 -19
rect 922 -55 1048 -53
rect 922 -89 934 -55
rect 968 -89 1048 -55
rect 922 -91 1048 -89
rect 922 -125 1008 -91
rect 1042 -125 1048 -91
rect 922 -127 1048 -125
rect 922 -161 934 -127
rect 968 -161 1048 -127
rect 922 -163 1048 -161
rect 922 -197 1008 -163
rect 1042 -197 1048 -163
rect 922 -199 1048 -197
rect 922 -233 934 -199
rect 968 -233 1048 -199
rect 922 -235 1048 -233
rect 922 -269 1008 -235
rect 1042 -269 1048 -235
rect 922 -271 1048 -269
rect 922 -305 934 -271
rect 968 -305 1048 -271
rect 922 -307 1048 -305
rect 922 -341 1008 -307
rect 1042 -341 1048 -307
rect 922 -343 1048 -341
rect 922 -377 934 -343
rect 968 -377 1048 -343
rect 922 -379 1048 -377
rect 922 -413 1008 -379
rect 1042 -413 1048 -379
rect 922 -415 1048 -413
rect 922 -449 934 -415
rect 968 -449 1048 -415
rect 922 -451 1048 -449
rect 922 -485 1008 -451
rect 1042 -485 1048 -451
rect 922 -487 1048 -485
rect 922 -521 934 -487
rect 968 -521 1048 -487
rect 922 -523 1048 -521
rect 922 -557 1008 -523
rect 1042 -557 1048 -523
rect 922 -559 1048 -557
rect 922 -593 934 -559
rect 968 -593 1048 -559
rect 922 -595 1048 -593
rect 922 -629 1008 -595
rect 1042 -629 1048 -595
rect 922 -631 1048 -629
rect 922 -665 934 -631
rect 968 -665 1048 -631
rect 922 -667 1048 -665
rect 922 -701 1008 -667
rect 1042 -701 1048 -667
rect 922 -703 1048 -701
rect 922 -737 934 -703
rect 968 -737 1048 -703
rect 922 -739 1048 -737
rect 922 -773 1008 -739
rect 1042 -773 1048 -739
rect 922 -775 1048 -773
rect 922 -809 934 -775
rect 968 -809 1048 -775
rect 922 -811 1048 -809
rect 922 -845 1008 -811
rect 1042 -845 1048 -811
rect 922 -847 1048 -845
rect 922 -881 934 -847
rect 968 -881 1048 -847
rect 922 -883 1048 -881
rect 922 -917 1008 -883
rect 1042 -917 1048 -883
rect 922 -919 1048 -917
rect 922 -953 934 -919
rect 968 -953 1048 -919
rect 922 -955 1048 -953
rect 922 -989 1008 -955
rect 1042 -989 1048 -955
rect 922 -991 1048 -989
rect 922 -1025 934 -991
rect 968 -1025 1048 -991
rect 922 -1027 1048 -1025
rect 922 -1061 1008 -1027
rect 1042 -1061 1048 -1027
rect 922 -1063 1048 -1061
rect 922 -1097 934 -1063
rect 968 -1097 1048 -1063
rect 922 -1099 1048 -1097
rect 922 -1133 1008 -1099
rect 1042 -1133 1048 -1099
rect 922 -1135 1048 -1133
rect 922 -1169 934 -1135
rect 968 -1169 1048 -1135
rect 922 -1171 1048 -1169
rect 922 -1205 1008 -1171
rect 1042 -1205 1048 -1171
rect 922 -1207 1048 -1205
rect 922 -1241 934 -1207
rect 968 -1241 1048 -1207
rect 922 -1243 1048 -1241
rect 922 -1277 1008 -1243
rect 1042 -1277 1048 -1243
rect 922 -1279 1048 -1277
rect 922 -1313 934 -1279
rect 968 -1313 1048 -1279
rect 922 -1315 1048 -1313
rect 922 -1349 1008 -1315
rect 1042 -1349 1048 -1315
rect 922 -1351 1048 -1349
rect 922 -1385 934 -1351
rect 968 -1385 1048 -1351
rect 922 -1387 1048 -1385
rect 922 -1421 1008 -1387
rect 1042 -1421 1048 -1387
rect 922 -1423 1048 -1421
rect 922 -1457 934 -1423
rect 968 -1457 1048 -1423
rect 922 -1459 1048 -1457
rect 922 -1493 1008 -1459
rect 1042 -1493 1048 -1459
rect 922 -1495 1048 -1493
rect 922 -1529 934 -1495
rect 968 -1529 1048 -1495
rect 922 -1531 1048 -1529
rect 922 -1565 1008 -1531
rect 1042 -1565 1048 -1531
rect 922 -1567 1048 -1565
rect 922 -1601 934 -1567
rect 968 -1601 1048 -1567
rect 922 -1603 1048 -1601
rect 922 -1637 1008 -1603
rect 1042 -1637 1048 -1603
rect 922 -1639 1048 -1637
rect 922 -1673 934 -1639
rect 968 -1673 1048 -1639
rect 922 -1675 1048 -1673
rect 922 -1709 1008 -1675
rect 1042 -1709 1048 -1675
rect 922 -1711 1048 -1709
rect 922 -1745 934 -1711
rect 968 -1745 1048 -1711
rect 922 -1747 1048 -1745
rect 922 -1781 1008 -1747
rect 1042 -1781 1048 -1747
rect 922 -1783 1048 -1781
rect 922 -1817 934 -1783
rect 968 -1817 1048 -1783
rect 922 -1819 1048 -1817
rect 922 -1853 1008 -1819
rect 1042 -1853 1048 -1819
rect 922 -1855 1048 -1853
rect 922 -1889 934 -1855
rect 968 -1889 1048 -1855
rect 922 -1891 1048 -1889
rect 922 -1925 1008 -1891
rect 1042 -1925 1048 -1891
rect 922 -1927 1048 -1925
rect 922 -1961 934 -1927
rect 968 -1961 1048 -1927
rect 922 -1963 1048 -1961
rect 922 -1997 1008 -1963
rect 1042 -1997 1048 -1963
rect 922 -1999 1048 -1997
rect 922 -2033 934 -1999
rect 968 -2033 1048 -1999
rect 922 -2035 1048 -2033
rect 922 -2069 1008 -2035
rect 1042 -2069 1048 -2035
rect 922 -2071 1048 -2069
rect 922 -2105 934 -2071
rect 968 -2105 1048 -2071
rect 922 -2107 1048 -2105
rect 922 -2141 1008 -2107
rect 1042 -2141 1048 -2107
rect 922 -2143 1048 -2141
rect 922 -2177 934 -2143
rect 968 -2177 1048 -2143
rect 922 -2179 1048 -2177
rect 922 -2213 1008 -2179
rect 1042 -2213 1048 -2179
rect 922 -2215 1048 -2213
rect 922 -2249 934 -2215
rect 968 -2249 1048 -2215
rect 922 -2251 1048 -2249
rect 922 -2285 1008 -2251
rect 1042 -2285 1048 -2251
rect 922 -2287 1048 -2285
rect 922 -2321 934 -2287
rect 968 -2321 1048 -2287
rect 922 -2323 1048 -2321
rect 922 -2357 1008 -2323
rect 1042 -2357 1048 -2323
rect 922 -2359 1048 -2357
rect 922 -2393 934 -2359
rect 968 -2393 1048 -2359
rect 922 -2395 1048 -2393
rect 922 -2429 1008 -2395
rect 1042 -2429 1048 -2395
rect 922 -2431 1048 -2429
rect 922 -2465 934 -2431
rect 968 -2465 1048 -2431
rect 922 -2467 1048 -2465
rect 922 -2501 1008 -2467
rect 1042 -2501 1048 -2467
rect 922 -2503 1048 -2501
rect 922 -2537 934 -2503
rect 968 -2537 1048 -2503
rect 922 -2539 1048 -2537
rect 922 -2573 1008 -2539
rect 1042 -2573 1048 -2539
rect 922 -2575 1048 -2573
rect 922 -2609 934 -2575
rect 968 -2609 1048 -2575
rect 922 -2611 1048 -2609
rect 922 -2645 1008 -2611
rect 1042 -2645 1048 -2611
rect 922 -2647 1048 -2645
rect 922 -2681 934 -2647
rect 968 -2681 1048 -2647
rect 922 -2683 1048 -2681
rect 922 -2717 1008 -2683
rect 1042 -2717 1048 -2683
rect 922 -2719 1048 -2717
rect 922 -2753 934 -2719
rect 968 -2753 1048 -2719
rect 922 -2755 1048 -2753
rect 922 -2789 1008 -2755
rect 1042 -2789 1048 -2755
rect 922 -2791 1048 -2789
rect 922 -2825 934 -2791
rect 968 -2825 1048 -2791
rect 922 -2827 1048 -2825
rect 922 -2861 1008 -2827
rect 1042 -2861 1048 -2827
rect 922 -2863 1048 -2861
rect 922 -2897 934 -2863
rect 968 -2897 1048 -2863
rect 922 -2899 1048 -2897
rect 922 -2933 1008 -2899
rect 1042 -2933 1048 -2899
rect 922 -2935 1048 -2933
rect 922 -2969 934 -2935
rect 968 -2969 1048 -2935
rect 922 -2971 1048 -2969
rect 922 -3005 1008 -2971
rect 1042 -3005 1048 -2971
rect 922 -3007 1048 -3005
rect 922 -3041 934 -3007
rect 968 -3041 1048 -3007
rect 922 -3043 1048 -3041
rect 922 -3077 1008 -3043
rect 1042 -3077 1048 -3043
rect 922 -3079 1048 -3077
rect 922 -3113 934 -3079
rect 968 -3113 1048 -3079
rect 922 -3115 1048 -3113
rect 922 -3149 1008 -3115
rect 1042 -3149 1048 -3115
rect 922 -3151 1048 -3149
rect 922 -3185 934 -3151
rect 968 -3185 1048 -3151
rect 922 -3187 1048 -3185
rect 922 -3221 1008 -3187
rect 1042 -3221 1048 -3187
rect 922 -3223 1048 -3221
rect 922 -3257 934 -3223
rect 968 -3257 1048 -3223
rect 922 -3259 1048 -3257
rect 922 -3293 1008 -3259
rect 1042 -3293 1048 -3259
rect 922 -3295 1048 -3293
rect 922 -3329 934 -3295
rect 968 -3329 1048 -3295
rect 922 -3331 1048 -3329
rect 922 -3365 1008 -3331
rect 1042 -3365 1048 -3331
rect 922 -3367 1048 -3365
rect 922 -3401 934 -3367
rect 968 -3401 1048 -3367
rect 922 -3403 1048 -3401
rect 922 -3437 1008 -3403
rect 1042 -3437 1048 -3403
rect 922 -3439 1048 -3437
rect 922 -3473 934 -3439
rect 968 -3473 1048 -3439
rect 922 -3475 1048 -3473
rect 922 -3509 1008 -3475
rect 1042 -3509 1048 -3475
rect 922 -3511 1048 -3509
rect 922 -3545 934 -3511
rect 968 -3545 1048 -3511
rect 922 -3547 1048 -3545
rect 922 -3581 1008 -3547
rect 1042 -3581 1048 -3547
rect 922 -3583 1048 -3581
rect 922 -3617 934 -3583
rect 968 -3617 1048 -3583
rect 922 -3619 1048 -3617
rect 922 -3653 1008 -3619
rect 1042 -3653 1048 -3619
rect 922 -3655 1048 -3653
rect 922 -3689 934 -3655
rect 968 -3689 1048 -3655
rect 922 -3691 1048 -3689
rect 922 -3725 1008 -3691
rect 1042 -3725 1048 -3691
rect 922 -3727 1048 -3725
rect 922 -3761 934 -3727
rect 968 -3761 1048 -3727
rect 922 -3763 1048 -3761
rect 922 -3797 1008 -3763
rect 1042 -3797 1048 -3763
rect 922 -3799 1048 -3797
rect 922 -3833 934 -3799
rect 968 -3833 1048 -3799
rect 922 -3835 1048 -3833
rect 922 -3869 1008 -3835
rect 1042 -3869 1048 -3835
rect 922 -3871 1048 -3869
rect 922 -3905 934 -3871
rect 968 -3905 1048 -3871
rect 922 -3907 1048 -3905
rect 922 -3941 1008 -3907
rect 1042 -3941 1048 -3907
rect 922 -3943 1048 -3941
rect 922 -3977 934 -3943
rect 968 -3977 1048 -3943
rect 922 -3979 1048 -3977
rect 922 -4013 1008 -3979
rect 1042 -4013 1048 -3979
rect 922 -4015 1048 -4013
rect 922 -4049 934 -4015
rect 968 -4049 1048 -4015
rect 922 -4051 1048 -4049
rect 922 -4085 1008 -4051
rect 1042 -4085 1048 -4051
rect 922 -4087 1048 -4085
rect 922 -4121 934 -4087
rect 968 -4121 1048 -4087
rect 922 -4123 1048 -4121
rect 922 -4157 1008 -4123
rect 1042 -4157 1048 -4123
rect 922 -4159 1048 -4157
rect 922 -4193 934 -4159
rect 968 -4193 1048 -4159
rect 922 -4195 1048 -4193
rect 922 -4229 1008 -4195
rect 1042 -4229 1048 -4195
rect 922 -4231 1048 -4229
rect 922 -4265 934 -4231
rect 968 -4265 1048 -4231
rect 922 -4267 1048 -4265
rect 922 -4301 1008 -4267
rect 1042 -4301 1048 -4267
rect 922 -4303 1048 -4301
rect 922 -4337 934 -4303
rect 968 -4337 1048 -4303
rect 922 -4339 1048 -4337
rect 922 -4373 1008 -4339
rect 1042 -4373 1048 -4339
rect 922 -4375 1048 -4373
rect 922 -4409 934 -4375
rect 968 -4409 1048 -4375
rect 922 -4411 1048 -4409
rect 922 -4445 1008 -4411
rect 1042 -4445 1048 -4411
rect 922 -4447 1048 -4445
rect 922 -4481 934 -4447
rect 968 -4481 1048 -4447
rect 922 -4483 1048 -4481
rect 922 -4517 1008 -4483
rect 1042 -4517 1048 -4483
rect 922 -4519 1048 -4517
rect 922 -4553 934 -4519
rect 968 -4553 1048 -4519
rect 922 -4555 1048 -4553
rect 922 -4589 1008 -4555
rect 1042 -4589 1048 -4555
rect 922 -4591 1048 -4589
rect 922 -4625 934 -4591
rect 968 -4625 1048 -4591
rect 922 -4627 1048 -4625
rect 922 -4661 1008 -4627
rect 1042 -4661 1048 -4627
rect 922 -4663 1048 -4661
rect 922 -4697 934 -4663
rect 968 -4697 1048 -4663
rect 922 -4699 1048 -4697
rect 922 -4733 1008 -4699
rect 1042 -4733 1048 -4699
rect 922 -4735 1048 -4733
rect 922 -4769 934 -4735
rect 968 -4769 1048 -4735
rect 922 -4771 1048 -4769
rect 922 -4805 1008 -4771
rect 1042 -4805 1048 -4771
rect 922 -4807 1048 -4805
rect 922 -4841 934 -4807
rect 968 -4841 1048 -4807
rect 922 -4843 1048 -4841
rect 922 -4877 1008 -4843
rect 1042 -4877 1048 -4843
rect 922 -4879 1048 -4877
rect 922 -4913 934 -4879
rect 968 -4913 1048 -4879
rect 922 -4915 1048 -4913
rect 922 -4949 1008 -4915
rect 1042 -4949 1048 -4915
rect 922 -4951 1048 -4949
rect 922 -4985 934 -4951
rect 968 -4985 1048 -4951
rect 922 -4987 1048 -4985
rect 922 -5021 1008 -4987
rect 1042 -5021 1048 -4987
tri 1138 5000 1158 5020 se
rect 1158 5000 1306 5020
tri 1306 5000 1326 5020 sw
rect 1138 4985 1326 5000
rect 1138 -4985 1179 4985
rect 1285 -4985 1326 4985
rect 1138 -5000 1326 -4985
tri 1138 -5020 1158 -5000 ne
rect 1158 -5020 1306 -5000
tri 1306 -5020 1326 -5000 nw
rect 922 -5023 1048 -5021
rect 922 -5057 934 -5023
rect 968 -5057 1048 -5023
rect 1416 -5021 1422 5021
rect 1528 -5021 1540 5021
rect 1416 -5023 1540 -5021
tri 1048 -5057 1061 -5044 sw
tri 1403 -5057 1416 -5044 se
rect 1416 -5057 1494 -5023
rect 1528 -5057 1540 -5023
rect 922 -5084 1061 -5057
tri 1061 -5084 1088 -5057 sw
tri 1398 -5062 1403 -5057 se
rect 1403 -5062 1540 -5057
tri 1376 -5084 1398 -5062 se
rect 1398 -5084 1540 -5062
rect 922 -5090 1540 -5084
rect 922 -5124 1107 -5090
rect 1141 -5124 1179 -5090
rect 1213 -5124 1251 -5090
rect 1285 -5124 1323 -5090
rect 1357 -5124 1540 -5090
rect 922 -5188 1540 -5124
<< properties >>
string FIXED_BBOX 1024 -5106 1438 5106
string GDS_END 5365438
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io__analog.gds
string GDS_START 5241946
<< end >>
