magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -38 261 1234 582
<< pwell >>
rect 29 21 1171 203
rect 29 -17 63 21
<< scnmos >>
rect 107 47 137 177
rect 191 47 221 177
rect 275 47 305 177
rect 359 47 389 177
rect 443 47 473 177
rect 615 47 645 177
rect 699 47 729 177
rect 783 47 813 177
rect 979 47 1009 177
rect 1063 47 1093 177
<< scpmoshvt >>
rect 103 297 133 497
rect 187 297 217 497
rect 271 297 301 497
rect 355 297 385 497
rect 543 297 573 497
rect 627 297 657 497
rect 711 297 741 497
rect 863 297 893 497
rect 975 297 1005 497
rect 1059 297 1089 497
<< ndiff >>
rect 55 129 107 177
rect 55 95 63 129
rect 97 95 107 129
rect 55 47 107 95
rect 137 89 191 177
rect 137 55 147 89
rect 181 55 191 89
rect 137 47 191 55
rect 221 129 275 177
rect 221 95 231 129
rect 265 95 275 129
rect 221 47 275 95
rect 305 89 359 177
rect 305 55 315 89
rect 349 55 359 89
rect 305 47 359 55
rect 389 129 443 177
rect 389 95 399 129
rect 433 95 443 129
rect 389 47 443 95
rect 473 89 615 177
rect 473 55 493 89
rect 527 55 561 89
rect 595 55 615 89
rect 473 47 615 55
rect 645 129 699 177
rect 645 95 655 129
rect 689 95 699 129
rect 645 47 699 95
rect 729 89 783 177
rect 729 55 739 89
rect 773 55 783 89
rect 729 47 783 55
rect 813 169 869 177
rect 813 135 823 169
rect 857 135 869 169
rect 813 47 869 135
rect 923 169 979 177
rect 923 135 935 169
rect 969 135 979 169
rect 923 47 979 135
rect 1009 89 1063 177
rect 1009 55 1019 89
rect 1053 55 1063 89
rect 1009 47 1063 55
rect 1093 129 1145 177
rect 1093 95 1103 129
rect 1137 95 1145 129
rect 1093 47 1145 95
<< pdiff >>
rect 51 448 103 497
rect 51 414 59 448
rect 93 414 103 448
rect 51 380 103 414
rect 51 346 59 380
rect 93 346 103 380
rect 51 297 103 346
rect 133 489 187 497
rect 133 455 143 489
rect 177 455 187 489
rect 133 421 187 455
rect 133 387 143 421
rect 177 387 187 421
rect 133 297 187 387
rect 217 448 271 497
rect 217 414 227 448
rect 261 414 271 448
rect 217 380 271 414
rect 217 346 227 380
rect 261 346 271 380
rect 217 297 271 346
rect 301 489 355 497
rect 301 455 311 489
rect 345 455 355 489
rect 301 421 355 455
rect 301 387 311 421
rect 345 387 355 421
rect 301 297 355 387
rect 385 380 437 497
rect 385 346 395 380
rect 429 346 437 380
rect 385 297 437 346
rect 491 380 543 497
rect 491 346 499 380
rect 533 346 543 380
rect 491 297 543 346
rect 573 489 627 497
rect 573 455 583 489
rect 617 455 627 489
rect 573 421 627 455
rect 573 387 583 421
rect 617 387 627 421
rect 573 297 627 387
rect 657 448 711 497
rect 657 414 667 448
rect 701 414 711 448
rect 657 380 711 414
rect 657 346 667 380
rect 701 346 711 380
rect 657 297 711 346
rect 741 489 863 497
rect 741 387 751 489
rect 853 387 863 489
rect 741 297 863 387
rect 893 448 975 497
rect 893 414 917 448
rect 951 414 975 448
rect 893 380 975 414
rect 893 346 917 380
rect 951 346 975 380
rect 893 297 975 346
rect 1005 489 1059 497
rect 1005 455 1015 489
rect 1049 455 1059 489
rect 1005 421 1059 455
rect 1005 387 1015 421
rect 1049 387 1059 421
rect 1005 297 1059 387
rect 1089 448 1141 497
rect 1089 414 1099 448
rect 1133 414 1141 448
rect 1089 380 1141 414
rect 1089 346 1099 380
rect 1133 346 1141 380
rect 1089 297 1141 346
<< ndiffc >>
rect 63 95 97 129
rect 147 55 181 89
rect 231 95 265 129
rect 315 55 349 89
rect 399 95 433 129
rect 493 55 527 89
rect 561 55 595 89
rect 655 95 689 129
rect 739 55 773 89
rect 823 135 857 169
rect 935 135 969 169
rect 1019 55 1053 89
rect 1103 95 1137 129
<< pdiffc >>
rect 59 414 93 448
rect 59 346 93 380
rect 143 455 177 489
rect 143 387 177 421
rect 227 414 261 448
rect 227 346 261 380
rect 311 455 345 489
rect 311 387 345 421
rect 395 346 429 380
rect 499 346 533 380
rect 583 455 617 489
rect 583 387 617 421
rect 667 414 701 448
rect 667 346 701 380
rect 751 387 853 489
rect 917 414 951 448
rect 917 346 951 380
rect 1015 455 1049 489
rect 1015 387 1049 421
rect 1099 414 1133 448
rect 1099 346 1133 380
<< poly >>
rect 103 497 133 523
rect 187 497 217 523
rect 271 497 301 523
rect 355 497 385 523
rect 543 497 573 523
rect 627 497 657 523
rect 711 497 741 523
rect 863 497 893 523
rect 975 497 1005 523
rect 1059 497 1089 523
rect 103 259 133 297
rect 187 259 217 297
rect 271 259 301 297
rect 355 259 385 297
rect 543 259 573 297
rect 627 259 657 297
rect 711 259 741 297
rect 863 259 893 297
rect 87 249 221 259
rect 87 215 103 249
rect 137 215 171 249
rect 205 215 221 249
rect 87 205 221 215
rect 263 249 397 259
rect 263 215 279 249
rect 313 215 347 249
rect 381 215 397 249
rect 263 205 397 215
rect 443 249 657 259
rect 443 215 481 249
rect 515 215 549 249
rect 583 215 657 249
rect 443 205 657 215
rect 699 249 893 259
rect 699 215 715 249
rect 749 215 783 249
rect 817 215 893 249
rect 699 205 893 215
rect 975 259 1005 297
rect 1059 259 1089 297
rect 975 249 1151 259
rect 975 215 1033 249
rect 1067 215 1101 249
rect 1135 215 1151 249
rect 975 205 1151 215
rect 107 177 137 205
rect 191 177 221 205
rect 275 177 305 205
rect 359 177 389 205
rect 443 177 473 205
rect 615 177 645 205
rect 699 177 729 205
rect 783 177 813 205
rect 979 177 1009 205
rect 1063 177 1093 205
rect 107 21 137 47
rect 191 21 221 47
rect 275 21 305 47
rect 359 21 389 47
rect 443 21 473 47
rect 615 21 645 47
rect 699 21 729 47
rect 783 21 813 47
rect 979 21 1009 47
rect 1063 21 1093 47
<< polycont >>
rect 103 215 137 249
rect 171 215 205 249
rect 279 215 313 249
rect 347 215 381 249
rect 481 215 515 249
rect 549 215 583 249
rect 715 215 749 249
rect 783 215 817 249
rect 1033 215 1067 249
rect 1101 215 1135 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 17 448 93 493
rect 17 414 59 448
rect 17 380 93 414
rect 17 346 59 380
rect 127 489 193 527
rect 127 455 143 489
rect 177 455 193 489
rect 127 421 193 455
rect 127 387 143 421
rect 177 387 193 421
rect 127 379 193 387
rect 227 448 261 493
rect 227 380 261 414
rect 17 345 93 346
rect 295 489 633 493
rect 295 455 311 489
rect 345 459 583 489
rect 345 455 361 459
rect 295 421 361 455
rect 567 455 583 459
rect 617 455 633 489
rect 295 387 311 421
rect 345 387 361 421
rect 295 379 361 387
rect 395 380 445 425
rect 227 345 261 346
rect 429 346 445 380
rect 395 345 445 346
rect 17 297 445 345
rect 483 380 533 425
rect 483 346 499 380
rect 567 421 633 455
rect 567 387 583 421
rect 617 387 633 421
rect 567 379 633 387
rect 667 448 701 493
rect 667 380 701 414
rect 483 345 533 346
rect 735 489 869 527
rect 735 387 751 489
rect 853 387 869 489
rect 735 379 869 387
rect 903 448 965 493
rect 903 414 917 448
rect 951 414 965 448
rect 903 380 965 414
rect 667 345 701 346
rect 903 346 917 380
rect 951 346 965 380
rect 999 489 1065 527
rect 999 455 1015 489
rect 1049 455 1065 489
rect 999 421 1065 455
rect 999 387 1015 421
rect 1049 387 1065 421
rect 999 379 1065 387
rect 1099 448 1179 493
rect 1133 414 1179 448
rect 1099 380 1179 414
rect 903 345 965 346
rect 1133 346 1179 380
rect 1099 345 1179 346
rect 483 297 1179 345
rect 17 249 221 263
rect 17 215 103 249
rect 137 215 171 249
rect 205 215 221 249
rect 17 211 221 215
rect 255 249 431 263
rect 255 215 279 249
rect 313 215 347 249
rect 381 215 431 249
rect 255 211 431 215
rect 465 249 615 263
rect 465 215 481 249
rect 515 215 549 249
rect 583 215 615 249
rect 465 211 615 215
rect 673 249 877 263
rect 673 215 715 249
rect 749 215 783 249
rect 817 215 877 249
rect 673 211 877 215
rect 911 177 983 297
rect 1017 249 1179 263
rect 1017 215 1033 249
rect 1067 215 1101 249
rect 1135 215 1179 249
rect 1017 211 1179 215
rect 17 169 877 177
rect 17 135 823 169
rect 857 135 877 169
rect 17 131 877 135
rect 911 169 1179 177
rect 911 135 935 169
rect 969 135 1179 169
rect 911 131 1179 135
rect 17 129 97 131
rect 17 95 63 129
rect 231 129 265 131
rect 17 51 97 95
rect 131 89 197 97
rect 131 55 147 89
rect 181 55 197 89
rect 131 17 197 55
rect 399 129 433 131
rect 231 51 265 95
rect 299 89 365 97
rect 299 55 315 89
rect 349 55 365 89
rect 299 17 365 55
rect 655 129 689 131
rect 399 51 433 95
rect 467 89 621 97
rect 467 55 493 89
rect 527 55 561 89
rect 595 55 621 89
rect 467 17 621 55
rect 1103 129 1179 131
rect 655 51 689 95
rect 723 89 1069 97
rect 723 55 739 89
rect 773 55 1019 89
rect 1053 55 1069 89
rect 723 51 1069 55
rect 1137 95 1179 129
rect 1103 51 1179 95
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
flabel locali s 29 221 63 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 949 221 983 255 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 1133 221 1167 255 0 FreeSans 200 0 0 0 C1
port 5 nsew signal input
flabel locali s 1041 221 1075 255 0 FreeSans 200 0 0 0 C1
port 5 nsew signal input
flabel locali s 765 221 799 255 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 673 221 707 255 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 581 221 615 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 489 221 523 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 397 221 431 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 305 221 339 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 121 221 155 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 489 357 523 391 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 949 289 983 323 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 1133 425 1167 459 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 1133 357 1167 391 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 1133 85 1167 119 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 949 153 983 187 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional abutment
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 o311ai_2
rlabel metal1 s 0 -48 1196 48 1 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1196 592 1 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1196 544
string GDS_END 902188
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 891792
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 5.980 0.000 
<< end >>
