magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect 11776 2435 12131 3859
rect 11973 1496 12623 1911
rect 8626 697 9486 1429
<< pwell >>
rect 8774 1597 9446 1849
<< mvnmos >>
rect 8867 1623 8987 1823
rect 9043 1623 9163 1823
rect 9247 1623 9367 1823
<< mvpmos >>
rect 8867 763 8987 1363
rect 9043 763 9163 1363
rect 9247 763 9367 1363
<< mvndiff >>
rect 8800 1805 8867 1823
rect 8800 1771 8808 1805
rect 8842 1771 8867 1805
rect 8800 1737 8867 1771
rect 8800 1703 8808 1737
rect 8842 1703 8867 1737
rect 8800 1669 8867 1703
rect 8800 1635 8808 1669
rect 8842 1635 8867 1669
rect 8800 1623 8867 1635
rect 8987 1805 9043 1823
rect 8987 1771 8998 1805
rect 9032 1771 9043 1805
rect 8987 1737 9043 1771
rect 8987 1703 8998 1737
rect 9032 1703 9043 1737
rect 8987 1669 9043 1703
rect 8987 1635 8998 1669
rect 9032 1635 9043 1669
rect 8987 1623 9043 1635
rect 9163 1805 9247 1823
rect 9163 1771 9188 1805
rect 9222 1771 9247 1805
rect 9163 1737 9247 1771
rect 9163 1703 9188 1737
rect 9222 1703 9247 1737
rect 9163 1669 9247 1703
rect 9163 1635 9188 1669
rect 9222 1635 9247 1669
rect 9163 1623 9247 1635
rect 9367 1805 9420 1823
rect 9367 1771 9378 1805
rect 9412 1771 9420 1805
rect 9367 1737 9420 1771
rect 9367 1703 9378 1737
rect 9412 1703 9420 1737
rect 9367 1669 9420 1703
rect 9367 1635 9378 1669
rect 9412 1635 9420 1669
rect 9367 1623 9420 1635
<< mvpdiff >>
rect 8800 1351 8867 1363
rect 8800 1317 8808 1351
rect 8842 1317 8867 1351
rect 8800 1283 8867 1317
rect 8800 1249 8808 1283
rect 8842 1249 8867 1283
rect 8800 1215 8867 1249
rect 8800 1181 8808 1215
rect 8842 1181 8867 1215
rect 8800 1147 8867 1181
rect 8800 1113 8808 1147
rect 8842 1113 8867 1147
rect 8800 1079 8867 1113
rect 8800 1045 8808 1079
rect 8842 1045 8867 1079
rect 8800 1011 8867 1045
rect 8800 977 8808 1011
rect 8842 977 8867 1011
rect 8800 943 8867 977
rect 8800 909 8808 943
rect 8842 909 8867 943
rect 8800 875 8867 909
rect 8800 841 8808 875
rect 8842 841 8867 875
rect 8800 763 8867 841
rect 8987 763 9043 1363
rect 9163 1351 9247 1363
rect 9163 1317 9188 1351
rect 9222 1317 9247 1351
rect 9163 1283 9247 1317
rect 9163 1249 9188 1283
rect 9222 1249 9247 1283
rect 9163 1215 9247 1249
rect 9163 1181 9188 1215
rect 9222 1181 9247 1215
rect 9163 1147 9247 1181
rect 9163 1113 9188 1147
rect 9222 1113 9247 1147
rect 9163 1079 9247 1113
rect 9163 1045 9188 1079
rect 9222 1045 9247 1079
rect 9163 1011 9247 1045
rect 9163 977 9188 1011
rect 9222 977 9247 1011
rect 9163 943 9247 977
rect 9163 909 9188 943
rect 9222 909 9247 943
rect 9163 875 9247 909
rect 9163 841 9188 875
rect 9222 841 9247 875
rect 9163 763 9247 841
rect 9367 1351 9420 1363
rect 9367 1317 9378 1351
rect 9412 1317 9420 1351
rect 9367 1283 9420 1317
rect 9367 1249 9378 1283
rect 9412 1249 9420 1283
rect 9367 1215 9420 1249
rect 9367 1181 9378 1215
rect 9412 1181 9420 1215
rect 9367 1147 9420 1181
rect 9367 1113 9378 1147
rect 9412 1113 9420 1147
rect 9367 1079 9420 1113
rect 9367 1045 9378 1079
rect 9412 1045 9420 1079
rect 9367 1011 9420 1045
rect 9367 977 9378 1011
rect 9412 977 9420 1011
rect 9367 943 9420 977
rect 9367 909 9378 943
rect 9412 909 9420 943
rect 9367 875 9420 909
rect 9367 841 9378 875
rect 9412 841 9420 875
rect 9367 763 9420 841
<< mvndiffc >>
rect 8808 1771 8842 1805
rect 8808 1703 8842 1737
rect 8808 1635 8842 1669
rect 8998 1771 9032 1805
rect 8998 1703 9032 1737
rect 8998 1635 9032 1669
rect 9188 1771 9222 1805
rect 9188 1703 9222 1737
rect 9188 1635 9222 1669
rect 9378 1771 9412 1805
rect 9378 1703 9412 1737
rect 9378 1635 9412 1669
<< mvpdiffc >>
rect 8808 1317 8842 1351
rect 8808 1249 8842 1283
rect 8808 1181 8842 1215
rect 8808 1113 8842 1147
rect 8808 1045 8842 1079
rect 8808 977 8842 1011
rect 8808 909 8842 943
rect 8808 841 8842 875
rect 9188 1317 9222 1351
rect 9188 1249 9222 1283
rect 9188 1181 9222 1215
rect 9188 1113 9222 1147
rect 9188 1045 9222 1079
rect 9188 977 9222 1011
rect 9188 909 9222 943
rect 9188 841 9222 875
rect 9378 1317 9412 1351
rect 9378 1249 9412 1283
rect 9378 1181 9412 1215
rect 9378 1113 9412 1147
rect 9378 1045 9412 1079
rect 9378 977 9412 1011
rect 9378 909 9412 943
rect 9378 841 9412 875
<< mvnsubdiff >>
rect 8692 1339 8726 1363
rect 8692 1265 8726 1305
rect 8692 1191 8726 1231
rect 8692 1117 8726 1157
rect 8692 1043 8726 1083
rect 8692 969 8726 1009
rect 8692 895 8726 935
rect 8692 821 8726 861
rect 8692 763 8726 787
<< mvnsubdiffcont >>
rect 8692 1305 8726 1339
rect 8692 1231 8726 1265
rect 8692 1157 8726 1191
rect 8692 1083 8726 1117
rect 8692 1009 8726 1043
rect 8692 935 8726 969
rect 8692 861 8726 895
rect 8692 787 8726 821
<< poly >>
rect 8867 1823 8987 1849
rect 9043 1823 9163 1849
rect 9247 1823 9367 1849
rect 8867 1513 8987 1623
rect 8867 1479 8910 1513
rect 8944 1479 8987 1513
rect 8867 1445 8987 1479
rect 8867 1411 8910 1445
rect 8944 1411 8987 1445
rect 8867 1363 8987 1411
rect 9043 1513 9163 1623
rect 9043 1479 9086 1513
rect 9120 1479 9163 1513
rect 9043 1445 9163 1479
rect 9043 1411 9086 1445
rect 9120 1411 9163 1445
rect 9043 1363 9163 1411
rect 9247 1513 9367 1623
rect 9247 1479 9263 1513
rect 9297 1479 9367 1513
rect 10751 1511 10871 1519
rect 10927 1511 11047 1519
rect 11103 1511 11223 1519
rect 11279 1511 11399 1519
rect 11455 1511 11575 1519
rect 9247 1445 9367 1479
rect 9247 1411 9263 1445
rect 9297 1411 9367 1445
rect 9247 1363 9367 1411
rect 8867 737 8987 763
rect 9043 737 9163 763
rect 9247 737 9367 763
rect 9970 5 10026 71
<< polycont >>
rect 8910 1479 8944 1513
rect 8910 1411 8944 1445
rect 9086 1479 9120 1513
rect 9086 1411 9120 1445
rect 9263 1479 9297 1513
rect 9263 1411 9297 1445
<< locali >>
rect 9903 3477 10032 3691
rect 9903 3443 9904 3477
rect 9938 3443 9976 3477
rect 10010 3443 10032 3477
rect 10158 3477 10286 3691
rect 10192 3443 10230 3477
rect 10264 3443 10286 3477
rect 10459 3289 10497 3323
rect 8808 1805 8842 1813
rect 8808 1737 8842 1741
rect 8808 1669 8842 1703
rect 8808 1619 8842 1635
rect 8998 1805 9032 1821
rect 8998 1737 9032 1771
rect 8998 1669 9032 1703
rect 8998 1585 9032 1635
rect 9188 1805 9222 1813
rect 9188 1737 9222 1741
rect 9188 1669 9222 1703
rect 9188 1619 9222 1635
rect 9378 1805 9412 1821
rect 9378 1737 9412 1771
rect 9378 1669 9412 1703
rect 8808 1551 9313 1585
rect 8659 1339 8765 1363
rect 8659 1305 8692 1339
rect 8726 1305 8765 1339
rect 2562 1267 2603 1301
rect 2637 1267 2678 1301
rect 2712 1267 2753 1301
rect 2787 1267 2828 1301
rect 2862 1267 2903 1301
rect 2937 1267 2978 1301
rect 3012 1267 3053 1301
rect 3087 1267 3128 1301
rect 3162 1267 3203 1301
rect 3237 1267 3278 1301
rect 3312 1267 3354 1301
rect 3388 1267 3430 1301
rect 3464 1267 3506 1301
rect 8659 1265 8765 1305
rect 8659 1231 8692 1265
rect 8726 1231 8765 1265
rect 8659 1191 8765 1231
rect 8659 1157 8692 1191
rect 8726 1157 8765 1191
rect 8659 1117 8765 1157
rect 8659 1083 8692 1117
rect 8726 1083 8765 1117
rect 8659 1043 8765 1083
rect 8659 1009 8692 1043
rect 8726 1009 8765 1043
rect 8659 969 8765 1009
rect 8659 935 8692 969
rect 8726 935 8765 969
rect 8659 895 8765 935
rect 8659 861 8692 895
rect 8726 861 8765 895
rect 8659 821 8765 861
rect 8808 1351 8842 1551
rect 9247 1513 9313 1551
rect 9378 1523 9412 1635
rect 8894 1479 8910 1513
rect 8944 1479 8960 1513
rect 8894 1445 8960 1479
rect 8894 1441 8910 1445
rect 8944 1441 8960 1445
rect 9070 1479 9086 1513
rect 9120 1479 9136 1513
rect 9070 1445 9136 1479
rect 9070 1441 9086 1445
rect 8944 1411 8948 1441
rect 8910 1407 8948 1411
rect 9083 1411 9086 1441
rect 9120 1441 9136 1445
rect 9247 1479 9263 1513
rect 9297 1479 9313 1513
rect 9397 1489 9435 1523
rect 9247 1445 9313 1479
rect 9120 1411 9121 1441
rect 9083 1407 9121 1411
rect 9247 1411 9263 1445
rect 9297 1411 9313 1445
rect 8808 1283 8842 1317
rect 8808 1215 8842 1249
rect 8808 1147 8842 1181
rect 9159 1351 9265 1367
rect 9159 1317 9188 1351
rect 9222 1317 9265 1351
rect 9159 1283 9265 1317
rect 9159 1249 9188 1283
rect 9222 1249 9265 1283
rect 9159 1215 9265 1249
rect 9159 1181 9188 1215
rect 9222 1181 9265 1215
rect 9159 1147 9265 1181
rect 8842 1112 8880 1146
rect 9159 1113 9188 1147
rect 9222 1113 9265 1147
rect 8808 1079 8842 1112
rect 8808 1011 8842 1045
rect 8808 943 8842 977
rect 8808 875 8842 909
rect 8808 825 8842 841
rect 9159 1079 9265 1113
rect 9159 1045 9188 1079
rect 9222 1045 9265 1079
rect 9159 1011 9265 1045
rect 9159 977 9188 1011
rect 9222 977 9265 1011
rect 9159 943 9265 977
rect 9159 909 9188 943
rect 9222 909 9265 943
rect 9159 875 9265 909
rect 9159 841 9188 875
rect 9222 841 9265 875
rect 8659 796 8692 821
rect 8726 796 8765 821
rect 8726 787 8731 796
rect 8693 762 8731 787
rect 9159 821 9265 841
rect 9378 1351 9412 1489
rect 9378 1283 9412 1317
rect 9378 1215 9412 1249
rect 9378 1147 9412 1181
rect 9378 1079 9412 1113
rect 9378 1011 9412 1045
rect 9378 943 9412 977
rect 10086 961 10168 965
rect 10084 927 10122 961
rect 10156 927 10168 961
rect 9378 875 9412 909
rect 9378 825 9412 841
rect 9193 787 9231 821
rect 6259 52 6297 86
rect 10086 55 10168 927
rect 9970 21 10026 55
rect 11351 -92 11385 73
<< viali >>
rect 9904 3443 9938 3477
rect 9976 3443 10010 3477
rect 10158 3443 10192 3477
rect 10230 3443 10264 3477
rect 10425 3289 10459 3323
rect 10497 3289 10531 3323
rect 8808 1813 8842 1847
rect 8808 1771 8842 1775
rect 8808 1741 8842 1771
rect 9188 1813 9222 1847
rect 9188 1771 9222 1775
rect 9188 1741 9222 1771
rect 2528 1267 2562 1301
rect 2603 1267 2637 1301
rect 2678 1267 2712 1301
rect 2753 1267 2787 1301
rect 2828 1267 2862 1301
rect 2903 1267 2937 1301
rect 2978 1267 3012 1301
rect 3053 1267 3087 1301
rect 3128 1267 3162 1301
rect 3203 1267 3237 1301
rect 3278 1267 3312 1301
rect 3354 1267 3388 1301
rect 3430 1267 3464 1301
rect 3506 1267 3540 1301
rect 8876 1407 8910 1441
rect 8948 1407 8982 1441
rect 9049 1407 9083 1441
rect 9363 1489 9397 1523
rect 9435 1489 9469 1523
rect 9121 1407 9155 1441
rect 8808 1113 8842 1146
rect 8808 1112 8842 1113
rect 8880 1112 8914 1146
rect 8659 787 8692 796
rect 8692 787 8693 796
rect 8659 762 8693 787
rect 8731 762 8765 796
rect 10050 927 10084 961
rect 10122 927 10156 961
rect 9159 787 9193 821
rect 9231 787 9265 821
rect 6225 52 6259 86
rect 6297 52 6331 86
<< metal1 >>
rect 0 3511 11256 3657
rect 9584 3477 10276 3483
rect 9636 3443 9904 3477
rect 9938 3443 9976 3477
rect 10010 3443 10158 3477
rect 10192 3443 10230 3477
rect 10264 3443 10276 3477
rect 9636 3437 10276 3443
rect 9584 3413 9636 3425
tri 9636 3412 9661 3437 nw
rect 9584 3355 9636 3361
rect 9829 3283 9835 3335
rect 9887 3283 9899 3335
rect 9951 3323 10697 3335
rect 9951 3289 10425 3323
rect 10459 3289 10497 3323
rect 10531 3289 10697 3323
rect 9951 3283 10697 3289
tri 7324 3093 7386 3155 se
rect 7386 3103 8662 3155
tri 7386 3093 7396 3103 nw
tri 7310 3079 7324 3093 se
rect 7324 3079 7372 3093
tri 7372 3079 7386 3093 nw
rect 6705 3027 6711 3079
rect 6763 3027 6775 3079
rect 6827 3027 7320 3079
tri 7320 3027 7372 3079 nw
rect 11435 3027 11441 3079
rect 11493 3027 11505 3079
rect 11557 3027 11563 3079
rect 0 2919 9580 2999
tri 9580 2919 9660 2999 sw
tri 10631 2919 10711 2999 se
rect 10711 2919 11256 2999
rect 0 2841 11256 2919
rect 0 2797 847 2841
rect 1066 2797 11256 2841
tri 9550 2772 9575 2797 ne
rect 9575 2772 9627 2797
tri 9627 2772 9652 2797 nw
rect 9576 2770 9626 2771
rect 9575 2734 9627 2770
rect 9576 2733 9626 2734
rect 9575 2689 9627 2732
tri 9627 2689 9652 2714 sw
rect 9575 2637 9759 2689
rect 9811 2637 9823 2689
rect 9875 2637 9881 2689
rect 11435 2557 11441 2609
rect 11493 2557 11505 2609
rect 11557 2557 11563 2609
rect 0 2428 9600 2473
tri 9600 2428 9645 2473 sw
tri 9811 2428 9856 2473 se
rect 9856 2428 11256 2473
rect 0 2271 11256 2428
rect 0 1859 11776 1989
tri 8777 1847 8789 1859 ne
rect 8789 1847 9228 1859
tri 8789 1834 8802 1847 ne
rect 8802 1813 8808 1847
rect 8842 1813 9188 1847
rect 9222 1813 9228 1847
tri 9228 1834 9253 1859 nw
rect 8802 1775 9228 1813
rect 8802 1741 8808 1775
rect 8842 1741 9188 1775
rect 9222 1741 9228 1775
rect 8802 1729 9228 1741
rect 9285 1779 9426 1831
rect 9428 1830 9464 1831
rect 9427 1780 9465 1830
rect 9428 1779 9464 1780
rect 9466 1779 9514 1831
rect 9566 1779 9578 1831
rect 9630 1779 9637 1831
tri 9637 1779 9689 1831 sw
rect 9753 1779 9759 1831
rect 9811 1779 9823 1831
rect 9875 1779 9881 1831
rect 6560 1656 6711 1708
rect 6763 1656 6775 1708
rect 6827 1656 7292 1708
tri 9260 1675 9285 1700 se
rect 9285 1675 9337 1779
tri 9337 1754 9362 1779 nw
tri 9615 1754 9640 1779 ne
rect 9640 1754 9689 1779
tri 9640 1705 9689 1754 ne
tri 9689 1711 9757 1779 sw
tri 9804 1754 9829 1779 ne
rect 9829 1754 9881 1779
rect 9830 1752 9880 1753
rect 9830 1715 9880 1716
tri 9826 1711 9829 1714 se
rect 9829 1711 9881 1714
rect 9689 1705 9757 1711
tri 9689 1700 9694 1705 ne
rect 9694 1700 9757 1705
tri 9337 1675 9362 1700 sw
tri 9694 1675 9719 1700 ne
rect 9719 1689 9757 1700
tri 9757 1689 9779 1711 sw
tri 9804 1689 9826 1711 se
rect 9826 1689 9881 1711
rect 9719 1675 9881 1689
rect 6907 1607 7010 1628
tri 7010 1607 7031 1628 sw
rect 8628 1623 8634 1675
rect 8686 1623 8698 1675
rect 8750 1623 9363 1675
rect 9365 1674 9401 1675
rect 9364 1624 9402 1674
rect 9365 1623 9401 1624
rect 9403 1623 9514 1675
rect 9566 1623 9578 1675
rect 9630 1623 9636 1675
tri 9719 1637 9757 1675 ne
rect 9757 1637 9881 1675
tri 9804 1623 9818 1637 ne
rect 9818 1623 9881 1637
tri 9404 1607 9420 1623 ne
rect 9420 1607 9481 1623
rect 6907 1576 7031 1607
tri 6988 1533 7031 1576 ne
tri 7031 1533 7105 1607 sw
tri 9420 1598 9429 1607 ne
rect 9429 1598 9481 1607
tri 9481 1598 9506 1623 nw
tri 9818 1612 9829 1623 ne
rect 9430 1596 9480 1597
rect 9430 1559 9480 1560
tri 9404 1533 9429 1558 se
rect 9429 1533 9481 1558
tri 9481 1533 9506 1558 sw
tri 9804 1533 9829 1558 se
rect 9829 1533 9881 1623
tri 7031 1523 7041 1533 ne
rect 7041 1523 9561 1533
tri 7041 1489 7075 1523 ne
rect 7075 1489 9363 1523
rect 9397 1489 9435 1523
rect 9469 1489 9561 1523
tri 7075 1481 7083 1489 ne
rect 7083 1481 9561 1489
rect 9562 1482 9563 1532
rect 9599 1482 9600 1532
rect 9601 1481 9881 1533
rect 1880 1373 3684 1479
rect 8864 1441 8994 1447
rect 8864 1407 8876 1441
rect 8910 1407 8948 1441
rect 8982 1407 8994 1441
rect 8864 1401 8994 1407
rect 9037 1441 9167 1447
rect 9037 1407 9049 1441
rect 9083 1407 9121 1441
rect 9155 1407 9167 1441
rect 9037 1401 9167 1407
rect 40 1349 3684 1373
rect 40 1243 2367 1349
rect 2516 1258 2522 1310
rect 2574 1258 2588 1310
rect 2640 1258 2654 1310
rect 2706 1301 2720 1310
rect 2772 1301 2786 1310
rect 2838 1301 2853 1310
rect 2905 1301 2920 1310
rect 2972 1301 2987 1310
rect 3039 1301 3054 1310
rect 3106 1307 3112 1310
rect 3106 1301 3552 1307
rect 2712 1267 2720 1301
rect 2972 1267 2978 1301
rect 3039 1267 3053 1301
rect 3106 1267 3128 1301
rect 3162 1267 3203 1301
rect 3237 1267 3278 1301
rect 3312 1267 3354 1301
rect 3388 1267 3430 1301
rect 3464 1267 3506 1301
rect 3540 1267 3552 1301
rect 2706 1258 2720 1267
rect 2772 1258 2786 1267
rect 2838 1258 2853 1267
rect 2905 1258 2920 1267
rect 2972 1258 2987 1267
rect 3039 1258 3054 1267
rect 3106 1261 3552 1267
rect 3106 1258 3112 1261
rect 3726 1243 11776 1373
rect 6835 1170 6904 1211
rect 8479 1180 8667 1215
rect 8479 1170 8480 1180
tri 8480 1170 8490 1180 nw
tri 8479 1169 8480 1170 nw
tri 8554 1146 8560 1152 se
rect 8560 1146 8926 1152
tri 8549 1141 8554 1146 se
rect 8554 1141 8808 1146
tri 7635 1125 7651 1141 se
rect 7651 1125 8808 1141
rect 6256 1073 6262 1125
rect 6314 1073 6326 1125
rect 6378 1112 7255 1125
tri 7255 1112 7268 1125 sw
tri 7622 1112 7635 1125 se
rect 7635 1112 8808 1125
rect 8842 1112 8880 1146
rect 8914 1112 8926 1146
rect 6378 1096 7268 1112
tri 7268 1096 7284 1112 sw
tri 7606 1096 7622 1112 se
rect 7622 1106 8926 1112
rect 7622 1096 8570 1106
rect 6378 1073 7284 1096
tri 7233 1022 7284 1073 ne
tri 7284 1022 7358 1096 sw
tri 7589 1079 7606 1096 se
rect 7606 1089 8570 1096
tri 8570 1089 8587 1106 nw
rect 7606 1079 7651 1089
tri 7651 1079 7661 1089 nw
tri 9188 1079 9195 1086 se
tri 7532 1022 7589 1079 se
rect 7589 1022 7594 1079
tri 7594 1022 7651 1079 nw
tri 9186 1077 9188 1079 se
rect 9188 1077 9195 1079
tri 8587 1027 8637 1077 se
rect 8637 1034 9195 1077
rect 8637 1027 8661 1034
tri 8661 1027 8668 1034 nw
tri 7284 970 7336 1022 ne
rect 7336 970 7542 1022
tri 7542 970 7594 1022 nw
rect 8172 975 8178 1027
rect 8230 975 8242 1027
rect 8294 975 8609 1027
tri 8609 975 8661 1027 nw
rect 8628 876 8634 928
rect 8686 876 8698 928
rect 8750 876 8756 928
rect 9508 921 9514 973
rect 9566 921 9578 973
rect 9630 961 10168 973
rect 9630 927 10050 961
rect 10084 927 10122 961
rect 10156 927 10168 961
rect 9630 921 10168 927
rect 83 843 11776 848
rect 83 791 2667 843
rect 2719 791 2750 843
rect 2802 791 2833 843
rect 2885 791 2917 843
rect 2969 821 11776 843
rect 2969 796 9159 821
rect 2969 791 8659 796
rect 83 775 8659 791
rect 83 723 2667 775
rect 2719 723 2750 775
rect 2802 723 2833 775
rect 2885 723 2917 775
rect 2969 762 8659 775
rect 8693 762 8731 796
rect 8765 787 9159 796
rect 9193 787 9231 821
rect 9265 787 11776 821
rect 8765 762 11776 787
rect 2969 723 11776 762
rect 83 707 11776 723
rect 83 655 2667 707
rect 2719 655 2750 707
rect 2802 655 2833 707
rect 2885 655 2917 707
rect 2969 655 11776 707
rect 83 646 11776 655
rect 8808 493 8844 574
rect 8172 406 8178 458
rect 8230 406 8242 458
rect 8294 406 8300 458
rect 266 120 11776 322
rect 6213 86 6262 92
rect 6314 86 6326 92
rect 6213 52 6225 86
rect 6259 52 6262 86
rect 6213 40 6262 52
rect 6314 40 6326 52
rect 6378 40 6384 92
rect 8567 40 8612 92
<< rmetal1 >>
rect 9575 2771 9627 2772
rect 9575 2770 9576 2771
rect 9626 2770 9627 2771
rect 9575 2733 9576 2734
rect 9626 2733 9627 2734
rect 9575 2732 9627 2733
rect 9426 1830 9428 1831
rect 9464 1830 9466 1831
rect 9426 1780 9427 1830
rect 9465 1780 9466 1830
rect 9426 1779 9428 1780
rect 9464 1779 9466 1780
rect 9829 1753 9881 1754
rect 9829 1752 9830 1753
rect 9880 1752 9881 1753
rect 9829 1715 9830 1716
rect 9880 1715 9881 1716
rect 9829 1714 9881 1715
rect 9363 1674 9365 1675
rect 9401 1674 9403 1675
rect 9363 1624 9364 1674
rect 9402 1624 9403 1674
rect 9363 1623 9365 1624
rect 9401 1623 9403 1624
rect 9429 1597 9481 1598
rect 9429 1596 9430 1597
rect 9480 1596 9481 1597
rect 9429 1559 9430 1560
rect 9480 1559 9481 1560
rect 9429 1558 9481 1559
rect 9561 1532 9563 1533
rect 9561 1482 9562 1532
rect 9561 1481 9563 1482
rect 9599 1532 9601 1533
rect 9600 1482 9601 1532
rect 9599 1481 9601 1482
<< via1 >>
rect 9584 3425 9636 3477
rect 9584 3361 9636 3413
rect 9835 3283 9887 3335
rect 9899 3283 9951 3335
rect 6711 3027 6763 3079
rect 6775 3027 6827 3079
rect 11441 3027 11493 3079
rect 11505 3027 11557 3079
rect 9759 2637 9811 2689
rect 9823 2637 9875 2689
rect 11441 2557 11493 2609
rect 11505 2557 11557 2609
rect 9514 1779 9566 1831
rect 9578 1779 9630 1831
rect 9759 1779 9811 1831
rect 9823 1779 9875 1831
rect 6711 1656 6763 1708
rect 6775 1656 6827 1708
rect 8634 1623 8686 1675
rect 8698 1623 8750 1675
rect 9514 1623 9566 1675
rect 9578 1623 9630 1675
rect 2522 1301 2574 1310
rect 2522 1267 2528 1301
rect 2528 1267 2562 1301
rect 2562 1267 2574 1301
rect 2522 1258 2574 1267
rect 2588 1301 2640 1310
rect 2588 1267 2603 1301
rect 2603 1267 2637 1301
rect 2637 1267 2640 1301
rect 2588 1258 2640 1267
rect 2654 1301 2706 1310
rect 2720 1301 2772 1310
rect 2786 1301 2838 1310
rect 2853 1301 2905 1310
rect 2920 1301 2972 1310
rect 2987 1301 3039 1310
rect 3054 1301 3106 1310
rect 2654 1267 2678 1301
rect 2678 1267 2706 1301
rect 2720 1267 2753 1301
rect 2753 1267 2772 1301
rect 2786 1267 2787 1301
rect 2787 1267 2828 1301
rect 2828 1267 2838 1301
rect 2853 1267 2862 1301
rect 2862 1267 2903 1301
rect 2903 1267 2905 1301
rect 2920 1267 2937 1301
rect 2937 1267 2972 1301
rect 2987 1267 3012 1301
rect 3012 1267 3039 1301
rect 3054 1267 3087 1301
rect 3087 1267 3106 1301
rect 2654 1258 2706 1267
rect 2720 1258 2772 1267
rect 2786 1258 2838 1267
rect 2853 1258 2905 1267
rect 2920 1258 2972 1267
rect 2987 1258 3039 1267
rect 3054 1258 3106 1267
rect 6262 1073 6314 1125
rect 6326 1073 6378 1125
rect 8178 975 8230 1027
rect 8242 975 8294 1027
rect 8634 876 8686 928
rect 8698 876 8750 928
rect 9514 921 9566 973
rect 9578 921 9630 973
rect 2667 791 2719 843
rect 2750 791 2802 843
rect 2833 791 2885 843
rect 2917 791 2969 843
rect 2667 723 2719 775
rect 2750 723 2802 775
rect 2833 723 2885 775
rect 2917 723 2969 775
rect 2667 655 2719 707
rect 2750 655 2802 707
rect 2833 655 2885 707
rect 2917 655 2969 707
rect 8178 406 8230 458
rect 8242 406 8294 458
rect 6262 86 6314 92
rect 6326 86 6378 92
rect 6262 52 6297 86
rect 6297 52 6314 86
rect 6326 52 6331 86
rect 6331 52 6378 86
rect 6262 40 6314 52
rect 6326 40 6378 52
<< metal2 >>
rect 9584 3477 9636 3483
rect 9584 3413 9636 3425
tri 8577 3079 8601 3103 ne
rect 8601 3079 8653 3103
rect 6705 3027 6711 3079
rect 6763 3027 6775 3079
rect 6827 3027 6833 3079
tri 8601 3027 8653 3079 ne
rect 6705 1708 6757 3027
tri 6757 3002 6782 3027 nw
tri 6757 1708 6782 1733 sw
rect 6705 1656 6711 1708
rect 6763 1656 6775 1708
rect 6827 1656 6833 1708
rect 8628 1623 8634 1675
rect 8686 1623 8698 1675
rect 8750 1623 8756 1675
rect 2516 1258 2522 1310
rect 2574 1258 2588 1310
rect 2640 1258 2654 1310
rect 2706 1258 2720 1310
rect 2772 1258 2786 1310
rect 2838 1258 2853 1310
rect 2905 1258 2920 1310
rect 2972 1258 2987 1310
rect 3039 1258 3054 1310
rect 3106 1258 3112 1310
rect 2656 843 2979 1258
rect 2656 791 2667 843
rect 2719 791 2750 843
rect 2802 791 2833 843
rect 2885 791 2917 843
rect 2969 791 2979 843
rect 2656 775 2979 791
rect 2656 723 2667 775
rect 2719 723 2750 775
rect 2802 723 2833 775
rect 2885 723 2917 775
rect 2969 723 2979 775
rect 2656 707 2979 723
rect 2656 655 2667 707
rect 2719 655 2750 707
rect 2802 655 2833 707
rect 2885 655 2917 707
rect 2969 655 2979 707
rect 2656 650 2979 655
rect 6256 1073 6262 1125
rect 6314 1073 6326 1125
rect 6378 1073 6384 1125
rect 6256 92 6327 1073
tri 6327 1048 6352 1073 nw
rect 8172 975 8178 1027
rect 8230 975 8242 1027
rect 8294 975 8300 1027
tri 8208 973 8210 975 ne
rect 8210 973 8300 975
tri 8210 950 8233 973 ne
tri 8208 458 8233 483 se
rect 8233 458 8300 973
rect 8628 928 8692 1623
tri 8692 1598 8717 1623 nw
rect 8796 1006 8848 3027
tri 9559 1831 9584 1856 se
rect 9584 1831 9636 3361
rect 9829 3283 9835 3335
rect 9887 3283 9899 3335
rect 9951 3283 9957 3335
rect 9664 3107 9722 3159
tri 9804 2689 9829 2714 se
rect 9829 2689 9881 3283
tri 9881 3258 9906 3283 nw
rect 9753 2637 9759 2689
rect 9811 2637 9823 2689
rect 9875 2637 9881 2689
tri 9804 2612 9829 2637 ne
tri 9804 1831 9829 1856 se
rect 9829 1831 9881 2637
rect 9508 1779 9514 1831
rect 9566 1779 9578 1831
rect 9630 1779 9636 1831
rect 9753 1779 9759 1831
rect 9811 1779 9823 1831
rect 9875 1779 9881 1831
rect 11435 3027 11441 3079
rect 11493 3027 11505 3079
rect 11557 3027 11563 3079
rect 11435 2609 11563 3027
rect 11435 2557 11441 2609
rect 11493 2557 11505 2609
rect 11557 2557 11563 2609
rect 9508 1623 9514 1675
rect 9566 1623 9578 1675
rect 9630 1623 9636 1675
rect 9195 1034 9242 1086
rect 9508 973 9636 1623
tri 8692 928 8717 953 sw
rect 8628 876 8634 928
rect 8686 876 8698 928
rect 8750 876 8756 928
rect 9508 921 9514 973
rect 9566 921 9578 973
rect 9630 921 9636 973
rect 8172 406 8178 458
rect 8230 406 8242 458
rect 8294 406 8300 458
tri 6327 92 6352 117 sw
rect 6256 40 6262 92
rect 6314 40 6326 92
rect 6378 40 6384 92
rect 11435 40 11563 2557
use sky130_fd_io__gpio_ovtv2_pdpredrvr_pbias  sky130_fd_io__gpio_ovtv2_pdpredrvr_pbias_0
timestamp 1704896540
transform -1 0 20068 0 1 -2980
box 7295 2861 20071 6839
use sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_nr2  sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_nr2_0
timestamp 1704896540
transform -1 0 11035 0 -1 1911
box -727 369 2877 1910
use sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_nr3  sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_nr3_0
timestamp 1704896540
transform -1 0 11256 0 1 1909
box -827 -420 4208 1950
use sky130_fd_io__tk_em1o_cdns_5595914180880  sky130_fd_io__tk_em1o_cdns_5595914180880_0
timestamp 1704896540
transform 0 1 9429 1 0 1506
box 0 0 1 1
use sky130_fd_io__tk_em1o_cdns_5595914180880  sky130_fd_io__tk_em1o_cdns_5595914180880_1
timestamp 1704896540
transform 0 1 9829 -1 0 1806
box 0 0 1 1
use sky130_fd_io__tk_em1o_cdns_5595914180880  sky130_fd_io__tk_em1o_cdns_5595914180880_2
timestamp 1704896540
transform 1 0 9509 0 1 1481
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_5595914180882  sky130_fd_io__tk_em1s_cdns_5595914180882_0
timestamp 1704896540
transform -1 0 9455 0 -1 1675
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_5595914180882  sky130_fd_io__tk_em1s_cdns_5595914180882_1
timestamp 1704896540
transform 0 -1 9627 1 0 2680
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_5595914180882  sky130_fd_io__tk_em1s_cdns_5595914180882_2
timestamp 1704896540
transform -1 0 9518 0 1 1779
box 0 0 1 1
use sky130_fd_pr__model__nfet_highvoltage__example_55959141808139  sky130_fd_pr__model__nfet_highvoltage__example_55959141808139_0
timestamp 1704896540
transform 1 0 8867 0 1 1623
box -15 0 311 1
use sky130_fd_pr__model__nfet_highvoltage__example_55959141808183  sky130_fd_pr__model__nfet_highvoltage__example_55959141808183_0
timestamp 1704896540
transform 1 0 9247 0 1 1623
box -15 0 121 1
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808141  sky130_fd_pr__model__pfet_highvoltage__example_55959141808141_0
timestamp 1704896540
transform 1 0 8867 0 -1 1363
box -15 0 -14 1
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808141  sky130_fd_pr__model__pfet_highvoltage__example_55959141808141_1
timestamp 1704896540
transform -1 0 9163 0 -1 1363
box -15 0 -14 1
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808184  sky130_fd_pr__model__pfet_highvoltage__example_55959141808184_0
timestamp 1704896540
transform 1 0 9247 0 -1 1363
box -15 0 121 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1704896540
transform 1 0 10158 0 1 3443
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_1
timestamp 1704896540
transform 1 0 9904 0 1 3443
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_2
timestamp 1704896540
transform 1 0 10425 0 1 3289
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_3
timestamp 1704896540
transform 1 0 9159 0 -1 821
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_4
timestamp 1704896540
transform 1 0 9049 0 -1 1441
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_5
timestamp 1704896540
transform 1 0 8876 0 -1 1441
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_6
timestamp 1704896540
transform 0 1 9188 1 0 1741
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_7
timestamp 1704896540
transform 0 1 8808 1 0 1741
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_8
timestamp 1704896540
transform 1 0 8808 0 -1 1146
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_9
timestamp 1704896540
transform 1 0 6225 0 1 52
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_10
timestamp 1704896540
transform 1 0 9363 0 -1 1523
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_11
timestamp 1704896540
transform 1 0 8659 0 -1 796
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_12
timestamp 1704896540
transform -1 0 10156 0 1 927
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_0
timestamp 1704896540
transform 1 0 9508 0 1 1779
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_1
timestamp 1704896540
transform 0 -1 9636 -1 0 3483
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_2
timestamp 1704896540
transform 1 0 9829 0 1 3283
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_3
timestamp 1704896540
transform -1 0 9881 0 1 2637
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_4
timestamp 1704896540
transform -1 0 9881 0 1 1779
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_5
timestamp 1704896540
transform 1 0 8172 0 1 975
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_6
timestamp 1704896540
transform 1 0 6256 0 1 40
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_7
timestamp 1704896540
transform 1 0 6256 0 1 1073
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_8
timestamp 1704896540
transform 1 0 8172 0 1 406
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_9
timestamp 1704896540
transform 1 0 8628 0 1 876
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_10
timestamp 1704896540
transform 1 0 8628 0 1 1623
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_11
timestamp 1704896540
transform 1 0 9508 0 1 921
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_12
timestamp 1704896540
transform 1 0 9508 0 1 1623
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_13
timestamp 1704896540
transform 1 0 6705 0 1 3027
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_14
timestamp 1704896540
transform 1 0 6705 0 1 1656
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_0
timestamp 1704896540
transform 0 1 8894 1 0 1395
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_1
timestamp 1704896540
transform 0 1 9070 1 0 1395
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_2
timestamp 1704896540
transform 0 1 9247 1 0 1395
box 0 0 1 1
<< labels >>
flabel metal2 s 9195 1034 9242 1086 3 FreeSans 300 180 0 0 PD_H[2]
port 1 nsew
flabel metal2 s 9664 3107 9722 3159 7 FreeSans 300 180 0 0 PD_H[3]
port 2 nsew
flabel metal1 s 8879 1401 8927 1447 3 FreeSans 200 90 0 0 EN_CMOS_B
port 4 nsew
flabel metal1 s 11216 2271 11256 2473 7 FreeSans 300 180 0 0 VGND_IO
port 5 nsew
flabel metal1 s 11216 2797 11256 2999 7 FreeSans 300 180 0 0 VCC_IO
port 6 nsew
flabel metal1 s 11216 3511 11256 3657 7 FreeSans 300 180 0 0 VCC_IO
port 6 nsew
flabel metal1 s 11235 2372 11235 2372 7 FreeSans 300 180 0 0 VGND_IO
flabel metal1 s 11736 646 11776 848 7 FreeSans 300 180 0 0 VCC_IO
port 6 nsew
flabel metal1 s 11736 120 11776 322 7 FreeSans 300 180 0 0 VGND_IO
port 5 nsew
flabel metal1 s 11736 1243 11776 1373 7 FreeSans 300 180 0 0 VGND_IO
port 5 nsew
flabel metal1 s 11216 1859 11256 1989 7 FreeSans 300 180 0 0 VGND_IO
port 5 nsew
flabel metal1 s 8567 40 8612 92 8 FreeSans 300 180 0 0 DRVLO_H_N
port 7 nsew
flabel metal1 s 9121 1401 9167 1447 7 FreeSans 300 180 0 0 SLOW_H
port 8 nsew
flabel metal1 s 0 2271 40 2473 3 FreeSans 300 180 0 0 VGND_IO
port 5 nsew
flabel metal1 s 0 1859 40 1989 3 FreeSans 300 180 0 0 VGND_IO
port 5 nsew
flabel metal1 s 43 1243 83 1373 3 FreeSans 300 180 0 0 VGND_IO
port 5 nsew
flabel metal1 s 83 646 123 848 3 FreeSans 300 180 0 0 VCC_IO
port 6 nsew
flabel metal1 s 276 120 316 322 3 FreeSans 300 180 0 0 VGND_IO
port 5 nsew
flabel metal1 s 0 2797 40 2999 3 FreeSans 300 180 0 0 VCC_IO
port 6 nsew
flabel metal1 s 0 3511 40 3657 7 FreeSans 300 180 0 0 VCC_IO
port 6 nsew
flabel metal1 s 6835 1170 6904 1211 3 FreeSans 520 0 0 0 DRVHI_H
port 9 nsew
flabel metal1 s 8808 493 8844 574 3 FreeSans 520 0 0 0 NSW_EN
port 10 nsew
flabel metal1 s 6560 1656 6593 1702 3 FreeSans 240 0 0 0 PDEN_H_N
port 11 nsew
flabel comment s 8277 742 8277 742 0 FreeSans 300 0 0 0 VCC_IO
flabel comment s 8253 210 8253 210 0 FreeSans 300 0 0 0 VGND_IO
flabel comment s 7705 3061 7705 3061 0 FreeSans 300 0 0 0 PDEN_H_N
flabel comment s 8813 3706 8813 3706 0 FreeSans 300 90 0 0 PDEN_H_N
flabel comment s 8812 2082 8812 2082 0 FreeSans 300 90 0 0 PDEN_H_N
flabel comment s 8698 1667 8698 1667 0 FreeSans 300 0 0 0 PBIAS
flabel comment s 6897 1611 6897 1611 0 FreeSans 300 0 0 0 EN_FAST_H_N
flabel comment s 9463 1511 9463 1511 0 FreeSans 300 0 0 0 EN_FAST_H_N
flabel comment s 8310 1126 8310 1126 0 FreeSans 300 0 0 0 EN_FAST_H
flabel comment s 6333 1097 6333 1097 0 FreeSans 300 0 0 0 EN_FAST_H
flabel comment s 9956 1467 9956 1467 0 FreeSans 300 0 0 0 PBIAS
flabel comment s 9841 2135 9841 2135 0 FreeSans 300 90 0 0 EN_FAST2_N0
flabel comment s 9565 1662 9565 1662 0 FreeSans 300 0 0 0 EN_FAST_N1
flabel comment s 9546 2130 9546 2130 0 FreeSans 300 90 0 0 EN_FAST2_N1
<< properties >>
string GDS_END 67930392
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 67912300
<< end >>
