magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< dnwell >>
rect 1846 1716 94204 77780
<< nwell >>
rect 1762 77696 94288 77864
rect 1762 1800 1930 77696
rect 94120 1800 94288 77696
rect 1762 1632 94288 1800
<< nsubdiff >>
rect 2157 77797 2207 77821
rect 2157 77763 2165 77797
rect 2199 77763 2207 77797
rect 2157 77739 2207 77763
rect 2493 77797 2543 77821
rect 2493 77763 2501 77797
rect 2535 77763 2543 77797
rect 2493 77739 2543 77763
rect 2829 77797 2879 77821
rect 2829 77763 2837 77797
rect 2871 77763 2879 77797
rect 2829 77739 2879 77763
rect 3165 77797 3215 77821
rect 3165 77763 3173 77797
rect 3207 77763 3215 77797
rect 3165 77739 3215 77763
rect 3501 77797 3551 77821
rect 3501 77763 3509 77797
rect 3543 77763 3551 77797
rect 3501 77739 3551 77763
rect 3837 77797 3887 77821
rect 3837 77763 3845 77797
rect 3879 77763 3887 77797
rect 3837 77739 3887 77763
rect 4173 77797 4223 77821
rect 4173 77763 4181 77797
rect 4215 77763 4223 77797
rect 4173 77739 4223 77763
rect 4509 77797 4559 77821
rect 4509 77763 4517 77797
rect 4551 77763 4559 77797
rect 4509 77739 4559 77763
rect 4845 77797 4895 77821
rect 4845 77763 4853 77797
rect 4887 77763 4895 77797
rect 4845 77739 4895 77763
rect 5181 77797 5231 77821
rect 5181 77763 5189 77797
rect 5223 77763 5231 77797
rect 5181 77739 5231 77763
rect 5517 77797 5567 77821
rect 5517 77763 5525 77797
rect 5559 77763 5567 77797
rect 5517 77739 5567 77763
rect 5853 77797 5903 77821
rect 5853 77763 5861 77797
rect 5895 77763 5903 77797
rect 5853 77739 5903 77763
rect 6189 77797 6239 77821
rect 6189 77763 6197 77797
rect 6231 77763 6239 77797
rect 6189 77739 6239 77763
rect 6525 77797 6575 77821
rect 6525 77763 6533 77797
rect 6567 77763 6575 77797
rect 6525 77739 6575 77763
rect 6861 77797 6911 77821
rect 6861 77763 6869 77797
rect 6903 77763 6911 77797
rect 6861 77739 6911 77763
rect 7197 77797 7247 77821
rect 7197 77763 7205 77797
rect 7239 77763 7247 77797
rect 7197 77739 7247 77763
rect 7533 77797 7583 77821
rect 7533 77763 7541 77797
rect 7575 77763 7583 77797
rect 7533 77739 7583 77763
rect 7869 77797 7919 77821
rect 7869 77763 7877 77797
rect 7911 77763 7919 77797
rect 7869 77739 7919 77763
rect 8205 77797 8255 77821
rect 8205 77763 8213 77797
rect 8247 77763 8255 77797
rect 8205 77739 8255 77763
rect 8541 77797 8591 77821
rect 8541 77763 8549 77797
rect 8583 77763 8591 77797
rect 8541 77739 8591 77763
rect 8877 77797 8927 77821
rect 8877 77763 8885 77797
rect 8919 77763 8927 77797
rect 8877 77739 8927 77763
rect 9213 77797 9263 77821
rect 9213 77763 9221 77797
rect 9255 77763 9263 77797
rect 9213 77739 9263 77763
rect 9549 77797 9599 77821
rect 9549 77763 9557 77797
rect 9591 77763 9599 77797
rect 9549 77739 9599 77763
rect 9885 77797 9935 77821
rect 9885 77763 9893 77797
rect 9927 77763 9935 77797
rect 9885 77739 9935 77763
rect 10221 77797 10271 77821
rect 10221 77763 10229 77797
rect 10263 77763 10271 77797
rect 10221 77739 10271 77763
rect 10557 77797 10607 77821
rect 10557 77763 10565 77797
rect 10599 77763 10607 77797
rect 10557 77739 10607 77763
rect 10893 77797 10943 77821
rect 10893 77763 10901 77797
rect 10935 77763 10943 77797
rect 10893 77739 10943 77763
rect 11229 77797 11279 77821
rect 11229 77763 11237 77797
rect 11271 77763 11279 77797
rect 11229 77739 11279 77763
rect 11565 77797 11615 77821
rect 11565 77763 11573 77797
rect 11607 77763 11615 77797
rect 11565 77739 11615 77763
rect 11901 77797 11951 77821
rect 11901 77763 11909 77797
rect 11943 77763 11951 77797
rect 11901 77739 11951 77763
rect 12237 77797 12287 77821
rect 12237 77763 12245 77797
rect 12279 77763 12287 77797
rect 12237 77739 12287 77763
rect 12573 77797 12623 77821
rect 12573 77763 12581 77797
rect 12615 77763 12623 77797
rect 12573 77739 12623 77763
rect 12909 77797 12959 77821
rect 12909 77763 12917 77797
rect 12951 77763 12959 77797
rect 12909 77739 12959 77763
rect 13245 77797 13295 77821
rect 13245 77763 13253 77797
rect 13287 77763 13295 77797
rect 13245 77739 13295 77763
rect 13581 77797 13631 77821
rect 13581 77763 13589 77797
rect 13623 77763 13631 77797
rect 13581 77739 13631 77763
rect 13917 77797 13967 77821
rect 13917 77763 13925 77797
rect 13959 77763 13967 77797
rect 13917 77739 13967 77763
rect 14253 77797 14303 77821
rect 14253 77763 14261 77797
rect 14295 77763 14303 77797
rect 14253 77739 14303 77763
rect 14589 77797 14639 77821
rect 14589 77763 14597 77797
rect 14631 77763 14639 77797
rect 14589 77739 14639 77763
rect 14925 77797 14975 77821
rect 14925 77763 14933 77797
rect 14967 77763 14975 77797
rect 14925 77739 14975 77763
rect 15261 77797 15311 77821
rect 15261 77763 15269 77797
rect 15303 77763 15311 77797
rect 15261 77739 15311 77763
rect 15597 77797 15647 77821
rect 15597 77763 15605 77797
rect 15639 77763 15647 77797
rect 15597 77739 15647 77763
rect 15933 77797 15983 77821
rect 15933 77763 15941 77797
rect 15975 77763 15983 77797
rect 15933 77739 15983 77763
rect 16269 77797 16319 77821
rect 16269 77763 16277 77797
rect 16311 77763 16319 77797
rect 16269 77739 16319 77763
rect 16605 77797 16655 77821
rect 16605 77763 16613 77797
rect 16647 77763 16655 77797
rect 16605 77739 16655 77763
rect 16941 77797 16991 77821
rect 16941 77763 16949 77797
rect 16983 77763 16991 77797
rect 16941 77739 16991 77763
rect 17277 77797 17327 77821
rect 17277 77763 17285 77797
rect 17319 77763 17327 77797
rect 17277 77739 17327 77763
rect 17613 77797 17663 77821
rect 17613 77763 17621 77797
rect 17655 77763 17663 77797
rect 17613 77739 17663 77763
rect 17949 77797 17999 77821
rect 17949 77763 17957 77797
rect 17991 77763 17999 77797
rect 17949 77739 17999 77763
rect 18285 77797 18335 77821
rect 18285 77763 18293 77797
rect 18327 77763 18335 77797
rect 18285 77739 18335 77763
rect 18621 77797 18671 77821
rect 18621 77763 18629 77797
rect 18663 77763 18671 77797
rect 18621 77739 18671 77763
rect 18957 77797 19007 77821
rect 18957 77763 18965 77797
rect 18999 77763 19007 77797
rect 18957 77739 19007 77763
rect 19293 77797 19343 77821
rect 19293 77763 19301 77797
rect 19335 77763 19343 77797
rect 19293 77739 19343 77763
rect 19629 77797 19679 77821
rect 19629 77763 19637 77797
rect 19671 77763 19679 77797
rect 19629 77739 19679 77763
rect 19965 77797 20015 77821
rect 19965 77763 19973 77797
rect 20007 77763 20015 77797
rect 19965 77739 20015 77763
rect 20301 77797 20351 77821
rect 20301 77763 20309 77797
rect 20343 77763 20351 77797
rect 20301 77739 20351 77763
rect 20637 77797 20687 77821
rect 20637 77763 20645 77797
rect 20679 77763 20687 77797
rect 20637 77739 20687 77763
rect 20973 77797 21023 77821
rect 20973 77763 20981 77797
rect 21015 77763 21023 77797
rect 20973 77739 21023 77763
rect 21309 77797 21359 77821
rect 21309 77763 21317 77797
rect 21351 77763 21359 77797
rect 21309 77739 21359 77763
rect 21645 77797 21695 77821
rect 21645 77763 21653 77797
rect 21687 77763 21695 77797
rect 21645 77739 21695 77763
rect 21981 77797 22031 77821
rect 21981 77763 21989 77797
rect 22023 77763 22031 77797
rect 21981 77739 22031 77763
rect 22317 77797 22367 77821
rect 22317 77763 22325 77797
rect 22359 77763 22367 77797
rect 22317 77739 22367 77763
rect 22653 77797 22703 77821
rect 22653 77763 22661 77797
rect 22695 77763 22703 77797
rect 22653 77739 22703 77763
rect 22989 77797 23039 77821
rect 22989 77763 22997 77797
rect 23031 77763 23039 77797
rect 22989 77739 23039 77763
rect 23325 77797 23375 77821
rect 23325 77763 23333 77797
rect 23367 77763 23375 77797
rect 23325 77739 23375 77763
rect 23661 77797 23711 77821
rect 23661 77763 23669 77797
rect 23703 77763 23711 77797
rect 23661 77739 23711 77763
rect 23997 77797 24047 77821
rect 23997 77763 24005 77797
rect 24039 77763 24047 77797
rect 23997 77739 24047 77763
rect 24333 77797 24383 77821
rect 24333 77763 24341 77797
rect 24375 77763 24383 77797
rect 24333 77739 24383 77763
rect 24669 77797 24719 77821
rect 24669 77763 24677 77797
rect 24711 77763 24719 77797
rect 24669 77739 24719 77763
rect 25005 77797 25055 77821
rect 25005 77763 25013 77797
rect 25047 77763 25055 77797
rect 25005 77739 25055 77763
rect 25341 77797 25391 77821
rect 25341 77763 25349 77797
rect 25383 77763 25391 77797
rect 25341 77739 25391 77763
rect 25677 77797 25727 77821
rect 25677 77763 25685 77797
rect 25719 77763 25727 77797
rect 25677 77739 25727 77763
rect 26013 77797 26063 77821
rect 26013 77763 26021 77797
rect 26055 77763 26063 77797
rect 26013 77739 26063 77763
rect 26349 77797 26399 77821
rect 26349 77763 26357 77797
rect 26391 77763 26399 77797
rect 26349 77739 26399 77763
rect 26685 77797 26735 77821
rect 26685 77763 26693 77797
rect 26727 77763 26735 77797
rect 26685 77739 26735 77763
rect 27021 77797 27071 77821
rect 27021 77763 27029 77797
rect 27063 77763 27071 77797
rect 27021 77739 27071 77763
rect 27357 77797 27407 77821
rect 27357 77763 27365 77797
rect 27399 77763 27407 77797
rect 27357 77739 27407 77763
rect 27693 77797 27743 77821
rect 27693 77763 27701 77797
rect 27735 77763 27743 77797
rect 27693 77739 27743 77763
rect 28029 77797 28079 77821
rect 28029 77763 28037 77797
rect 28071 77763 28079 77797
rect 28029 77739 28079 77763
rect 28365 77797 28415 77821
rect 28365 77763 28373 77797
rect 28407 77763 28415 77797
rect 28365 77739 28415 77763
rect 28701 77797 28751 77821
rect 28701 77763 28709 77797
rect 28743 77763 28751 77797
rect 28701 77739 28751 77763
rect 29037 77797 29087 77821
rect 29037 77763 29045 77797
rect 29079 77763 29087 77797
rect 29037 77739 29087 77763
rect 29373 77797 29423 77821
rect 29373 77763 29381 77797
rect 29415 77763 29423 77797
rect 29373 77739 29423 77763
rect 29709 77797 29759 77821
rect 29709 77763 29717 77797
rect 29751 77763 29759 77797
rect 29709 77739 29759 77763
rect 30045 77797 30095 77821
rect 30045 77763 30053 77797
rect 30087 77763 30095 77797
rect 30045 77739 30095 77763
rect 30381 77797 30431 77821
rect 30381 77763 30389 77797
rect 30423 77763 30431 77797
rect 30381 77739 30431 77763
rect 30717 77797 30767 77821
rect 30717 77763 30725 77797
rect 30759 77763 30767 77797
rect 30717 77739 30767 77763
rect 31053 77797 31103 77821
rect 31053 77763 31061 77797
rect 31095 77763 31103 77797
rect 31053 77739 31103 77763
rect 31389 77797 31439 77821
rect 31389 77763 31397 77797
rect 31431 77763 31439 77797
rect 31389 77739 31439 77763
rect 31725 77797 31775 77821
rect 31725 77763 31733 77797
rect 31767 77763 31775 77797
rect 31725 77739 31775 77763
rect 32061 77797 32111 77821
rect 32061 77763 32069 77797
rect 32103 77763 32111 77797
rect 32061 77739 32111 77763
rect 32397 77797 32447 77821
rect 32397 77763 32405 77797
rect 32439 77763 32447 77797
rect 32397 77739 32447 77763
rect 32733 77797 32783 77821
rect 32733 77763 32741 77797
rect 32775 77763 32783 77797
rect 32733 77739 32783 77763
rect 33069 77797 33119 77821
rect 33069 77763 33077 77797
rect 33111 77763 33119 77797
rect 33069 77739 33119 77763
rect 33405 77797 33455 77821
rect 33405 77763 33413 77797
rect 33447 77763 33455 77797
rect 33405 77739 33455 77763
rect 33741 77797 33791 77821
rect 33741 77763 33749 77797
rect 33783 77763 33791 77797
rect 33741 77739 33791 77763
rect 34077 77797 34127 77821
rect 34077 77763 34085 77797
rect 34119 77763 34127 77797
rect 34077 77739 34127 77763
rect 34413 77797 34463 77821
rect 34413 77763 34421 77797
rect 34455 77763 34463 77797
rect 34413 77739 34463 77763
rect 34749 77797 34799 77821
rect 34749 77763 34757 77797
rect 34791 77763 34799 77797
rect 34749 77739 34799 77763
rect 35085 77797 35135 77821
rect 35085 77763 35093 77797
rect 35127 77763 35135 77797
rect 35085 77739 35135 77763
rect 35421 77797 35471 77821
rect 35421 77763 35429 77797
rect 35463 77763 35471 77797
rect 35421 77739 35471 77763
rect 35757 77797 35807 77821
rect 35757 77763 35765 77797
rect 35799 77763 35807 77797
rect 35757 77739 35807 77763
rect 36093 77797 36143 77821
rect 36093 77763 36101 77797
rect 36135 77763 36143 77797
rect 36093 77739 36143 77763
rect 36429 77797 36479 77821
rect 36429 77763 36437 77797
rect 36471 77763 36479 77797
rect 36429 77739 36479 77763
rect 36765 77797 36815 77821
rect 36765 77763 36773 77797
rect 36807 77763 36815 77797
rect 36765 77739 36815 77763
rect 37101 77797 37151 77821
rect 37101 77763 37109 77797
rect 37143 77763 37151 77797
rect 37101 77739 37151 77763
rect 37437 77797 37487 77821
rect 37437 77763 37445 77797
rect 37479 77763 37487 77797
rect 37437 77739 37487 77763
rect 37773 77797 37823 77821
rect 37773 77763 37781 77797
rect 37815 77763 37823 77797
rect 37773 77739 37823 77763
rect 38109 77797 38159 77821
rect 38109 77763 38117 77797
rect 38151 77763 38159 77797
rect 38109 77739 38159 77763
rect 38445 77797 38495 77821
rect 38445 77763 38453 77797
rect 38487 77763 38495 77797
rect 38445 77739 38495 77763
rect 38781 77797 38831 77821
rect 38781 77763 38789 77797
rect 38823 77763 38831 77797
rect 38781 77739 38831 77763
rect 39117 77797 39167 77821
rect 39117 77763 39125 77797
rect 39159 77763 39167 77797
rect 39117 77739 39167 77763
rect 39453 77797 39503 77821
rect 39453 77763 39461 77797
rect 39495 77763 39503 77797
rect 39453 77739 39503 77763
rect 39789 77797 39839 77821
rect 39789 77763 39797 77797
rect 39831 77763 39839 77797
rect 39789 77739 39839 77763
rect 40125 77797 40175 77821
rect 40125 77763 40133 77797
rect 40167 77763 40175 77797
rect 40125 77739 40175 77763
rect 40461 77797 40511 77821
rect 40461 77763 40469 77797
rect 40503 77763 40511 77797
rect 40461 77739 40511 77763
rect 40797 77797 40847 77821
rect 40797 77763 40805 77797
rect 40839 77763 40847 77797
rect 40797 77739 40847 77763
rect 41133 77797 41183 77821
rect 41133 77763 41141 77797
rect 41175 77763 41183 77797
rect 41133 77739 41183 77763
rect 41469 77797 41519 77821
rect 41469 77763 41477 77797
rect 41511 77763 41519 77797
rect 41469 77739 41519 77763
rect 41805 77797 41855 77821
rect 41805 77763 41813 77797
rect 41847 77763 41855 77797
rect 41805 77739 41855 77763
rect 42141 77797 42191 77821
rect 42141 77763 42149 77797
rect 42183 77763 42191 77797
rect 42141 77739 42191 77763
rect 42477 77797 42527 77821
rect 42477 77763 42485 77797
rect 42519 77763 42527 77797
rect 42477 77739 42527 77763
rect 42813 77797 42863 77821
rect 42813 77763 42821 77797
rect 42855 77763 42863 77797
rect 42813 77739 42863 77763
rect 43149 77797 43199 77821
rect 43149 77763 43157 77797
rect 43191 77763 43199 77797
rect 43149 77739 43199 77763
rect 43485 77797 43535 77821
rect 43485 77763 43493 77797
rect 43527 77763 43535 77797
rect 43485 77739 43535 77763
rect 43821 77797 43871 77821
rect 43821 77763 43829 77797
rect 43863 77763 43871 77797
rect 43821 77739 43871 77763
rect 44157 77797 44207 77821
rect 44157 77763 44165 77797
rect 44199 77763 44207 77797
rect 44157 77739 44207 77763
rect 44493 77797 44543 77821
rect 44493 77763 44501 77797
rect 44535 77763 44543 77797
rect 44493 77739 44543 77763
rect 44829 77797 44879 77821
rect 44829 77763 44837 77797
rect 44871 77763 44879 77797
rect 44829 77739 44879 77763
rect 45165 77797 45215 77821
rect 45165 77763 45173 77797
rect 45207 77763 45215 77797
rect 45165 77739 45215 77763
rect 45501 77797 45551 77821
rect 45501 77763 45509 77797
rect 45543 77763 45551 77797
rect 45501 77739 45551 77763
rect 45837 77797 45887 77821
rect 45837 77763 45845 77797
rect 45879 77763 45887 77797
rect 45837 77739 45887 77763
rect 46173 77797 46223 77821
rect 46173 77763 46181 77797
rect 46215 77763 46223 77797
rect 46173 77739 46223 77763
rect 46509 77797 46559 77821
rect 46509 77763 46517 77797
rect 46551 77763 46559 77797
rect 46509 77739 46559 77763
rect 46845 77797 46895 77821
rect 46845 77763 46853 77797
rect 46887 77763 46895 77797
rect 46845 77739 46895 77763
rect 47181 77797 47231 77821
rect 47181 77763 47189 77797
rect 47223 77763 47231 77797
rect 47181 77739 47231 77763
rect 47517 77797 47567 77821
rect 47517 77763 47525 77797
rect 47559 77763 47567 77797
rect 47517 77739 47567 77763
rect 47853 77797 47903 77821
rect 47853 77763 47861 77797
rect 47895 77763 47903 77797
rect 47853 77739 47903 77763
rect 48189 77797 48239 77821
rect 48189 77763 48197 77797
rect 48231 77763 48239 77797
rect 48189 77739 48239 77763
rect 48525 77797 48575 77821
rect 48525 77763 48533 77797
rect 48567 77763 48575 77797
rect 48525 77739 48575 77763
rect 48861 77797 48911 77821
rect 48861 77763 48869 77797
rect 48903 77763 48911 77797
rect 48861 77739 48911 77763
rect 49197 77797 49247 77821
rect 49197 77763 49205 77797
rect 49239 77763 49247 77797
rect 49197 77739 49247 77763
rect 49533 77797 49583 77821
rect 49533 77763 49541 77797
rect 49575 77763 49583 77797
rect 49533 77739 49583 77763
rect 49869 77797 49919 77821
rect 49869 77763 49877 77797
rect 49911 77763 49919 77797
rect 49869 77739 49919 77763
rect 50205 77797 50255 77821
rect 50205 77763 50213 77797
rect 50247 77763 50255 77797
rect 50205 77739 50255 77763
rect 50541 77797 50591 77821
rect 50541 77763 50549 77797
rect 50583 77763 50591 77797
rect 50541 77739 50591 77763
rect 50877 77797 50927 77821
rect 50877 77763 50885 77797
rect 50919 77763 50927 77797
rect 50877 77739 50927 77763
rect 51213 77797 51263 77821
rect 51213 77763 51221 77797
rect 51255 77763 51263 77797
rect 51213 77739 51263 77763
rect 51549 77797 51599 77821
rect 51549 77763 51557 77797
rect 51591 77763 51599 77797
rect 51549 77739 51599 77763
rect 51885 77797 51935 77821
rect 51885 77763 51893 77797
rect 51927 77763 51935 77797
rect 51885 77739 51935 77763
rect 52221 77797 52271 77821
rect 52221 77763 52229 77797
rect 52263 77763 52271 77797
rect 52221 77739 52271 77763
rect 52557 77797 52607 77821
rect 52557 77763 52565 77797
rect 52599 77763 52607 77797
rect 52557 77739 52607 77763
rect 52893 77797 52943 77821
rect 52893 77763 52901 77797
rect 52935 77763 52943 77797
rect 52893 77739 52943 77763
rect 53229 77797 53279 77821
rect 53229 77763 53237 77797
rect 53271 77763 53279 77797
rect 53229 77739 53279 77763
rect 53565 77797 53615 77821
rect 53565 77763 53573 77797
rect 53607 77763 53615 77797
rect 53565 77739 53615 77763
rect 53901 77797 53951 77821
rect 53901 77763 53909 77797
rect 53943 77763 53951 77797
rect 53901 77739 53951 77763
rect 54237 77797 54287 77821
rect 54237 77763 54245 77797
rect 54279 77763 54287 77797
rect 54237 77739 54287 77763
rect 54573 77797 54623 77821
rect 54573 77763 54581 77797
rect 54615 77763 54623 77797
rect 54573 77739 54623 77763
rect 54909 77797 54959 77821
rect 54909 77763 54917 77797
rect 54951 77763 54959 77797
rect 54909 77739 54959 77763
rect 55245 77797 55295 77821
rect 55245 77763 55253 77797
rect 55287 77763 55295 77797
rect 55245 77739 55295 77763
rect 55581 77797 55631 77821
rect 55581 77763 55589 77797
rect 55623 77763 55631 77797
rect 55581 77739 55631 77763
rect 55917 77797 55967 77821
rect 55917 77763 55925 77797
rect 55959 77763 55967 77797
rect 55917 77739 55967 77763
rect 56253 77797 56303 77821
rect 56253 77763 56261 77797
rect 56295 77763 56303 77797
rect 56253 77739 56303 77763
rect 56589 77797 56639 77821
rect 56589 77763 56597 77797
rect 56631 77763 56639 77797
rect 56589 77739 56639 77763
rect 56925 77797 56975 77821
rect 56925 77763 56933 77797
rect 56967 77763 56975 77797
rect 56925 77739 56975 77763
rect 57261 77797 57311 77821
rect 57261 77763 57269 77797
rect 57303 77763 57311 77797
rect 57261 77739 57311 77763
rect 57597 77797 57647 77821
rect 57597 77763 57605 77797
rect 57639 77763 57647 77797
rect 57597 77739 57647 77763
rect 57933 77797 57983 77821
rect 57933 77763 57941 77797
rect 57975 77763 57983 77797
rect 57933 77739 57983 77763
rect 58269 77797 58319 77821
rect 58269 77763 58277 77797
rect 58311 77763 58319 77797
rect 58269 77739 58319 77763
rect 58605 77797 58655 77821
rect 58605 77763 58613 77797
rect 58647 77763 58655 77797
rect 58605 77739 58655 77763
rect 58941 77797 58991 77821
rect 58941 77763 58949 77797
rect 58983 77763 58991 77797
rect 58941 77739 58991 77763
rect 59277 77797 59327 77821
rect 59277 77763 59285 77797
rect 59319 77763 59327 77797
rect 59277 77739 59327 77763
rect 59613 77797 59663 77821
rect 59613 77763 59621 77797
rect 59655 77763 59663 77797
rect 59613 77739 59663 77763
rect 59949 77797 59999 77821
rect 59949 77763 59957 77797
rect 59991 77763 59999 77797
rect 59949 77739 59999 77763
rect 60285 77797 60335 77821
rect 60285 77763 60293 77797
rect 60327 77763 60335 77797
rect 60285 77739 60335 77763
rect 60621 77797 60671 77821
rect 60621 77763 60629 77797
rect 60663 77763 60671 77797
rect 60621 77739 60671 77763
rect 60957 77797 61007 77821
rect 60957 77763 60965 77797
rect 60999 77763 61007 77797
rect 60957 77739 61007 77763
rect 61293 77797 61343 77821
rect 61293 77763 61301 77797
rect 61335 77763 61343 77797
rect 61293 77739 61343 77763
rect 61629 77797 61679 77821
rect 61629 77763 61637 77797
rect 61671 77763 61679 77797
rect 61629 77739 61679 77763
rect 61965 77797 62015 77821
rect 61965 77763 61973 77797
rect 62007 77763 62015 77797
rect 61965 77739 62015 77763
rect 62301 77797 62351 77821
rect 62301 77763 62309 77797
rect 62343 77763 62351 77797
rect 62301 77739 62351 77763
rect 62637 77797 62687 77821
rect 62637 77763 62645 77797
rect 62679 77763 62687 77797
rect 62637 77739 62687 77763
rect 62973 77797 63023 77821
rect 62973 77763 62981 77797
rect 63015 77763 63023 77797
rect 62973 77739 63023 77763
rect 63309 77797 63359 77821
rect 63309 77763 63317 77797
rect 63351 77763 63359 77797
rect 63309 77739 63359 77763
rect 63645 77797 63695 77821
rect 63645 77763 63653 77797
rect 63687 77763 63695 77797
rect 63645 77739 63695 77763
rect 63981 77797 64031 77821
rect 63981 77763 63989 77797
rect 64023 77763 64031 77797
rect 63981 77739 64031 77763
rect 64317 77797 64367 77821
rect 64317 77763 64325 77797
rect 64359 77763 64367 77797
rect 64317 77739 64367 77763
rect 64653 77797 64703 77821
rect 64653 77763 64661 77797
rect 64695 77763 64703 77797
rect 64653 77739 64703 77763
rect 64989 77797 65039 77821
rect 64989 77763 64997 77797
rect 65031 77763 65039 77797
rect 64989 77739 65039 77763
rect 65325 77797 65375 77821
rect 65325 77763 65333 77797
rect 65367 77763 65375 77797
rect 65325 77739 65375 77763
rect 65661 77797 65711 77821
rect 65661 77763 65669 77797
rect 65703 77763 65711 77797
rect 65661 77739 65711 77763
rect 65997 77797 66047 77821
rect 65997 77763 66005 77797
rect 66039 77763 66047 77797
rect 65997 77739 66047 77763
rect 66333 77797 66383 77821
rect 66333 77763 66341 77797
rect 66375 77763 66383 77797
rect 66333 77739 66383 77763
rect 66669 77797 66719 77821
rect 66669 77763 66677 77797
rect 66711 77763 66719 77797
rect 66669 77739 66719 77763
rect 67005 77797 67055 77821
rect 67005 77763 67013 77797
rect 67047 77763 67055 77797
rect 67005 77739 67055 77763
rect 67341 77797 67391 77821
rect 67341 77763 67349 77797
rect 67383 77763 67391 77797
rect 67341 77739 67391 77763
rect 67677 77797 67727 77821
rect 67677 77763 67685 77797
rect 67719 77763 67727 77797
rect 67677 77739 67727 77763
rect 68013 77797 68063 77821
rect 68013 77763 68021 77797
rect 68055 77763 68063 77797
rect 68013 77739 68063 77763
rect 68349 77797 68399 77821
rect 68349 77763 68357 77797
rect 68391 77763 68399 77797
rect 68349 77739 68399 77763
rect 68685 77797 68735 77821
rect 68685 77763 68693 77797
rect 68727 77763 68735 77797
rect 68685 77739 68735 77763
rect 69021 77797 69071 77821
rect 69021 77763 69029 77797
rect 69063 77763 69071 77797
rect 69021 77739 69071 77763
rect 69357 77797 69407 77821
rect 69357 77763 69365 77797
rect 69399 77763 69407 77797
rect 69357 77739 69407 77763
rect 69693 77797 69743 77821
rect 69693 77763 69701 77797
rect 69735 77763 69743 77797
rect 69693 77739 69743 77763
rect 70029 77797 70079 77821
rect 70029 77763 70037 77797
rect 70071 77763 70079 77797
rect 70029 77739 70079 77763
rect 70365 77797 70415 77821
rect 70365 77763 70373 77797
rect 70407 77763 70415 77797
rect 70365 77739 70415 77763
rect 70701 77797 70751 77821
rect 70701 77763 70709 77797
rect 70743 77763 70751 77797
rect 70701 77739 70751 77763
rect 71037 77797 71087 77821
rect 71037 77763 71045 77797
rect 71079 77763 71087 77797
rect 71037 77739 71087 77763
rect 71373 77797 71423 77821
rect 71373 77763 71381 77797
rect 71415 77763 71423 77797
rect 71373 77739 71423 77763
rect 71709 77797 71759 77821
rect 71709 77763 71717 77797
rect 71751 77763 71759 77797
rect 71709 77739 71759 77763
rect 72045 77797 72095 77821
rect 72045 77763 72053 77797
rect 72087 77763 72095 77797
rect 72045 77739 72095 77763
rect 72381 77797 72431 77821
rect 72381 77763 72389 77797
rect 72423 77763 72431 77797
rect 72381 77739 72431 77763
rect 72717 77797 72767 77821
rect 72717 77763 72725 77797
rect 72759 77763 72767 77797
rect 72717 77739 72767 77763
rect 73053 77797 73103 77821
rect 73053 77763 73061 77797
rect 73095 77763 73103 77797
rect 73053 77739 73103 77763
rect 73389 77797 73439 77821
rect 73389 77763 73397 77797
rect 73431 77763 73439 77797
rect 73389 77739 73439 77763
rect 73725 77797 73775 77821
rect 73725 77763 73733 77797
rect 73767 77763 73775 77797
rect 73725 77739 73775 77763
rect 74061 77797 74111 77821
rect 74061 77763 74069 77797
rect 74103 77763 74111 77797
rect 74061 77739 74111 77763
rect 74397 77797 74447 77821
rect 74397 77763 74405 77797
rect 74439 77763 74447 77797
rect 74397 77739 74447 77763
rect 74733 77797 74783 77821
rect 74733 77763 74741 77797
rect 74775 77763 74783 77797
rect 74733 77739 74783 77763
rect 75069 77797 75119 77821
rect 75069 77763 75077 77797
rect 75111 77763 75119 77797
rect 75069 77739 75119 77763
rect 75405 77797 75455 77821
rect 75405 77763 75413 77797
rect 75447 77763 75455 77797
rect 75405 77739 75455 77763
rect 75741 77797 75791 77821
rect 75741 77763 75749 77797
rect 75783 77763 75791 77797
rect 75741 77739 75791 77763
rect 76077 77797 76127 77821
rect 76077 77763 76085 77797
rect 76119 77763 76127 77797
rect 76077 77739 76127 77763
rect 76413 77797 76463 77821
rect 76413 77763 76421 77797
rect 76455 77763 76463 77797
rect 76413 77739 76463 77763
rect 76749 77797 76799 77821
rect 76749 77763 76757 77797
rect 76791 77763 76799 77797
rect 76749 77739 76799 77763
rect 77085 77797 77135 77821
rect 77085 77763 77093 77797
rect 77127 77763 77135 77797
rect 77085 77739 77135 77763
rect 77421 77797 77471 77821
rect 77421 77763 77429 77797
rect 77463 77763 77471 77797
rect 77421 77739 77471 77763
rect 77757 77797 77807 77821
rect 77757 77763 77765 77797
rect 77799 77763 77807 77797
rect 77757 77739 77807 77763
rect 78093 77797 78143 77821
rect 78093 77763 78101 77797
rect 78135 77763 78143 77797
rect 78093 77739 78143 77763
rect 78429 77797 78479 77821
rect 78429 77763 78437 77797
rect 78471 77763 78479 77797
rect 78429 77739 78479 77763
rect 78765 77797 78815 77821
rect 78765 77763 78773 77797
rect 78807 77763 78815 77797
rect 78765 77739 78815 77763
rect 79101 77797 79151 77821
rect 79101 77763 79109 77797
rect 79143 77763 79151 77797
rect 79101 77739 79151 77763
rect 79437 77797 79487 77821
rect 79437 77763 79445 77797
rect 79479 77763 79487 77797
rect 79437 77739 79487 77763
rect 79773 77797 79823 77821
rect 79773 77763 79781 77797
rect 79815 77763 79823 77797
rect 79773 77739 79823 77763
rect 80109 77797 80159 77821
rect 80109 77763 80117 77797
rect 80151 77763 80159 77797
rect 80109 77739 80159 77763
rect 80445 77797 80495 77821
rect 80445 77763 80453 77797
rect 80487 77763 80495 77797
rect 80445 77739 80495 77763
rect 80781 77797 80831 77821
rect 80781 77763 80789 77797
rect 80823 77763 80831 77797
rect 80781 77739 80831 77763
rect 81117 77797 81167 77821
rect 81117 77763 81125 77797
rect 81159 77763 81167 77797
rect 81117 77739 81167 77763
rect 81453 77797 81503 77821
rect 81453 77763 81461 77797
rect 81495 77763 81503 77797
rect 81453 77739 81503 77763
rect 81789 77797 81839 77821
rect 81789 77763 81797 77797
rect 81831 77763 81839 77797
rect 81789 77739 81839 77763
rect 82125 77797 82175 77821
rect 82125 77763 82133 77797
rect 82167 77763 82175 77797
rect 82125 77739 82175 77763
rect 82461 77797 82511 77821
rect 82461 77763 82469 77797
rect 82503 77763 82511 77797
rect 82461 77739 82511 77763
rect 82797 77797 82847 77821
rect 82797 77763 82805 77797
rect 82839 77763 82847 77797
rect 82797 77739 82847 77763
rect 83133 77797 83183 77821
rect 83133 77763 83141 77797
rect 83175 77763 83183 77797
rect 83133 77739 83183 77763
rect 83469 77797 83519 77821
rect 83469 77763 83477 77797
rect 83511 77763 83519 77797
rect 83469 77739 83519 77763
rect 83805 77797 83855 77821
rect 83805 77763 83813 77797
rect 83847 77763 83855 77797
rect 83805 77739 83855 77763
rect 84141 77797 84191 77821
rect 84141 77763 84149 77797
rect 84183 77763 84191 77797
rect 84141 77739 84191 77763
rect 84477 77797 84527 77821
rect 84477 77763 84485 77797
rect 84519 77763 84527 77797
rect 84477 77739 84527 77763
rect 84813 77797 84863 77821
rect 84813 77763 84821 77797
rect 84855 77763 84863 77797
rect 84813 77739 84863 77763
rect 85149 77797 85199 77821
rect 85149 77763 85157 77797
rect 85191 77763 85199 77797
rect 85149 77739 85199 77763
rect 85485 77797 85535 77821
rect 85485 77763 85493 77797
rect 85527 77763 85535 77797
rect 85485 77739 85535 77763
rect 85821 77797 85871 77821
rect 85821 77763 85829 77797
rect 85863 77763 85871 77797
rect 85821 77739 85871 77763
rect 86157 77797 86207 77821
rect 86157 77763 86165 77797
rect 86199 77763 86207 77797
rect 86157 77739 86207 77763
rect 86493 77797 86543 77821
rect 86493 77763 86501 77797
rect 86535 77763 86543 77797
rect 86493 77739 86543 77763
rect 86829 77797 86879 77821
rect 86829 77763 86837 77797
rect 86871 77763 86879 77797
rect 86829 77739 86879 77763
rect 87165 77797 87215 77821
rect 87165 77763 87173 77797
rect 87207 77763 87215 77797
rect 87165 77739 87215 77763
rect 87501 77797 87551 77821
rect 87501 77763 87509 77797
rect 87543 77763 87551 77797
rect 87501 77739 87551 77763
rect 87837 77797 87887 77821
rect 87837 77763 87845 77797
rect 87879 77763 87887 77797
rect 87837 77739 87887 77763
rect 88173 77797 88223 77821
rect 88173 77763 88181 77797
rect 88215 77763 88223 77797
rect 88173 77739 88223 77763
rect 88509 77797 88559 77821
rect 88509 77763 88517 77797
rect 88551 77763 88559 77797
rect 88509 77739 88559 77763
rect 88845 77797 88895 77821
rect 88845 77763 88853 77797
rect 88887 77763 88895 77797
rect 88845 77739 88895 77763
rect 89181 77797 89231 77821
rect 89181 77763 89189 77797
rect 89223 77763 89231 77797
rect 89181 77739 89231 77763
rect 89517 77797 89567 77821
rect 89517 77763 89525 77797
rect 89559 77763 89567 77797
rect 89517 77739 89567 77763
rect 89853 77797 89903 77821
rect 89853 77763 89861 77797
rect 89895 77763 89903 77797
rect 89853 77739 89903 77763
rect 90189 77797 90239 77821
rect 90189 77763 90197 77797
rect 90231 77763 90239 77797
rect 90189 77739 90239 77763
rect 90525 77797 90575 77821
rect 90525 77763 90533 77797
rect 90567 77763 90575 77797
rect 90525 77739 90575 77763
rect 90861 77797 90911 77821
rect 90861 77763 90869 77797
rect 90903 77763 90911 77797
rect 90861 77739 90911 77763
rect 91197 77797 91247 77821
rect 91197 77763 91205 77797
rect 91239 77763 91247 77797
rect 91197 77739 91247 77763
rect 91533 77797 91583 77821
rect 91533 77763 91541 77797
rect 91575 77763 91583 77797
rect 91533 77739 91583 77763
rect 91869 77797 91919 77821
rect 91869 77763 91877 77797
rect 91911 77763 91919 77797
rect 91869 77739 91919 77763
rect 92205 77797 92255 77821
rect 92205 77763 92213 77797
rect 92247 77763 92255 77797
rect 92205 77739 92255 77763
rect 92541 77797 92591 77821
rect 92541 77763 92549 77797
rect 92583 77763 92591 77797
rect 92541 77739 92591 77763
rect 92877 77797 92927 77821
rect 92877 77763 92885 77797
rect 92919 77763 92927 77797
rect 92877 77739 92927 77763
rect 93213 77797 93263 77821
rect 93213 77763 93221 77797
rect 93255 77763 93263 77797
rect 93213 77739 93263 77763
rect 93549 77797 93599 77821
rect 93549 77763 93557 77797
rect 93591 77763 93599 77797
rect 93549 77739 93599 77763
rect 1821 77333 1871 77357
rect 1821 77299 1829 77333
rect 1863 77299 1871 77333
rect 1821 77275 1871 77299
rect 94179 77333 94229 77357
rect 94179 77299 94187 77333
rect 94221 77299 94229 77333
rect 94179 77275 94229 77299
rect 1821 76997 1871 77021
rect 1821 76963 1829 76997
rect 1863 76963 1871 76997
rect 1821 76939 1871 76963
rect 94179 76997 94229 77021
rect 94179 76963 94187 76997
rect 94221 76963 94229 76997
rect 94179 76939 94229 76963
rect 1821 76661 1871 76685
rect 1821 76627 1829 76661
rect 1863 76627 1871 76661
rect 1821 76603 1871 76627
rect 94179 76661 94229 76685
rect 94179 76627 94187 76661
rect 94221 76627 94229 76661
rect 94179 76603 94229 76627
rect 1821 76325 1871 76349
rect 1821 76291 1829 76325
rect 1863 76291 1871 76325
rect 1821 76267 1871 76291
rect 94179 76325 94229 76349
rect 94179 76291 94187 76325
rect 94221 76291 94229 76325
rect 94179 76267 94229 76291
rect 1821 75989 1871 76013
rect 1821 75955 1829 75989
rect 1863 75955 1871 75989
rect 1821 75931 1871 75955
rect 94179 75989 94229 76013
rect 94179 75955 94187 75989
rect 94221 75955 94229 75989
rect 94179 75931 94229 75955
rect 1821 75653 1871 75677
rect 1821 75619 1829 75653
rect 1863 75619 1871 75653
rect 1821 75595 1871 75619
rect 94179 75653 94229 75677
rect 94179 75619 94187 75653
rect 94221 75619 94229 75653
rect 94179 75595 94229 75619
rect 1821 75317 1871 75341
rect 1821 75283 1829 75317
rect 1863 75283 1871 75317
rect 1821 75259 1871 75283
rect 94179 75317 94229 75341
rect 94179 75283 94187 75317
rect 94221 75283 94229 75317
rect 94179 75259 94229 75283
rect 1821 74981 1871 75005
rect 1821 74947 1829 74981
rect 1863 74947 1871 74981
rect 1821 74923 1871 74947
rect 94179 74981 94229 75005
rect 94179 74947 94187 74981
rect 94221 74947 94229 74981
rect 94179 74923 94229 74947
rect 1821 74645 1871 74669
rect 1821 74611 1829 74645
rect 1863 74611 1871 74645
rect 1821 74587 1871 74611
rect 94179 74645 94229 74669
rect 94179 74611 94187 74645
rect 94221 74611 94229 74645
rect 94179 74587 94229 74611
rect 1821 74309 1871 74333
rect 1821 74275 1829 74309
rect 1863 74275 1871 74309
rect 1821 74251 1871 74275
rect 94179 74309 94229 74333
rect 94179 74275 94187 74309
rect 94221 74275 94229 74309
rect 94179 74251 94229 74275
rect 1821 73973 1871 73997
rect 1821 73939 1829 73973
rect 1863 73939 1871 73973
rect 1821 73915 1871 73939
rect 94179 73973 94229 73997
rect 94179 73939 94187 73973
rect 94221 73939 94229 73973
rect 94179 73915 94229 73939
rect 1821 73637 1871 73661
rect 1821 73603 1829 73637
rect 1863 73603 1871 73637
rect 1821 73579 1871 73603
rect 94179 73637 94229 73661
rect 94179 73603 94187 73637
rect 94221 73603 94229 73637
rect 94179 73579 94229 73603
rect 1821 73301 1871 73325
rect 1821 73267 1829 73301
rect 1863 73267 1871 73301
rect 1821 73243 1871 73267
rect 94179 73301 94229 73325
rect 94179 73267 94187 73301
rect 94221 73267 94229 73301
rect 94179 73243 94229 73267
rect 1821 72965 1871 72989
rect 1821 72931 1829 72965
rect 1863 72931 1871 72965
rect 1821 72907 1871 72931
rect 94179 72965 94229 72989
rect 94179 72931 94187 72965
rect 94221 72931 94229 72965
rect 94179 72907 94229 72931
rect 1821 72629 1871 72653
rect 1821 72595 1829 72629
rect 1863 72595 1871 72629
rect 1821 72571 1871 72595
rect 94179 72629 94229 72653
rect 94179 72595 94187 72629
rect 94221 72595 94229 72629
rect 94179 72571 94229 72595
rect 1821 72293 1871 72317
rect 1821 72259 1829 72293
rect 1863 72259 1871 72293
rect 1821 72235 1871 72259
rect 94179 72293 94229 72317
rect 94179 72259 94187 72293
rect 94221 72259 94229 72293
rect 94179 72235 94229 72259
rect 1821 71957 1871 71981
rect 1821 71923 1829 71957
rect 1863 71923 1871 71957
rect 1821 71899 1871 71923
rect 94179 71957 94229 71981
rect 94179 71923 94187 71957
rect 94221 71923 94229 71957
rect 94179 71899 94229 71923
rect 1821 71621 1871 71645
rect 1821 71587 1829 71621
rect 1863 71587 1871 71621
rect 1821 71563 1871 71587
rect 94179 71621 94229 71645
rect 94179 71587 94187 71621
rect 94221 71587 94229 71621
rect 94179 71563 94229 71587
rect 1821 71285 1871 71309
rect 1821 71251 1829 71285
rect 1863 71251 1871 71285
rect 1821 71227 1871 71251
rect 94179 71285 94229 71309
rect 94179 71251 94187 71285
rect 94221 71251 94229 71285
rect 94179 71227 94229 71251
rect 1821 70949 1871 70973
rect 1821 70915 1829 70949
rect 1863 70915 1871 70949
rect 1821 70891 1871 70915
rect 94179 70949 94229 70973
rect 94179 70915 94187 70949
rect 94221 70915 94229 70949
rect 94179 70891 94229 70915
rect 1821 70613 1871 70637
rect 1821 70579 1829 70613
rect 1863 70579 1871 70613
rect 1821 70555 1871 70579
rect 94179 70613 94229 70637
rect 94179 70579 94187 70613
rect 94221 70579 94229 70613
rect 94179 70555 94229 70579
rect 1821 70277 1871 70301
rect 1821 70243 1829 70277
rect 1863 70243 1871 70277
rect 1821 70219 1871 70243
rect 94179 70277 94229 70301
rect 94179 70243 94187 70277
rect 94221 70243 94229 70277
rect 94179 70219 94229 70243
rect 1821 69941 1871 69965
rect 1821 69907 1829 69941
rect 1863 69907 1871 69941
rect 1821 69883 1871 69907
rect 94179 69941 94229 69965
rect 94179 69907 94187 69941
rect 94221 69907 94229 69941
rect 94179 69883 94229 69907
rect 1821 69605 1871 69629
rect 1821 69571 1829 69605
rect 1863 69571 1871 69605
rect 1821 69547 1871 69571
rect 94179 69605 94229 69629
rect 94179 69571 94187 69605
rect 94221 69571 94229 69605
rect 94179 69547 94229 69571
rect 1821 69269 1871 69293
rect 1821 69235 1829 69269
rect 1863 69235 1871 69269
rect 1821 69211 1871 69235
rect 94179 69269 94229 69293
rect 94179 69235 94187 69269
rect 94221 69235 94229 69269
rect 94179 69211 94229 69235
rect 1821 68933 1871 68957
rect 1821 68899 1829 68933
rect 1863 68899 1871 68933
rect 1821 68875 1871 68899
rect 94179 68933 94229 68957
rect 94179 68899 94187 68933
rect 94221 68899 94229 68933
rect 94179 68875 94229 68899
rect 1821 68597 1871 68621
rect 1821 68563 1829 68597
rect 1863 68563 1871 68597
rect 1821 68539 1871 68563
rect 94179 68597 94229 68621
rect 94179 68563 94187 68597
rect 94221 68563 94229 68597
rect 94179 68539 94229 68563
rect 1821 68261 1871 68285
rect 1821 68227 1829 68261
rect 1863 68227 1871 68261
rect 1821 68203 1871 68227
rect 94179 68261 94229 68285
rect 94179 68227 94187 68261
rect 94221 68227 94229 68261
rect 94179 68203 94229 68227
rect 1821 67925 1871 67949
rect 1821 67891 1829 67925
rect 1863 67891 1871 67925
rect 1821 67867 1871 67891
rect 94179 67925 94229 67949
rect 94179 67891 94187 67925
rect 94221 67891 94229 67925
rect 94179 67867 94229 67891
rect 1821 67589 1871 67613
rect 1821 67555 1829 67589
rect 1863 67555 1871 67589
rect 1821 67531 1871 67555
rect 94179 67589 94229 67613
rect 94179 67555 94187 67589
rect 94221 67555 94229 67589
rect 94179 67531 94229 67555
rect 1821 67253 1871 67277
rect 1821 67219 1829 67253
rect 1863 67219 1871 67253
rect 1821 67195 1871 67219
rect 94179 67253 94229 67277
rect 94179 67219 94187 67253
rect 94221 67219 94229 67253
rect 94179 67195 94229 67219
rect 1821 66917 1871 66941
rect 1821 66883 1829 66917
rect 1863 66883 1871 66917
rect 1821 66859 1871 66883
rect 94179 66917 94229 66941
rect 94179 66883 94187 66917
rect 94221 66883 94229 66917
rect 94179 66859 94229 66883
rect 1821 66581 1871 66605
rect 1821 66547 1829 66581
rect 1863 66547 1871 66581
rect 1821 66523 1871 66547
rect 94179 66581 94229 66605
rect 94179 66547 94187 66581
rect 94221 66547 94229 66581
rect 94179 66523 94229 66547
rect 1821 66245 1871 66269
rect 1821 66211 1829 66245
rect 1863 66211 1871 66245
rect 1821 66187 1871 66211
rect 94179 66245 94229 66269
rect 94179 66211 94187 66245
rect 94221 66211 94229 66245
rect 94179 66187 94229 66211
rect 1821 65909 1871 65933
rect 1821 65875 1829 65909
rect 1863 65875 1871 65909
rect 1821 65851 1871 65875
rect 94179 65909 94229 65933
rect 94179 65875 94187 65909
rect 94221 65875 94229 65909
rect 94179 65851 94229 65875
rect 1821 65573 1871 65597
rect 1821 65539 1829 65573
rect 1863 65539 1871 65573
rect 1821 65515 1871 65539
rect 94179 65573 94229 65597
rect 94179 65539 94187 65573
rect 94221 65539 94229 65573
rect 94179 65515 94229 65539
rect 1821 65237 1871 65261
rect 1821 65203 1829 65237
rect 1863 65203 1871 65237
rect 1821 65179 1871 65203
rect 94179 65237 94229 65261
rect 94179 65203 94187 65237
rect 94221 65203 94229 65237
rect 94179 65179 94229 65203
rect 1821 64901 1871 64925
rect 1821 64867 1829 64901
rect 1863 64867 1871 64901
rect 1821 64843 1871 64867
rect 94179 64901 94229 64925
rect 94179 64867 94187 64901
rect 94221 64867 94229 64901
rect 94179 64843 94229 64867
rect 1821 64565 1871 64589
rect 1821 64531 1829 64565
rect 1863 64531 1871 64565
rect 1821 64507 1871 64531
rect 94179 64565 94229 64589
rect 94179 64531 94187 64565
rect 94221 64531 94229 64565
rect 94179 64507 94229 64531
rect 1821 64229 1871 64253
rect 1821 64195 1829 64229
rect 1863 64195 1871 64229
rect 1821 64171 1871 64195
rect 94179 64229 94229 64253
rect 94179 64195 94187 64229
rect 94221 64195 94229 64229
rect 94179 64171 94229 64195
rect 1821 63893 1871 63917
rect 1821 63859 1829 63893
rect 1863 63859 1871 63893
rect 1821 63835 1871 63859
rect 94179 63893 94229 63917
rect 94179 63859 94187 63893
rect 94221 63859 94229 63893
rect 94179 63835 94229 63859
rect 1821 63557 1871 63581
rect 1821 63523 1829 63557
rect 1863 63523 1871 63557
rect 1821 63499 1871 63523
rect 94179 63557 94229 63581
rect 94179 63523 94187 63557
rect 94221 63523 94229 63557
rect 94179 63499 94229 63523
rect 1821 63221 1871 63245
rect 1821 63187 1829 63221
rect 1863 63187 1871 63221
rect 1821 63163 1871 63187
rect 94179 63221 94229 63245
rect 94179 63187 94187 63221
rect 94221 63187 94229 63221
rect 94179 63163 94229 63187
rect 1821 62885 1871 62909
rect 1821 62851 1829 62885
rect 1863 62851 1871 62885
rect 1821 62827 1871 62851
rect 94179 62885 94229 62909
rect 94179 62851 94187 62885
rect 94221 62851 94229 62885
rect 94179 62827 94229 62851
rect 1821 62549 1871 62573
rect 1821 62515 1829 62549
rect 1863 62515 1871 62549
rect 1821 62491 1871 62515
rect 94179 62549 94229 62573
rect 94179 62515 94187 62549
rect 94221 62515 94229 62549
rect 94179 62491 94229 62515
rect 1821 62213 1871 62237
rect 1821 62179 1829 62213
rect 1863 62179 1871 62213
rect 1821 62155 1871 62179
rect 94179 62213 94229 62237
rect 94179 62179 94187 62213
rect 94221 62179 94229 62213
rect 94179 62155 94229 62179
rect 1821 61877 1871 61901
rect 1821 61843 1829 61877
rect 1863 61843 1871 61877
rect 1821 61819 1871 61843
rect 94179 61877 94229 61901
rect 94179 61843 94187 61877
rect 94221 61843 94229 61877
rect 94179 61819 94229 61843
rect 1821 61541 1871 61565
rect 1821 61507 1829 61541
rect 1863 61507 1871 61541
rect 1821 61483 1871 61507
rect 94179 61541 94229 61565
rect 94179 61507 94187 61541
rect 94221 61507 94229 61541
rect 94179 61483 94229 61507
rect 1821 61205 1871 61229
rect 1821 61171 1829 61205
rect 1863 61171 1871 61205
rect 1821 61147 1871 61171
rect 94179 61205 94229 61229
rect 94179 61171 94187 61205
rect 94221 61171 94229 61205
rect 94179 61147 94229 61171
rect 1821 60869 1871 60893
rect 1821 60835 1829 60869
rect 1863 60835 1871 60869
rect 1821 60811 1871 60835
rect 94179 60869 94229 60893
rect 94179 60835 94187 60869
rect 94221 60835 94229 60869
rect 94179 60811 94229 60835
rect 1821 60533 1871 60557
rect 1821 60499 1829 60533
rect 1863 60499 1871 60533
rect 1821 60475 1871 60499
rect 94179 60533 94229 60557
rect 94179 60499 94187 60533
rect 94221 60499 94229 60533
rect 94179 60475 94229 60499
rect 1821 60197 1871 60221
rect 1821 60163 1829 60197
rect 1863 60163 1871 60197
rect 1821 60139 1871 60163
rect 94179 60197 94229 60221
rect 94179 60163 94187 60197
rect 94221 60163 94229 60197
rect 94179 60139 94229 60163
rect 1821 59861 1871 59885
rect 1821 59827 1829 59861
rect 1863 59827 1871 59861
rect 1821 59803 1871 59827
rect 94179 59861 94229 59885
rect 94179 59827 94187 59861
rect 94221 59827 94229 59861
rect 94179 59803 94229 59827
rect 1821 59525 1871 59549
rect 1821 59491 1829 59525
rect 1863 59491 1871 59525
rect 1821 59467 1871 59491
rect 94179 59525 94229 59549
rect 94179 59491 94187 59525
rect 94221 59491 94229 59525
rect 94179 59467 94229 59491
rect 1821 59189 1871 59213
rect 1821 59155 1829 59189
rect 1863 59155 1871 59189
rect 1821 59131 1871 59155
rect 94179 59189 94229 59213
rect 94179 59155 94187 59189
rect 94221 59155 94229 59189
rect 94179 59131 94229 59155
rect 1821 58853 1871 58877
rect 1821 58819 1829 58853
rect 1863 58819 1871 58853
rect 1821 58795 1871 58819
rect 94179 58853 94229 58877
rect 94179 58819 94187 58853
rect 94221 58819 94229 58853
rect 94179 58795 94229 58819
rect 1821 58517 1871 58541
rect 1821 58483 1829 58517
rect 1863 58483 1871 58517
rect 1821 58459 1871 58483
rect 94179 58517 94229 58541
rect 94179 58483 94187 58517
rect 94221 58483 94229 58517
rect 94179 58459 94229 58483
rect 1821 58181 1871 58205
rect 1821 58147 1829 58181
rect 1863 58147 1871 58181
rect 1821 58123 1871 58147
rect 94179 58181 94229 58205
rect 94179 58147 94187 58181
rect 94221 58147 94229 58181
rect 94179 58123 94229 58147
rect 1821 57845 1871 57869
rect 1821 57811 1829 57845
rect 1863 57811 1871 57845
rect 1821 57787 1871 57811
rect 94179 57845 94229 57869
rect 94179 57811 94187 57845
rect 94221 57811 94229 57845
rect 94179 57787 94229 57811
rect 1821 57509 1871 57533
rect 1821 57475 1829 57509
rect 1863 57475 1871 57509
rect 1821 57451 1871 57475
rect 94179 57509 94229 57533
rect 94179 57475 94187 57509
rect 94221 57475 94229 57509
rect 94179 57451 94229 57475
rect 1821 57173 1871 57197
rect 1821 57139 1829 57173
rect 1863 57139 1871 57173
rect 1821 57115 1871 57139
rect 94179 57173 94229 57197
rect 94179 57139 94187 57173
rect 94221 57139 94229 57173
rect 94179 57115 94229 57139
rect 1821 56837 1871 56861
rect 1821 56803 1829 56837
rect 1863 56803 1871 56837
rect 1821 56779 1871 56803
rect 94179 56837 94229 56861
rect 94179 56803 94187 56837
rect 94221 56803 94229 56837
rect 94179 56779 94229 56803
rect 1821 56501 1871 56525
rect 1821 56467 1829 56501
rect 1863 56467 1871 56501
rect 1821 56443 1871 56467
rect 94179 56501 94229 56525
rect 94179 56467 94187 56501
rect 94221 56467 94229 56501
rect 94179 56443 94229 56467
rect 1821 56165 1871 56189
rect 1821 56131 1829 56165
rect 1863 56131 1871 56165
rect 1821 56107 1871 56131
rect 94179 56165 94229 56189
rect 94179 56131 94187 56165
rect 94221 56131 94229 56165
rect 94179 56107 94229 56131
rect 1821 55829 1871 55853
rect 1821 55795 1829 55829
rect 1863 55795 1871 55829
rect 1821 55771 1871 55795
rect 94179 55829 94229 55853
rect 94179 55795 94187 55829
rect 94221 55795 94229 55829
rect 94179 55771 94229 55795
rect 1821 55493 1871 55517
rect 1821 55459 1829 55493
rect 1863 55459 1871 55493
rect 1821 55435 1871 55459
rect 94179 55493 94229 55517
rect 94179 55459 94187 55493
rect 94221 55459 94229 55493
rect 94179 55435 94229 55459
rect 1821 55157 1871 55181
rect 1821 55123 1829 55157
rect 1863 55123 1871 55157
rect 1821 55099 1871 55123
rect 94179 55157 94229 55181
rect 94179 55123 94187 55157
rect 94221 55123 94229 55157
rect 94179 55099 94229 55123
rect 1821 54821 1871 54845
rect 1821 54787 1829 54821
rect 1863 54787 1871 54821
rect 1821 54763 1871 54787
rect 94179 54821 94229 54845
rect 94179 54787 94187 54821
rect 94221 54787 94229 54821
rect 94179 54763 94229 54787
rect 1821 54485 1871 54509
rect 1821 54451 1829 54485
rect 1863 54451 1871 54485
rect 1821 54427 1871 54451
rect 94179 54485 94229 54509
rect 94179 54451 94187 54485
rect 94221 54451 94229 54485
rect 94179 54427 94229 54451
rect 1821 54149 1871 54173
rect 1821 54115 1829 54149
rect 1863 54115 1871 54149
rect 1821 54091 1871 54115
rect 94179 54149 94229 54173
rect 94179 54115 94187 54149
rect 94221 54115 94229 54149
rect 94179 54091 94229 54115
rect 1821 53813 1871 53837
rect 1821 53779 1829 53813
rect 1863 53779 1871 53813
rect 1821 53755 1871 53779
rect 94179 53813 94229 53837
rect 94179 53779 94187 53813
rect 94221 53779 94229 53813
rect 94179 53755 94229 53779
rect 1821 53477 1871 53501
rect 1821 53443 1829 53477
rect 1863 53443 1871 53477
rect 1821 53419 1871 53443
rect 94179 53477 94229 53501
rect 94179 53443 94187 53477
rect 94221 53443 94229 53477
rect 94179 53419 94229 53443
rect 1821 53141 1871 53165
rect 1821 53107 1829 53141
rect 1863 53107 1871 53141
rect 1821 53083 1871 53107
rect 94179 53141 94229 53165
rect 94179 53107 94187 53141
rect 94221 53107 94229 53141
rect 94179 53083 94229 53107
rect 1821 52805 1871 52829
rect 1821 52771 1829 52805
rect 1863 52771 1871 52805
rect 1821 52747 1871 52771
rect 94179 52805 94229 52829
rect 94179 52771 94187 52805
rect 94221 52771 94229 52805
rect 94179 52747 94229 52771
rect 1821 52469 1871 52493
rect 1821 52435 1829 52469
rect 1863 52435 1871 52469
rect 1821 52411 1871 52435
rect 94179 52469 94229 52493
rect 94179 52435 94187 52469
rect 94221 52435 94229 52469
rect 94179 52411 94229 52435
rect 1821 52133 1871 52157
rect 1821 52099 1829 52133
rect 1863 52099 1871 52133
rect 1821 52075 1871 52099
rect 94179 52133 94229 52157
rect 94179 52099 94187 52133
rect 94221 52099 94229 52133
rect 94179 52075 94229 52099
rect 1821 51797 1871 51821
rect 1821 51763 1829 51797
rect 1863 51763 1871 51797
rect 1821 51739 1871 51763
rect 94179 51797 94229 51821
rect 94179 51763 94187 51797
rect 94221 51763 94229 51797
rect 94179 51739 94229 51763
rect 1821 51461 1871 51485
rect 1821 51427 1829 51461
rect 1863 51427 1871 51461
rect 1821 51403 1871 51427
rect 94179 51461 94229 51485
rect 94179 51427 94187 51461
rect 94221 51427 94229 51461
rect 94179 51403 94229 51427
rect 1821 51125 1871 51149
rect 1821 51091 1829 51125
rect 1863 51091 1871 51125
rect 1821 51067 1871 51091
rect 94179 51125 94229 51149
rect 94179 51091 94187 51125
rect 94221 51091 94229 51125
rect 94179 51067 94229 51091
rect 1821 50789 1871 50813
rect 1821 50755 1829 50789
rect 1863 50755 1871 50789
rect 1821 50731 1871 50755
rect 94179 50789 94229 50813
rect 94179 50755 94187 50789
rect 94221 50755 94229 50789
rect 94179 50731 94229 50755
rect 1821 50453 1871 50477
rect 1821 50419 1829 50453
rect 1863 50419 1871 50453
rect 1821 50395 1871 50419
rect 94179 50453 94229 50477
rect 94179 50419 94187 50453
rect 94221 50419 94229 50453
rect 94179 50395 94229 50419
rect 1821 50117 1871 50141
rect 1821 50083 1829 50117
rect 1863 50083 1871 50117
rect 1821 50059 1871 50083
rect 94179 50117 94229 50141
rect 94179 50083 94187 50117
rect 94221 50083 94229 50117
rect 94179 50059 94229 50083
rect 1821 49781 1871 49805
rect 1821 49747 1829 49781
rect 1863 49747 1871 49781
rect 1821 49723 1871 49747
rect 94179 49781 94229 49805
rect 94179 49747 94187 49781
rect 94221 49747 94229 49781
rect 94179 49723 94229 49747
rect 1821 49445 1871 49469
rect 1821 49411 1829 49445
rect 1863 49411 1871 49445
rect 1821 49387 1871 49411
rect 94179 49445 94229 49469
rect 94179 49411 94187 49445
rect 94221 49411 94229 49445
rect 94179 49387 94229 49411
rect 1821 49109 1871 49133
rect 1821 49075 1829 49109
rect 1863 49075 1871 49109
rect 1821 49051 1871 49075
rect 94179 49109 94229 49133
rect 94179 49075 94187 49109
rect 94221 49075 94229 49109
rect 94179 49051 94229 49075
rect 1821 48773 1871 48797
rect 1821 48739 1829 48773
rect 1863 48739 1871 48773
rect 1821 48715 1871 48739
rect 94179 48773 94229 48797
rect 94179 48739 94187 48773
rect 94221 48739 94229 48773
rect 94179 48715 94229 48739
rect 1821 48437 1871 48461
rect 1821 48403 1829 48437
rect 1863 48403 1871 48437
rect 1821 48379 1871 48403
rect 94179 48437 94229 48461
rect 94179 48403 94187 48437
rect 94221 48403 94229 48437
rect 94179 48379 94229 48403
rect 1821 48101 1871 48125
rect 1821 48067 1829 48101
rect 1863 48067 1871 48101
rect 1821 48043 1871 48067
rect 94179 48101 94229 48125
rect 94179 48067 94187 48101
rect 94221 48067 94229 48101
rect 94179 48043 94229 48067
rect 1821 47765 1871 47789
rect 1821 47731 1829 47765
rect 1863 47731 1871 47765
rect 1821 47707 1871 47731
rect 94179 47765 94229 47789
rect 94179 47731 94187 47765
rect 94221 47731 94229 47765
rect 94179 47707 94229 47731
rect 1821 47429 1871 47453
rect 1821 47395 1829 47429
rect 1863 47395 1871 47429
rect 1821 47371 1871 47395
rect 94179 47429 94229 47453
rect 94179 47395 94187 47429
rect 94221 47395 94229 47429
rect 94179 47371 94229 47395
rect 1821 47093 1871 47117
rect 1821 47059 1829 47093
rect 1863 47059 1871 47093
rect 1821 47035 1871 47059
rect 94179 47093 94229 47117
rect 94179 47059 94187 47093
rect 94221 47059 94229 47093
rect 94179 47035 94229 47059
rect 1821 46757 1871 46781
rect 1821 46723 1829 46757
rect 1863 46723 1871 46757
rect 1821 46699 1871 46723
rect 94179 46757 94229 46781
rect 94179 46723 94187 46757
rect 94221 46723 94229 46757
rect 94179 46699 94229 46723
rect 1821 46421 1871 46445
rect 1821 46387 1829 46421
rect 1863 46387 1871 46421
rect 1821 46363 1871 46387
rect 94179 46421 94229 46445
rect 94179 46387 94187 46421
rect 94221 46387 94229 46421
rect 94179 46363 94229 46387
rect 1821 46085 1871 46109
rect 1821 46051 1829 46085
rect 1863 46051 1871 46085
rect 1821 46027 1871 46051
rect 94179 46085 94229 46109
rect 94179 46051 94187 46085
rect 94221 46051 94229 46085
rect 94179 46027 94229 46051
rect 1821 45749 1871 45773
rect 1821 45715 1829 45749
rect 1863 45715 1871 45749
rect 1821 45691 1871 45715
rect 94179 45749 94229 45773
rect 94179 45715 94187 45749
rect 94221 45715 94229 45749
rect 94179 45691 94229 45715
rect 1821 45413 1871 45437
rect 1821 45379 1829 45413
rect 1863 45379 1871 45413
rect 1821 45355 1871 45379
rect 94179 45413 94229 45437
rect 94179 45379 94187 45413
rect 94221 45379 94229 45413
rect 94179 45355 94229 45379
rect 1821 45077 1871 45101
rect 1821 45043 1829 45077
rect 1863 45043 1871 45077
rect 1821 45019 1871 45043
rect 94179 45077 94229 45101
rect 94179 45043 94187 45077
rect 94221 45043 94229 45077
rect 94179 45019 94229 45043
rect 1821 44741 1871 44765
rect 1821 44707 1829 44741
rect 1863 44707 1871 44741
rect 1821 44683 1871 44707
rect 94179 44741 94229 44765
rect 94179 44707 94187 44741
rect 94221 44707 94229 44741
rect 94179 44683 94229 44707
rect 1821 44405 1871 44429
rect 1821 44371 1829 44405
rect 1863 44371 1871 44405
rect 1821 44347 1871 44371
rect 94179 44405 94229 44429
rect 94179 44371 94187 44405
rect 94221 44371 94229 44405
rect 94179 44347 94229 44371
rect 1821 44069 1871 44093
rect 1821 44035 1829 44069
rect 1863 44035 1871 44069
rect 1821 44011 1871 44035
rect 94179 44069 94229 44093
rect 94179 44035 94187 44069
rect 94221 44035 94229 44069
rect 94179 44011 94229 44035
rect 1821 43733 1871 43757
rect 1821 43699 1829 43733
rect 1863 43699 1871 43733
rect 1821 43675 1871 43699
rect 94179 43733 94229 43757
rect 94179 43699 94187 43733
rect 94221 43699 94229 43733
rect 94179 43675 94229 43699
rect 1821 43397 1871 43421
rect 1821 43363 1829 43397
rect 1863 43363 1871 43397
rect 1821 43339 1871 43363
rect 94179 43397 94229 43421
rect 94179 43363 94187 43397
rect 94221 43363 94229 43397
rect 94179 43339 94229 43363
rect 1821 43061 1871 43085
rect 1821 43027 1829 43061
rect 1863 43027 1871 43061
rect 1821 43003 1871 43027
rect 94179 43061 94229 43085
rect 94179 43027 94187 43061
rect 94221 43027 94229 43061
rect 94179 43003 94229 43027
rect 1821 42725 1871 42749
rect 1821 42691 1829 42725
rect 1863 42691 1871 42725
rect 1821 42667 1871 42691
rect 94179 42725 94229 42749
rect 94179 42691 94187 42725
rect 94221 42691 94229 42725
rect 94179 42667 94229 42691
rect 1821 42389 1871 42413
rect 1821 42355 1829 42389
rect 1863 42355 1871 42389
rect 1821 42331 1871 42355
rect 94179 42389 94229 42413
rect 94179 42355 94187 42389
rect 94221 42355 94229 42389
rect 94179 42331 94229 42355
rect 1821 42053 1871 42077
rect 1821 42019 1829 42053
rect 1863 42019 1871 42053
rect 1821 41995 1871 42019
rect 94179 42053 94229 42077
rect 94179 42019 94187 42053
rect 94221 42019 94229 42053
rect 94179 41995 94229 42019
rect 1821 41717 1871 41741
rect 1821 41683 1829 41717
rect 1863 41683 1871 41717
rect 1821 41659 1871 41683
rect 94179 41717 94229 41741
rect 94179 41683 94187 41717
rect 94221 41683 94229 41717
rect 94179 41659 94229 41683
rect 1821 41381 1871 41405
rect 1821 41347 1829 41381
rect 1863 41347 1871 41381
rect 1821 41323 1871 41347
rect 94179 41381 94229 41405
rect 94179 41347 94187 41381
rect 94221 41347 94229 41381
rect 94179 41323 94229 41347
rect 1821 41045 1871 41069
rect 1821 41011 1829 41045
rect 1863 41011 1871 41045
rect 1821 40987 1871 41011
rect 94179 41045 94229 41069
rect 94179 41011 94187 41045
rect 94221 41011 94229 41045
rect 94179 40987 94229 41011
rect 1821 40709 1871 40733
rect 1821 40675 1829 40709
rect 1863 40675 1871 40709
rect 1821 40651 1871 40675
rect 94179 40709 94229 40733
rect 94179 40675 94187 40709
rect 94221 40675 94229 40709
rect 94179 40651 94229 40675
rect 1821 40373 1871 40397
rect 1821 40339 1829 40373
rect 1863 40339 1871 40373
rect 1821 40315 1871 40339
rect 94179 40373 94229 40397
rect 94179 40339 94187 40373
rect 94221 40339 94229 40373
rect 94179 40315 94229 40339
rect 1821 40037 1871 40061
rect 1821 40003 1829 40037
rect 1863 40003 1871 40037
rect 1821 39979 1871 40003
rect 94179 40037 94229 40061
rect 94179 40003 94187 40037
rect 94221 40003 94229 40037
rect 94179 39979 94229 40003
rect 1821 39701 1871 39725
rect 1821 39667 1829 39701
rect 1863 39667 1871 39701
rect 1821 39643 1871 39667
rect 94179 39701 94229 39725
rect 94179 39667 94187 39701
rect 94221 39667 94229 39701
rect 94179 39643 94229 39667
rect 1821 39365 1871 39389
rect 1821 39331 1829 39365
rect 1863 39331 1871 39365
rect 1821 39307 1871 39331
rect 94179 39365 94229 39389
rect 94179 39331 94187 39365
rect 94221 39331 94229 39365
rect 94179 39307 94229 39331
rect 1821 39029 1871 39053
rect 1821 38995 1829 39029
rect 1863 38995 1871 39029
rect 1821 38971 1871 38995
rect 94179 39029 94229 39053
rect 94179 38995 94187 39029
rect 94221 38995 94229 39029
rect 94179 38971 94229 38995
rect 1821 38693 1871 38717
rect 1821 38659 1829 38693
rect 1863 38659 1871 38693
rect 1821 38635 1871 38659
rect 94179 38693 94229 38717
rect 94179 38659 94187 38693
rect 94221 38659 94229 38693
rect 94179 38635 94229 38659
rect 1821 38357 1871 38381
rect 1821 38323 1829 38357
rect 1863 38323 1871 38357
rect 1821 38299 1871 38323
rect 94179 38357 94229 38381
rect 94179 38323 94187 38357
rect 94221 38323 94229 38357
rect 94179 38299 94229 38323
rect 1821 38021 1871 38045
rect 1821 37987 1829 38021
rect 1863 37987 1871 38021
rect 1821 37963 1871 37987
rect 94179 38021 94229 38045
rect 94179 37987 94187 38021
rect 94221 37987 94229 38021
rect 94179 37963 94229 37987
rect 1821 37685 1871 37709
rect 1821 37651 1829 37685
rect 1863 37651 1871 37685
rect 1821 37627 1871 37651
rect 94179 37685 94229 37709
rect 94179 37651 94187 37685
rect 94221 37651 94229 37685
rect 94179 37627 94229 37651
rect 1821 37349 1871 37373
rect 1821 37315 1829 37349
rect 1863 37315 1871 37349
rect 1821 37291 1871 37315
rect 94179 37349 94229 37373
rect 94179 37315 94187 37349
rect 94221 37315 94229 37349
rect 94179 37291 94229 37315
rect 1821 37013 1871 37037
rect 1821 36979 1829 37013
rect 1863 36979 1871 37013
rect 1821 36955 1871 36979
rect 94179 37013 94229 37037
rect 94179 36979 94187 37013
rect 94221 36979 94229 37013
rect 94179 36955 94229 36979
rect 1821 36677 1871 36701
rect 1821 36643 1829 36677
rect 1863 36643 1871 36677
rect 1821 36619 1871 36643
rect 94179 36677 94229 36701
rect 94179 36643 94187 36677
rect 94221 36643 94229 36677
rect 94179 36619 94229 36643
rect 1821 36341 1871 36365
rect 1821 36307 1829 36341
rect 1863 36307 1871 36341
rect 1821 36283 1871 36307
rect 94179 36341 94229 36365
rect 94179 36307 94187 36341
rect 94221 36307 94229 36341
rect 94179 36283 94229 36307
rect 1821 36005 1871 36029
rect 1821 35971 1829 36005
rect 1863 35971 1871 36005
rect 1821 35947 1871 35971
rect 94179 36005 94229 36029
rect 94179 35971 94187 36005
rect 94221 35971 94229 36005
rect 94179 35947 94229 35971
rect 1821 35669 1871 35693
rect 1821 35635 1829 35669
rect 1863 35635 1871 35669
rect 1821 35611 1871 35635
rect 94179 35669 94229 35693
rect 94179 35635 94187 35669
rect 94221 35635 94229 35669
rect 94179 35611 94229 35635
rect 1821 35333 1871 35357
rect 1821 35299 1829 35333
rect 1863 35299 1871 35333
rect 1821 35275 1871 35299
rect 94179 35333 94229 35357
rect 94179 35299 94187 35333
rect 94221 35299 94229 35333
rect 94179 35275 94229 35299
rect 1821 34997 1871 35021
rect 1821 34963 1829 34997
rect 1863 34963 1871 34997
rect 1821 34939 1871 34963
rect 94179 34997 94229 35021
rect 94179 34963 94187 34997
rect 94221 34963 94229 34997
rect 94179 34939 94229 34963
rect 1821 34661 1871 34685
rect 1821 34627 1829 34661
rect 1863 34627 1871 34661
rect 1821 34603 1871 34627
rect 94179 34661 94229 34685
rect 94179 34627 94187 34661
rect 94221 34627 94229 34661
rect 94179 34603 94229 34627
rect 1821 34325 1871 34349
rect 1821 34291 1829 34325
rect 1863 34291 1871 34325
rect 1821 34267 1871 34291
rect 94179 34325 94229 34349
rect 94179 34291 94187 34325
rect 94221 34291 94229 34325
rect 94179 34267 94229 34291
rect 1821 33989 1871 34013
rect 1821 33955 1829 33989
rect 1863 33955 1871 33989
rect 1821 33931 1871 33955
rect 94179 33989 94229 34013
rect 94179 33955 94187 33989
rect 94221 33955 94229 33989
rect 94179 33931 94229 33955
rect 1821 33653 1871 33677
rect 1821 33619 1829 33653
rect 1863 33619 1871 33653
rect 1821 33595 1871 33619
rect 94179 33653 94229 33677
rect 94179 33619 94187 33653
rect 94221 33619 94229 33653
rect 94179 33595 94229 33619
rect 1821 33317 1871 33341
rect 1821 33283 1829 33317
rect 1863 33283 1871 33317
rect 1821 33259 1871 33283
rect 94179 33317 94229 33341
rect 94179 33283 94187 33317
rect 94221 33283 94229 33317
rect 94179 33259 94229 33283
rect 1821 32981 1871 33005
rect 1821 32947 1829 32981
rect 1863 32947 1871 32981
rect 1821 32923 1871 32947
rect 94179 32981 94229 33005
rect 94179 32947 94187 32981
rect 94221 32947 94229 32981
rect 94179 32923 94229 32947
rect 1821 32645 1871 32669
rect 1821 32611 1829 32645
rect 1863 32611 1871 32645
rect 1821 32587 1871 32611
rect 94179 32645 94229 32669
rect 94179 32611 94187 32645
rect 94221 32611 94229 32645
rect 94179 32587 94229 32611
rect 1821 32309 1871 32333
rect 1821 32275 1829 32309
rect 1863 32275 1871 32309
rect 1821 32251 1871 32275
rect 94179 32309 94229 32333
rect 94179 32275 94187 32309
rect 94221 32275 94229 32309
rect 94179 32251 94229 32275
rect 1821 31973 1871 31997
rect 1821 31939 1829 31973
rect 1863 31939 1871 31973
rect 1821 31915 1871 31939
rect 94179 31973 94229 31997
rect 94179 31939 94187 31973
rect 94221 31939 94229 31973
rect 94179 31915 94229 31939
rect 1821 31637 1871 31661
rect 1821 31603 1829 31637
rect 1863 31603 1871 31637
rect 1821 31579 1871 31603
rect 94179 31637 94229 31661
rect 94179 31603 94187 31637
rect 94221 31603 94229 31637
rect 94179 31579 94229 31603
rect 1821 31301 1871 31325
rect 1821 31267 1829 31301
rect 1863 31267 1871 31301
rect 1821 31243 1871 31267
rect 94179 31301 94229 31325
rect 94179 31267 94187 31301
rect 94221 31267 94229 31301
rect 94179 31243 94229 31267
rect 1821 30965 1871 30989
rect 1821 30931 1829 30965
rect 1863 30931 1871 30965
rect 1821 30907 1871 30931
rect 94179 30965 94229 30989
rect 94179 30931 94187 30965
rect 94221 30931 94229 30965
rect 94179 30907 94229 30931
rect 1821 30629 1871 30653
rect 1821 30595 1829 30629
rect 1863 30595 1871 30629
rect 1821 30571 1871 30595
rect 94179 30629 94229 30653
rect 94179 30595 94187 30629
rect 94221 30595 94229 30629
rect 94179 30571 94229 30595
rect 1821 30293 1871 30317
rect 1821 30259 1829 30293
rect 1863 30259 1871 30293
rect 1821 30235 1871 30259
rect 94179 30293 94229 30317
rect 94179 30259 94187 30293
rect 94221 30259 94229 30293
rect 94179 30235 94229 30259
rect 1821 29957 1871 29981
rect 1821 29923 1829 29957
rect 1863 29923 1871 29957
rect 1821 29899 1871 29923
rect 94179 29957 94229 29981
rect 94179 29923 94187 29957
rect 94221 29923 94229 29957
rect 94179 29899 94229 29923
rect 1821 29621 1871 29645
rect 1821 29587 1829 29621
rect 1863 29587 1871 29621
rect 1821 29563 1871 29587
rect 94179 29621 94229 29645
rect 94179 29587 94187 29621
rect 94221 29587 94229 29621
rect 94179 29563 94229 29587
rect 1821 29285 1871 29309
rect 1821 29251 1829 29285
rect 1863 29251 1871 29285
rect 1821 29227 1871 29251
rect 94179 29285 94229 29309
rect 94179 29251 94187 29285
rect 94221 29251 94229 29285
rect 94179 29227 94229 29251
rect 1821 28949 1871 28973
rect 1821 28915 1829 28949
rect 1863 28915 1871 28949
rect 1821 28891 1871 28915
rect 94179 28949 94229 28973
rect 94179 28915 94187 28949
rect 94221 28915 94229 28949
rect 94179 28891 94229 28915
rect 1821 28613 1871 28637
rect 1821 28579 1829 28613
rect 1863 28579 1871 28613
rect 1821 28555 1871 28579
rect 94179 28613 94229 28637
rect 94179 28579 94187 28613
rect 94221 28579 94229 28613
rect 94179 28555 94229 28579
rect 1821 28277 1871 28301
rect 1821 28243 1829 28277
rect 1863 28243 1871 28277
rect 1821 28219 1871 28243
rect 94179 28277 94229 28301
rect 94179 28243 94187 28277
rect 94221 28243 94229 28277
rect 94179 28219 94229 28243
rect 1821 27941 1871 27965
rect 1821 27907 1829 27941
rect 1863 27907 1871 27941
rect 1821 27883 1871 27907
rect 94179 27941 94229 27965
rect 94179 27907 94187 27941
rect 94221 27907 94229 27941
rect 94179 27883 94229 27907
rect 1821 27605 1871 27629
rect 1821 27571 1829 27605
rect 1863 27571 1871 27605
rect 1821 27547 1871 27571
rect 94179 27605 94229 27629
rect 94179 27571 94187 27605
rect 94221 27571 94229 27605
rect 94179 27547 94229 27571
rect 1821 27269 1871 27293
rect 1821 27235 1829 27269
rect 1863 27235 1871 27269
rect 1821 27211 1871 27235
rect 94179 27269 94229 27293
rect 94179 27235 94187 27269
rect 94221 27235 94229 27269
rect 94179 27211 94229 27235
rect 1821 26933 1871 26957
rect 1821 26899 1829 26933
rect 1863 26899 1871 26933
rect 1821 26875 1871 26899
rect 94179 26933 94229 26957
rect 94179 26899 94187 26933
rect 94221 26899 94229 26933
rect 94179 26875 94229 26899
rect 1821 26597 1871 26621
rect 1821 26563 1829 26597
rect 1863 26563 1871 26597
rect 1821 26539 1871 26563
rect 94179 26597 94229 26621
rect 94179 26563 94187 26597
rect 94221 26563 94229 26597
rect 94179 26539 94229 26563
rect 1821 26261 1871 26285
rect 1821 26227 1829 26261
rect 1863 26227 1871 26261
rect 1821 26203 1871 26227
rect 94179 26261 94229 26285
rect 94179 26227 94187 26261
rect 94221 26227 94229 26261
rect 94179 26203 94229 26227
rect 1821 25925 1871 25949
rect 1821 25891 1829 25925
rect 1863 25891 1871 25925
rect 1821 25867 1871 25891
rect 94179 25925 94229 25949
rect 94179 25891 94187 25925
rect 94221 25891 94229 25925
rect 94179 25867 94229 25891
rect 1821 25589 1871 25613
rect 1821 25555 1829 25589
rect 1863 25555 1871 25589
rect 1821 25531 1871 25555
rect 94179 25589 94229 25613
rect 94179 25555 94187 25589
rect 94221 25555 94229 25589
rect 94179 25531 94229 25555
rect 1821 25253 1871 25277
rect 1821 25219 1829 25253
rect 1863 25219 1871 25253
rect 1821 25195 1871 25219
rect 94179 25253 94229 25277
rect 94179 25219 94187 25253
rect 94221 25219 94229 25253
rect 94179 25195 94229 25219
rect 1821 24917 1871 24941
rect 1821 24883 1829 24917
rect 1863 24883 1871 24917
rect 1821 24859 1871 24883
rect 94179 24917 94229 24941
rect 94179 24883 94187 24917
rect 94221 24883 94229 24917
rect 94179 24859 94229 24883
rect 1821 24581 1871 24605
rect 1821 24547 1829 24581
rect 1863 24547 1871 24581
rect 1821 24523 1871 24547
rect 94179 24581 94229 24605
rect 94179 24547 94187 24581
rect 94221 24547 94229 24581
rect 94179 24523 94229 24547
rect 1821 24245 1871 24269
rect 1821 24211 1829 24245
rect 1863 24211 1871 24245
rect 1821 24187 1871 24211
rect 94179 24245 94229 24269
rect 94179 24211 94187 24245
rect 94221 24211 94229 24245
rect 94179 24187 94229 24211
rect 1821 23909 1871 23933
rect 1821 23875 1829 23909
rect 1863 23875 1871 23909
rect 1821 23851 1871 23875
rect 94179 23909 94229 23933
rect 94179 23875 94187 23909
rect 94221 23875 94229 23909
rect 94179 23851 94229 23875
rect 1821 23573 1871 23597
rect 1821 23539 1829 23573
rect 1863 23539 1871 23573
rect 1821 23515 1871 23539
rect 94179 23573 94229 23597
rect 94179 23539 94187 23573
rect 94221 23539 94229 23573
rect 94179 23515 94229 23539
rect 1821 23237 1871 23261
rect 1821 23203 1829 23237
rect 1863 23203 1871 23237
rect 1821 23179 1871 23203
rect 94179 23237 94229 23261
rect 94179 23203 94187 23237
rect 94221 23203 94229 23237
rect 94179 23179 94229 23203
rect 1821 22901 1871 22925
rect 1821 22867 1829 22901
rect 1863 22867 1871 22901
rect 1821 22843 1871 22867
rect 94179 22901 94229 22925
rect 94179 22867 94187 22901
rect 94221 22867 94229 22901
rect 94179 22843 94229 22867
rect 1821 22565 1871 22589
rect 1821 22531 1829 22565
rect 1863 22531 1871 22565
rect 1821 22507 1871 22531
rect 94179 22565 94229 22589
rect 94179 22531 94187 22565
rect 94221 22531 94229 22565
rect 94179 22507 94229 22531
rect 1821 22229 1871 22253
rect 1821 22195 1829 22229
rect 1863 22195 1871 22229
rect 1821 22171 1871 22195
rect 94179 22229 94229 22253
rect 94179 22195 94187 22229
rect 94221 22195 94229 22229
rect 94179 22171 94229 22195
rect 1821 21893 1871 21917
rect 1821 21859 1829 21893
rect 1863 21859 1871 21893
rect 1821 21835 1871 21859
rect 94179 21893 94229 21917
rect 94179 21859 94187 21893
rect 94221 21859 94229 21893
rect 94179 21835 94229 21859
rect 1821 21557 1871 21581
rect 1821 21523 1829 21557
rect 1863 21523 1871 21557
rect 1821 21499 1871 21523
rect 94179 21557 94229 21581
rect 94179 21523 94187 21557
rect 94221 21523 94229 21557
rect 94179 21499 94229 21523
rect 1821 21221 1871 21245
rect 1821 21187 1829 21221
rect 1863 21187 1871 21221
rect 1821 21163 1871 21187
rect 94179 21221 94229 21245
rect 94179 21187 94187 21221
rect 94221 21187 94229 21221
rect 94179 21163 94229 21187
rect 1821 20885 1871 20909
rect 1821 20851 1829 20885
rect 1863 20851 1871 20885
rect 1821 20827 1871 20851
rect 94179 20885 94229 20909
rect 94179 20851 94187 20885
rect 94221 20851 94229 20885
rect 94179 20827 94229 20851
rect 1821 20549 1871 20573
rect 1821 20515 1829 20549
rect 1863 20515 1871 20549
rect 1821 20491 1871 20515
rect 94179 20549 94229 20573
rect 94179 20515 94187 20549
rect 94221 20515 94229 20549
rect 94179 20491 94229 20515
rect 1821 20213 1871 20237
rect 1821 20179 1829 20213
rect 1863 20179 1871 20213
rect 1821 20155 1871 20179
rect 94179 20213 94229 20237
rect 94179 20179 94187 20213
rect 94221 20179 94229 20213
rect 94179 20155 94229 20179
rect 1821 19877 1871 19901
rect 1821 19843 1829 19877
rect 1863 19843 1871 19877
rect 1821 19819 1871 19843
rect 94179 19877 94229 19901
rect 94179 19843 94187 19877
rect 94221 19843 94229 19877
rect 94179 19819 94229 19843
rect 1821 19541 1871 19565
rect 1821 19507 1829 19541
rect 1863 19507 1871 19541
rect 1821 19483 1871 19507
rect 94179 19541 94229 19565
rect 94179 19507 94187 19541
rect 94221 19507 94229 19541
rect 94179 19483 94229 19507
rect 1821 19205 1871 19229
rect 1821 19171 1829 19205
rect 1863 19171 1871 19205
rect 1821 19147 1871 19171
rect 94179 19205 94229 19229
rect 94179 19171 94187 19205
rect 94221 19171 94229 19205
rect 94179 19147 94229 19171
rect 1821 18869 1871 18893
rect 1821 18835 1829 18869
rect 1863 18835 1871 18869
rect 1821 18811 1871 18835
rect 94179 18869 94229 18893
rect 94179 18835 94187 18869
rect 94221 18835 94229 18869
rect 94179 18811 94229 18835
rect 1821 18533 1871 18557
rect 1821 18499 1829 18533
rect 1863 18499 1871 18533
rect 1821 18475 1871 18499
rect 94179 18533 94229 18557
rect 94179 18499 94187 18533
rect 94221 18499 94229 18533
rect 94179 18475 94229 18499
rect 1821 18197 1871 18221
rect 1821 18163 1829 18197
rect 1863 18163 1871 18197
rect 1821 18139 1871 18163
rect 94179 18197 94229 18221
rect 94179 18163 94187 18197
rect 94221 18163 94229 18197
rect 94179 18139 94229 18163
rect 1821 17861 1871 17885
rect 1821 17827 1829 17861
rect 1863 17827 1871 17861
rect 1821 17803 1871 17827
rect 94179 17861 94229 17885
rect 94179 17827 94187 17861
rect 94221 17827 94229 17861
rect 94179 17803 94229 17827
rect 1821 17525 1871 17549
rect 1821 17491 1829 17525
rect 1863 17491 1871 17525
rect 1821 17467 1871 17491
rect 94179 17525 94229 17549
rect 94179 17491 94187 17525
rect 94221 17491 94229 17525
rect 94179 17467 94229 17491
rect 1821 17189 1871 17213
rect 1821 17155 1829 17189
rect 1863 17155 1871 17189
rect 1821 17131 1871 17155
rect 94179 17189 94229 17213
rect 94179 17155 94187 17189
rect 94221 17155 94229 17189
rect 94179 17131 94229 17155
rect 1821 16853 1871 16877
rect 1821 16819 1829 16853
rect 1863 16819 1871 16853
rect 1821 16795 1871 16819
rect 94179 16853 94229 16877
rect 94179 16819 94187 16853
rect 94221 16819 94229 16853
rect 94179 16795 94229 16819
rect 1821 16517 1871 16541
rect 1821 16483 1829 16517
rect 1863 16483 1871 16517
rect 1821 16459 1871 16483
rect 94179 16517 94229 16541
rect 94179 16483 94187 16517
rect 94221 16483 94229 16517
rect 94179 16459 94229 16483
rect 1821 16181 1871 16205
rect 1821 16147 1829 16181
rect 1863 16147 1871 16181
rect 1821 16123 1871 16147
rect 94179 16181 94229 16205
rect 94179 16147 94187 16181
rect 94221 16147 94229 16181
rect 94179 16123 94229 16147
rect 1821 15845 1871 15869
rect 1821 15811 1829 15845
rect 1863 15811 1871 15845
rect 1821 15787 1871 15811
rect 94179 15845 94229 15869
rect 94179 15811 94187 15845
rect 94221 15811 94229 15845
rect 94179 15787 94229 15811
rect 1821 15509 1871 15533
rect 1821 15475 1829 15509
rect 1863 15475 1871 15509
rect 1821 15451 1871 15475
rect 94179 15509 94229 15533
rect 94179 15475 94187 15509
rect 94221 15475 94229 15509
rect 94179 15451 94229 15475
rect 1821 15173 1871 15197
rect 1821 15139 1829 15173
rect 1863 15139 1871 15173
rect 1821 15115 1871 15139
rect 94179 15173 94229 15197
rect 94179 15139 94187 15173
rect 94221 15139 94229 15173
rect 94179 15115 94229 15139
rect 1821 14837 1871 14861
rect 1821 14803 1829 14837
rect 1863 14803 1871 14837
rect 1821 14779 1871 14803
rect 94179 14837 94229 14861
rect 94179 14803 94187 14837
rect 94221 14803 94229 14837
rect 94179 14779 94229 14803
rect 1821 14501 1871 14525
rect 1821 14467 1829 14501
rect 1863 14467 1871 14501
rect 1821 14443 1871 14467
rect 94179 14501 94229 14525
rect 94179 14467 94187 14501
rect 94221 14467 94229 14501
rect 94179 14443 94229 14467
rect 1821 14165 1871 14189
rect 1821 14131 1829 14165
rect 1863 14131 1871 14165
rect 1821 14107 1871 14131
rect 94179 14165 94229 14189
rect 94179 14131 94187 14165
rect 94221 14131 94229 14165
rect 94179 14107 94229 14131
rect 1821 13829 1871 13853
rect 1821 13795 1829 13829
rect 1863 13795 1871 13829
rect 1821 13771 1871 13795
rect 94179 13829 94229 13853
rect 94179 13795 94187 13829
rect 94221 13795 94229 13829
rect 94179 13771 94229 13795
rect 1821 13493 1871 13517
rect 1821 13459 1829 13493
rect 1863 13459 1871 13493
rect 1821 13435 1871 13459
rect 94179 13493 94229 13517
rect 94179 13459 94187 13493
rect 94221 13459 94229 13493
rect 94179 13435 94229 13459
rect 1821 13157 1871 13181
rect 1821 13123 1829 13157
rect 1863 13123 1871 13157
rect 1821 13099 1871 13123
rect 94179 13157 94229 13181
rect 94179 13123 94187 13157
rect 94221 13123 94229 13157
rect 94179 13099 94229 13123
rect 1821 12821 1871 12845
rect 1821 12787 1829 12821
rect 1863 12787 1871 12821
rect 1821 12763 1871 12787
rect 94179 12821 94229 12845
rect 94179 12787 94187 12821
rect 94221 12787 94229 12821
rect 94179 12763 94229 12787
rect 1821 12485 1871 12509
rect 1821 12451 1829 12485
rect 1863 12451 1871 12485
rect 1821 12427 1871 12451
rect 94179 12485 94229 12509
rect 94179 12451 94187 12485
rect 94221 12451 94229 12485
rect 94179 12427 94229 12451
rect 1821 12149 1871 12173
rect 1821 12115 1829 12149
rect 1863 12115 1871 12149
rect 1821 12091 1871 12115
rect 94179 12149 94229 12173
rect 94179 12115 94187 12149
rect 94221 12115 94229 12149
rect 94179 12091 94229 12115
rect 1821 11813 1871 11837
rect 1821 11779 1829 11813
rect 1863 11779 1871 11813
rect 1821 11755 1871 11779
rect 94179 11813 94229 11837
rect 94179 11779 94187 11813
rect 94221 11779 94229 11813
rect 94179 11755 94229 11779
rect 1821 11477 1871 11501
rect 1821 11443 1829 11477
rect 1863 11443 1871 11477
rect 1821 11419 1871 11443
rect 94179 11477 94229 11501
rect 94179 11443 94187 11477
rect 94221 11443 94229 11477
rect 94179 11419 94229 11443
rect 1821 11141 1871 11165
rect 1821 11107 1829 11141
rect 1863 11107 1871 11141
rect 1821 11083 1871 11107
rect 94179 11141 94229 11165
rect 94179 11107 94187 11141
rect 94221 11107 94229 11141
rect 94179 11083 94229 11107
rect 1821 10805 1871 10829
rect 1821 10771 1829 10805
rect 1863 10771 1871 10805
rect 1821 10747 1871 10771
rect 94179 10805 94229 10829
rect 94179 10771 94187 10805
rect 94221 10771 94229 10805
rect 94179 10747 94229 10771
rect 1821 10469 1871 10493
rect 1821 10435 1829 10469
rect 1863 10435 1871 10469
rect 1821 10411 1871 10435
rect 94179 10469 94229 10493
rect 94179 10435 94187 10469
rect 94221 10435 94229 10469
rect 94179 10411 94229 10435
rect 1821 10133 1871 10157
rect 1821 10099 1829 10133
rect 1863 10099 1871 10133
rect 1821 10075 1871 10099
rect 94179 10133 94229 10157
rect 94179 10099 94187 10133
rect 94221 10099 94229 10133
rect 94179 10075 94229 10099
rect 1821 9797 1871 9821
rect 1821 9763 1829 9797
rect 1863 9763 1871 9797
rect 1821 9739 1871 9763
rect 94179 9797 94229 9821
rect 94179 9763 94187 9797
rect 94221 9763 94229 9797
rect 94179 9739 94229 9763
rect 1821 9461 1871 9485
rect 1821 9427 1829 9461
rect 1863 9427 1871 9461
rect 1821 9403 1871 9427
rect 94179 9461 94229 9485
rect 94179 9427 94187 9461
rect 94221 9427 94229 9461
rect 94179 9403 94229 9427
rect 1821 9125 1871 9149
rect 1821 9091 1829 9125
rect 1863 9091 1871 9125
rect 1821 9067 1871 9091
rect 94179 9125 94229 9149
rect 94179 9091 94187 9125
rect 94221 9091 94229 9125
rect 94179 9067 94229 9091
rect 1821 8789 1871 8813
rect 1821 8755 1829 8789
rect 1863 8755 1871 8789
rect 1821 8731 1871 8755
rect 94179 8789 94229 8813
rect 94179 8755 94187 8789
rect 94221 8755 94229 8789
rect 94179 8731 94229 8755
rect 1821 8453 1871 8477
rect 1821 8419 1829 8453
rect 1863 8419 1871 8453
rect 1821 8395 1871 8419
rect 94179 8453 94229 8477
rect 94179 8419 94187 8453
rect 94221 8419 94229 8453
rect 94179 8395 94229 8419
rect 1821 8117 1871 8141
rect 1821 8083 1829 8117
rect 1863 8083 1871 8117
rect 1821 8059 1871 8083
rect 94179 8117 94229 8141
rect 94179 8083 94187 8117
rect 94221 8083 94229 8117
rect 94179 8059 94229 8083
rect 1821 7781 1871 7805
rect 1821 7747 1829 7781
rect 1863 7747 1871 7781
rect 1821 7723 1871 7747
rect 94179 7781 94229 7805
rect 94179 7747 94187 7781
rect 94221 7747 94229 7781
rect 94179 7723 94229 7747
rect 1821 7445 1871 7469
rect 1821 7411 1829 7445
rect 1863 7411 1871 7445
rect 1821 7387 1871 7411
rect 94179 7445 94229 7469
rect 94179 7411 94187 7445
rect 94221 7411 94229 7445
rect 94179 7387 94229 7411
rect 1821 7109 1871 7133
rect 1821 7075 1829 7109
rect 1863 7075 1871 7109
rect 1821 7051 1871 7075
rect 94179 7109 94229 7133
rect 94179 7075 94187 7109
rect 94221 7075 94229 7109
rect 94179 7051 94229 7075
rect 1821 6773 1871 6797
rect 1821 6739 1829 6773
rect 1863 6739 1871 6773
rect 1821 6715 1871 6739
rect 94179 6773 94229 6797
rect 94179 6739 94187 6773
rect 94221 6739 94229 6773
rect 94179 6715 94229 6739
rect 1821 6437 1871 6461
rect 1821 6403 1829 6437
rect 1863 6403 1871 6437
rect 1821 6379 1871 6403
rect 94179 6437 94229 6461
rect 94179 6403 94187 6437
rect 94221 6403 94229 6437
rect 94179 6379 94229 6403
rect 1821 6101 1871 6125
rect 1821 6067 1829 6101
rect 1863 6067 1871 6101
rect 1821 6043 1871 6067
rect 94179 6101 94229 6125
rect 94179 6067 94187 6101
rect 94221 6067 94229 6101
rect 94179 6043 94229 6067
rect 1821 5765 1871 5789
rect 1821 5731 1829 5765
rect 1863 5731 1871 5765
rect 1821 5707 1871 5731
rect 94179 5765 94229 5789
rect 94179 5731 94187 5765
rect 94221 5731 94229 5765
rect 94179 5707 94229 5731
rect 1821 5429 1871 5453
rect 1821 5395 1829 5429
rect 1863 5395 1871 5429
rect 1821 5371 1871 5395
rect 94179 5429 94229 5453
rect 94179 5395 94187 5429
rect 94221 5395 94229 5429
rect 94179 5371 94229 5395
rect 1821 5093 1871 5117
rect 1821 5059 1829 5093
rect 1863 5059 1871 5093
rect 1821 5035 1871 5059
rect 94179 5093 94229 5117
rect 94179 5059 94187 5093
rect 94221 5059 94229 5093
rect 94179 5035 94229 5059
rect 1821 4757 1871 4781
rect 1821 4723 1829 4757
rect 1863 4723 1871 4757
rect 1821 4699 1871 4723
rect 94179 4757 94229 4781
rect 94179 4723 94187 4757
rect 94221 4723 94229 4757
rect 94179 4699 94229 4723
rect 1821 4421 1871 4445
rect 1821 4387 1829 4421
rect 1863 4387 1871 4421
rect 1821 4363 1871 4387
rect 94179 4421 94229 4445
rect 94179 4387 94187 4421
rect 94221 4387 94229 4421
rect 94179 4363 94229 4387
rect 1821 4085 1871 4109
rect 1821 4051 1829 4085
rect 1863 4051 1871 4085
rect 1821 4027 1871 4051
rect 94179 4085 94229 4109
rect 94179 4051 94187 4085
rect 94221 4051 94229 4085
rect 94179 4027 94229 4051
rect 1821 3749 1871 3773
rect 1821 3715 1829 3749
rect 1863 3715 1871 3749
rect 1821 3691 1871 3715
rect 94179 3749 94229 3773
rect 94179 3715 94187 3749
rect 94221 3715 94229 3749
rect 94179 3691 94229 3715
rect 1821 3413 1871 3437
rect 1821 3379 1829 3413
rect 1863 3379 1871 3413
rect 1821 3355 1871 3379
rect 94179 3413 94229 3437
rect 94179 3379 94187 3413
rect 94221 3379 94229 3413
rect 94179 3355 94229 3379
rect 1821 3077 1871 3101
rect 1821 3043 1829 3077
rect 1863 3043 1871 3077
rect 1821 3019 1871 3043
rect 94179 3077 94229 3101
rect 94179 3043 94187 3077
rect 94221 3043 94229 3077
rect 94179 3019 94229 3043
rect 1821 2741 1871 2765
rect 1821 2707 1829 2741
rect 1863 2707 1871 2741
rect 1821 2683 1871 2707
rect 94179 2741 94229 2765
rect 94179 2707 94187 2741
rect 94221 2707 94229 2741
rect 94179 2683 94229 2707
rect 1821 2405 1871 2429
rect 1821 2371 1829 2405
rect 1863 2371 1871 2405
rect 1821 2347 1871 2371
rect 94179 2405 94229 2429
rect 94179 2371 94187 2405
rect 94221 2371 94229 2405
rect 94179 2347 94229 2371
rect 1821 2069 1871 2093
rect 1821 2035 1829 2069
rect 1863 2035 1871 2069
rect 1821 2011 1871 2035
rect 94179 2069 94229 2093
rect 94179 2035 94187 2069
rect 94221 2035 94229 2069
rect 94179 2011 94229 2035
rect 2157 1733 2207 1757
rect 2157 1699 2165 1733
rect 2199 1699 2207 1733
rect 2157 1675 2207 1699
rect 2493 1733 2543 1757
rect 2493 1699 2501 1733
rect 2535 1699 2543 1733
rect 2493 1675 2543 1699
rect 2829 1733 2879 1757
rect 2829 1699 2837 1733
rect 2871 1699 2879 1733
rect 2829 1675 2879 1699
rect 3165 1733 3215 1757
rect 3165 1699 3173 1733
rect 3207 1699 3215 1733
rect 3165 1675 3215 1699
rect 3501 1733 3551 1757
rect 3501 1699 3509 1733
rect 3543 1699 3551 1733
rect 3501 1675 3551 1699
rect 3837 1733 3887 1757
rect 3837 1699 3845 1733
rect 3879 1699 3887 1733
rect 3837 1675 3887 1699
rect 4173 1733 4223 1757
rect 4173 1699 4181 1733
rect 4215 1699 4223 1733
rect 4173 1675 4223 1699
rect 4509 1733 4559 1757
rect 4509 1699 4517 1733
rect 4551 1699 4559 1733
rect 4509 1675 4559 1699
rect 4845 1733 4895 1757
rect 4845 1699 4853 1733
rect 4887 1699 4895 1733
rect 4845 1675 4895 1699
rect 5181 1733 5231 1757
rect 5181 1699 5189 1733
rect 5223 1699 5231 1733
rect 5181 1675 5231 1699
rect 5517 1733 5567 1757
rect 5517 1699 5525 1733
rect 5559 1699 5567 1733
rect 5517 1675 5567 1699
rect 5853 1733 5903 1757
rect 5853 1699 5861 1733
rect 5895 1699 5903 1733
rect 5853 1675 5903 1699
rect 6189 1733 6239 1757
rect 6189 1699 6197 1733
rect 6231 1699 6239 1733
rect 6189 1675 6239 1699
rect 6525 1733 6575 1757
rect 6525 1699 6533 1733
rect 6567 1699 6575 1733
rect 6525 1675 6575 1699
rect 6861 1733 6911 1757
rect 6861 1699 6869 1733
rect 6903 1699 6911 1733
rect 6861 1675 6911 1699
rect 7197 1733 7247 1757
rect 7197 1699 7205 1733
rect 7239 1699 7247 1733
rect 7197 1675 7247 1699
rect 7533 1733 7583 1757
rect 7533 1699 7541 1733
rect 7575 1699 7583 1733
rect 7533 1675 7583 1699
rect 7869 1733 7919 1757
rect 7869 1699 7877 1733
rect 7911 1699 7919 1733
rect 7869 1675 7919 1699
rect 8205 1733 8255 1757
rect 8205 1699 8213 1733
rect 8247 1699 8255 1733
rect 8205 1675 8255 1699
rect 8541 1733 8591 1757
rect 8541 1699 8549 1733
rect 8583 1699 8591 1733
rect 8541 1675 8591 1699
rect 8877 1733 8927 1757
rect 8877 1699 8885 1733
rect 8919 1699 8927 1733
rect 8877 1675 8927 1699
rect 9213 1733 9263 1757
rect 9213 1699 9221 1733
rect 9255 1699 9263 1733
rect 9213 1675 9263 1699
rect 9549 1733 9599 1757
rect 9549 1699 9557 1733
rect 9591 1699 9599 1733
rect 9549 1675 9599 1699
rect 9885 1733 9935 1757
rect 9885 1699 9893 1733
rect 9927 1699 9935 1733
rect 9885 1675 9935 1699
rect 10221 1733 10271 1757
rect 10221 1699 10229 1733
rect 10263 1699 10271 1733
rect 10221 1675 10271 1699
rect 10557 1733 10607 1757
rect 10557 1699 10565 1733
rect 10599 1699 10607 1733
rect 10557 1675 10607 1699
rect 10893 1733 10943 1757
rect 10893 1699 10901 1733
rect 10935 1699 10943 1733
rect 10893 1675 10943 1699
rect 11229 1733 11279 1757
rect 11229 1699 11237 1733
rect 11271 1699 11279 1733
rect 11229 1675 11279 1699
rect 11565 1733 11615 1757
rect 11565 1699 11573 1733
rect 11607 1699 11615 1733
rect 11565 1675 11615 1699
rect 11901 1733 11951 1757
rect 11901 1699 11909 1733
rect 11943 1699 11951 1733
rect 11901 1675 11951 1699
rect 12237 1733 12287 1757
rect 12237 1699 12245 1733
rect 12279 1699 12287 1733
rect 12237 1675 12287 1699
rect 12573 1733 12623 1757
rect 12573 1699 12581 1733
rect 12615 1699 12623 1733
rect 12573 1675 12623 1699
rect 12909 1733 12959 1757
rect 12909 1699 12917 1733
rect 12951 1699 12959 1733
rect 12909 1675 12959 1699
rect 13245 1733 13295 1757
rect 13245 1699 13253 1733
rect 13287 1699 13295 1733
rect 13245 1675 13295 1699
rect 13581 1733 13631 1757
rect 13581 1699 13589 1733
rect 13623 1699 13631 1733
rect 13581 1675 13631 1699
rect 13917 1733 13967 1757
rect 13917 1699 13925 1733
rect 13959 1699 13967 1733
rect 13917 1675 13967 1699
rect 14253 1733 14303 1757
rect 14253 1699 14261 1733
rect 14295 1699 14303 1733
rect 14253 1675 14303 1699
rect 14589 1733 14639 1757
rect 14589 1699 14597 1733
rect 14631 1699 14639 1733
rect 14589 1675 14639 1699
rect 14925 1733 14975 1757
rect 14925 1699 14933 1733
rect 14967 1699 14975 1733
rect 14925 1675 14975 1699
rect 15261 1733 15311 1757
rect 15261 1699 15269 1733
rect 15303 1699 15311 1733
rect 15261 1675 15311 1699
rect 15597 1733 15647 1757
rect 15597 1699 15605 1733
rect 15639 1699 15647 1733
rect 15597 1675 15647 1699
rect 15933 1733 15983 1757
rect 15933 1699 15941 1733
rect 15975 1699 15983 1733
rect 15933 1675 15983 1699
rect 16269 1733 16319 1757
rect 16269 1699 16277 1733
rect 16311 1699 16319 1733
rect 16269 1675 16319 1699
rect 16605 1733 16655 1757
rect 16605 1699 16613 1733
rect 16647 1699 16655 1733
rect 16605 1675 16655 1699
rect 16941 1733 16991 1757
rect 16941 1699 16949 1733
rect 16983 1699 16991 1733
rect 16941 1675 16991 1699
rect 17277 1733 17327 1757
rect 17277 1699 17285 1733
rect 17319 1699 17327 1733
rect 17277 1675 17327 1699
rect 17613 1733 17663 1757
rect 17613 1699 17621 1733
rect 17655 1699 17663 1733
rect 17613 1675 17663 1699
rect 17949 1733 17999 1757
rect 17949 1699 17957 1733
rect 17991 1699 17999 1733
rect 17949 1675 17999 1699
rect 18285 1733 18335 1757
rect 18285 1699 18293 1733
rect 18327 1699 18335 1733
rect 18285 1675 18335 1699
rect 18621 1733 18671 1757
rect 18621 1699 18629 1733
rect 18663 1699 18671 1733
rect 18621 1675 18671 1699
rect 18957 1733 19007 1757
rect 18957 1699 18965 1733
rect 18999 1699 19007 1733
rect 18957 1675 19007 1699
rect 19293 1733 19343 1757
rect 19293 1699 19301 1733
rect 19335 1699 19343 1733
rect 19293 1675 19343 1699
rect 19629 1733 19679 1757
rect 19629 1699 19637 1733
rect 19671 1699 19679 1733
rect 19629 1675 19679 1699
rect 19965 1733 20015 1757
rect 19965 1699 19973 1733
rect 20007 1699 20015 1733
rect 19965 1675 20015 1699
rect 20301 1733 20351 1757
rect 20301 1699 20309 1733
rect 20343 1699 20351 1733
rect 20301 1675 20351 1699
rect 20637 1733 20687 1757
rect 20637 1699 20645 1733
rect 20679 1699 20687 1733
rect 20637 1675 20687 1699
rect 20973 1733 21023 1757
rect 20973 1699 20981 1733
rect 21015 1699 21023 1733
rect 20973 1675 21023 1699
rect 21309 1733 21359 1757
rect 21309 1699 21317 1733
rect 21351 1699 21359 1733
rect 21309 1675 21359 1699
rect 21645 1733 21695 1757
rect 21645 1699 21653 1733
rect 21687 1699 21695 1733
rect 21645 1675 21695 1699
rect 21981 1733 22031 1757
rect 21981 1699 21989 1733
rect 22023 1699 22031 1733
rect 21981 1675 22031 1699
rect 22317 1733 22367 1757
rect 22317 1699 22325 1733
rect 22359 1699 22367 1733
rect 22317 1675 22367 1699
rect 22653 1733 22703 1757
rect 22653 1699 22661 1733
rect 22695 1699 22703 1733
rect 22653 1675 22703 1699
rect 22989 1733 23039 1757
rect 22989 1699 22997 1733
rect 23031 1699 23039 1733
rect 22989 1675 23039 1699
rect 23325 1733 23375 1757
rect 23325 1699 23333 1733
rect 23367 1699 23375 1733
rect 23325 1675 23375 1699
rect 23661 1733 23711 1757
rect 23661 1699 23669 1733
rect 23703 1699 23711 1733
rect 23661 1675 23711 1699
rect 23997 1733 24047 1757
rect 23997 1699 24005 1733
rect 24039 1699 24047 1733
rect 23997 1675 24047 1699
rect 24333 1733 24383 1757
rect 24333 1699 24341 1733
rect 24375 1699 24383 1733
rect 24333 1675 24383 1699
rect 24669 1733 24719 1757
rect 24669 1699 24677 1733
rect 24711 1699 24719 1733
rect 24669 1675 24719 1699
rect 25005 1733 25055 1757
rect 25005 1699 25013 1733
rect 25047 1699 25055 1733
rect 25005 1675 25055 1699
rect 25341 1733 25391 1757
rect 25341 1699 25349 1733
rect 25383 1699 25391 1733
rect 25341 1675 25391 1699
rect 25677 1733 25727 1757
rect 25677 1699 25685 1733
rect 25719 1699 25727 1733
rect 25677 1675 25727 1699
rect 26013 1733 26063 1757
rect 26013 1699 26021 1733
rect 26055 1699 26063 1733
rect 26013 1675 26063 1699
rect 26349 1733 26399 1757
rect 26349 1699 26357 1733
rect 26391 1699 26399 1733
rect 26349 1675 26399 1699
rect 26685 1733 26735 1757
rect 26685 1699 26693 1733
rect 26727 1699 26735 1733
rect 26685 1675 26735 1699
rect 27021 1733 27071 1757
rect 27021 1699 27029 1733
rect 27063 1699 27071 1733
rect 27021 1675 27071 1699
rect 27357 1733 27407 1757
rect 27357 1699 27365 1733
rect 27399 1699 27407 1733
rect 27357 1675 27407 1699
rect 27693 1733 27743 1757
rect 27693 1699 27701 1733
rect 27735 1699 27743 1733
rect 27693 1675 27743 1699
rect 28029 1733 28079 1757
rect 28029 1699 28037 1733
rect 28071 1699 28079 1733
rect 28029 1675 28079 1699
rect 28365 1733 28415 1757
rect 28365 1699 28373 1733
rect 28407 1699 28415 1733
rect 28365 1675 28415 1699
rect 28701 1733 28751 1757
rect 28701 1699 28709 1733
rect 28743 1699 28751 1733
rect 28701 1675 28751 1699
rect 29037 1733 29087 1757
rect 29037 1699 29045 1733
rect 29079 1699 29087 1733
rect 29037 1675 29087 1699
rect 29373 1733 29423 1757
rect 29373 1699 29381 1733
rect 29415 1699 29423 1733
rect 29373 1675 29423 1699
rect 29709 1733 29759 1757
rect 29709 1699 29717 1733
rect 29751 1699 29759 1733
rect 29709 1675 29759 1699
rect 30045 1733 30095 1757
rect 30045 1699 30053 1733
rect 30087 1699 30095 1733
rect 30045 1675 30095 1699
rect 30381 1733 30431 1757
rect 30381 1699 30389 1733
rect 30423 1699 30431 1733
rect 30381 1675 30431 1699
rect 30717 1733 30767 1757
rect 30717 1699 30725 1733
rect 30759 1699 30767 1733
rect 30717 1675 30767 1699
rect 31053 1733 31103 1757
rect 31053 1699 31061 1733
rect 31095 1699 31103 1733
rect 31053 1675 31103 1699
rect 31389 1733 31439 1757
rect 31389 1699 31397 1733
rect 31431 1699 31439 1733
rect 31389 1675 31439 1699
rect 31725 1733 31775 1757
rect 31725 1699 31733 1733
rect 31767 1699 31775 1733
rect 31725 1675 31775 1699
rect 32061 1733 32111 1757
rect 32061 1699 32069 1733
rect 32103 1699 32111 1733
rect 32061 1675 32111 1699
rect 32397 1733 32447 1757
rect 32397 1699 32405 1733
rect 32439 1699 32447 1733
rect 32397 1675 32447 1699
rect 32733 1733 32783 1757
rect 32733 1699 32741 1733
rect 32775 1699 32783 1733
rect 32733 1675 32783 1699
rect 33069 1733 33119 1757
rect 33069 1699 33077 1733
rect 33111 1699 33119 1733
rect 33069 1675 33119 1699
rect 33405 1733 33455 1757
rect 33405 1699 33413 1733
rect 33447 1699 33455 1733
rect 33405 1675 33455 1699
rect 33741 1733 33791 1757
rect 33741 1699 33749 1733
rect 33783 1699 33791 1733
rect 33741 1675 33791 1699
rect 34077 1733 34127 1757
rect 34077 1699 34085 1733
rect 34119 1699 34127 1733
rect 34077 1675 34127 1699
rect 34413 1733 34463 1757
rect 34413 1699 34421 1733
rect 34455 1699 34463 1733
rect 34413 1675 34463 1699
rect 34749 1733 34799 1757
rect 34749 1699 34757 1733
rect 34791 1699 34799 1733
rect 34749 1675 34799 1699
rect 35085 1733 35135 1757
rect 35085 1699 35093 1733
rect 35127 1699 35135 1733
rect 35085 1675 35135 1699
rect 35421 1733 35471 1757
rect 35421 1699 35429 1733
rect 35463 1699 35471 1733
rect 35421 1675 35471 1699
rect 35757 1733 35807 1757
rect 35757 1699 35765 1733
rect 35799 1699 35807 1733
rect 35757 1675 35807 1699
rect 36093 1733 36143 1757
rect 36093 1699 36101 1733
rect 36135 1699 36143 1733
rect 36093 1675 36143 1699
rect 36429 1733 36479 1757
rect 36429 1699 36437 1733
rect 36471 1699 36479 1733
rect 36429 1675 36479 1699
rect 36765 1733 36815 1757
rect 36765 1699 36773 1733
rect 36807 1699 36815 1733
rect 36765 1675 36815 1699
rect 37101 1733 37151 1757
rect 37101 1699 37109 1733
rect 37143 1699 37151 1733
rect 37101 1675 37151 1699
rect 37437 1733 37487 1757
rect 37437 1699 37445 1733
rect 37479 1699 37487 1733
rect 37437 1675 37487 1699
rect 37773 1733 37823 1757
rect 37773 1699 37781 1733
rect 37815 1699 37823 1733
rect 37773 1675 37823 1699
rect 38109 1733 38159 1757
rect 38109 1699 38117 1733
rect 38151 1699 38159 1733
rect 38109 1675 38159 1699
rect 38445 1733 38495 1757
rect 38445 1699 38453 1733
rect 38487 1699 38495 1733
rect 38445 1675 38495 1699
rect 38781 1733 38831 1757
rect 38781 1699 38789 1733
rect 38823 1699 38831 1733
rect 38781 1675 38831 1699
rect 39117 1733 39167 1757
rect 39117 1699 39125 1733
rect 39159 1699 39167 1733
rect 39117 1675 39167 1699
rect 39453 1733 39503 1757
rect 39453 1699 39461 1733
rect 39495 1699 39503 1733
rect 39453 1675 39503 1699
rect 39789 1733 39839 1757
rect 39789 1699 39797 1733
rect 39831 1699 39839 1733
rect 39789 1675 39839 1699
rect 40125 1733 40175 1757
rect 40125 1699 40133 1733
rect 40167 1699 40175 1733
rect 40125 1675 40175 1699
rect 40461 1733 40511 1757
rect 40461 1699 40469 1733
rect 40503 1699 40511 1733
rect 40461 1675 40511 1699
rect 40797 1733 40847 1757
rect 40797 1699 40805 1733
rect 40839 1699 40847 1733
rect 40797 1675 40847 1699
rect 41133 1733 41183 1757
rect 41133 1699 41141 1733
rect 41175 1699 41183 1733
rect 41133 1675 41183 1699
rect 41469 1733 41519 1757
rect 41469 1699 41477 1733
rect 41511 1699 41519 1733
rect 41469 1675 41519 1699
rect 41805 1733 41855 1757
rect 41805 1699 41813 1733
rect 41847 1699 41855 1733
rect 41805 1675 41855 1699
rect 42141 1733 42191 1757
rect 42141 1699 42149 1733
rect 42183 1699 42191 1733
rect 42141 1675 42191 1699
rect 42477 1733 42527 1757
rect 42477 1699 42485 1733
rect 42519 1699 42527 1733
rect 42477 1675 42527 1699
rect 42813 1733 42863 1757
rect 42813 1699 42821 1733
rect 42855 1699 42863 1733
rect 42813 1675 42863 1699
rect 43149 1733 43199 1757
rect 43149 1699 43157 1733
rect 43191 1699 43199 1733
rect 43149 1675 43199 1699
rect 43485 1733 43535 1757
rect 43485 1699 43493 1733
rect 43527 1699 43535 1733
rect 43485 1675 43535 1699
rect 43821 1733 43871 1757
rect 43821 1699 43829 1733
rect 43863 1699 43871 1733
rect 43821 1675 43871 1699
rect 44157 1733 44207 1757
rect 44157 1699 44165 1733
rect 44199 1699 44207 1733
rect 44157 1675 44207 1699
rect 44493 1733 44543 1757
rect 44493 1699 44501 1733
rect 44535 1699 44543 1733
rect 44493 1675 44543 1699
rect 44829 1733 44879 1757
rect 44829 1699 44837 1733
rect 44871 1699 44879 1733
rect 44829 1675 44879 1699
rect 45165 1733 45215 1757
rect 45165 1699 45173 1733
rect 45207 1699 45215 1733
rect 45165 1675 45215 1699
rect 45501 1733 45551 1757
rect 45501 1699 45509 1733
rect 45543 1699 45551 1733
rect 45501 1675 45551 1699
rect 45837 1733 45887 1757
rect 45837 1699 45845 1733
rect 45879 1699 45887 1733
rect 45837 1675 45887 1699
rect 46173 1733 46223 1757
rect 46173 1699 46181 1733
rect 46215 1699 46223 1733
rect 46173 1675 46223 1699
rect 46509 1733 46559 1757
rect 46509 1699 46517 1733
rect 46551 1699 46559 1733
rect 46509 1675 46559 1699
rect 46845 1733 46895 1757
rect 46845 1699 46853 1733
rect 46887 1699 46895 1733
rect 46845 1675 46895 1699
rect 47181 1733 47231 1757
rect 47181 1699 47189 1733
rect 47223 1699 47231 1733
rect 47181 1675 47231 1699
rect 47517 1733 47567 1757
rect 47517 1699 47525 1733
rect 47559 1699 47567 1733
rect 47517 1675 47567 1699
rect 47853 1733 47903 1757
rect 47853 1699 47861 1733
rect 47895 1699 47903 1733
rect 47853 1675 47903 1699
rect 48189 1733 48239 1757
rect 48189 1699 48197 1733
rect 48231 1699 48239 1733
rect 48189 1675 48239 1699
rect 48525 1733 48575 1757
rect 48525 1699 48533 1733
rect 48567 1699 48575 1733
rect 48525 1675 48575 1699
rect 48861 1733 48911 1757
rect 48861 1699 48869 1733
rect 48903 1699 48911 1733
rect 48861 1675 48911 1699
rect 49197 1733 49247 1757
rect 49197 1699 49205 1733
rect 49239 1699 49247 1733
rect 49197 1675 49247 1699
rect 49533 1733 49583 1757
rect 49533 1699 49541 1733
rect 49575 1699 49583 1733
rect 49533 1675 49583 1699
rect 49869 1733 49919 1757
rect 49869 1699 49877 1733
rect 49911 1699 49919 1733
rect 49869 1675 49919 1699
rect 50205 1733 50255 1757
rect 50205 1699 50213 1733
rect 50247 1699 50255 1733
rect 50205 1675 50255 1699
rect 50541 1733 50591 1757
rect 50541 1699 50549 1733
rect 50583 1699 50591 1733
rect 50541 1675 50591 1699
rect 50877 1733 50927 1757
rect 50877 1699 50885 1733
rect 50919 1699 50927 1733
rect 50877 1675 50927 1699
rect 51213 1733 51263 1757
rect 51213 1699 51221 1733
rect 51255 1699 51263 1733
rect 51213 1675 51263 1699
rect 51549 1733 51599 1757
rect 51549 1699 51557 1733
rect 51591 1699 51599 1733
rect 51549 1675 51599 1699
rect 51885 1733 51935 1757
rect 51885 1699 51893 1733
rect 51927 1699 51935 1733
rect 51885 1675 51935 1699
rect 52221 1733 52271 1757
rect 52221 1699 52229 1733
rect 52263 1699 52271 1733
rect 52221 1675 52271 1699
rect 52557 1733 52607 1757
rect 52557 1699 52565 1733
rect 52599 1699 52607 1733
rect 52557 1675 52607 1699
rect 52893 1733 52943 1757
rect 52893 1699 52901 1733
rect 52935 1699 52943 1733
rect 52893 1675 52943 1699
rect 53229 1733 53279 1757
rect 53229 1699 53237 1733
rect 53271 1699 53279 1733
rect 53229 1675 53279 1699
rect 53565 1733 53615 1757
rect 53565 1699 53573 1733
rect 53607 1699 53615 1733
rect 53565 1675 53615 1699
rect 53901 1733 53951 1757
rect 53901 1699 53909 1733
rect 53943 1699 53951 1733
rect 53901 1675 53951 1699
rect 54237 1733 54287 1757
rect 54237 1699 54245 1733
rect 54279 1699 54287 1733
rect 54237 1675 54287 1699
rect 54573 1733 54623 1757
rect 54573 1699 54581 1733
rect 54615 1699 54623 1733
rect 54573 1675 54623 1699
rect 54909 1733 54959 1757
rect 54909 1699 54917 1733
rect 54951 1699 54959 1733
rect 54909 1675 54959 1699
rect 55245 1733 55295 1757
rect 55245 1699 55253 1733
rect 55287 1699 55295 1733
rect 55245 1675 55295 1699
rect 55581 1733 55631 1757
rect 55581 1699 55589 1733
rect 55623 1699 55631 1733
rect 55581 1675 55631 1699
rect 55917 1733 55967 1757
rect 55917 1699 55925 1733
rect 55959 1699 55967 1733
rect 55917 1675 55967 1699
rect 56253 1733 56303 1757
rect 56253 1699 56261 1733
rect 56295 1699 56303 1733
rect 56253 1675 56303 1699
rect 56589 1733 56639 1757
rect 56589 1699 56597 1733
rect 56631 1699 56639 1733
rect 56589 1675 56639 1699
rect 56925 1733 56975 1757
rect 56925 1699 56933 1733
rect 56967 1699 56975 1733
rect 56925 1675 56975 1699
rect 57261 1733 57311 1757
rect 57261 1699 57269 1733
rect 57303 1699 57311 1733
rect 57261 1675 57311 1699
rect 57597 1733 57647 1757
rect 57597 1699 57605 1733
rect 57639 1699 57647 1733
rect 57597 1675 57647 1699
rect 57933 1733 57983 1757
rect 57933 1699 57941 1733
rect 57975 1699 57983 1733
rect 57933 1675 57983 1699
rect 58269 1733 58319 1757
rect 58269 1699 58277 1733
rect 58311 1699 58319 1733
rect 58269 1675 58319 1699
rect 58605 1733 58655 1757
rect 58605 1699 58613 1733
rect 58647 1699 58655 1733
rect 58605 1675 58655 1699
rect 58941 1733 58991 1757
rect 58941 1699 58949 1733
rect 58983 1699 58991 1733
rect 58941 1675 58991 1699
rect 59277 1733 59327 1757
rect 59277 1699 59285 1733
rect 59319 1699 59327 1733
rect 59277 1675 59327 1699
rect 59613 1733 59663 1757
rect 59613 1699 59621 1733
rect 59655 1699 59663 1733
rect 59613 1675 59663 1699
rect 59949 1733 59999 1757
rect 59949 1699 59957 1733
rect 59991 1699 59999 1733
rect 59949 1675 59999 1699
rect 60285 1733 60335 1757
rect 60285 1699 60293 1733
rect 60327 1699 60335 1733
rect 60285 1675 60335 1699
rect 60621 1733 60671 1757
rect 60621 1699 60629 1733
rect 60663 1699 60671 1733
rect 60621 1675 60671 1699
rect 60957 1733 61007 1757
rect 60957 1699 60965 1733
rect 60999 1699 61007 1733
rect 60957 1675 61007 1699
rect 61293 1733 61343 1757
rect 61293 1699 61301 1733
rect 61335 1699 61343 1733
rect 61293 1675 61343 1699
rect 61629 1733 61679 1757
rect 61629 1699 61637 1733
rect 61671 1699 61679 1733
rect 61629 1675 61679 1699
rect 61965 1733 62015 1757
rect 61965 1699 61973 1733
rect 62007 1699 62015 1733
rect 61965 1675 62015 1699
rect 62301 1733 62351 1757
rect 62301 1699 62309 1733
rect 62343 1699 62351 1733
rect 62301 1675 62351 1699
rect 62637 1733 62687 1757
rect 62637 1699 62645 1733
rect 62679 1699 62687 1733
rect 62637 1675 62687 1699
rect 62973 1733 63023 1757
rect 62973 1699 62981 1733
rect 63015 1699 63023 1733
rect 62973 1675 63023 1699
rect 63309 1733 63359 1757
rect 63309 1699 63317 1733
rect 63351 1699 63359 1733
rect 63309 1675 63359 1699
rect 63645 1733 63695 1757
rect 63645 1699 63653 1733
rect 63687 1699 63695 1733
rect 63645 1675 63695 1699
rect 63981 1733 64031 1757
rect 63981 1699 63989 1733
rect 64023 1699 64031 1733
rect 63981 1675 64031 1699
rect 64317 1733 64367 1757
rect 64317 1699 64325 1733
rect 64359 1699 64367 1733
rect 64317 1675 64367 1699
rect 64653 1733 64703 1757
rect 64653 1699 64661 1733
rect 64695 1699 64703 1733
rect 64653 1675 64703 1699
rect 64989 1733 65039 1757
rect 64989 1699 64997 1733
rect 65031 1699 65039 1733
rect 64989 1675 65039 1699
rect 65325 1733 65375 1757
rect 65325 1699 65333 1733
rect 65367 1699 65375 1733
rect 65325 1675 65375 1699
rect 65661 1733 65711 1757
rect 65661 1699 65669 1733
rect 65703 1699 65711 1733
rect 65661 1675 65711 1699
rect 65997 1733 66047 1757
rect 65997 1699 66005 1733
rect 66039 1699 66047 1733
rect 65997 1675 66047 1699
rect 66333 1733 66383 1757
rect 66333 1699 66341 1733
rect 66375 1699 66383 1733
rect 66333 1675 66383 1699
rect 66669 1733 66719 1757
rect 66669 1699 66677 1733
rect 66711 1699 66719 1733
rect 66669 1675 66719 1699
rect 67005 1733 67055 1757
rect 67005 1699 67013 1733
rect 67047 1699 67055 1733
rect 67005 1675 67055 1699
rect 67341 1733 67391 1757
rect 67341 1699 67349 1733
rect 67383 1699 67391 1733
rect 67341 1675 67391 1699
rect 67677 1733 67727 1757
rect 67677 1699 67685 1733
rect 67719 1699 67727 1733
rect 67677 1675 67727 1699
rect 68013 1733 68063 1757
rect 68013 1699 68021 1733
rect 68055 1699 68063 1733
rect 68013 1675 68063 1699
rect 68349 1733 68399 1757
rect 68349 1699 68357 1733
rect 68391 1699 68399 1733
rect 68349 1675 68399 1699
rect 68685 1733 68735 1757
rect 68685 1699 68693 1733
rect 68727 1699 68735 1733
rect 68685 1675 68735 1699
rect 69021 1733 69071 1757
rect 69021 1699 69029 1733
rect 69063 1699 69071 1733
rect 69021 1675 69071 1699
rect 69357 1733 69407 1757
rect 69357 1699 69365 1733
rect 69399 1699 69407 1733
rect 69357 1675 69407 1699
rect 69693 1733 69743 1757
rect 69693 1699 69701 1733
rect 69735 1699 69743 1733
rect 69693 1675 69743 1699
rect 70029 1733 70079 1757
rect 70029 1699 70037 1733
rect 70071 1699 70079 1733
rect 70029 1675 70079 1699
rect 70365 1733 70415 1757
rect 70365 1699 70373 1733
rect 70407 1699 70415 1733
rect 70365 1675 70415 1699
rect 70701 1733 70751 1757
rect 70701 1699 70709 1733
rect 70743 1699 70751 1733
rect 70701 1675 70751 1699
rect 71037 1733 71087 1757
rect 71037 1699 71045 1733
rect 71079 1699 71087 1733
rect 71037 1675 71087 1699
rect 71373 1733 71423 1757
rect 71373 1699 71381 1733
rect 71415 1699 71423 1733
rect 71373 1675 71423 1699
rect 71709 1733 71759 1757
rect 71709 1699 71717 1733
rect 71751 1699 71759 1733
rect 71709 1675 71759 1699
rect 72045 1733 72095 1757
rect 72045 1699 72053 1733
rect 72087 1699 72095 1733
rect 72045 1675 72095 1699
rect 72381 1733 72431 1757
rect 72381 1699 72389 1733
rect 72423 1699 72431 1733
rect 72381 1675 72431 1699
rect 72717 1733 72767 1757
rect 72717 1699 72725 1733
rect 72759 1699 72767 1733
rect 72717 1675 72767 1699
rect 73053 1733 73103 1757
rect 73053 1699 73061 1733
rect 73095 1699 73103 1733
rect 73053 1675 73103 1699
rect 73389 1733 73439 1757
rect 73389 1699 73397 1733
rect 73431 1699 73439 1733
rect 73389 1675 73439 1699
rect 73725 1733 73775 1757
rect 73725 1699 73733 1733
rect 73767 1699 73775 1733
rect 73725 1675 73775 1699
rect 74061 1733 74111 1757
rect 74061 1699 74069 1733
rect 74103 1699 74111 1733
rect 74061 1675 74111 1699
rect 74397 1733 74447 1757
rect 74397 1699 74405 1733
rect 74439 1699 74447 1733
rect 74397 1675 74447 1699
rect 74733 1733 74783 1757
rect 74733 1699 74741 1733
rect 74775 1699 74783 1733
rect 74733 1675 74783 1699
rect 75069 1733 75119 1757
rect 75069 1699 75077 1733
rect 75111 1699 75119 1733
rect 75069 1675 75119 1699
rect 75405 1733 75455 1757
rect 75405 1699 75413 1733
rect 75447 1699 75455 1733
rect 75405 1675 75455 1699
rect 75741 1733 75791 1757
rect 75741 1699 75749 1733
rect 75783 1699 75791 1733
rect 75741 1675 75791 1699
rect 76077 1733 76127 1757
rect 76077 1699 76085 1733
rect 76119 1699 76127 1733
rect 76077 1675 76127 1699
rect 76413 1733 76463 1757
rect 76413 1699 76421 1733
rect 76455 1699 76463 1733
rect 76413 1675 76463 1699
rect 76749 1733 76799 1757
rect 76749 1699 76757 1733
rect 76791 1699 76799 1733
rect 76749 1675 76799 1699
rect 77085 1733 77135 1757
rect 77085 1699 77093 1733
rect 77127 1699 77135 1733
rect 77085 1675 77135 1699
rect 77421 1733 77471 1757
rect 77421 1699 77429 1733
rect 77463 1699 77471 1733
rect 77421 1675 77471 1699
rect 77757 1733 77807 1757
rect 77757 1699 77765 1733
rect 77799 1699 77807 1733
rect 77757 1675 77807 1699
rect 78093 1733 78143 1757
rect 78093 1699 78101 1733
rect 78135 1699 78143 1733
rect 78093 1675 78143 1699
rect 78429 1733 78479 1757
rect 78429 1699 78437 1733
rect 78471 1699 78479 1733
rect 78429 1675 78479 1699
rect 78765 1733 78815 1757
rect 78765 1699 78773 1733
rect 78807 1699 78815 1733
rect 78765 1675 78815 1699
rect 79101 1733 79151 1757
rect 79101 1699 79109 1733
rect 79143 1699 79151 1733
rect 79101 1675 79151 1699
rect 79437 1733 79487 1757
rect 79437 1699 79445 1733
rect 79479 1699 79487 1733
rect 79437 1675 79487 1699
rect 79773 1733 79823 1757
rect 79773 1699 79781 1733
rect 79815 1699 79823 1733
rect 79773 1675 79823 1699
rect 80109 1733 80159 1757
rect 80109 1699 80117 1733
rect 80151 1699 80159 1733
rect 80109 1675 80159 1699
rect 80445 1733 80495 1757
rect 80445 1699 80453 1733
rect 80487 1699 80495 1733
rect 80445 1675 80495 1699
rect 80781 1733 80831 1757
rect 80781 1699 80789 1733
rect 80823 1699 80831 1733
rect 80781 1675 80831 1699
rect 81117 1733 81167 1757
rect 81117 1699 81125 1733
rect 81159 1699 81167 1733
rect 81117 1675 81167 1699
rect 81453 1733 81503 1757
rect 81453 1699 81461 1733
rect 81495 1699 81503 1733
rect 81453 1675 81503 1699
rect 81789 1733 81839 1757
rect 81789 1699 81797 1733
rect 81831 1699 81839 1733
rect 81789 1675 81839 1699
rect 82125 1733 82175 1757
rect 82125 1699 82133 1733
rect 82167 1699 82175 1733
rect 82125 1675 82175 1699
rect 82461 1733 82511 1757
rect 82461 1699 82469 1733
rect 82503 1699 82511 1733
rect 82461 1675 82511 1699
rect 82797 1733 82847 1757
rect 82797 1699 82805 1733
rect 82839 1699 82847 1733
rect 82797 1675 82847 1699
rect 83133 1733 83183 1757
rect 83133 1699 83141 1733
rect 83175 1699 83183 1733
rect 83133 1675 83183 1699
rect 83469 1733 83519 1757
rect 83469 1699 83477 1733
rect 83511 1699 83519 1733
rect 83469 1675 83519 1699
rect 83805 1733 83855 1757
rect 83805 1699 83813 1733
rect 83847 1699 83855 1733
rect 83805 1675 83855 1699
rect 84141 1733 84191 1757
rect 84141 1699 84149 1733
rect 84183 1699 84191 1733
rect 84141 1675 84191 1699
rect 84477 1733 84527 1757
rect 84477 1699 84485 1733
rect 84519 1699 84527 1733
rect 84477 1675 84527 1699
rect 84813 1733 84863 1757
rect 84813 1699 84821 1733
rect 84855 1699 84863 1733
rect 84813 1675 84863 1699
rect 85149 1733 85199 1757
rect 85149 1699 85157 1733
rect 85191 1699 85199 1733
rect 85149 1675 85199 1699
rect 85485 1733 85535 1757
rect 85485 1699 85493 1733
rect 85527 1699 85535 1733
rect 85485 1675 85535 1699
rect 85821 1733 85871 1757
rect 85821 1699 85829 1733
rect 85863 1699 85871 1733
rect 85821 1675 85871 1699
rect 86157 1733 86207 1757
rect 86157 1699 86165 1733
rect 86199 1699 86207 1733
rect 86157 1675 86207 1699
rect 86493 1733 86543 1757
rect 86493 1699 86501 1733
rect 86535 1699 86543 1733
rect 86493 1675 86543 1699
rect 86829 1733 86879 1757
rect 86829 1699 86837 1733
rect 86871 1699 86879 1733
rect 86829 1675 86879 1699
rect 87165 1733 87215 1757
rect 87165 1699 87173 1733
rect 87207 1699 87215 1733
rect 87165 1675 87215 1699
rect 87501 1733 87551 1757
rect 87501 1699 87509 1733
rect 87543 1699 87551 1733
rect 87501 1675 87551 1699
rect 87837 1733 87887 1757
rect 87837 1699 87845 1733
rect 87879 1699 87887 1733
rect 87837 1675 87887 1699
rect 88173 1733 88223 1757
rect 88173 1699 88181 1733
rect 88215 1699 88223 1733
rect 88173 1675 88223 1699
rect 88509 1733 88559 1757
rect 88509 1699 88517 1733
rect 88551 1699 88559 1733
rect 88509 1675 88559 1699
rect 88845 1733 88895 1757
rect 88845 1699 88853 1733
rect 88887 1699 88895 1733
rect 88845 1675 88895 1699
rect 89181 1733 89231 1757
rect 89181 1699 89189 1733
rect 89223 1699 89231 1733
rect 89181 1675 89231 1699
rect 89517 1733 89567 1757
rect 89517 1699 89525 1733
rect 89559 1699 89567 1733
rect 89517 1675 89567 1699
rect 89853 1733 89903 1757
rect 89853 1699 89861 1733
rect 89895 1699 89903 1733
rect 89853 1675 89903 1699
rect 90189 1733 90239 1757
rect 90189 1699 90197 1733
rect 90231 1699 90239 1733
rect 90189 1675 90239 1699
rect 90525 1733 90575 1757
rect 90525 1699 90533 1733
rect 90567 1699 90575 1733
rect 90525 1675 90575 1699
rect 90861 1733 90911 1757
rect 90861 1699 90869 1733
rect 90903 1699 90911 1733
rect 90861 1675 90911 1699
rect 91197 1733 91247 1757
rect 91197 1699 91205 1733
rect 91239 1699 91247 1733
rect 91197 1675 91247 1699
rect 91533 1733 91583 1757
rect 91533 1699 91541 1733
rect 91575 1699 91583 1733
rect 91533 1675 91583 1699
rect 91869 1733 91919 1757
rect 91869 1699 91877 1733
rect 91911 1699 91919 1733
rect 91869 1675 91919 1699
rect 92205 1733 92255 1757
rect 92205 1699 92213 1733
rect 92247 1699 92255 1733
rect 92205 1675 92255 1699
rect 92541 1733 92591 1757
rect 92541 1699 92549 1733
rect 92583 1699 92591 1733
rect 92541 1675 92591 1699
rect 92877 1733 92927 1757
rect 92877 1699 92885 1733
rect 92919 1699 92927 1733
rect 92877 1675 92927 1699
rect 93213 1733 93263 1757
rect 93213 1699 93221 1733
rect 93255 1699 93263 1733
rect 93213 1675 93263 1699
rect 93549 1733 93599 1757
rect 93549 1699 93557 1733
rect 93591 1699 93599 1733
rect 93549 1675 93599 1699
<< nsubdiffcont >>
rect 2165 77763 2199 77797
rect 2501 77763 2535 77797
rect 2837 77763 2871 77797
rect 3173 77763 3207 77797
rect 3509 77763 3543 77797
rect 3845 77763 3879 77797
rect 4181 77763 4215 77797
rect 4517 77763 4551 77797
rect 4853 77763 4887 77797
rect 5189 77763 5223 77797
rect 5525 77763 5559 77797
rect 5861 77763 5895 77797
rect 6197 77763 6231 77797
rect 6533 77763 6567 77797
rect 6869 77763 6903 77797
rect 7205 77763 7239 77797
rect 7541 77763 7575 77797
rect 7877 77763 7911 77797
rect 8213 77763 8247 77797
rect 8549 77763 8583 77797
rect 8885 77763 8919 77797
rect 9221 77763 9255 77797
rect 9557 77763 9591 77797
rect 9893 77763 9927 77797
rect 10229 77763 10263 77797
rect 10565 77763 10599 77797
rect 10901 77763 10935 77797
rect 11237 77763 11271 77797
rect 11573 77763 11607 77797
rect 11909 77763 11943 77797
rect 12245 77763 12279 77797
rect 12581 77763 12615 77797
rect 12917 77763 12951 77797
rect 13253 77763 13287 77797
rect 13589 77763 13623 77797
rect 13925 77763 13959 77797
rect 14261 77763 14295 77797
rect 14597 77763 14631 77797
rect 14933 77763 14967 77797
rect 15269 77763 15303 77797
rect 15605 77763 15639 77797
rect 15941 77763 15975 77797
rect 16277 77763 16311 77797
rect 16613 77763 16647 77797
rect 16949 77763 16983 77797
rect 17285 77763 17319 77797
rect 17621 77763 17655 77797
rect 17957 77763 17991 77797
rect 18293 77763 18327 77797
rect 18629 77763 18663 77797
rect 18965 77763 18999 77797
rect 19301 77763 19335 77797
rect 19637 77763 19671 77797
rect 19973 77763 20007 77797
rect 20309 77763 20343 77797
rect 20645 77763 20679 77797
rect 20981 77763 21015 77797
rect 21317 77763 21351 77797
rect 21653 77763 21687 77797
rect 21989 77763 22023 77797
rect 22325 77763 22359 77797
rect 22661 77763 22695 77797
rect 22997 77763 23031 77797
rect 23333 77763 23367 77797
rect 23669 77763 23703 77797
rect 24005 77763 24039 77797
rect 24341 77763 24375 77797
rect 24677 77763 24711 77797
rect 25013 77763 25047 77797
rect 25349 77763 25383 77797
rect 25685 77763 25719 77797
rect 26021 77763 26055 77797
rect 26357 77763 26391 77797
rect 26693 77763 26727 77797
rect 27029 77763 27063 77797
rect 27365 77763 27399 77797
rect 27701 77763 27735 77797
rect 28037 77763 28071 77797
rect 28373 77763 28407 77797
rect 28709 77763 28743 77797
rect 29045 77763 29079 77797
rect 29381 77763 29415 77797
rect 29717 77763 29751 77797
rect 30053 77763 30087 77797
rect 30389 77763 30423 77797
rect 30725 77763 30759 77797
rect 31061 77763 31095 77797
rect 31397 77763 31431 77797
rect 31733 77763 31767 77797
rect 32069 77763 32103 77797
rect 32405 77763 32439 77797
rect 32741 77763 32775 77797
rect 33077 77763 33111 77797
rect 33413 77763 33447 77797
rect 33749 77763 33783 77797
rect 34085 77763 34119 77797
rect 34421 77763 34455 77797
rect 34757 77763 34791 77797
rect 35093 77763 35127 77797
rect 35429 77763 35463 77797
rect 35765 77763 35799 77797
rect 36101 77763 36135 77797
rect 36437 77763 36471 77797
rect 36773 77763 36807 77797
rect 37109 77763 37143 77797
rect 37445 77763 37479 77797
rect 37781 77763 37815 77797
rect 38117 77763 38151 77797
rect 38453 77763 38487 77797
rect 38789 77763 38823 77797
rect 39125 77763 39159 77797
rect 39461 77763 39495 77797
rect 39797 77763 39831 77797
rect 40133 77763 40167 77797
rect 40469 77763 40503 77797
rect 40805 77763 40839 77797
rect 41141 77763 41175 77797
rect 41477 77763 41511 77797
rect 41813 77763 41847 77797
rect 42149 77763 42183 77797
rect 42485 77763 42519 77797
rect 42821 77763 42855 77797
rect 43157 77763 43191 77797
rect 43493 77763 43527 77797
rect 43829 77763 43863 77797
rect 44165 77763 44199 77797
rect 44501 77763 44535 77797
rect 44837 77763 44871 77797
rect 45173 77763 45207 77797
rect 45509 77763 45543 77797
rect 45845 77763 45879 77797
rect 46181 77763 46215 77797
rect 46517 77763 46551 77797
rect 46853 77763 46887 77797
rect 47189 77763 47223 77797
rect 47525 77763 47559 77797
rect 47861 77763 47895 77797
rect 48197 77763 48231 77797
rect 48533 77763 48567 77797
rect 48869 77763 48903 77797
rect 49205 77763 49239 77797
rect 49541 77763 49575 77797
rect 49877 77763 49911 77797
rect 50213 77763 50247 77797
rect 50549 77763 50583 77797
rect 50885 77763 50919 77797
rect 51221 77763 51255 77797
rect 51557 77763 51591 77797
rect 51893 77763 51927 77797
rect 52229 77763 52263 77797
rect 52565 77763 52599 77797
rect 52901 77763 52935 77797
rect 53237 77763 53271 77797
rect 53573 77763 53607 77797
rect 53909 77763 53943 77797
rect 54245 77763 54279 77797
rect 54581 77763 54615 77797
rect 54917 77763 54951 77797
rect 55253 77763 55287 77797
rect 55589 77763 55623 77797
rect 55925 77763 55959 77797
rect 56261 77763 56295 77797
rect 56597 77763 56631 77797
rect 56933 77763 56967 77797
rect 57269 77763 57303 77797
rect 57605 77763 57639 77797
rect 57941 77763 57975 77797
rect 58277 77763 58311 77797
rect 58613 77763 58647 77797
rect 58949 77763 58983 77797
rect 59285 77763 59319 77797
rect 59621 77763 59655 77797
rect 59957 77763 59991 77797
rect 60293 77763 60327 77797
rect 60629 77763 60663 77797
rect 60965 77763 60999 77797
rect 61301 77763 61335 77797
rect 61637 77763 61671 77797
rect 61973 77763 62007 77797
rect 62309 77763 62343 77797
rect 62645 77763 62679 77797
rect 62981 77763 63015 77797
rect 63317 77763 63351 77797
rect 63653 77763 63687 77797
rect 63989 77763 64023 77797
rect 64325 77763 64359 77797
rect 64661 77763 64695 77797
rect 64997 77763 65031 77797
rect 65333 77763 65367 77797
rect 65669 77763 65703 77797
rect 66005 77763 66039 77797
rect 66341 77763 66375 77797
rect 66677 77763 66711 77797
rect 67013 77763 67047 77797
rect 67349 77763 67383 77797
rect 67685 77763 67719 77797
rect 68021 77763 68055 77797
rect 68357 77763 68391 77797
rect 68693 77763 68727 77797
rect 69029 77763 69063 77797
rect 69365 77763 69399 77797
rect 69701 77763 69735 77797
rect 70037 77763 70071 77797
rect 70373 77763 70407 77797
rect 70709 77763 70743 77797
rect 71045 77763 71079 77797
rect 71381 77763 71415 77797
rect 71717 77763 71751 77797
rect 72053 77763 72087 77797
rect 72389 77763 72423 77797
rect 72725 77763 72759 77797
rect 73061 77763 73095 77797
rect 73397 77763 73431 77797
rect 73733 77763 73767 77797
rect 74069 77763 74103 77797
rect 74405 77763 74439 77797
rect 74741 77763 74775 77797
rect 75077 77763 75111 77797
rect 75413 77763 75447 77797
rect 75749 77763 75783 77797
rect 76085 77763 76119 77797
rect 76421 77763 76455 77797
rect 76757 77763 76791 77797
rect 77093 77763 77127 77797
rect 77429 77763 77463 77797
rect 77765 77763 77799 77797
rect 78101 77763 78135 77797
rect 78437 77763 78471 77797
rect 78773 77763 78807 77797
rect 79109 77763 79143 77797
rect 79445 77763 79479 77797
rect 79781 77763 79815 77797
rect 80117 77763 80151 77797
rect 80453 77763 80487 77797
rect 80789 77763 80823 77797
rect 81125 77763 81159 77797
rect 81461 77763 81495 77797
rect 81797 77763 81831 77797
rect 82133 77763 82167 77797
rect 82469 77763 82503 77797
rect 82805 77763 82839 77797
rect 83141 77763 83175 77797
rect 83477 77763 83511 77797
rect 83813 77763 83847 77797
rect 84149 77763 84183 77797
rect 84485 77763 84519 77797
rect 84821 77763 84855 77797
rect 85157 77763 85191 77797
rect 85493 77763 85527 77797
rect 85829 77763 85863 77797
rect 86165 77763 86199 77797
rect 86501 77763 86535 77797
rect 86837 77763 86871 77797
rect 87173 77763 87207 77797
rect 87509 77763 87543 77797
rect 87845 77763 87879 77797
rect 88181 77763 88215 77797
rect 88517 77763 88551 77797
rect 88853 77763 88887 77797
rect 89189 77763 89223 77797
rect 89525 77763 89559 77797
rect 89861 77763 89895 77797
rect 90197 77763 90231 77797
rect 90533 77763 90567 77797
rect 90869 77763 90903 77797
rect 91205 77763 91239 77797
rect 91541 77763 91575 77797
rect 91877 77763 91911 77797
rect 92213 77763 92247 77797
rect 92549 77763 92583 77797
rect 92885 77763 92919 77797
rect 93221 77763 93255 77797
rect 93557 77763 93591 77797
rect 1829 77299 1863 77333
rect 94187 77299 94221 77333
rect 1829 76963 1863 76997
rect 94187 76963 94221 76997
rect 1829 76627 1863 76661
rect 94187 76627 94221 76661
rect 1829 76291 1863 76325
rect 94187 76291 94221 76325
rect 1829 75955 1863 75989
rect 94187 75955 94221 75989
rect 1829 75619 1863 75653
rect 94187 75619 94221 75653
rect 1829 75283 1863 75317
rect 94187 75283 94221 75317
rect 1829 74947 1863 74981
rect 94187 74947 94221 74981
rect 1829 74611 1863 74645
rect 94187 74611 94221 74645
rect 1829 74275 1863 74309
rect 94187 74275 94221 74309
rect 1829 73939 1863 73973
rect 94187 73939 94221 73973
rect 1829 73603 1863 73637
rect 94187 73603 94221 73637
rect 1829 73267 1863 73301
rect 94187 73267 94221 73301
rect 1829 72931 1863 72965
rect 94187 72931 94221 72965
rect 1829 72595 1863 72629
rect 94187 72595 94221 72629
rect 1829 72259 1863 72293
rect 94187 72259 94221 72293
rect 1829 71923 1863 71957
rect 94187 71923 94221 71957
rect 1829 71587 1863 71621
rect 94187 71587 94221 71621
rect 1829 71251 1863 71285
rect 94187 71251 94221 71285
rect 1829 70915 1863 70949
rect 94187 70915 94221 70949
rect 1829 70579 1863 70613
rect 94187 70579 94221 70613
rect 1829 70243 1863 70277
rect 94187 70243 94221 70277
rect 1829 69907 1863 69941
rect 94187 69907 94221 69941
rect 1829 69571 1863 69605
rect 94187 69571 94221 69605
rect 1829 69235 1863 69269
rect 94187 69235 94221 69269
rect 1829 68899 1863 68933
rect 94187 68899 94221 68933
rect 1829 68563 1863 68597
rect 94187 68563 94221 68597
rect 1829 68227 1863 68261
rect 94187 68227 94221 68261
rect 1829 67891 1863 67925
rect 94187 67891 94221 67925
rect 1829 67555 1863 67589
rect 94187 67555 94221 67589
rect 1829 67219 1863 67253
rect 94187 67219 94221 67253
rect 1829 66883 1863 66917
rect 94187 66883 94221 66917
rect 1829 66547 1863 66581
rect 94187 66547 94221 66581
rect 1829 66211 1863 66245
rect 94187 66211 94221 66245
rect 1829 65875 1863 65909
rect 94187 65875 94221 65909
rect 1829 65539 1863 65573
rect 94187 65539 94221 65573
rect 1829 65203 1863 65237
rect 94187 65203 94221 65237
rect 1829 64867 1863 64901
rect 94187 64867 94221 64901
rect 1829 64531 1863 64565
rect 94187 64531 94221 64565
rect 1829 64195 1863 64229
rect 94187 64195 94221 64229
rect 1829 63859 1863 63893
rect 94187 63859 94221 63893
rect 1829 63523 1863 63557
rect 94187 63523 94221 63557
rect 1829 63187 1863 63221
rect 94187 63187 94221 63221
rect 1829 62851 1863 62885
rect 94187 62851 94221 62885
rect 1829 62515 1863 62549
rect 94187 62515 94221 62549
rect 1829 62179 1863 62213
rect 94187 62179 94221 62213
rect 1829 61843 1863 61877
rect 94187 61843 94221 61877
rect 1829 61507 1863 61541
rect 94187 61507 94221 61541
rect 1829 61171 1863 61205
rect 94187 61171 94221 61205
rect 1829 60835 1863 60869
rect 94187 60835 94221 60869
rect 1829 60499 1863 60533
rect 94187 60499 94221 60533
rect 1829 60163 1863 60197
rect 94187 60163 94221 60197
rect 1829 59827 1863 59861
rect 94187 59827 94221 59861
rect 1829 59491 1863 59525
rect 94187 59491 94221 59525
rect 1829 59155 1863 59189
rect 94187 59155 94221 59189
rect 1829 58819 1863 58853
rect 94187 58819 94221 58853
rect 1829 58483 1863 58517
rect 94187 58483 94221 58517
rect 1829 58147 1863 58181
rect 94187 58147 94221 58181
rect 1829 57811 1863 57845
rect 94187 57811 94221 57845
rect 1829 57475 1863 57509
rect 94187 57475 94221 57509
rect 1829 57139 1863 57173
rect 94187 57139 94221 57173
rect 1829 56803 1863 56837
rect 94187 56803 94221 56837
rect 1829 56467 1863 56501
rect 94187 56467 94221 56501
rect 1829 56131 1863 56165
rect 94187 56131 94221 56165
rect 1829 55795 1863 55829
rect 94187 55795 94221 55829
rect 1829 55459 1863 55493
rect 94187 55459 94221 55493
rect 1829 55123 1863 55157
rect 94187 55123 94221 55157
rect 1829 54787 1863 54821
rect 94187 54787 94221 54821
rect 1829 54451 1863 54485
rect 94187 54451 94221 54485
rect 1829 54115 1863 54149
rect 94187 54115 94221 54149
rect 1829 53779 1863 53813
rect 94187 53779 94221 53813
rect 1829 53443 1863 53477
rect 94187 53443 94221 53477
rect 1829 53107 1863 53141
rect 94187 53107 94221 53141
rect 1829 52771 1863 52805
rect 94187 52771 94221 52805
rect 1829 52435 1863 52469
rect 94187 52435 94221 52469
rect 1829 52099 1863 52133
rect 94187 52099 94221 52133
rect 1829 51763 1863 51797
rect 94187 51763 94221 51797
rect 1829 51427 1863 51461
rect 94187 51427 94221 51461
rect 1829 51091 1863 51125
rect 94187 51091 94221 51125
rect 1829 50755 1863 50789
rect 94187 50755 94221 50789
rect 1829 50419 1863 50453
rect 94187 50419 94221 50453
rect 1829 50083 1863 50117
rect 94187 50083 94221 50117
rect 1829 49747 1863 49781
rect 94187 49747 94221 49781
rect 1829 49411 1863 49445
rect 94187 49411 94221 49445
rect 1829 49075 1863 49109
rect 94187 49075 94221 49109
rect 1829 48739 1863 48773
rect 94187 48739 94221 48773
rect 1829 48403 1863 48437
rect 94187 48403 94221 48437
rect 1829 48067 1863 48101
rect 94187 48067 94221 48101
rect 1829 47731 1863 47765
rect 94187 47731 94221 47765
rect 1829 47395 1863 47429
rect 94187 47395 94221 47429
rect 1829 47059 1863 47093
rect 94187 47059 94221 47093
rect 1829 46723 1863 46757
rect 94187 46723 94221 46757
rect 1829 46387 1863 46421
rect 94187 46387 94221 46421
rect 1829 46051 1863 46085
rect 94187 46051 94221 46085
rect 1829 45715 1863 45749
rect 94187 45715 94221 45749
rect 1829 45379 1863 45413
rect 94187 45379 94221 45413
rect 1829 45043 1863 45077
rect 94187 45043 94221 45077
rect 1829 44707 1863 44741
rect 94187 44707 94221 44741
rect 1829 44371 1863 44405
rect 94187 44371 94221 44405
rect 1829 44035 1863 44069
rect 94187 44035 94221 44069
rect 1829 43699 1863 43733
rect 94187 43699 94221 43733
rect 1829 43363 1863 43397
rect 94187 43363 94221 43397
rect 1829 43027 1863 43061
rect 94187 43027 94221 43061
rect 1829 42691 1863 42725
rect 94187 42691 94221 42725
rect 1829 42355 1863 42389
rect 94187 42355 94221 42389
rect 1829 42019 1863 42053
rect 94187 42019 94221 42053
rect 1829 41683 1863 41717
rect 94187 41683 94221 41717
rect 1829 41347 1863 41381
rect 94187 41347 94221 41381
rect 1829 41011 1863 41045
rect 94187 41011 94221 41045
rect 1829 40675 1863 40709
rect 94187 40675 94221 40709
rect 1829 40339 1863 40373
rect 94187 40339 94221 40373
rect 1829 40003 1863 40037
rect 94187 40003 94221 40037
rect 1829 39667 1863 39701
rect 94187 39667 94221 39701
rect 1829 39331 1863 39365
rect 94187 39331 94221 39365
rect 1829 38995 1863 39029
rect 94187 38995 94221 39029
rect 1829 38659 1863 38693
rect 94187 38659 94221 38693
rect 1829 38323 1863 38357
rect 94187 38323 94221 38357
rect 1829 37987 1863 38021
rect 94187 37987 94221 38021
rect 1829 37651 1863 37685
rect 94187 37651 94221 37685
rect 1829 37315 1863 37349
rect 94187 37315 94221 37349
rect 1829 36979 1863 37013
rect 94187 36979 94221 37013
rect 1829 36643 1863 36677
rect 94187 36643 94221 36677
rect 1829 36307 1863 36341
rect 94187 36307 94221 36341
rect 1829 35971 1863 36005
rect 94187 35971 94221 36005
rect 1829 35635 1863 35669
rect 94187 35635 94221 35669
rect 1829 35299 1863 35333
rect 94187 35299 94221 35333
rect 1829 34963 1863 34997
rect 94187 34963 94221 34997
rect 1829 34627 1863 34661
rect 94187 34627 94221 34661
rect 1829 34291 1863 34325
rect 94187 34291 94221 34325
rect 1829 33955 1863 33989
rect 94187 33955 94221 33989
rect 1829 33619 1863 33653
rect 94187 33619 94221 33653
rect 1829 33283 1863 33317
rect 94187 33283 94221 33317
rect 1829 32947 1863 32981
rect 94187 32947 94221 32981
rect 1829 32611 1863 32645
rect 94187 32611 94221 32645
rect 1829 32275 1863 32309
rect 94187 32275 94221 32309
rect 1829 31939 1863 31973
rect 94187 31939 94221 31973
rect 1829 31603 1863 31637
rect 94187 31603 94221 31637
rect 1829 31267 1863 31301
rect 94187 31267 94221 31301
rect 1829 30931 1863 30965
rect 94187 30931 94221 30965
rect 1829 30595 1863 30629
rect 94187 30595 94221 30629
rect 1829 30259 1863 30293
rect 94187 30259 94221 30293
rect 1829 29923 1863 29957
rect 94187 29923 94221 29957
rect 1829 29587 1863 29621
rect 94187 29587 94221 29621
rect 1829 29251 1863 29285
rect 94187 29251 94221 29285
rect 1829 28915 1863 28949
rect 94187 28915 94221 28949
rect 1829 28579 1863 28613
rect 94187 28579 94221 28613
rect 1829 28243 1863 28277
rect 94187 28243 94221 28277
rect 1829 27907 1863 27941
rect 94187 27907 94221 27941
rect 1829 27571 1863 27605
rect 94187 27571 94221 27605
rect 1829 27235 1863 27269
rect 94187 27235 94221 27269
rect 1829 26899 1863 26933
rect 94187 26899 94221 26933
rect 1829 26563 1863 26597
rect 94187 26563 94221 26597
rect 1829 26227 1863 26261
rect 94187 26227 94221 26261
rect 1829 25891 1863 25925
rect 94187 25891 94221 25925
rect 1829 25555 1863 25589
rect 94187 25555 94221 25589
rect 1829 25219 1863 25253
rect 94187 25219 94221 25253
rect 1829 24883 1863 24917
rect 94187 24883 94221 24917
rect 1829 24547 1863 24581
rect 94187 24547 94221 24581
rect 1829 24211 1863 24245
rect 94187 24211 94221 24245
rect 1829 23875 1863 23909
rect 94187 23875 94221 23909
rect 1829 23539 1863 23573
rect 94187 23539 94221 23573
rect 1829 23203 1863 23237
rect 94187 23203 94221 23237
rect 1829 22867 1863 22901
rect 94187 22867 94221 22901
rect 1829 22531 1863 22565
rect 94187 22531 94221 22565
rect 1829 22195 1863 22229
rect 94187 22195 94221 22229
rect 1829 21859 1863 21893
rect 94187 21859 94221 21893
rect 1829 21523 1863 21557
rect 94187 21523 94221 21557
rect 1829 21187 1863 21221
rect 94187 21187 94221 21221
rect 1829 20851 1863 20885
rect 94187 20851 94221 20885
rect 1829 20515 1863 20549
rect 94187 20515 94221 20549
rect 1829 20179 1863 20213
rect 94187 20179 94221 20213
rect 1829 19843 1863 19877
rect 94187 19843 94221 19877
rect 1829 19507 1863 19541
rect 94187 19507 94221 19541
rect 1829 19171 1863 19205
rect 94187 19171 94221 19205
rect 1829 18835 1863 18869
rect 94187 18835 94221 18869
rect 1829 18499 1863 18533
rect 94187 18499 94221 18533
rect 1829 18163 1863 18197
rect 94187 18163 94221 18197
rect 1829 17827 1863 17861
rect 94187 17827 94221 17861
rect 1829 17491 1863 17525
rect 94187 17491 94221 17525
rect 1829 17155 1863 17189
rect 94187 17155 94221 17189
rect 1829 16819 1863 16853
rect 94187 16819 94221 16853
rect 1829 16483 1863 16517
rect 94187 16483 94221 16517
rect 1829 16147 1863 16181
rect 94187 16147 94221 16181
rect 1829 15811 1863 15845
rect 94187 15811 94221 15845
rect 1829 15475 1863 15509
rect 94187 15475 94221 15509
rect 1829 15139 1863 15173
rect 94187 15139 94221 15173
rect 1829 14803 1863 14837
rect 94187 14803 94221 14837
rect 1829 14467 1863 14501
rect 94187 14467 94221 14501
rect 1829 14131 1863 14165
rect 94187 14131 94221 14165
rect 1829 13795 1863 13829
rect 94187 13795 94221 13829
rect 1829 13459 1863 13493
rect 94187 13459 94221 13493
rect 1829 13123 1863 13157
rect 94187 13123 94221 13157
rect 1829 12787 1863 12821
rect 94187 12787 94221 12821
rect 1829 12451 1863 12485
rect 94187 12451 94221 12485
rect 1829 12115 1863 12149
rect 94187 12115 94221 12149
rect 1829 11779 1863 11813
rect 94187 11779 94221 11813
rect 1829 11443 1863 11477
rect 94187 11443 94221 11477
rect 1829 11107 1863 11141
rect 94187 11107 94221 11141
rect 1829 10771 1863 10805
rect 94187 10771 94221 10805
rect 1829 10435 1863 10469
rect 94187 10435 94221 10469
rect 1829 10099 1863 10133
rect 94187 10099 94221 10133
rect 1829 9763 1863 9797
rect 94187 9763 94221 9797
rect 1829 9427 1863 9461
rect 94187 9427 94221 9461
rect 1829 9091 1863 9125
rect 94187 9091 94221 9125
rect 1829 8755 1863 8789
rect 94187 8755 94221 8789
rect 1829 8419 1863 8453
rect 94187 8419 94221 8453
rect 1829 8083 1863 8117
rect 94187 8083 94221 8117
rect 1829 7747 1863 7781
rect 94187 7747 94221 7781
rect 1829 7411 1863 7445
rect 94187 7411 94221 7445
rect 1829 7075 1863 7109
rect 94187 7075 94221 7109
rect 1829 6739 1863 6773
rect 94187 6739 94221 6773
rect 1829 6403 1863 6437
rect 94187 6403 94221 6437
rect 1829 6067 1863 6101
rect 94187 6067 94221 6101
rect 1829 5731 1863 5765
rect 94187 5731 94221 5765
rect 1829 5395 1863 5429
rect 94187 5395 94221 5429
rect 1829 5059 1863 5093
rect 94187 5059 94221 5093
rect 1829 4723 1863 4757
rect 94187 4723 94221 4757
rect 1829 4387 1863 4421
rect 94187 4387 94221 4421
rect 1829 4051 1863 4085
rect 94187 4051 94221 4085
rect 1829 3715 1863 3749
rect 94187 3715 94221 3749
rect 1829 3379 1863 3413
rect 94187 3379 94221 3413
rect 1829 3043 1863 3077
rect 94187 3043 94221 3077
rect 1829 2707 1863 2741
rect 94187 2707 94221 2741
rect 1829 2371 1863 2405
rect 94187 2371 94221 2405
rect 1829 2035 1863 2069
rect 94187 2035 94221 2069
rect 2165 1699 2199 1733
rect 2501 1699 2535 1733
rect 2837 1699 2871 1733
rect 3173 1699 3207 1733
rect 3509 1699 3543 1733
rect 3845 1699 3879 1733
rect 4181 1699 4215 1733
rect 4517 1699 4551 1733
rect 4853 1699 4887 1733
rect 5189 1699 5223 1733
rect 5525 1699 5559 1733
rect 5861 1699 5895 1733
rect 6197 1699 6231 1733
rect 6533 1699 6567 1733
rect 6869 1699 6903 1733
rect 7205 1699 7239 1733
rect 7541 1699 7575 1733
rect 7877 1699 7911 1733
rect 8213 1699 8247 1733
rect 8549 1699 8583 1733
rect 8885 1699 8919 1733
rect 9221 1699 9255 1733
rect 9557 1699 9591 1733
rect 9893 1699 9927 1733
rect 10229 1699 10263 1733
rect 10565 1699 10599 1733
rect 10901 1699 10935 1733
rect 11237 1699 11271 1733
rect 11573 1699 11607 1733
rect 11909 1699 11943 1733
rect 12245 1699 12279 1733
rect 12581 1699 12615 1733
rect 12917 1699 12951 1733
rect 13253 1699 13287 1733
rect 13589 1699 13623 1733
rect 13925 1699 13959 1733
rect 14261 1699 14295 1733
rect 14597 1699 14631 1733
rect 14933 1699 14967 1733
rect 15269 1699 15303 1733
rect 15605 1699 15639 1733
rect 15941 1699 15975 1733
rect 16277 1699 16311 1733
rect 16613 1699 16647 1733
rect 16949 1699 16983 1733
rect 17285 1699 17319 1733
rect 17621 1699 17655 1733
rect 17957 1699 17991 1733
rect 18293 1699 18327 1733
rect 18629 1699 18663 1733
rect 18965 1699 18999 1733
rect 19301 1699 19335 1733
rect 19637 1699 19671 1733
rect 19973 1699 20007 1733
rect 20309 1699 20343 1733
rect 20645 1699 20679 1733
rect 20981 1699 21015 1733
rect 21317 1699 21351 1733
rect 21653 1699 21687 1733
rect 21989 1699 22023 1733
rect 22325 1699 22359 1733
rect 22661 1699 22695 1733
rect 22997 1699 23031 1733
rect 23333 1699 23367 1733
rect 23669 1699 23703 1733
rect 24005 1699 24039 1733
rect 24341 1699 24375 1733
rect 24677 1699 24711 1733
rect 25013 1699 25047 1733
rect 25349 1699 25383 1733
rect 25685 1699 25719 1733
rect 26021 1699 26055 1733
rect 26357 1699 26391 1733
rect 26693 1699 26727 1733
rect 27029 1699 27063 1733
rect 27365 1699 27399 1733
rect 27701 1699 27735 1733
rect 28037 1699 28071 1733
rect 28373 1699 28407 1733
rect 28709 1699 28743 1733
rect 29045 1699 29079 1733
rect 29381 1699 29415 1733
rect 29717 1699 29751 1733
rect 30053 1699 30087 1733
rect 30389 1699 30423 1733
rect 30725 1699 30759 1733
rect 31061 1699 31095 1733
rect 31397 1699 31431 1733
rect 31733 1699 31767 1733
rect 32069 1699 32103 1733
rect 32405 1699 32439 1733
rect 32741 1699 32775 1733
rect 33077 1699 33111 1733
rect 33413 1699 33447 1733
rect 33749 1699 33783 1733
rect 34085 1699 34119 1733
rect 34421 1699 34455 1733
rect 34757 1699 34791 1733
rect 35093 1699 35127 1733
rect 35429 1699 35463 1733
rect 35765 1699 35799 1733
rect 36101 1699 36135 1733
rect 36437 1699 36471 1733
rect 36773 1699 36807 1733
rect 37109 1699 37143 1733
rect 37445 1699 37479 1733
rect 37781 1699 37815 1733
rect 38117 1699 38151 1733
rect 38453 1699 38487 1733
rect 38789 1699 38823 1733
rect 39125 1699 39159 1733
rect 39461 1699 39495 1733
rect 39797 1699 39831 1733
rect 40133 1699 40167 1733
rect 40469 1699 40503 1733
rect 40805 1699 40839 1733
rect 41141 1699 41175 1733
rect 41477 1699 41511 1733
rect 41813 1699 41847 1733
rect 42149 1699 42183 1733
rect 42485 1699 42519 1733
rect 42821 1699 42855 1733
rect 43157 1699 43191 1733
rect 43493 1699 43527 1733
rect 43829 1699 43863 1733
rect 44165 1699 44199 1733
rect 44501 1699 44535 1733
rect 44837 1699 44871 1733
rect 45173 1699 45207 1733
rect 45509 1699 45543 1733
rect 45845 1699 45879 1733
rect 46181 1699 46215 1733
rect 46517 1699 46551 1733
rect 46853 1699 46887 1733
rect 47189 1699 47223 1733
rect 47525 1699 47559 1733
rect 47861 1699 47895 1733
rect 48197 1699 48231 1733
rect 48533 1699 48567 1733
rect 48869 1699 48903 1733
rect 49205 1699 49239 1733
rect 49541 1699 49575 1733
rect 49877 1699 49911 1733
rect 50213 1699 50247 1733
rect 50549 1699 50583 1733
rect 50885 1699 50919 1733
rect 51221 1699 51255 1733
rect 51557 1699 51591 1733
rect 51893 1699 51927 1733
rect 52229 1699 52263 1733
rect 52565 1699 52599 1733
rect 52901 1699 52935 1733
rect 53237 1699 53271 1733
rect 53573 1699 53607 1733
rect 53909 1699 53943 1733
rect 54245 1699 54279 1733
rect 54581 1699 54615 1733
rect 54917 1699 54951 1733
rect 55253 1699 55287 1733
rect 55589 1699 55623 1733
rect 55925 1699 55959 1733
rect 56261 1699 56295 1733
rect 56597 1699 56631 1733
rect 56933 1699 56967 1733
rect 57269 1699 57303 1733
rect 57605 1699 57639 1733
rect 57941 1699 57975 1733
rect 58277 1699 58311 1733
rect 58613 1699 58647 1733
rect 58949 1699 58983 1733
rect 59285 1699 59319 1733
rect 59621 1699 59655 1733
rect 59957 1699 59991 1733
rect 60293 1699 60327 1733
rect 60629 1699 60663 1733
rect 60965 1699 60999 1733
rect 61301 1699 61335 1733
rect 61637 1699 61671 1733
rect 61973 1699 62007 1733
rect 62309 1699 62343 1733
rect 62645 1699 62679 1733
rect 62981 1699 63015 1733
rect 63317 1699 63351 1733
rect 63653 1699 63687 1733
rect 63989 1699 64023 1733
rect 64325 1699 64359 1733
rect 64661 1699 64695 1733
rect 64997 1699 65031 1733
rect 65333 1699 65367 1733
rect 65669 1699 65703 1733
rect 66005 1699 66039 1733
rect 66341 1699 66375 1733
rect 66677 1699 66711 1733
rect 67013 1699 67047 1733
rect 67349 1699 67383 1733
rect 67685 1699 67719 1733
rect 68021 1699 68055 1733
rect 68357 1699 68391 1733
rect 68693 1699 68727 1733
rect 69029 1699 69063 1733
rect 69365 1699 69399 1733
rect 69701 1699 69735 1733
rect 70037 1699 70071 1733
rect 70373 1699 70407 1733
rect 70709 1699 70743 1733
rect 71045 1699 71079 1733
rect 71381 1699 71415 1733
rect 71717 1699 71751 1733
rect 72053 1699 72087 1733
rect 72389 1699 72423 1733
rect 72725 1699 72759 1733
rect 73061 1699 73095 1733
rect 73397 1699 73431 1733
rect 73733 1699 73767 1733
rect 74069 1699 74103 1733
rect 74405 1699 74439 1733
rect 74741 1699 74775 1733
rect 75077 1699 75111 1733
rect 75413 1699 75447 1733
rect 75749 1699 75783 1733
rect 76085 1699 76119 1733
rect 76421 1699 76455 1733
rect 76757 1699 76791 1733
rect 77093 1699 77127 1733
rect 77429 1699 77463 1733
rect 77765 1699 77799 1733
rect 78101 1699 78135 1733
rect 78437 1699 78471 1733
rect 78773 1699 78807 1733
rect 79109 1699 79143 1733
rect 79445 1699 79479 1733
rect 79781 1699 79815 1733
rect 80117 1699 80151 1733
rect 80453 1699 80487 1733
rect 80789 1699 80823 1733
rect 81125 1699 81159 1733
rect 81461 1699 81495 1733
rect 81797 1699 81831 1733
rect 82133 1699 82167 1733
rect 82469 1699 82503 1733
rect 82805 1699 82839 1733
rect 83141 1699 83175 1733
rect 83477 1699 83511 1733
rect 83813 1699 83847 1733
rect 84149 1699 84183 1733
rect 84485 1699 84519 1733
rect 84821 1699 84855 1733
rect 85157 1699 85191 1733
rect 85493 1699 85527 1733
rect 85829 1699 85863 1733
rect 86165 1699 86199 1733
rect 86501 1699 86535 1733
rect 86837 1699 86871 1733
rect 87173 1699 87207 1733
rect 87509 1699 87543 1733
rect 87845 1699 87879 1733
rect 88181 1699 88215 1733
rect 88517 1699 88551 1733
rect 88853 1699 88887 1733
rect 89189 1699 89223 1733
rect 89525 1699 89559 1733
rect 89861 1699 89895 1733
rect 90197 1699 90231 1733
rect 90533 1699 90567 1733
rect 90869 1699 90903 1733
rect 91205 1699 91239 1733
rect 91541 1699 91575 1733
rect 91877 1699 91911 1733
rect 92213 1699 92247 1733
rect 92549 1699 92583 1733
rect 92885 1699 92919 1733
rect 93221 1699 93255 1733
rect 93557 1699 93591 1733
<< locali >>
rect 2165 77797 2199 77813
rect 2165 77747 2199 77763
rect 2501 77797 2535 77813
rect 2501 77747 2535 77763
rect 2837 77797 2871 77813
rect 2837 77747 2871 77763
rect 3173 77797 3207 77813
rect 3173 77747 3207 77763
rect 3509 77797 3543 77813
rect 3509 77747 3543 77763
rect 3845 77797 3879 77813
rect 3845 77747 3879 77763
rect 4181 77797 4215 77813
rect 4181 77747 4215 77763
rect 4517 77797 4551 77813
rect 4517 77747 4551 77763
rect 4853 77797 4887 77813
rect 4853 77747 4887 77763
rect 5189 77797 5223 77813
rect 5189 77747 5223 77763
rect 5525 77797 5559 77813
rect 5525 77747 5559 77763
rect 5861 77797 5895 77813
rect 5861 77747 5895 77763
rect 6197 77797 6231 77813
rect 6197 77747 6231 77763
rect 6533 77797 6567 77813
rect 6533 77747 6567 77763
rect 6869 77797 6903 77813
rect 6869 77747 6903 77763
rect 7205 77797 7239 77813
rect 7205 77747 7239 77763
rect 7541 77797 7575 77813
rect 7541 77747 7575 77763
rect 7877 77797 7911 77813
rect 7877 77747 7911 77763
rect 8213 77797 8247 77813
rect 8213 77747 8247 77763
rect 8549 77797 8583 77813
rect 8549 77747 8583 77763
rect 8885 77797 8919 77813
rect 8885 77747 8919 77763
rect 9221 77797 9255 77813
rect 9221 77747 9255 77763
rect 9557 77797 9591 77813
rect 9557 77747 9591 77763
rect 9893 77797 9927 77813
rect 9893 77747 9927 77763
rect 10229 77797 10263 77813
rect 10229 77747 10263 77763
rect 10565 77797 10599 77813
rect 10565 77747 10599 77763
rect 10901 77797 10935 77813
rect 10901 77747 10935 77763
rect 11237 77797 11271 77813
rect 11237 77747 11271 77763
rect 11573 77797 11607 77813
rect 11573 77747 11607 77763
rect 11909 77797 11943 77813
rect 11909 77747 11943 77763
rect 12245 77797 12279 77813
rect 12245 77747 12279 77763
rect 12581 77797 12615 77813
rect 12581 77747 12615 77763
rect 12917 77797 12951 77813
rect 12917 77747 12951 77763
rect 13253 77797 13287 77813
rect 13253 77747 13287 77763
rect 13589 77797 13623 77813
rect 13589 77747 13623 77763
rect 13925 77797 13959 77813
rect 13925 77747 13959 77763
rect 14261 77797 14295 77813
rect 14261 77747 14295 77763
rect 14597 77797 14631 77813
rect 14597 77747 14631 77763
rect 14933 77797 14967 77813
rect 14933 77747 14967 77763
rect 15269 77797 15303 77813
rect 15269 77747 15303 77763
rect 15605 77797 15639 77813
rect 15605 77747 15639 77763
rect 15941 77797 15975 77813
rect 15941 77747 15975 77763
rect 16277 77797 16311 77813
rect 16277 77747 16311 77763
rect 16613 77797 16647 77813
rect 16613 77747 16647 77763
rect 16949 77797 16983 77813
rect 16949 77747 16983 77763
rect 17285 77797 17319 77813
rect 17285 77747 17319 77763
rect 17621 77797 17655 77813
rect 17621 77747 17655 77763
rect 17957 77797 17991 77813
rect 17957 77747 17991 77763
rect 18293 77797 18327 77813
rect 18293 77747 18327 77763
rect 18629 77797 18663 77813
rect 18629 77747 18663 77763
rect 18965 77797 18999 77813
rect 18965 77747 18999 77763
rect 19301 77797 19335 77813
rect 19301 77747 19335 77763
rect 19637 77797 19671 77813
rect 19637 77747 19671 77763
rect 19973 77797 20007 77813
rect 19973 77747 20007 77763
rect 20309 77797 20343 77813
rect 20309 77747 20343 77763
rect 20645 77797 20679 77813
rect 20645 77747 20679 77763
rect 20981 77797 21015 77813
rect 20981 77747 21015 77763
rect 21317 77797 21351 77813
rect 21317 77747 21351 77763
rect 21653 77797 21687 77813
rect 21653 77747 21687 77763
rect 21989 77797 22023 77813
rect 21989 77747 22023 77763
rect 22325 77797 22359 77813
rect 22325 77747 22359 77763
rect 22661 77797 22695 77813
rect 22661 77747 22695 77763
rect 22997 77797 23031 77813
rect 22997 77747 23031 77763
rect 23333 77797 23367 77813
rect 23333 77747 23367 77763
rect 23669 77797 23703 77813
rect 23669 77747 23703 77763
rect 24005 77797 24039 77813
rect 24005 77747 24039 77763
rect 24341 77797 24375 77813
rect 24341 77747 24375 77763
rect 24677 77797 24711 77813
rect 24677 77747 24711 77763
rect 25013 77797 25047 77813
rect 25013 77747 25047 77763
rect 25349 77797 25383 77813
rect 25349 77747 25383 77763
rect 25685 77797 25719 77813
rect 25685 77747 25719 77763
rect 26021 77797 26055 77813
rect 26021 77747 26055 77763
rect 26357 77797 26391 77813
rect 26357 77747 26391 77763
rect 26693 77797 26727 77813
rect 26693 77747 26727 77763
rect 27029 77797 27063 77813
rect 27029 77747 27063 77763
rect 27365 77797 27399 77813
rect 27365 77747 27399 77763
rect 27701 77797 27735 77813
rect 27701 77747 27735 77763
rect 28037 77797 28071 77813
rect 28037 77747 28071 77763
rect 28373 77797 28407 77813
rect 28373 77747 28407 77763
rect 28709 77797 28743 77813
rect 28709 77747 28743 77763
rect 29045 77797 29079 77813
rect 29045 77747 29079 77763
rect 29381 77797 29415 77813
rect 29381 77747 29415 77763
rect 29717 77797 29751 77813
rect 29717 77747 29751 77763
rect 30053 77797 30087 77813
rect 30053 77747 30087 77763
rect 30389 77797 30423 77813
rect 30389 77747 30423 77763
rect 30725 77797 30759 77813
rect 30725 77747 30759 77763
rect 31061 77797 31095 77813
rect 31061 77747 31095 77763
rect 31397 77797 31431 77813
rect 31397 77747 31431 77763
rect 31733 77797 31767 77813
rect 31733 77747 31767 77763
rect 32069 77797 32103 77813
rect 32069 77747 32103 77763
rect 32405 77797 32439 77813
rect 32405 77747 32439 77763
rect 32741 77797 32775 77813
rect 32741 77747 32775 77763
rect 33077 77797 33111 77813
rect 33077 77747 33111 77763
rect 33413 77797 33447 77813
rect 33413 77747 33447 77763
rect 33749 77797 33783 77813
rect 33749 77747 33783 77763
rect 34085 77797 34119 77813
rect 34085 77747 34119 77763
rect 34421 77797 34455 77813
rect 34421 77747 34455 77763
rect 34757 77797 34791 77813
rect 34757 77747 34791 77763
rect 35093 77797 35127 77813
rect 35093 77747 35127 77763
rect 35429 77797 35463 77813
rect 35429 77747 35463 77763
rect 35765 77797 35799 77813
rect 35765 77747 35799 77763
rect 36101 77797 36135 77813
rect 36101 77747 36135 77763
rect 36437 77797 36471 77813
rect 36437 77747 36471 77763
rect 36773 77797 36807 77813
rect 36773 77747 36807 77763
rect 37109 77797 37143 77813
rect 37109 77747 37143 77763
rect 37445 77797 37479 77813
rect 37445 77747 37479 77763
rect 37781 77797 37815 77813
rect 37781 77747 37815 77763
rect 38117 77797 38151 77813
rect 38117 77747 38151 77763
rect 38453 77797 38487 77813
rect 38453 77747 38487 77763
rect 38789 77797 38823 77813
rect 38789 77747 38823 77763
rect 39125 77797 39159 77813
rect 39125 77747 39159 77763
rect 39461 77797 39495 77813
rect 39461 77747 39495 77763
rect 39797 77797 39831 77813
rect 39797 77747 39831 77763
rect 40133 77797 40167 77813
rect 40133 77747 40167 77763
rect 40469 77797 40503 77813
rect 40469 77747 40503 77763
rect 40805 77797 40839 77813
rect 40805 77747 40839 77763
rect 41141 77797 41175 77813
rect 41141 77747 41175 77763
rect 41477 77797 41511 77813
rect 41477 77747 41511 77763
rect 41813 77797 41847 77813
rect 41813 77747 41847 77763
rect 42149 77797 42183 77813
rect 42149 77747 42183 77763
rect 42485 77797 42519 77813
rect 42485 77747 42519 77763
rect 42821 77797 42855 77813
rect 42821 77747 42855 77763
rect 43157 77797 43191 77813
rect 43157 77747 43191 77763
rect 43493 77797 43527 77813
rect 43493 77747 43527 77763
rect 43829 77797 43863 77813
rect 43829 77747 43863 77763
rect 44165 77797 44199 77813
rect 44165 77747 44199 77763
rect 44501 77797 44535 77813
rect 44501 77747 44535 77763
rect 44837 77797 44871 77813
rect 44837 77747 44871 77763
rect 45173 77797 45207 77813
rect 45173 77747 45207 77763
rect 45509 77797 45543 77813
rect 45509 77747 45543 77763
rect 45845 77797 45879 77813
rect 45845 77747 45879 77763
rect 46181 77797 46215 77813
rect 46181 77747 46215 77763
rect 46517 77797 46551 77813
rect 46517 77747 46551 77763
rect 46853 77797 46887 77813
rect 46853 77747 46887 77763
rect 47189 77797 47223 77813
rect 47189 77747 47223 77763
rect 47525 77797 47559 77813
rect 47525 77747 47559 77763
rect 47861 77797 47895 77813
rect 47861 77747 47895 77763
rect 48197 77797 48231 77813
rect 48197 77747 48231 77763
rect 48533 77797 48567 77813
rect 48533 77747 48567 77763
rect 48869 77797 48903 77813
rect 48869 77747 48903 77763
rect 49205 77797 49239 77813
rect 49205 77747 49239 77763
rect 49541 77797 49575 77813
rect 49541 77747 49575 77763
rect 49877 77797 49911 77813
rect 49877 77747 49911 77763
rect 50213 77797 50247 77813
rect 50213 77747 50247 77763
rect 50549 77797 50583 77813
rect 50549 77747 50583 77763
rect 50885 77797 50919 77813
rect 50885 77747 50919 77763
rect 51221 77797 51255 77813
rect 51221 77747 51255 77763
rect 51557 77797 51591 77813
rect 51557 77747 51591 77763
rect 51893 77797 51927 77813
rect 51893 77747 51927 77763
rect 52229 77797 52263 77813
rect 52229 77747 52263 77763
rect 52565 77797 52599 77813
rect 52565 77747 52599 77763
rect 52901 77797 52935 77813
rect 52901 77747 52935 77763
rect 53237 77797 53271 77813
rect 53237 77747 53271 77763
rect 53573 77797 53607 77813
rect 53573 77747 53607 77763
rect 53909 77797 53943 77813
rect 53909 77747 53943 77763
rect 54245 77797 54279 77813
rect 54245 77747 54279 77763
rect 54581 77797 54615 77813
rect 54581 77747 54615 77763
rect 54917 77797 54951 77813
rect 54917 77747 54951 77763
rect 55253 77797 55287 77813
rect 55253 77747 55287 77763
rect 55589 77797 55623 77813
rect 55589 77747 55623 77763
rect 55925 77797 55959 77813
rect 55925 77747 55959 77763
rect 56261 77797 56295 77813
rect 56261 77747 56295 77763
rect 56597 77797 56631 77813
rect 56597 77747 56631 77763
rect 56933 77797 56967 77813
rect 56933 77747 56967 77763
rect 57269 77797 57303 77813
rect 57269 77747 57303 77763
rect 57605 77797 57639 77813
rect 57605 77747 57639 77763
rect 57941 77797 57975 77813
rect 57941 77747 57975 77763
rect 58277 77797 58311 77813
rect 58277 77747 58311 77763
rect 58613 77797 58647 77813
rect 58613 77747 58647 77763
rect 58949 77797 58983 77813
rect 58949 77747 58983 77763
rect 59285 77797 59319 77813
rect 59285 77747 59319 77763
rect 59621 77797 59655 77813
rect 59621 77747 59655 77763
rect 59957 77797 59991 77813
rect 59957 77747 59991 77763
rect 60293 77797 60327 77813
rect 60293 77747 60327 77763
rect 60629 77797 60663 77813
rect 60629 77747 60663 77763
rect 60965 77797 60999 77813
rect 60965 77747 60999 77763
rect 61301 77797 61335 77813
rect 61301 77747 61335 77763
rect 61637 77797 61671 77813
rect 61637 77747 61671 77763
rect 61973 77797 62007 77813
rect 61973 77747 62007 77763
rect 62309 77797 62343 77813
rect 62309 77747 62343 77763
rect 62645 77797 62679 77813
rect 62645 77747 62679 77763
rect 62981 77797 63015 77813
rect 62981 77747 63015 77763
rect 63317 77797 63351 77813
rect 63317 77747 63351 77763
rect 63653 77797 63687 77813
rect 63653 77747 63687 77763
rect 63989 77797 64023 77813
rect 63989 77747 64023 77763
rect 64325 77797 64359 77813
rect 64325 77747 64359 77763
rect 64661 77797 64695 77813
rect 64661 77747 64695 77763
rect 64997 77797 65031 77813
rect 64997 77747 65031 77763
rect 65333 77797 65367 77813
rect 65333 77747 65367 77763
rect 65669 77797 65703 77813
rect 65669 77747 65703 77763
rect 66005 77797 66039 77813
rect 66005 77747 66039 77763
rect 66341 77797 66375 77813
rect 66341 77747 66375 77763
rect 66677 77797 66711 77813
rect 66677 77747 66711 77763
rect 67013 77797 67047 77813
rect 67013 77747 67047 77763
rect 67349 77797 67383 77813
rect 67349 77747 67383 77763
rect 67685 77797 67719 77813
rect 67685 77747 67719 77763
rect 68021 77797 68055 77813
rect 68021 77747 68055 77763
rect 68357 77797 68391 77813
rect 68357 77747 68391 77763
rect 68693 77797 68727 77813
rect 68693 77747 68727 77763
rect 69029 77797 69063 77813
rect 69029 77747 69063 77763
rect 69365 77797 69399 77813
rect 69365 77747 69399 77763
rect 69701 77797 69735 77813
rect 69701 77747 69735 77763
rect 70037 77797 70071 77813
rect 70037 77747 70071 77763
rect 70373 77797 70407 77813
rect 70373 77747 70407 77763
rect 70709 77797 70743 77813
rect 70709 77747 70743 77763
rect 71045 77797 71079 77813
rect 71045 77747 71079 77763
rect 71381 77797 71415 77813
rect 71381 77747 71415 77763
rect 71717 77797 71751 77813
rect 71717 77747 71751 77763
rect 72053 77797 72087 77813
rect 72053 77747 72087 77763
rect 72389 77797 72423 77813
rect 72389 77747 72423 77763
rect 72725 77797 72759 77813
rect 72725 77747 72759 77763
rect 73061 77797 73095 77813
rect 73061 77747 73095 77763
rect 73397 77797 73431 77813
rect 73397 77747 73431 77763
rect 73733 77797 73767 77813
rect 73733 77747 73767 77763
rect 74069 77797 74103 77813
rect 74069 77747 74103 77763
rect 74405 77797 74439 77813
rect 74405 77747 74439 77763
rect 74741 77797 74775 77813
rect 74741 77747 74775 77763
rect 75077 77797 75111 77813
rect 75077 77747 75111 77763
rect 75413 77797 75447 77813
rect 75413 77747 75447 77763
rect 75749 77797 75783 77813
rect 75749 77747 75783 77763
rect 76085 77797 76119 77813
rect 76085 77747 76119 77763
rect 76421 77797 76455 77813
rect 76421 77747 76455 77763
rect 76757 77797 76791 77813
rect 76757 77747 76791 77763
rect 77093 77797 77127 77813
rect 77093 77747 77127 77763
rect 77429 77797 77463 77813
rect 77429 77747 77463 77763
rect 77765 77797 77799 77813
rect 77765 77747 77799 77763
rect 78101 77797 78135 77813
rect 78101 77747 78135 77763
rect 78437 77797 78471 77813
rect 78437 77747 78471 77763
rect 78773 77797 78807 77813
rect 78773 77747 78807 77763
rect 79109 77797 79143 77813
rect 79109 77747 79143 77763
rect 79445 77797 79479 77813
rect 79445 77747 79479 77763
rect 79781 77797 79815 77813
rect 79781 77747 79815 77763
rect 80117 77797 80151 77813
rect 80117 77747 80151 77763
rect 80453 77797 80487 77813
rect 80453 77747 80487 77763
rect 80789 77797 80823 77813
rect 80789 77747 80823 77763
rect 81125 77797 81159 77813
rect 81125 77747 81159 77763
rect 81461 77797 81495 77813
rect 81461 77747 81495 77763
rect 81797 77797 81831 77813
rect 81797 77747 81831 77763
rect 82133 77797 82167 77813
rect 82133 77747 82167 77763
rect 82469 77797 82503 77813
rect 82469 77747 82503 77763
rect 82805 77797 82839 77813
rect 82805 77747 82839 77763
rect 83141 77797 83175 77813
rect 83141 77747 83175 77763
rect 83477 77797 83511 77813
rect 83477 77747 83511 77763
rect 83813 77797 83847 77813
rect 83813 77747 83847 77763
rect 84149 77797 84183 77813
rect 84149 77747 84183 77763
rect 84485 77797 84519 77813
rect 84485 77747 84519 77763
rect 84821 77797 84855 77813
rect 84821 77747 84855 77763
rect 85157 77797 85191 77813
rect 85157 77747 85191 77763
rect 85493 77797 85527 77813
rect 85493 77747 85527 77763
rect 85829 77797 85863 77813
rect 85829 77747 85863 77763
rect 86165 77797 86199 77813
rect 86165 77747 86199 77763
rect 86501 77797 86535 77813
rect 86501 77747 86535 77763
rect 86837 77797 86871 77813
rect 86837 77747 86871 77763
rect 87173 77797 87207 77813
rect 87173 77747 87207 77763
rect 87509 77797 87543 77813
rect 87509 77747 87543 77763
rect 87845 77797 87879 77813
rect 87845 77747 87879 77763
rect 88181 77797 88215 77813
rect 88181 77747 88215 77763
rect 88517 77797 88551 77813
rect 88517 77747 88551 77763
rect 88853 77797 88887 77813
rect 88853 77747 88887 77763
rect 89189 77797 89223 77813
rect 89189 77747 89223 77763
rect 89525 77797 89559 77813
rect 89525 77747 89559 77763
rect 89861 77797 89895 77813
rect 89861 77747 89895 77763
rect 90197 77797 90231 77813
rect 90197 77747 90231 77763
rect 90533 77797 90567 77813
rect 90533 77747 90567 77763
rect 90869 77797 90903 77813
rect 90869 77747 90903 77763
rect 91205 77797 91239 77813
rect 91205 77747 91239 77763
rect 91541 77797 91575 77813
rect 91541 77747 91575 77763
rect 91877 77797 91911 77813
rect 91877 77747 91911 77763
rect 92213 77797 92247 77813
rect 92213 77747 92247 77763
rect 92549 77797 92583 77813
rect 92549 77747 92583 77763
rect 92885 77797 92919 77813
rect 92885 77747 92919 77763
rect 93221 77797 93255 77813
rect 93221 77747 93255 77763
rect 93557 77797 93591 77813
rect 93557 77747 93591 77763
rect 1829 77333 1863 77349
rect 1829 77283 1863 77299
rect 94187 77333 94221 77349
rect 94187 77283 94221 77299
rect 1829 76997 1863 77013
rect 1829 76947 1863 76963
rect 94187 76997 94221 77013
rect 94187 76947 94221 76963
rect 1829 76661 1863 76677
rect 1829 76611 1863 76627
rect 94187 76661 94221 76677
rect 94187 76611 94221 76627
rect 1829 76325 1863 76341
rect 1829 76275 1863 76291
rect 94187 76325 94221 76341
rect 94187 76275 94221 76291
rect 1829 75989 1863 76005
rect 1829 75939 1863 75955
rect 94187 75989 94221 76005
rect 94187 75939 94221 75955
rect 1829 75653 1863 75669
rect 1829 75603 1863 75619
rect 94187 75653 94221 75669
rect 94187 75603 94221 75619
rect 1829 75317 1863 75333
rect 1829 75267 1863 75283
rect 94187 75317 94221 75333
rect 94187 75267 94221 75283
rect 1829 74981 1863 74997
rect 1829 74931 1863 74947
rect 94187 74981 94221 74997
rect 94187 74931 94221 74947
rect 1829 74645 1863 74661
rect 1829 74595 1863 74611
rect 94187 74645 94221 74661
rect 94187 74595 94221 74611
rect 1829 74309 1863 74325
rect 1829 74259 1863 74275
rect 94187 74309 94221 74325
rect 94187 74259 94221 74275
rect 1829 73973 1863 73989
rect 1829 73923 1863 73939
rect 94187 73973 94221 73989
rect 94187 73923 94221 73939
rect 1829 73637 1863 73653
rect 1829 73587 1863 73603
rect 94187 73637 94221 73653
rect 94187 73587 94221 73603
rect 1829 73301 1863 73317
rect 1829 73251 1863 73267
rect 94187 73301 94221 73317
rect 94187 73251 94221 73267
rect 1829 72965 1863 72981
rect 1829 72915 1863 72931
rect 94187 72965 94221 72981
rect 94187 72915 94221 72931
rect 1829 72629 1863 72645
rect 1829 72579 1863 72595
rect 94187 72629 94221 72645
rect 94187 72579 94221 72595
rect 1829 72293 1863 72309
rect 1829 72243 1863 72259
rect 94187 72293 94221 72309
rect 94187 72243 94221 72259
rect 1829 71957 1863 71973
rect 1829 71907 1863 71923
rect 94187 71957 94221 71973
rect 94187 71907 94221 71923
rect 1829 71621 1863 71637
rect 1829 71571 1863 71587
rect 94187 71621 94221 71637
rect 94187 71571 94221 71587
rect 1829 71285 1863 71301
rect 1829 71235 1863 71251
rect 94187 71285 94221 71301
rect 94187 71235 94221 71251
rect 1829 70949 1863 70965
rect 1829 70899 1863 70915
rect 94187 70949 94221 70965
rect 94187 70899 94221 70915
rect 1829 70613 1863 70629
rect 1829 70563 1863 70579
rect 94187 70613 94221 70629
rect 94187 70563 94221 70579
rect 1829 70277 1863 70293
rect 1829 70227 1863 70243
rect 94187 70277 94221 70293
rect 94187 70227 94221 70243
rect 1829 69941 1863 69957
rect 1829 69891 1863 69907
rect 94187 69941 94221 69957
rect 94187 69891 94221 69907
rect 1829 69605 1863 69621
rect 1829 69555 1863 69571
rect 94187 69605 94221 69621
rect 94187 69555 94221 69571
rect 1829 69269 1863 69285
rect 1829 69219 1863 69235
rect 94187 69269 94221 69285
rect 94187 69219 94221 69235
rect 1829 68933 1863 68949
rect 1829 68883 1863 68899
rect 94187 68933 94221 68949
rect 94187 68883 94221 68899
rect 1829 68597 1863 68613
rect 1829 68547 1863 68563
rect 94187 68597 94221 68613
rect 94187 68547 94221 68563
rect 1829 68261 1863 68277
rect 1829 68211 1863 68227
rect 94187 68261 94221 68277
rect 94187 68211 94221 68227
rect 1829 67925 1863 67941
rect 1829 67875 1863 67891
rect 94187 67925 94221 67941
rect 94187 67875 94221 67891
rect 1829 67589 1863 67605
rect 1829 67539 1863 67555
rect 94187 67589 94221 67605
rect 94187 67539 94221 67555
rect 1829 67253 1863 67269
rect 1829 67203 1863 67219
rect 94187 67253 94221 67269
rect 94187 67203 94221 67219
rect 1829 66917 1863 66933
rect 1829 66867 1863 66883
rect 94187 66917 94221 66933
rect 94187 66867 94221 66883
rect 1829 66581 1863 66597
rect 1829 66531 1863 66547
rect 94187 66581 94221 66597
rect 94187 66531 94221 66547
rect 1829 66245 1863 66261
rect 1829 66195 1863 66211
rect 94187 66245 94221 66261
rect 94187 66195 94221 66211
rect 1829 65909 1863 65925
rect 1829 65859 1863 65875
rect 94187 65909 94221 65925
rect 94187 65859 94221 65875
rect 1829 65573 1863 65589
rect 1829 65523 1863 65539
rect 94187 65573 94221 65589
rect 94187 65523 94221 65539
rect 1829 65237 1863 65253
rect 1829 65187 1863 65203
rect 94187 65237 94221 65253
rect 94187 65187 94221 65203
rect 1829 64901 1863 64917
rect 1829 64851 1863 64867
rect 94187 64901 94221 64917
rect 94187 64851 94221 64867
rect 1829 64565 1863 64581
rect 1829 64515 1863 64531
rect 94187 64565 94221 64581
rect 94187 64515 94221 64531
rect 1829 64229 1863 64245
rect 1829 64179 1863 64195
rect 94187 64229 94221 64245
rect 94187 64179 94221 64195
rect 1829 63893 1863 63909
rect 1829 63843 1863 63859
rect 94187 63893 94221 63909
rect 94187 63843 94221 63859
rect 1829 63557 1863 63573
rect 1829 63507 1863 63523
rect 94187 63557 94221 63573
rect 94187 63507 94221 63523
rect 1829 63221 1863 63237
rect 1829 63171 1863 63187
rect 94187 63221 94221 63237
rect 94187 63171 94221 63187
rect 1829 62885 1863 62901
rect 1829 62835 1863 62851
rect 94187 62885 94221 62901
rect 94187 62835 94221 62851
rect 1829 62549 1863 62565
rect 1829 62499 1863 62515
rect 94187 62549 94221 62565
rect 94187 62499 94221 62515
rect 1829 62213 1863 62229
rect 1829 62163 1863 62179
rect 94187 62213 94221 62229
rect 94187 62163 94221 62179
rect 1829 61877 1863 61893
rect 1829 61827 1863 61843
rect 94187 61877 94221 61893
rect 94187 61827 94221 61843
rect 1829 61541 1863 61557
rect 1829 61491 1863 61507
rect 94187 61541 94221 61557
rect 94187 61491 94221 61507
rect 1829 61205 1863 61221
rect 1829 61155 1863 61171
rect 94187 61205 94221 61221
rect 94187 61155 94221 61171
rect 1829 60869 1863 60885
rect 1829 60819 1863 60835
rect 94187 60869 94221 60885
rect 94187 60819 94221 60835
rect 1829 60533 1863 60549
rect 1829 60483 1863 60499
rect 94187 60533 94221 60549
rect 94187 60483 94221 60499
rect 1829 60197 1863 60213
rect 1829 60147 1863 60163
rect 94187 60197 94221 60213
rect 94187 60147 94221 60163
rect 1829 59861 1863 59877
rect 1829 59811 1863 59827
rect 94187 59861 94221 59877
rect 94187 59811 94221 59827
rect 1829 59525 1863 59541
rect 1829 59475 1863 59491
rect 94187 59525 94221 59541
rect 94187 59475 94221 59491
rect 1829 59189 1863 59205
rect 1829 59139 1863 59155
rect 94187 59189 94221 59205
rect 94187 59139 94221 59155
rect 1829 58853 1863 58869
rect 1829 58803 1863 58819
rect 94187 58853 94221 58869
rect 94187 58803 94221 58819
rect 1829 58517 1863 58533
rect 1829 58467 1863 58483
rect 94187 58517 94221 58533
rect 94187 58467 94221 58483
rect 1829 58181 1863 58197
rect 1829 58131 1863 58147
rect 94187 58181 94221 58197
rect 94187 58131 94221 58147
rect 1829 57845 1863 57861
rect 1829 57795 1863 57811
rect 94187 57845 94221 57861
rect 94187 57795 94221 57811
rect 1829 57509 1863 57525
rect 1829 57459 1863 57475
rect 94187 57509 94221 57525
rect 94187 57459 94221 57475
rect 1829 57173 1863 57189
rect 1829 57123 1863 57139
rect 94187 57173 94221 57189
rect 94187 57123 94221 57139
rect 1829 56837 1863 56853
rect 1829 56787 1863 56803
rect 94187 56837 94221 56853
rect 94187 56787 94221 56803
rect 1829 56501 1863 56517
rect 1829 56451 1863 56467
rect 94187 56501 94221 56517
rect 94187 56451 94221 56467
rect 1829 56165 1863 56181
rect 1829 56115 1863 56131
rect 94187 56165 94221 56181
rect 94187 56115 94221 56131
rect 1829 55829 1863 55845
rect 1829 55779 1863 55795
rect 94187 55829 94221 55845
rect 94187 55779 94221 55795
rect 1829 55493 1863 55509
rect 1829 55443 1863 55459
rect 94187 55493 94221 55509
rect 94187 55443 94221 55459
rect 1829 55157 1863 55173
rect 1829 55107 1863 55123
rect 94187 55157 94221 55173
rect 94187 55107 94221 55123
rect 1829 54821 1863 54837
rect 1829 54771 1863 54787
rect 94187 54821 94221 54837
rect 94187 54771 94221 54787
rect 1829 54485 1863 54501
rect 1829 54435 1863 54451
rect 94187 54485 94221 54501
rect 94187 54435 94221 54451
rect 1829 54149 1863 54165
rect 1829 54099 1863 54115
rect 94187 54149 94221 54165
rect 94187 54099 94221 54115
rect 1829 53813 1863 53829
rect 1829 53763 1863 53779
rect 94187 53813 94221 53829
rect 94187 53763 94221 53779
rect 1829 53477 1863 53493
rect 1829 53427 1863 53443
rect 94187 53477 94221 53493
rect 94187 53427 94221 53443
rect 1829 53141 1863 53157
rect 1829 53091 1863 53107
rect 94187 53141 94221 53157
rect 94187 53091 94221 53107
rect 1829 52805 1863 52821
rect 1829 52755 1863 52771
rect 94187 52805 94221 52821
rect 94187 52755 94221 52771
rect 1829 52469 1863 52485
rect 1829 52419 1863 52435
rect 94187 52469 94221 52485
rect 94187 52419 94221 52435
rect 1829 52133 1863 52149
rect 1829 52083 1863 52099
rect 94187 52133 94221 52149
rect 94187 52083 94221 52099
rect 1829 51797 1863 51813
rect 1829 51747 1863 51763
rect 94187 51797 94221 51813
rect 94187 51747 94221 51763
rect 1829 51461 1863 51477
rect 1829 51411 1863 51427
rect 94187 51461 94221 51477
rect 94187 51411 94221 51427
rect 1829 51125 1863 51141
rect 1829 51075 1863 51091
rect 94187 51125 94221 51141
rect 94187 51075 94221 51091
rect 1829 50789 1863 50805
rect 1829 50739 1863 50755
rect 94187 50789 94221 50805
rect 94187 50739 94221 50755
rect 1829 50453 1863 50469
rect 1829 50403 1863 50419
rect 94187 50453 94221 50469
rect 94187 50403 94221 50419
rect 1829 50117 1863 50133
rect 1829 50067 1863 50083
rect 94187 50117 94221 50133
rect 94187 50067 94221 50083
rect 1829 49781 1863 49797
rect 1829 49731 1863 49747
rect 94187 49781 94221 49797
rect 94187 49731 94221 49747
rect 1829 49445 1863 49461
rect 1829 49395 1863 49411
rect 94187 49445 94221 49461
rect 94187 49395 94221 49411
rect 1829 49109 1863 49125
rect 1829 49059 1863 49075
rect 94187 49109 94221 49125
rect 94187 49059 94221 49075
rect 1829 48773 1863 48789
rect 1829 48723 1863 48739
rect 94187 48773 94221 48789
rect 94187 48723 94221 48739
rect 1829 48437 1863 48453
rect 1829 48387 1863 48403
rect 94187 48437 94221 48453
rect 94187 48387 94221 48403
rect 1829 48101 1863 48117
rect 1829 48051 1863 48067
rect 94187 48101 94221 48117
rect 94187 48051 94221 48067
rect 1829 47765 1863 47781
rect 1829 47715 1863 47731
rect 94187 47765 94221 47781
rect 94187 47715 94221 47731
rect 1829 47429 1863 47445
rect 1829 47379 1863 47395
rect 94187 47429 94221 47445
rect 94187 47379 94221 47395
rect 1829 47093 1863 47109
rect 1829 47043 1863 47059
rect 94187 47093 94221 47109
rect 94187 47043 94221 47059
rect 1829 46757 1863 46773
rect 1829 46707 1863 46723
rect 94187 46757 94221 46773
rect 94187 46707 94221 46723
rect 1829 46421 1863 46437
rect 1829 46371 1863 46387
rect 94187 46421 94221 46437
rect 94187 46371 94221 46387
rect 1829 46085 1863 46101
rect 1829 46035 1863 46051
rect 94187 46085 94221 46101
rect 94187 46035 94221 46051
rect 1829 45749 1863 45765
rect 1829 45699 1863 45715
rect 94187 45749 94221 45765
rect 94187 45699 94221 45715
rect 1829 45413 1863 45429
rect 1829 45363 1863 45379
rect 94187 45413 94221 45429
rect 94187 45363 94221 45379
rect 1829 45077 1863 45093
rect 1829 45027 1863 45043
rect 94187 45077 94221 45093
rect 94187 45027 94221 45043
rect 1829 44741 1863 44757
rect 1829 44691 1863 44707
rect 94187 44741 94221 44757
rect 94187 44691 94221 44707
rect 1829 44405 1863 44421
rect 1829 44355 1863 44371
rect 94187 44405 94221 44421
rect 94187 44355 94221 44371
rect 1829 44069 1863 44085
rect 1829 44019 1863 44035
rect 94187 44069 94221 44085
rect 94187 44019 94221 44035
rect 1829 43733 1863 43749
rect 1829 43683 1863 43699
rect 94187 43733 94221 43749
rect 94187 43683 94221 43699
rect 1829 43397 1863 43413
rect 1829 43347 1863 43363
rect 94187 43397 94221 43413
rect 94187 43347 94221 43363
rect 1829 43061 1863 43077
rect 1829 43011 1863 43027
rect 94187 43061 94221 43077
rect 94187 43011 94221 43027
rect 1829 42725 1863 42741
rect 1829 42675 1863 42691
rect 94187 42725 94221 42741
rect 94187 42675 94221 42691
rect 1829 42389 1863 42405
rect 1829 42339 1863 42355
rect 94187 42389 94221 42405
rect 94187 42339 94221 42355
rect 1829 42053 1863 42069
rect 1829 42003 1863 42019
rect 94187 42053 94221 42069
rect 94187 42003 94221 42019
rect 1829 41717 1863 41733
rect 1829 41667 1863 41683
rect 94187 41717 94221 41733
rect 94187 41667 94221 41683
rect 1829 41381 1863 41397
rect 1829 41331 1863 41347
rect 94187 41381 94221 41397
rect 94187 41331 94221 41347
rect 1829 41045 1863 41061
rect 1829 40995 1863 41011
rect 94187 41045 94221 41061
rect 94187 40995 94221 41011
rect 1829 40709 1863 40725
rect 1829 40659 1863 40675
rect 94187 40709 94221 40725
rect 94187 40659 94221 40675
rect 1829 40373 1863 40389
rect 1829 40323 1863 40339
rect 94187 40373 94221 40389
rect 94187 40323 94221 40339
rect 1829 40037 1863 40053
rect 1829 39987 1863 40003
rect 94187 40037 94221 40053
rect 94187 39987 94221 40003
rect 1829 39701 1863 39717
rect 1829 39651 1863 39667
rect 94187 39701 94221 39717
rect 94187 39651 94221 39667
rect 1829 39365 1863 39381
rect 1829 39315 1863 39331
rect 94187 39365 94221 39381
rect 94187 39315 94221 39331
rect 1829 39029 1863 39045
rect 1829 38979 1863 38995
rect 94187 39029 94221 39045
rect 94187 38979 94221 38995
rect 1829 38693 1863 38709
rect 1829 38643 1863 38659
rect 94187 38693 94221 38709
rect 94187 38643 94221 38659
rect 1829 38357 1863 38373
rect 1829 38307 1863 38323
rect 94187 38357 94221 38373
rect 94187 38307 94221 38323
rect 1829 38021 1863 38037
rect 1829 37971 1863 37987
rect 94187 38021 94221 38037
rect 94187 37971 94221 37987
rect 1829 37685 1863 37701
rect 1829 37635 1863 37651
rect 94187 37685 94221 37701
rect 94187 37635 94221 37651
rect 1829 37349 1863 37365
rect 1829 37299 1863 37315
rect 94187 37349 94221 37365
rect 94187 37299 94221 37315
rect 1829 37013 1863 37029
rect 1829 36963 1863 36979
rect 94187 37013 94221 37029
rect 94187 36963 94221 36979
rect 1829 36677 1863 36693
rect 1829 36627 1863 36643
rect 94187 36677 94221 36693
rect 94187 36627 94221 36643
rect 1829 36341 1863 36357
rect 1829 36291 1863 36307
rect 94187 36341 94221 36357
rect 94187 36291 94221 36307
rect 1829 36005 1863 36021
rect 1829 35955 1863 35971
rect 94187 36005 94221 36021
rect 94187 35955 94221 35971
rect 1829 35669 1863 35685
rect 1829 35619 1863 35635
rect 94187 35669 94221 35685
rect 94187 35619 94221 35635
rect 1829 35333 1863 35349
rect 1829 35283 1863 35299
rect 94187 35333 94221 35349
rect 94187 35283 94221 35299
rect 1829 34997 1863 35013
rect 1829 34947 1863 34963
rect 94187 34997 94221 35013
rect 94187 34947 94221 34963
rect 1829 34661 1863 34677
rect 1829 34611 1863 34627
rect 94187 34661 94221 34677
rect 94187 34611 94221 34627
rect 1829 34325 1863 34341
rect 1829 34275 1863 34291
rect 94187 34325 94221 34341
rect 94187 34275 94221 34291
rect 1829 33989 1863 34005
rect 1829 33939 1863 33955
rect 94187 33989 94221 34005
rect 94187 33939 94221 33955
rect 1829 33653 1863 33669
rect 1829 33603 1863 33619
rect 94187 33653 94221 33669
rect 94187 33603 94221 33619
rect 1829 33317 1863 33333
rect 1829 33267 1863 33283
rect 94187 33317 94221 33333
rect 94187 33267 94221 33283
rect 1829 32981 1863 32997
rect 1829 32931 1863 32947
rect 94187 32981 94221 32997
rect 94187 32931 94221 32947
rect 1829 32645 1863 32661
rect 1829 32595 1863 32611
rect 94187 32645 94221 32661
rect 94187 32595 94221 32611
rect 1829 32309 1863 32325
rect 1829 32259 1863 32275
rect 94187 32309 94221 32325
rect 94187 32259 94221 32275
rect 1829 31973 1863 31989
rect 1829 31923 1863 31939
rect 94187 31973 94221 31989
rect 94187 31923 94221 31939
rect 1829 31637 1863 31653
rect 1829 31587 1863 31603
rect 94187 31637 94221 31653
rect 94187 31587 94221 31603
rect 1829 31301 1863 31317
rect 1829 31251 1863 31267
rect 94187 31301 94221 31317
rect 94187 31251 94221 31267
rect 1829 30965 1863 30981
rect 1829 30915 1863 30931
rect 94187 30965 94221 30981
rect 94187 30915 94221 30931
rect 1829 30629 1863 30645
rect 1829 30579 1863 30595
rect 94187 30629 94221 30645
rect 94187 30579 94221 30595
rect 1829 30293 1863 30309
rect 1829 30243 1863 30259
rect 94187 30293 94221 30309
rect 94187 30243 94221 30259
rect 1829 29957 1863 29973
rect 1829 29907 1863 29923
rect 94187 29957 94221 29973
rect 94187 29907 94221 29923
rect 1829 29621 1863 29637
rect 1829 29571 1863 29587
rect 94187 29621 94221 29637
rect 94187 29571 94221 29587
rect 1829 29285 1863 29301
rect 1829 29235 1863 29251
rect 94187 29285 94221 29301
rect 94187 29235 94221 29251
rect 1829 28949 1863 28965
rect 1829 28899 1863 28915
rect 94187 28949 94221 28965
rect 94187 28899 94221 28915
rect 1829 28613 1863 28629
rect 1829 28563 1863 28579
rect 94187 28613 94221 28629
rect 94187 28563 94221 28579
rect 1829 28277 1863 28293
rect 1829 28227 1863 28243
rect 94187 28277 94221 28293
rect 94187 28227 94221 28243
rect 1829 27941 1863 27957
rect 1829 27891 1863 27907
rect 94187 27941 94221 27957
rect 94187 27891 94221 27907
rect 1829 27605 1863 27621
rect 1829 27555 1863 27571
rect 94187 27605 94221 27621
rect 94187 27555 94221 27571
rect 1829 27269 1863 27285
rect 1829 27219 1863 27235
rect 94187 27269 94221 27285
rect 94187 27219 94221 27235
rect 1829 26933 1863 26949
rect 1829 26883 1863 26899
rect 94187 26933 94221 26949
rect 94187 26883 94221 26899
rect 1829 26597 1863 26613
rect 1829 26547 1863 26563
rect 94187 26597 94221 26613
rect 94187 26547 94221 26563
rect 1829 26261 1863 26277
rect 1829 26211 1863 26227
rect 94187 26261 94221 26277
rect 94187 26211 94221 26227
rect 1829 25925 1863 25941
rect 1829 25875 1863 25891
rect 94187 25925 94221 25941
rect 94187 25875 94221 25891
rect 1829 25589 1863 25605
rect 1829 25539 1863 25555
rect 94187 25589 94221 25605
rect 94187 25539 94221 25555
rect 1829 25253 1863 25269
rect 1829 25203 1863 25219
rect 94187 25253 94221 25269
rect 94187 25203 94221 25219
rect 1829 24917 1863 24933
rect 1829 24867 1863 24883
rect 94187 24917 94221 24933
rect 94187 24867 94221 24883
rect 1829 24581 1863 24597
rect 1829 24531 1863 24547
rect 94187 24581 94221 24597
rect 94187 24531 94221 24547
rect 1829 24245 1863 24261
rect 1829 24195 1863 24211
rect 94187 24245 94221 24261
rect 94187 24195 94221 24211
rect 1829 23909 1863 23925
rect 1829 23859 1863 23875
rect 94187 23909 94221 23925
rect 94187 23859 94221 23875
rect 1829 23573 1863 23589
rect 1829 23523 1863 23539
rect 94187 23573 94221 23589
rect 94187 23523 94221 23539
rect 1829 23237 1863 23253
rect 1829 23187 1863 23203
rect 94187 23237 94221 23253
rect 94187 23187 94221 23203
rect 1829 22901 1863 22917
rect 1829 22851 1863 22867
rect 94187 22901 94221 22917
rect 94187 22851 94221 22867
rect 1829 22565 1863 22581
rect 1829 22515 1863 22531
rect 94187 22565 94221 22581
rect 94187 22515 94221 22531
rect 1829 22229 1863 22245
rect 1829 22179 1863 22195
rect 94187 22229 94221 22245
rect 94187 22179 94221 22195
rect 1829 21893 1863 21909
rect 1829 21843 1863 21859
rect 94187 21893 94221 21909
rect 94187 21843 94221 21859
rect 1829 21557 1863 21573
rect 1829 21507 1863 21523
rect 94187 21557 94221 21573
rect 94187 21507 94221 21523
rect 1829 21221 1863 21237
rect 1829 21171 1863 21187
rect 94187 21221 94221 21237
rect 94187 21171 94221 21187
rect 1829 20885 1863 20901
rect 1829 20835 1863 20851
rect 94187 20885 94221 20901
rect 94187 20835 94221 20851
rect 1829 20549 1863 20565
rect 1829 20499 1863 20515
rect 94187 20549 94221 20565
rect 94187 20499 94221 20515
rect 1829 20213 1863 20229
rect 1829 20163 1863 20179
rect 94187 20213 94221 20229
rect 94187 20163 94221 20179
rect 1829 19877 1863 19893
rect 1829 19827 1863 19843
rect 94187 19877 94221 19893
rect 94187 19827 94221 19843
rect 1829 19541 1863 19557
rect 1829 19491 1863 19507
rect 94187 19541 94221 19557
rect 94187 19491 94221 19507
rect 1829 19205 1863 19221
rect 1829 19155 1863 19171
rect 94187 19205 94221 19221
rect 94187 19155 94221 19171
rect 1829 18869 1863 18885
rect 1829 18819 1863 18835
rect 94187 18869 94221 18885
rect 94187 18819 94221 18835
rect 1829 18533 1863 18549
rect 1829 18483 1863 18499
rect 94187 18533 94221 18549
rect 94187 18483 94221 18499
rect 1829 18197 1863 18213
rect 1829 18147 1863 18163
rect 94187 18197 94221 18213
rect 94187 18147 94221 18163
rect 1829 17861 1863 17877
rect 1829 17811 1863 17827
rect 94187 17861 94221 17877
rect 94187 17811 94221 17827
rect 1829 17525 1863 17541
rect 1829 17475 1863 17491
rect 94187 17525 94221 17541
rect 94187 17475 94221 17491
rect 1829 17189 1863 17205
rect 1829 17139 1863 17155
rect 94187 17189 94221 17205
rect 94187 17139 94221 17155
rect 1829 16853 1863 16869
rect 1829 16803 1863 16819
rect 94187 16853 94221 16869
rect 94187 16803 94221 16819
rect 1829 16517 1863 16533
rect 1829 16467 1863 16483
rect 94187 16517 94221 16533
rect 94187 16467 94221 16483
rect 1829 16181 1863 16197
rect 1829 16131 1863 16147
rect 94187 16181 94221 16197
rect 94187 16131 94221 16147
rect 1829 15845 1863 15861
rect 1829 15795 1863 15811
rect 94187 15845 94221 15861
rect 94187 15795 94221 15811
rect 1829 15509 1863 15525
rect 1829 15459 1863 15475
rect 94187 15509 94221 15525
rect 94187 15459 94221 15475
rect 1829 15173 1863 15189
rect 1829 15123 1863 15139
rect 94187 15173 94221 15189
rect 94187 15123 94221 15139
rect 1829 14837 1863 14853
rect 1829 14787 1863 14803
rect 94187 14837 94221 14853
rect 94187 14787 94221 14803
rect 1829 14501 1863 14517
rect 1829 14451 1863 14467
rect 94187 14501 94221 14517
rect 94187 14451 94221 14467
rect 1829 14165 1863 14181
rect 1829 14115 1863 14131
rect 94187 14165 94221 14181
rect 94187 14115 94221 14131
rect 1829 13829 1863 13845
rect 1829 13779 1863 13795
rect 94187 13829 94221 13845
rect 94187 13779 94221 13795
rect 1829 13493 1863 13509
rect 1829 13443 1863 13459
rect 94187 13493 94221 13509
rect 94187 13443 94221 13459
rect 1829 13157 1863 13173
rect 1829 13107 1863 13123
rect 94187 13157 94221 13173
rect 94187 13107 94221 13123
rect 1829 12821 1863 12837
rect 1829 12771 1863 12787
rect 94187 12821 94221 12837
rect 94187 12771 94221 12787
rect 1829 12485 1863 12501
rect 1829 12435 1863 12451
rect 94187 12485 94221 12501
rect 94187 12435 94221 12451
rect 1829 12149 1863 12165
rect 1829 12099 1863 12115
rect 94187 12149 94221 12165
rect 94187 12099 94221 12115
rect 1829 11813 1863 11829
rect 1829 11763 1863 11779
rect 94187 11813 94221 11829
rect 94187 11763 94221 11779
rect 1829 11477 1863 11493
rect 1829 11427 1863 11443
rect 94187 11477 94221 11493
rect 94187 11427 94221 11443
rect 1829 11141 1863 11157
rect 1829 11091 1863 11107
rect 94187 11141 94221 11157
rect 94187 11091 94221 11107
rect 1829 10805 1863 10821
rect 1829 10755 1863 10771
rect 94187 10805 94221 10821
rect 94187 10755 94221 10771
rect 1829 10469 1863 10485
rect 1829 10419 1863 10435
rect 94187 10469 94221 10485
rect 94187 10419 94221 10435
rect 1829 10133 1863 10149
rect 1829 10083 1863 10099
rect 94187 10133 94221 10149
rect 94187 10083 94221 10099
rect 1829 9797 1863 9813
rect 1829 9747 1863 9763
rect 94187 9797 94221 9813
rect 94187 9747 94221 9763
rect 1829 9461 1863 9477
rect 1829 9411 1863 9427
rect 94187 9461 94221 9477
rect 94187 9411 94221 9427
rect 1829 9125 1863 9141
rect 1829 9075 1863 9091
rect 94187 9125 94221 9141
rect 94187 9075 94221 9091
rect 1829 8789 1863 8805
rect 1829 8739 1863 8755
rect 94187 8789 94221 8805
rect 94187 8739 94221 8755
rect 1829 8453 1863 8469
rect 1829 8403 1863 8419
rect 94187 8453 94221 8469
rect 94187 8403 94221 8419
rect 1829 8117 1863 8133
rect 1829 8067 1863 8083
rect 94187 8117 94221 8133
rect 94187 8067 94221 8083
rect 1829 7781 1863 7797
rect 1829 7731 1863 7747
rect 94187 7781 94221 7797
rect 94187 7731 94221 7747
rect 1829 7445 1863 7461
rect 1829 7395 1863 7411
rect 94187 7445 94221 7461
rect 94187 7395 94221 7411
rect 1829 7109 1863 7125
rect 1829 7059 1863 7075
rect 94187 7109 94221 7125
rect 94187 7059 94221 7075
rect 1829 6773 1863 6789
rect 1829 6723 1863 6739
rect 94187 6773 94221 6789
rect 94187 6723 94221 6739
rect 1829 6437 1863 6453
rect 1829 6387 1863 6403
rect 94187 6437 94221 6453
rect 94187 6387 94221 6403
rect 1829 6101 1863 6117
rect 1829 6051 1863 6067
rect 94187 6101 94221 6117
rect 94187 6051 94221 6067
rect 1829 5765 1863 5781
rect 1829 5715 1863 5731
rect 94187 5765 94221 5781
rect 94187 5715 94221 5731
rect 1829 5429 1863 5445
rect 1829 5379 1863 5395
rect 94187 5429 94221 5445
rect 94187 5379 94221 5395
rect 1829 5093 1863 5109
rect 1829 5043 1863 5059
rect 94187 5093 94221 5109
rect 94187 5043 94221 5059
rect 1829 4757 1863 4773
rect 1829 4707 1863 4723
rect 94187 4757 94221 4773
rect 94187 4707 94221 4723
rect 1829 4421 1863 4437
rect 1829 4371 1863 4387
rect 94187 4421 94221 4437
rect 94187 4371 94221 4387
rect 1829 4085 1863 4101
rect 1829 4035 1863 4051
rect 94187 4085 94221 4101
rect 94187 4035 94221 4051
rect 1829 3749 1863 3765
rect 1829 3699 1863 3715
rect 94187 3749 94221 3765
rect 94187 3699 94221 3715
rect 1829 3413 1863 3429
rect 1829 3363 1863 3379
rect 94187 3413 94221 3429
rect 94187 3363 94221 3379
rect 1829 3077 1863 3093
rect 1829 3027 1863 3043
rect 94187 3077 94221 3093
rect 94187 3027 94221 3043
rect 1829 2741 1863 2757
rect 1829 2691 1863 2707
rect 94187 2741 94221 2757
rect 94187 2691 94221 2707
rect 1829 2405 1863 2421
rect 1829 2355 1863 2371
rect 94187 2405 94221 2421
rect 94187 2355 94221 2371
rect 1829 2069 1863 2085
rect 1829 2019 1863 2035
rect 94187 2069 94221 2085
rect 94187 2019 94221 2035
rect 2165 1733 2199 1749
rect 2165 1683 2199 1699
rect 2501 1733 2535 1749
rect 2501 1683 2535 1699
rect 2837 1733 2871 1749
rect 2837 1683 2871 1699
rect 3173 1733 3207 1749
rect 3173 1683 3207 1699
rect 3509 1733 3543 1749
rect 3509 1683 3543 1699
rect 3845 1733 3879 1749
rect 3845 1683 3879 1699
rect 4181 1733 4215 1749
rect 4181 1683 4215 1699
rect 4517 1733 4551 1749
rect 4517 1683 4551 1699
rect 4853 1733 4887 1749
rect 4853 1683 4887 1699
rect 5189 1733 5223 1749
rect 5189 1683 5223 1699
rect 5525 1733 5559 1749
rect 5525 1683 5559 1699
rect 5861 1733 5895 1749
rect 5861 1683 5895 1699
rect 6197 1733 6231 1749
rect 6197 1683 6231 1699
rect 6533 1733 6567 1749
rect 6533 1683 6567 1699
rect 6869 1733 6903 1749
rect 6869 1683 6903 1699
rect 7205 1733 7239 1749
rect 7205 1683 7239 1699
rect 7541 1733 7575 1749
rect 7541 1683 7575 1699
rect 7877 1733 7911 1749
rect 7877 1683 7911 1699
rect 8213 1733 8247 1749
rect 8213 1683 8247 1699
rect 8549 1733 8583 1749
rect 8549 1683 8583 1699
rect 8885 1733 8919 1749
rect 8885 1683 8919 1699
rect 9221 1733 9255 1749
rect 9221 1683 9255 1699
rect 9557 1733 9591 1749
rect 9557 1683 9591 1699
rect 9893 1733 9927 1749
rect 9893 1683 9927 1699
rect 10229 1733 10263 1749
rect 10229 1683 10263 1699
rect 10565 1733 10599 1749
rect 10565 1683 10599 1699
rect 10901 1733 10935 1749
rect 10901 1683 10935 1699
rect 11237 1733 11271 1749
rect 11237 1683 11271 1699
rect 11573 1733 11607 1749
rect 11573 1683 11607 1699
rect 11909 1733 11943 1749
rect 11909 1683 11943 1699
rect 12245 1733 12279 1749
rect 12245 1683 12279 1699
rect 12581 1733 12615 1749
rect 12581 1683 12615 1699
rect 12917 1733 12951 1749
rect 12917 1683 12951 1699
rect 13253 1733 13287 1749
rect 13253 1683 13287 1699
rect 13589 1733 13623 1749
rect 13589 1683 13623 1699
rect 13925 1733 13959 1749
rect 13925 1683 13959 1699
rect 14261 1733 14295 1749
rect 14261 1683 14295 1699
rect 14597 1733 14631 1749
rect 14597 1683 14631 1699
rect 14933 1733 14967 1749
rect 14933 1683 14967 1699
rect 15269 1733 15303 1749
rect 15269 1683 15303 1699
rect 15605 1733 15639 1749
rect 15605 1683 15639 1699
rect 15941 1733 15975 1749
rect 15941 1683 15975 1699
rect 16277 1733 16311 1749
rect 16277 1683 16311 1699
rect 16613 1733 16647 1749
rect 16613 1683 16647 1699
rect 16949 1733 16983 1749
rect 16949 1683 16983 1699
rect 17285 1733 17319 1749
rect 17285 1683 17319 1699
rect 17621 1733 17655 1749
rect 17621 1683 17655 1699
rect 17957 1733 17991 1749
rect 17957 1683 17991 1699
rect 18293 1733 18327 1749
rect 18293 1683 18327 1699
rect 18629 1733 18663 1749
rect 18629 1683 18663 1699
rect 18965 1733 18999 1749
rect 18965 1683 18999 1699
rect 19301 1733 19335 1749
rect 19301 1683 19335 1699
rect 19637 1733 19671 1749
rect 19637 1683 19671 1699
rect 19973 1733 20007 1749
rect 19973 1683 20007 1699
rect 20309 1733 20343 1749
rect 20309 1683 20343 1699
rect 20645 1733 20679 1749
rect 20645 1683 20679 1699
rect 20981 1733 21015 1749
rect 20981 1683 21015 1699
rect 21317 1733 21351 1749
rect 21317 1683 21351 1699
rect 21653 1733 21687 1749
rect 21653 1683 21687 1699
rect 21989 1733 22023 1749
rect 21989 1683 22023 1699
rect 22325 1733 22359 1749
rect 22325 1683 22359 1699
rect 22661 1733 22695 1749
rect 22661 1683 22695 1699
rect 22997 1733 23031 1749
rect 22997 1683 23031 1699
rect 23333 1733 23367 1749
rect 23333 1683 23367 1699
rect 23669 1733 23703 1749
rect 23669 1683 23703 1699
rect 24005 1733 24039 1749
rect 24005 1683 24039 1699
rect 24341 1733 24375 1749
rect 24341 1683 24375 1699
rect 24677 1733 24711 1749
rect 24677 1683 24711 1699
rect 25013 1733 25047 1749
rect 25013 1683 25047 1699
rect 25349 1733 25383 1749
rect 25349 1683 25383 1699
rect 25685 1733 25719 1749
rect 25685 1683 25719 1699
rect 26021 1733 26055 1749
rect 26021 1683 26055 1699
rect 26357 1733 26391 1749
rect 26357 1683 26391 1699
rect 26693 1733 26727 1749
rect 26693 1683 26727 1699
rect 27029 1733 27063 1749
rect 27029 1683 27063 1699
rect 27365 1733 27399 1749
rect 27365 1683 27399 1699
rect 27701 1733 27735 1749
rect 27701 1683 27735 1699
rect 28037 1733 28071 1749
rect 28037 1683 28071 1699
rect 28373 1733 28407 1749
rect 28373 1683 28407 1699
rect 28709 1733 28743 1749
rect 28709 1683 28743 1699
rect 29045 1733 29079 1749
rect 29045 1683 29079 1699
rect 29381 1733 29415 1749
rect 29381 1683 29415 1699
rect 29717 1733 29751 1749
rect 29717 1683 29751 1699
rect 30053 1733 30087 1749
rect 30053 1683 30087 1699
rect 30389 1733 30423 1749
rect 30389 1683 30423 1699
rect 30725 1733 30759 1749
rect 30725 1683 30759 1699
rect 31061 1733 31095 1749
rect 31061 1683 31095 1699
rect 31397 1733 31431 1749
rect 31397 1683 31431 1699
rect 31733 1733 31767 1749
rect 31733 1683 31767 1699
rect 32069 1733 32103 1749
rect 32069 1683 32103 1699
rect 32405 1733 32439 1749
rect 32405 1683 32439 1699
rect 32741 1733 32775 1749
rect 32741 1683 32775 1699
rect 33077 1733 33111 1749
rect 33077 1683 33111 1699
rect 33413 1733 33447 1749
rect 33413 1683 33447 1699
rect 33749 1733 33783 1749
rect 33749 1683 33783 1699
rect 34085 1733 34119 1749
rect 34085 1683 34119 1699
rect 34421 1733 34455 1749
rect 34421 1683 34455 1699
rect 34757 1733 34791 1749
rect 34757 1683 34791 1699
rect 35093 1733 35127 1749
rect 35093 1683 35127 1699
rect 35429 1733 35463 1749
rect 35429 1683 35463 1699
rect 35765 1733 35799 1749
rect 35765 1683 35799 1699
rect 36101 1733 36135 1749
rect 36101 1683 36135 1699
rect 36437 1733 36471 1749
rect 36437 1683 36471 1699
rect 36773 1733 36807 1749
rect 36773 1683 36807 1699
rect 37109 1733 37143 1749
rect 37109 1683 37143 1699
rect 37445 1733 37479 1749
rect 37445 1683 37479 1699
rect 37781 1733 37815 1749
rect 37781 1683 37815 1699
rect 38117 1733 38151 1749
rect 38117 1683 38151 1699
rect 38453 1733 38487 1749
rect 38453 1683 38487 1699
rect 38789 1733 38823 1749
rect 38789 1683 38823 1699
rect 39125 1733 39159 1749
rect 39125 1683 39159 1699
rect 39461 1733 39495 1749
rect 39461 1683 39495 1699
rect 39797 1733 39831 1749
rect 39797 1683 39831 1699
rect 40133 1733 40167 1749
rect 40133 1683 40167 1699
rect 40469 1733 40503 1749
rect 40469 1683 40503 1699
rect 40805 1733 40839 1749
rect 40805 1683 40839 1699
rect 41141 1733 41175 1749
rect 41141 1683 41175 1699
rect 41477 1733 41511 1749
rect 41477 1683 41511 1699
rect 41813 1733 41847 1749
rect 41813 1683 41847 1699
rect 42149 1733 42183 1749
rect 42149 1683 42183 1699
rect 42485 1733 42519 1749
rect 42485 1683 42519 1699
rect 42821 1733 42855 1749
rect 42821 1683 42855 1699
rect 43157 1733 43191 1749
rect 43157 1683 43191 1699
rect 43493 1733 43527 1749
rect 43493 1683 43527 1699
rect 43829 1733 43863 1749
rect 43829 1683 43863 1699
rect 44165 1733 44199 1749
rect 44165 1683 44199 1699
rect 44501 1733 44535 1749
rect 44501 1683 44535 1699
rect 44837 1733 44871 1749
rect 44837 1683 44871 1699
rect 45173 1733 45207 1749
rect 45173 1683 45207 1699
rect 45509 1733 45543 1749
rect 45509 1683 45543 1699
rect 45845 1733 45879 1749
rect 45845 1683 45879 1699
rect 46181 1733 46215 1749
rect 46181 1683 46215 1699
rect 46517 1733 46551 1749
rect 46517 1683 46551 1699
rect 46853 1733 46887 1749
rect 46853 1683 46887 1699
rect 47189 1733 47223 1749
rect 47189 1683 47223 1699
rect 47525 1733 47559 1749
rect 47525 1683 47559 1699
rect 47861 1733 47895 1749
rect 47861 1683 47895 1699
rect 48197 1733 48231 1749
rect 48197 1683 48231 1699
rect 48533 1733 48567 1749
rect 48533 1683 48567 1699
rect 48869 1733 48903 1749
rect 48869 1683 48903 1699
rect 49205 1733 49239 1749
rect 49205 1683 49239 1699
rect 49541 1733 49575 1749
rect 49541 1683 49575 1699
rect 49877 1733 49911 1749
rect 49877 1683 49911 1699
rect 50213 1733 50247 1749
rect 50213 1683 50247 1699
rect 50549 1733 50583 1749
rect 50549 1683 50583 1699
rect 50885 1733 50919 1749
rect 50885 1683 50919 1699
rect 51221 1733 51255 1749
rect 51221 1683 51255 1699
rect 51557 1733 51591 1749
rect 51557 1683 51591 1699
rect 51893 1733 51927 1749
rect 51893 1683 51927 1699
rect 52229 1733 52263 1749
rect 52229 1683 52263 1699
rect 52565 1733 52599 1749
rect 52565 1683 52599 1699
rect 52901 1733 52935 1749
rect 52901 1683 52935 1699
rect 53237 1733 53271 1749
rect 53237 1683 53271 1699
rect 53573 1733 53607 1749
rect 53573 1683 53607 1699
rect 53909 1733 53943 1749
rect 53909 1683 53943 1699
rect 54245 1733 54279 1749
rect 54245 1683 54279 1699
rect 54581 1733 54615 1749
rect 54581 1683 54615 1699
rect 54917 1733 54951 1749
rect 54917 1683 54951 1699
rect 55253 1733 55287 1749
rect 55253 1683 55287 1699
rect 55589 1733 55623 1749
rect 55589 1683 55623 1699
rect 55925 1733 55959 1749
rect 55925 1683 55959 1699
rect 56261 1733 56295 1749
rect 56261 1683 56295 1699
rect 56597 1733 56631 1749
rect 56597 1683 56631 1699
rect 56933 1733 56967 1749
rect 56933 1683 56967 1699
rect 57269 1733 57303 1749
rect 57269 1683 57303 1699
rect 57605 1733 57639 1749
rect 57605 1683 57639 1699
rect 57941 1733 57975 1749
rect 57941 1683 57975 1699
rect 58277 1733 58311 1749
rect 58277 1683 58311 1699
rect 58613 1733 58647 1749
rect 58613 1683 58647 1699
rect 58949 1733 58983 1749
rect 58949 1683 58983 1699
rect 59285 1733 59319 1749
rect 59285 1683 59319 1699
rect 59621 1733 59655 1749
rect 59621 1683 59655 1699
rect 59957 1733 59991 1749
rect 59957 1683 59991 1699
rect 60293 1733 60327 1749
rect 60293 1683 60327 1699
rect 60629 1733 60663 1749
rect 60629 1683 60663 1699
rect 60965 1733 60999 1749
rect 60965 1683 60999 1699
rect 61301 1733 61335 1749
rect 61301 1683 61335 1699
rect 61637 1733 61671 1749
rect 61637 1683 61671 1699
rect 61973 1733 62007 1749
rect 61973 1683 62007 1699
rect 62309 1733 62343 1749
rect 62309 1683 62343 1699
rect 62645 1733 62679 1749
rect 62645 1683 62679 1699
rect 62981 1733 63015 1749
rect 62981 1683 63015 1699
rect 63317 1733 63351 1749
rect 63317 1683 63351 1699
rect 63653 1733 63687 1749
rect 63653 1683 63687 1699
rect 63989 1733 64023 1749
rect 63989 1683 64023 1699
rect 64325 1733 64359 1749
rect 64325 1683 64359 1699
rect 64661 1733 64695 1749
rect 64661 1683 64695 1699
rect 64997 1733 65031 1749
rect 64997 1683 65031 1699
rect 65333 1733 65367 1749
rect 65333 1683 65367 1699
rect 65669 1733 65703 1749
rect 65669 1683 65703 1699
rect 66005 1733 66039 1749
rect 66005 1683 66039 1699
rect 66341 1733 66375 1749
rect 66341 1683 66375 1699
rect 66677 1733 66711 1749
rect 66677 1683 66711 1699
rect 67013 1733 67047 1749
rect 67013 1683 67047 1699
rect 67349 1733 67383 1749
rect 67349 1683 67383 1699
rect 67685 1733 67719 1749
rect 67685 1683 67719 1699
rect 68021 1733 68055 1749
rect 68021 1683 68055 1699
rect 68357 1733 68391 1749
rect 68357 1683 68391 1699
rect 68693 1733 68727 1749
rect 68693 1683 68727 1699
rect 69029 1733 69063 1749
rect 69029 1683 69063 1699
rect 69365 1733 69399 1749
rect 69365 1683 69399 1699
rect 69701 1733 69735 1749
rect 69701 1683 69735 1699
rect 70037 1733 70071 1749
rect 70037 1683 70071 1699
rect 70373 1733 70407 1749
rect 70373 1683 70407 1699
rect 70709 1733 70743 1749
rect 70709 1683 70743 1699
rect 71045 1733 71079 1749
rect 71045 1683 71079 1699
rect 71381 1733 71415 1749
rect 71381 1683 71415 1699
rect 71717 1733 71751 1749
rect 71717 1683 71751 1699
rect 72053 1733 72087 1749
rect 72053 1683 72087 1699
rect 72389 1733 72423 1749
rect 72389 1683 72423 1699
rect 72725 1733 72759 1749
rect 72725 1683 72759 1699
rect 73061 1733 73095 1749
rect 73061 1683 73095 1699
rect 73397 1733 73431 1749
rect 73397 1683 73431 1699
rect 73733 1733 73767 1749
rect 73733 1683 73767 1699
rect 74069 1733 74103 1749
rect 74069 1683 74103 1699
rect 74405 1733 74439 1749
rect 74405 1683 74439 1699
rect 74741 1733 74775 1749
rect 74741 1683 74775 1699
rect 75077 1733 75111 1749
rect 75077 1683 75111 1699
rect 75413 1733 75447 1749
rect 75413 1683 75447 1699
rect 75749 1733 75783 1749
rect 75749 1683 75783 1699
rect 76085 1733 76119 1749
rect 76085 1683 76119 1699
rect 76421 1733 76455 1749
rect 76421 1683 76455 1699
rect 76757 1733 76791 1749
rect 76757 1683 76791 1699
rect 77093 1733 77127 1749
rect 77093 1683 77127 1699
rect 77429 1733 77463 1749
rect 77429 1683 77463 1699
rect 77765 1733 77799 1749
rect 77765 1683 77799 1699
rect 78101 1733 78135 1749
rect 78101 1683 78135 1699
rect 78437 1733 78471 1749
rect 78437 1683 78471 1699
rect 78773 1733 78807 1749
rect 78773 1683 78807 1699
rect 79109 1733 79143 1749
rect 79109 1683 79143 1699
rect 79445 1733 79479 1749
rect 79445 1683 79479 1699
rect 79781 1733 79815 1749
rect 79781 1683 79815 1699
rect 80117 1733 80151 1749
rect 80117 1683 80151 1699
rect 80453 1733 80487 1749
rect 80453 1683 80487 1699
rect 80789 1733 80823 1749
rect 80789 1683 80823 1699
rect 81125 1733 81159 1749
rect 81125 1683 81159 1699
rect 81461 1733 81495 1749
rect 81461 1683 81495 1699
rect 81797 1733 81831 1749
rect 81797 1683 81831 1699
rect 82133 1733 82167 1749
rect 82133 1683 82167 1699
rect 82469 1733 82503 1749
rect 82469 1683 82503 1699
rect 82805 1733 82839 1749
rect 82805 1683 82839 1699
rect 83141 1733 83175 1749
rect 83141 1683 83175 1699
rect 83477 1733 83511 1749
rect 83477 1683 83511 1699
rect 83813 1733 83847 1749
rect 83813 1683 83847 1699
rect 84149 1733 84183 1749
rect 84149 1683 84183 1699
rect 84485 1733 84519 1749
rect 84485 1683 84519 1699
rect 84821 1733 84855 1749
rect 84821 1683 84855 1699
rect 85157 1733 85191 1749
rect 85157 1683 85191 1699
rect 85493 1733 85527 1749
rect 85493 1683 85527 1699
rect 85829 1733 85863 1749
rect 85829 1683 85863 1699
rect 86165 1733 86199 1749
rect 86165 1683 86199 1699
rect 86501 1733 86535 1749
rect 86501 1683 86535 1699
rect 86837 1733 86871 1749
rect 86837 1683 86871 1699
rect 87173 1733 87207 1749
rect 87173 1683 87207 1699
rect 87509 1733 87543 1749
rect 87509 1683 87543 1699
rect 87845 1733 87879 1749
rect 87845 1683 87879 1699
rect 88181 1733 88215 1749
rect 88181 1683 88215 1699
rect 88517 1733 88551 1749
rect 88517 1683 88551 1699
rect 88853 1733 88887 1749
rect 88853 1683 88887 1699
rect 89189 1733 89223 1749
rect 89189 1683 89223 1699
rect 89525 1733 89559 1749
rect 89525 1683 89559 1699
rect 89861 1733 89895 1749
rect 89861 1683 89895 1699
rect 90197 1733 90231 1749
rect 90197 1683 90231 1699
rect 90533 1733 90567 1749
rect 90533 1683 90567 1699
rect 90869 1733 90903 1749
rect 90869 1683 90903 1699
rect 91205 1733 91239 1749
rect 91205 1683 91239 1699
rect 91541 1733 91575 1749
rect 91541 1683 91575 1699
rect 91877 1733 91911 1749
rect 91877 1683 91911 1699
rect 92213 1733 92247 1749
rect 92213 1683 92247 1699
rect 92549 1733 92583 1749
rect 92549 1683 92583 1699
rect 92885 1733 92919 1749
rect 92885 1683 92919 1699
rect 93221 1733 93255 1749
rect 93221 1683 93255 1699
rect 93557 1733 93591 1749
rect 93557 1683 93591 1699
<< viali >>
rect 2165 77763 2199 77797
rect 2501 77763 2535 77797
rect 2837 77763 2871 77797
rect 3173 77763 3207 77797
rect 3509 77763 3543 77797
rect 3845 77763 3879 77797
rect 4181 77763 4215 77797
rect 4517 77763 4551 77797
rect 4853 77763 4887 77797
rect 5189 77763 5223 77797
rect 5525 77763 5559 77797
rect 5861 77763 5895 77797
rect 6197 77763 6231 77797
rect 6533 77763 6567 77797
rect 6869 77763 6903 77797
rect 7205 77763 7239 77797
rect 7541 77763 7575 77797
rect 7877 77763 7911 77797
rect 8213 77763 8247 77797
rect 8549 77763 8583 77797
rect 8885 77763 8919 77797
rect 9221 77763 9255 77797
rect 9557 77763 9591 77797
rect 9893 77763 9927 77797
rect 10229 77763 10263 77797
rect 10565 77763 10599 77797
rect 10901 77763 10935 77797
rect 11237 77763 11271 77797
rect 11573 77763 11607 77797
rect 11909 77763 11943 77797
rect 12245 77763 12279 77797
rect 12581 77763 12615 77797
rect 12917 77763 12951 77797
rect 13253 77763 13287 77797
rect 13589 77763 13623 77797
rect 13925 77763 13959 77797
rect 14261 77763 14295 77797
rect 14597 77763 14631 77797
rect 14933 77763 14967 77797
rect 15269 77763 15303 77797
rect 15605 77763 15639 77797
rect 15941 77763 15975 77797
rect 16277 77763 16311 77797
rect 16613 77763 16647 77797
rect 16949 77763 16983 77797
rect 17285 77763 17319 77797
rect 17621 77763 17655 77797
rect 17957 77763 17991 77797
rect 18293 77763 18327 77797
rect 18629 77763 18663 77797
rect 18965 77763 18999 77797
rect 19301 77763 19335 77797
rect 19637 77763 19671 77797
rect 19973 77763 20007 77797
rect 20309 77763 20343 77797
rect 20645 77763 20679 77797
rect 20981 77763 21015 77797
rect 21317 77763 21351 77797
rect 21653 77763 21687 77797
rect 21989 77763 22023 77797
rect 22325 77763 22359 77797
rect 22661 77763 22695 77797
rect 22997 77763 23031 77797
rect 23333 77763 23367 77797
rect 23669 77763 23703 77797
rect 24005 77763 24039 77797
rect 24341 77763 24375 77797
rect 24677 77763 24711 77797
rect 25013 77763 25047 77797
rect 25349 77763 25383 77797
rect 25685 77763 25719 77797
rect 26021 77763 26055 77797
rect 26357 77763 26391 77797
rect 26693 77763 26727 77797
rect 27029 77763 27063 77797
rect 27365 77763 27399 77797
rect 27701 77763 27735 77797
rect 28037 77763 28071 77797
rect 28373 77763 28407 77797
rect 28709 77763 28743 77797
rect 29045 77763 29079 77797
rect 29381 77763 29415 77797
rect 29717 77763 29751 77797
rect 30053 77763 30087 77797
rect 30389 77763 30423 77797
rect 30725 77763 30759 77797
rect 31061 77763 31095 77797
rect 31397 77763 31431 77797
rect 31733 77763 31767 77797
rect 32069 77763 32103 77797
rect 32405 77763 32439 77797
rect 32741 77763 32775 77797
rect 33077 77763 33111 77797
rect 33413 77763 33447 77797
rect 33749 77763 33783 77797
rect 34085 77763 34119 77797
rect 34421 77763 34455 77797
rect 34757 77763 34791 77797
rect 35093 77763 35127 77797
rect 35429 77763 35463 77797
rect 35765 77763 35799 77797
rect 36101 77763 36135 77797
rect 36437 77763 36471 77797
rect 36773 77763 36807 77797
rect 37109 77763 37143 77797
rect 37445 77763 37479 77797
rect 37781 77763 37815 77797
rect 38117 77763 38151 77797
rect 38453 77763 38487 77797
rect 38789 77763 38823 77797
rect 39125 77763 39159 77797
rect 39461 77763 39495 77797
rect 39797 77763 39831 77797
rect 40133 77763 40167 77797
rect 40469 77763 40503 77797
rect 40805 77763 40839 77797
rect 41141 77763 41175 77797
rect 41477 77763 41511 77797
rect 41813 77763 41847 77797
rect 42149 77763 42183 77797
rect 42485 77763 42519 77797
rect 42821 77763 42855 77797
rect 43157 77763 43191 77797
rect 43493 77763 43527 77797
rect 43829 77763 43863 77797
rect 44165 77763 44199 77797
rect 44501 77763 44535 77797
rect 44837 77763 44871 77797
rect 45173 77763 45207 77797
rect 45509 77763 45543 77797
rect 45845 77763 45879 77797
rect 46181 77763 46215 77797
rect 46517 77763 46551 77797
rect 46853 77763 46887 77797
rect 47189 77763 47223 77797
rect 47525 77763 47559 77797
rect 47861 77763 47895 77797
rect 48197 77763 48231 77797
rect 48533 77763 48567 77797
rect 48869 77763 48903 77797
rect 49205 77763 49239 77797
rect 49541 77763 49575 77797
rect 49877 77763 49911 77797
rect 50213 77763 50247 77797
rect 50549 77763 50583 77797
rect 50885 77763 50919 77797
rect 51221 77763 51255 77797
rect 51557 77763 51591 77797
rect 51893 77763 51927 77797
rect 52229 77763 52263 77797
rect 52565 77763 52599 77797
rect 52901 77763 52935 77797
rect 53237 77763 53271 77797
rect 53573 77763 53607 77797
rect 53909 77763 53943 77797
rect 54245 77763 54279 77797
rect 54581 77763 54615 77797
rect 54917 77763 54951 77797
rect 55253 77763 55287 77797
rect 55589 77763 55623 77797
rect 55925 77763 55959 77797
rect 56261 77763 56295 77797
rect 56597 77763 56631 77797
rect 56933 77763 56967 77797
rect 57269 77763 57303 77797
rect 57605 77763 57639 77797
rect 57941 77763 57975 77797
rect 58277 77763 58311 77797
rect 58613 77763 58647 77797
rect 58949 77763 58983 77797
rect 59285 77763 59319 77797
rect 59621 77763 59655 77797
rect 59957 77763 59991 77797
rect 60293 77763 60327 77797
rect 60629 77763 60663 77797
rect 60965 77763 60999 77797
rect 61301 77763 61335 77797
rect 61637 77763 61671 77797
rect 61973 77763 62007 77797
rect 62309 77763 62343 77797
rect 62645 77763 62679 77797
rect 62981 77763 63015 77797
rect 63317 77763 63351 77797
rect 63653 77763 63687 77797
rect 63989 77763 64023 77797
rect 64325 77763 64359 77797
rect 64661 77763 64695 77797
rect 64997 77763 65031 77797
rect 65333 77763 65367 77797
rect 65669 77763 65703 77797
rect 66005 77763 66039 77797
rect 66341 77763 66375 77797
rect 66677 77763 66711 77797
rect 67013 77763 67047 77797
rect 67349 77763 67383 77797
rect 67685 77763 67719 77797
rect 68021 77763 68055 77797
rect 68357 77763 68391 77797
rect 68693 77763 68727 77797
rect 69029 77763 69063 77797
rect 69365 77763 69399 77797
rect 69701 77763 69735 77797
rect 70037 77763 70071 77797
rect 70373 77763 70407 77797
rect 70709 77763 70743 77797
rect 71045 77763 71079 77797
rect 71381 77763 71415 77797
rect 71717 77763 71751 77797
rect 72053 77763 72087 77797
rect 72389 77763 72423 77797
rect 72725 77763 72759 77797
rect 73061 77763 73095 77797
rect 73397 77763 73431 77797
rect 73733 77763 73767 77797
rect 74069 77763 74103 77797
rect 74405 77763 74439 77797
rect 74741 77763 74775 77797
rect 75077 77763 75111 77797
rect 75413 77763 75447 77797
rect 75749 77763 75783 77797
rect 76085 77763 76119 77797
rect 76421 77763 76455 77797
rect 76757 77763 76791 77797
rect 77093 77763 77127 77797
rect 77429 77763 77463 77797
rect 77765 77763 77799 77797
rect 78101 77763 78135 77797
rect 78437 77763 78471 77797
rect 78773 77763 78807 77797
rect 79109 77763 79143 77797
rect 79445 77763 79479 77797
rect 79781 77763 79815 77797
rect 80117 77763 80151 77797
rect 80453 77763 80487 77797
rect 80789 77763 80823 77797
rect 81125 77763 81159 77797
rect 81461 77763 81495 77797
rect 81797 77763 81831 77797
rect 82133 77763 82167 77797
rect 82469 77763 82503 77797
rect 82805 77763 82839 77797
rect 83141 77763 83175 77797
rect 83477 77763 83511 77797
rect 83813 77763 83847 77797
rect 84149 77763 84183 77797
rect 84485 77763 84519 77797
rect 84821 77763 84855 77797
rect 85157 77763 85191 77797
rect 85493 77763 85527 77797
rect 85829 77763 85863 77797
rect 86165 77763 86199 77797
rect 86501 77763 86535 77797
rect 86837 77763 86871 77797
rect 87173 77763 87207 77797
rect 87509 77763 87543 77797
rect 87845 77763 87879 77797
rect 88181 77763 88215 77797
rect 88517 77763 88551 77797
rect 88853 77763 88887 77797
rect 89189 77763 89223 77797
rect 89525 77763 89559 77797
rect 89861 77763 89895 77797
rect 90197 77763 90231 77797
rect 90533 77763 90567 77797
rect 90869 77763 90903 77797
rect 91205 77763 91239 77797
rect 91541 77763 91575 77797
rect 91877 77763 91911 77797
rect 92213 77763 92247 77797
rect 92549 77763 92583 77797
rect 92885 77763 92919 77797
rect 93221 77763 93255 77797
rect 93557 77763 93591 77797
rect 1829 77299 1863 77333
rect 94187 77299 94221 77333
rect 1829 76963 1863 76997
rect 94187 76963 94221 76997
rect 1829 76627 1863 76661
rect 94187 76627 94221 76661
rect 1829 76291 1863 76325
rect 94187 76291 94221 76325
rect 1829 75955 1863 75989
rect 94187 75955 94221 75989
rect 1829 75619 1863 75653
rect 94187 75619 94221 75653
rect 1829 75283 1863 75317
rect 94187 75283 94221 75317
rect 1829 74947 1863 74981
rect 94187 74947 94221 74981
rect 1829 74611 1863 74645
rect 94187 74611 94221 74645
rect 1829 74275 1863 74309
rect 94187 74275 94221 74309
rect 1829 73939 1863 73973
rect 94187 73939 94221 73973
rect 1829 73603 1863 73637
rect 94187 73603 94221 73637
rect 1829 73267 1863 73301
rect 94187 73267 94221 73301
rect 1829 72931 1863 72965
rect 94187 72931 94221 72965
rect 1829 72595 1863 72629
rect 94187 72595 94221 72629
rect 1829 72259 1863 72293
rect 94187 72259 94221 72293
rect 1829 71923 1863 71957
rect 94187 71923 94221 71957
rect 1829 71587 1863 71621
rect 94187 71587 94221 71621
rect 1829 71251 1863 71285
rect 94187 71251 94221 71285
rect 1829 70915 1863 70949
rect 94187 70915 94221 70949
rect 1829 70579 1863 70613
rect 94187 70579 94221 70613
rect 1829 70243 1863 70277
rect 94187 70243 94221 70277
rect 1829 69907 1863 69941
rect 94187 69907 94221 69941
rect 1829 69571 1863 69605
rect 94187 69571 94221 69605
rect 1829 69235 1863 69269
rect 94187 69235 94221 69269
rect 1829 68899 1863 68933
rect 94187 68899 94221 68933
rect 1829 68563 1863 68597
rect 94187 68563 94221 68597
rect 1829 68227 1863 68261
rect 94187 68227 94221 68261
rect 1829 67891 1863 67925
rect 94187 67891 94221 67925
rect 1829 67555 1863 67589
rect 94187 67555 94221 67589
rect 1829 67219 1863 67253
rect 94187 67219 94221 67253
rect 1829 66883 1863 66917
rect 94187 66883 94221 66917
rect 1829 66547 1863 66581
rect 94187 66547 94221 66581
rect 1829 66211 1863 66245
rect 94187 66211 94221 66245
rect 1829 65875 1863 65909
rect 94187 65875 94221 65909
rect 1829 65539 1863 65573
rect 94187 65539 94221 65573
rect 1829 65203 1863 65237
rect 94187 65203 94221 65237
rect 1829 64867 1863 64901
rect 94187 64867 94221 64901
rect 1829 64531 1863 64565
rect 94187 64531 94221 64565
rect 1829 64195 1863 64229
rect 94187 64195 94221 64229
rect 1829 63859 1863 63893
rect 94187 63859 94221 63893
rect 1829 63523 1863 63557
rect 94187 63523 94221 63557
rect 1829 63187 1863 63221
rect 94187 63187 94221 63221
rect 1829 62851 1863 62885
rect 94187 62851 94221 62885
rect 1829 62515 1863 62549
rect 94187 62515 94221 62549
rect 1829 62179 1863 62213
rect 94187 62179 94221 62213
rect 1829 61843 1863 61877
rect 94187 61843 94221 61877
rect 1829 61507 1863 61541
rect 94187 61507 94221 61541
rect 1829 61171 1863 61205
rect 94187 61171 94221 61205
rect 1829 60835 1863 60869
rect 94187 60835 94221 60869
rect 1829 60499 1863 60533
rect 94187 60499 94221 60533
rect 1829 60163 1863 60197
rect 94187 60163 94221 60197
rect 1829 59827 1863 59861
rect 94187 59827 94221 59861
rect 1829 59491 1863 59525
rect 94187 59491 94221 59525
rect 1829 59155 1863 59189
rect 94187 59155 94221 59189
rect 1829 58819 1863 58853
rect 94187 58819 94221 58853
rect 1829 58483 1863 58517
rect 94187 58483 94221 58517
rect 1829 58147 1863 58181
rect 94187 58147 94221 58181
rect 1829 57811 1863 57845
rect 94187 57811 94221 57845
rect 1829 57475 1863 57509
rect 94187 57475 94221 57509
rect 1829 57139 1863 57173
rect 94187 57139 94221 57173
rect 1829 56803 1863 56837
rect 94187 56803 94221 56837
rect 1829 56467 1863 56501
rect 94187 56467 94221 56501
rect 1829 56131 1863 56165
rect 94187 56131 94221 56165
rect 1829 55795 1863 55829
rect 94187 55795 94221 55829
rect 1829 55459 1863 55493
rect 94187 55459 94221 55493
rect 1829 55123 1863 55157
rect 94187 55123 94221 55157
rect 1829 54787 1863 54821
rect 94187 54787 94221 54821
rect 1829 54451 1863 54485
rect 94187 54451 94221 54485
rect 1829 54115 1863 54149
rect 94187 54115 94221 54149
rect 1829 53779 1863 53813
rect 94187 53779 94221 53813
rect 1829 53443 1863 53477
rect 94187 53443 94221 53477
rect 1829 53107 1863 53141
rect 94187 53107 94221 53141
rect 1829 52771 1863 52805
rect 94187 52771 94221 52805
rect 1829 52435 1863 52469
rect 94187 52435 94221 52469
rect 1829 52099 1863 52133
rect 94187 52099 94221 52133
rect 1829 51763 1863 51797
rect 94187 51763 94221 51797
rect 1829 51427 1863 51461
rect 94187 51427 94221 51461
rect 1829 51091 1863 51125
rect 94187 51091 94221 51125
rect 1829 50755 1863 50789
rect 94187 50755 94221 50789
rect 1829 50419 1863 50453
rect 94187 50419 94221 50453
rect 1829 50083 1863 50117
rect 94187 50083 94221 50117
rect 1829 49747 1863 49781
rect 94187 49747 94221 49781
rect 1829 49411 1863 49445
rect 94187 49411 94221 49445
rect 1829 49075 1863 49109
rect 94187 49075 94221 49109
rect 1829 48739 1863 48773
rect 94187 48739 94221 48773
rect 1829 48403 1863 48437
rect 94187 48403 94221 48437
rect 1829 48067 1863 48101
rect 94187 48067 94221 48101
rect 1829 47731 1863 47765
rect 94187 47731 94221 47765
rect 1829 47395 1863 47429
rect 94187 47395 94221 47429
rect 1829 47059 1863 47093
rect 94187 47059 94221 47093
rect 1829 46723 1863 46757
rect 94187 46723 94221 46757
rect 1829 46387 1863 46421
rect 94187 46387 94221 46421
rect 1829 46051 1863 46085
rect 94187 46051 94221 46085
rect 1829 45715 1863 45749
rect 94187 45715 94221 45749
rect 1829 45379 1863 45413
rect 94187 45379 94221 45413
rect 1829 45043 1863 45077
rect 94187 45043 94221 45077
rect 1829 44707 1863 44741
rect 94187 44707 94221 44741
rect 1829 44371 1863 44405
rect 94187 44371 94221 44405
rect 1829 44035 1863 44069
rect 94187 44035 94221 44069
rect 1829 43699 1863 43733
rect 94187 43699 94221 43733
rect 1829 43363 1863 43397
rect 94187 43363 94221 43397
rect 1829 43027 1863 43061
rect 94187 43027 94221 43061
rect 1829 42691 1863 42725
rect 94187 42691 94221 42725
rect 1829 42355 1863 42389
rect 94187 42355 94221 42389
rect 1829 42019 1863 42053
rect 94187 42019 94221 42053
rect 1829 41683 1863 41717
rect 94187 41683 94221 41717
rect 1829 41347 1863 41381
rect 94187 41347 94221 41381
rect 1829 41011 1863 41045
rect 94187 41011 94221 41045
rect 1829 40675 1863 40709
rect 94187 40675 94221 40709
rect 1829 40339 1863 40373
rect 94187 40339 94221 40373
rect 1829 40003 1863 40037
rect 94187 40003 94221 40037
rect 1829 39667 1863 39701
rect 94187 39667 94221 39701
rect 1829 39331 1863 39365
rect 94187 39331 94221 39365
rect 1829 38995 1863 39029
rect 94187 38995 94221 39029
rect 1829 38659 1863 38693
rect 94187 38659 94221 38693
rect 1829 38323 1863 38357
rect 94187 38323 94221 38357
rect 1829 37987 1863 38021
rect 94187 37987 94221 38021
rect 1829 37651 1863 37685
rect 94187 37651 94221 37685
rect 1829 37315 1863 37349
rect 94187 37315 94221 37349
rect 1829 36979 1863 37013
rect 94187 36979 94221 37013
rect 1829 36643 1863 36677
rect 94187 36643 94221 36677
rect 1829 36307 1863 36341
rect 94187 36307 94221 36341
rect 1829 35971 1863 36005
rect 94187 35971 94221 36005
rect 1829 35635 1863 35669
rect 94187 35635 94221 35669
rect 1829 35299 1863 35333
rect 94187 35299 94221 35333
rect 1829 34963 1863 34997
rect 94187 34963 94221 34997
rect 1829 34627 1863 34661
rect 94187 34627 94221 34661
rect 1829 34291 1863 34325
rect 94187 34291 94221 34325
rect 1829 33955 1863 33989
rect 94187 33955 94221 33989
rect 1829 33619 1863 33653
rect 94187 33619 94221 33653
rect 1829 33283 1863 33317
rect 94187 33283 94221 33317
rect 1829 32947 1863 32981
rect 94187 32947 94221 32981
rect 1829 32611 1863 32645
rect 94187 32611 94221 32645
rect 1829 32275 1863 32309
rect 94187 32275 94221 32309
rect 1829 31939 1863 31973
rect 94187 31939 94221 31973
rect 1829 31603 1863 31637
rect 94187 31603 94221 31637
rect 1829 31267 1863 31301
rect 94187 31267 94221 31301
rect 1829 30931 1863 30965
rect 94187 30931 94221 30965
rect 1829 30595 1863 30629
rect 94187 30595 94221 30629
rect 1829 30259 1863 30293
rect 94187 30259 94221 30293
rect 1829 29923 1863 29957
rect 94187 29923 94221 29957
rect 1829 29587 1863 29621
rect 94187 29587 94221 29621
rect 1829 29251 1863 29285
rect 94187 29251 94221 29285
rect 1829 28915 1863 28949
rect 94187 28915 94221 28949
rect 1829 28579 1863 28613
rect 94187 28579 94221 28613
rect 1829 28243 1863 28277
rect 94187 28243 94221 28277
rect 1829 27907 1863 27941
rect 94187 27907 94221 27941
rect 1829 27571 1863 27605
rect 94187 27571 94221 27605
rect 1829 27235 1863 27269
rect 94187 27235 94221 27269
rect 1829 26899 1863 26933
rect 94187 26899 94221 26933
rect 1829 26563 1863 26597
rect 94187 26563 94221 26597
rect 1829 26227 1863 26261
rect 94187 26227 94221 26261
rect 1829 25891 1863 25925
rect 94187 25891 94221 25925
rect 1829 25555 1863 25589
rect 94187 25555 94221 25589
rect 1829 25219 1863 25253
rect 94187 25219 94221 25253
rect 1829 24883 1863 24917
rect 94187 24883 94221 24917
rect 1829 24547 1863 24581
rect 94187 24547 94221 24581
rect 1829 24211 1863 24245
rect 94187 24211 94221 24245
rect 1829 23875 1863 23909
rect 94187 23875 94221 23909
rect 1829 23539 1863 23573
rect 94187 23539 94221 23573
rect 1829 23203 1863 23237
rect 94187 23203 94221 23237
rect 1829 22867 1863 22901
rect 94187 22867 94221 22901
rect 1829 22531 1863 22565
rect 94187 22531 94221 22565
rect 1829 22195 1863 22229
rect 94187 22195 94221 22229
rect 1829 21859 1863 21893
rect 94187 21859 94221 21893
rect 1829 21523 1863 21557
rect 94187 21523 94221 21557
rect 1829 21187 1863 21221
rect 94187 21187 94221 21221
rect 1829 20851 1863 20885
rect 94187 20851 94221 20885
rect 1829 20515 1863 20549
rect 94187 20515 94221 20549
rect 1829 20179 1863 20213
rect 94187 20179 94221 20213
rect 1829 19843 1863 19877
rect 94187 19843 94221 19877
rect 1829 19507 1863 19541
rect 94187 19507 94221 19541
rect 1829 19171 1863 19205
rect 94187 19171 94221 19205
rect 1829 18835 1863 18869
rect 94187 18835 94221 18869
rect 1829 18499 1863 18533
rect 94187 18499 94221 18533
rect 1829 18163 1863 18197
rect 94187 18163 94221 18197
rect 1829 17827 1863 17861
rect 94187 17827 94221 17861
rect 1829 17491 1863 17525
rect 94187 17491 94221 17525
rect 1829 17155 1863 17189
rect 94187 17155 94221 17189
rect 1829 16819 1863 16853
rect 94187 16819 94221 16853
rect 1829 16483 1863 16517
rect 94187 16483 94221 16517
rect 1829 16147 1863 16181
rect 94187 16147 94221 16181
rect 1829 15811 1863 15845
rect 94187 15811 94221 15845
rect 1829 15475 1863 15509
rect 94187 15475 94221 15509
rect 1829 15139 1863 15173
rect 94187 15139 94221 15173
rect 1829 14803 1863 14837
rect 94187 14803 94221 14837
rect 1829 14467 1863 14501
rect 94187 14467 94221 14501
rect 1829 14131 1863 14165
rect 94187 14131 94221 14165
rect 1829 13795 1863 13829
rect 94187 13795 94221 13829
rect 1829 13459 1863 13493
rect 94187 13459 94221 13493
rect 1829 13123 1863 13157
rect 94187 13123 94221 13157
rect 1829 12787 1863 12821
rect 94187 12787 94221 12821
rect 1829 12451 1863 12485
rect 94187 12451 94221 12485
rect 1829 12115 1863 12149
rect 94187 12115 94221 12149
rect 1829 11779 1863 11813
rect 94187 11779 94221 11813
rect 1829 11443 1863 11477
rect 94187 11443 94221 11477
rect 1829 11107 1863 11141
rect 94187 11107 94221 11141
rect 1829 10771 1863 10805
rect 94187 10771 94221 10805
rect 1829 10435 1863 10469
rect 94187 10435 94221 10469
rect 1829 10099 1863 10133
rect 94187 10099 94221 10133
rect 1829 9763 1863 9797
rect 94187 9763 94221 9797
rect 1829 9427 1863 9461
rect 94187 9427 94221 9461
rect 1829 9091 1863 9125
rect 94187 9091 94221 9125
rect 1829 8755 1863 8789
rect 94187 8755 94221 8789
rect 1829 8419 1863 8453
rect 94187 8419 94221 8453
rect 1829 8083 1863 8117
rect 94187 8083 94221 8117
rect 1829 7747 1863 7781
rect 94187 7747 94221 7781
rect 1829 7411 1863 7445
rect 94187 7411 94221 7445
rect 1829 7075 1863 7109
rect 94187 7075 94221 7109
rect 1829 6739 1863 6773
rect 94187 6739 94221 6773
rect 1829 6403 1863 6437
rect 94187 6403 94221 6437
rect 1829 6067 1863 6101
rect 94187 6067 94221 6101
rect 1829 5731 1863 5765
rect 94187 5731 94221 5765
rect 1829 5395 1863 5429
rect 94187 5395 94221 5429
rect 1829 5059 1863 5093
rect 94187 5059 94221 5093
rect 1829 4723 1863 4757
rect 94187 4723 94221 4757
rect 1829 4387 1863 4421
rect 94187 4387 94221 4421
rect 1829 4051 1863 4085
rect 94187 4051 94221 4085
rect 1829 3715 1863 3749
rect 94187 3715 94221 3749
rect 1829 3379 1863 3413
rect 94187 3379 94221 3413
rect 1829 3043 1863 3077
rect 94187 3043 94221 3077
rect 1829 2707 1863 2741
rect 94187 2707 94221 2741
rect 1829 2371 1863 2405
rect 94187 2371 94221 2405
rect 1829 2035 1863 2069
rect 94187 2035 94221 2069
rect 2165 1699 2199 1733
rect 2501 1699 2535 1733
rect 2837 1699 2871 1733
rect 3173 1699 3207 1733
rect 3509 1699 3543 1733
rect 3845 1699 3879 1733
rect 4181 1699 4215 1733
rect 4517 1699 4551 1733
rect 4853 1699 4887 1733
rect 5189 1699 5223 1733
rect 5525 1699 5559 1733
rect 5861 1699 5895 1733
rect 6197 1699 6231 1733
rect 6533 1699 6567 1733
rect 6869 1699 6903 1733
rect 7205 1699 7239 1733
rect 7541 1699 7575 1733
rect 7877 1699 7911 1733
rect 8213 1699 8247 1733
rect 8549 1699 8583 1733
rect 8885 1699 8919 1733
rect 9221 1699 9255 1733
rect 9557 1699 9591 1733
rect 9893 1699 9927 1733
rect 10229 1699 10263 1733
rect 10565 1699 10599 1733
rect 10901 1699 10935 1733
rect 11237 1699 11271 1733
rect 11573 1699 11607 1733
rect 11909 1699 11943 1733
rect 12245 1699 12279 1733
rect 12581 1699 12615 1733
rect 12917 1699 12951 1733
rect 13253 1699 13287 1733
rect 13589 1699 13623 1733
rect 13925 1699 13959 1733
rect 14261 1699 14295 1733
rect 14597 1699 14631 1733
rect 14933 1699 14967 1733
rect 15269 1699 15303 1733
rect 15605 1699 15639 1733
rect 15941 1699 15975 1733
rect 16277 1699 16311 1733
rect 16613 1699 16647 1733
rect 16949 1699 16983 1733
rect 17285 1699 17319 1733
rect 17621 1699 17655 1733
rect 17957 1699 17991 1733
rect 18293 1699 18327 1733
rect 18629 1699 18663 1733
rect 18965 1699 18999 1733
rect 19301 1699 19335 1733
rect 19637 1699 19671 1733
rect 19973 1699 20007 1733
rect 20309 1699 20343 1733
rect 20645 1699 20679 1733
rect 20981 1699 21015 1733
rect 21317 1699 21351 1733
rect 21653 1699 21687 1733
rect 21989 1699 22023 1733
rect 22325 1699 22359 1733
rect 22661 1699 22695 1733
rect 22997 1699 23031 1733
rect 23333 1699 23367 1733
rect 23669 1699 23703 1733
rect 24005 1699 24039 1733
rect 24341 1699 24375 1733
rect 24677 1699 24711 1733
rect 25013 1699 25047 1733
rect 25349 1699 25383 1733
rect 25685 1699 25719 1733
rect 26021 1699 26055 1733
rect 26357 1699 26391 1733
rect 26693 1699 26727 1733
rect 27029 1699 27063 1733
rect 27365 1699 27399 1733
rect 27701 1699 27735 1733
rect 28037 1699 28071 1733
rect 28373 1699 28407 1733
rect 28709 1699 28743 1733
rect 29045 1699 29079 1733
rect 29381 1699 29415 1733
rect 29717 1699 29751 1733
rect 30053 1699 30087 1733
rect 30389 1699 30423 1733
rect 30725 1699 30759 1733
rect 31061 1699 31095 1733
rect 31397 1699 31431 1733
rect 31733 1699 31767 1733
rect 32069 1699 32103 1733
rect 32405 1699 32439 1733
rect 32741 1699 32775 1733
rect 33077 1699 33111 1733
rect 33413 1699 33447 1733
rect 33749 1699 33783 1733
rect 34085 1699 34119 1733
rect 34421 1699 34455 1733
rect 34757 1699 34791 1733
rect 35093 1699 35127 1733
rect 35429 1699 35463 1733
rect 35765 1699 35799 1733
rect 36101 1699 36135 1733
rect 36437 1699 36471 1733
rect 36773 1699 36807 1733
rect 37109 1699 37143 1733
rect 37445 1699 37479 1733
rect 37781 1699 37815 1733
rect 38117 1699 38151 1733
rect 38453 1699 38487 1733
rect 38789 1699 38823 1733
rect 39125 1699 39159 1733
rect 39461 1699 39495 1733
rect 39797 1699 39831 1733
rect 40133 1699 40167 1733
rect 40469 1699 40503 1733
rect 40805 1699 40839 1733
rect 41141 1699 41175 1733
rect 41477 1699 41511 1733
rect 41813 1699 41847 1733
rect 42149 1699 42183 1733
rect 42485 1699 42519 1733
rect 42821 1699 42855 1733
rect 43157 1699 43191 1733
rect 43493 1699 43527 1733
rect 43829 1699 43863 1733
rect 44165 1699 44199 1733
rect 44501 1699 44535 1733
rect 44837 1699 44871 1733
rect 45173 1699 45207 1733
rect 45509 1699 45543 1733
rect 45845 1699 45879 1733
rect 46181 1699 46215 1733
rect 46517 1699 46551 1733
rect 46853 1699 46887 1733
rect 47189 1699 47223 1733
rect 47525 1699 47559 1733
rect 47861 1699 47895 1733
rect 48197 1699 48231 1733
rect 48533 1699 48567 1733
rect 48869 1699 48903 1733
rect 49205 1699 49239 1733
rect 49541 1699 49575 1733
rect 49877 1699 49911 1733
rect 50213 1699 50247 1733
rect 50549 1699 50583 1733
rect 50885 1699 50919 1733
rect 51221 1699 51255 1733
rect 51557 1699 51591 1733
rect 51893 1699 51927 1733
rect 52229 1699 52263 1733
rect 52565 1699 52599 1733
rect 52901 1699 52935 1733
rect 53237 1699 53271 1733
rect 53573 1699 53607 1733
rect 53909 1699 53943 1733
rect 54245 1699 54279 1733
rect 54581 1699 54615 1733
rect 54917 1699 54951 1733
rect 55253 1699 55287 1733
rect 55589 1699 55623 1733
rect 55925 1699 55959 1733
rect 56261 1699 56295 1733
rect 56597 1699 56631 1733
rect 56933 1699 56967 1733
rect 57269 1699 57303 1733
rect 57605 1699 57639 1733
rect 57941 1699 57975 1733
rect 58277 1699 58311 1733
rect 58613 1699 58647 1733
rect 58949 1699 58983 1733
rect 59285 1699 59319 1733
rect 59621 1699 59655 1733
rect 59957 1699 59991 1733
rect 60293 1699 60327 1733
rect 60629 1699 60663 1733
rect 60965 1699 60999 1733
rect 61301 1699 61335 1733
rect 61637 1699 61671 1733
rect 61973 1699 62007 1733
rect 62309 1699 62343 1733
rect 62645 1699 62679 1733
rect 62981 1699 63015 1733
rect 63317 1699 63351 1733
rect 63653 1699 63687 1733
rect 63989 1699 64023 1733
rect 64325 1699 64359 1733
rect 64661 1699 64695 1733
rect 64997 1699 65031 1733
rect 65333 1699 65367 1733
rect 65669 1699 65703 1733
rect 66005 1699 66039 1733
rect 66341 1699 66375 1733
rect 66677 1699 66711 1733
rect 67013 1699 67047 1733
rect 67349 1699 67383 1733
rect 67685 1699 67719 1733
rect 68021 1699 68055 1733
rect 68357 1699 68391 1733
rect 68693 1699 68727 1733
rect 69029 1699 69063 1733
rect 69365 1699 69399 1733
rect 69701 1699 69735 1733
rect 70037 1699 70071 1733
rect 70373 1699 70407 1733
rect 70709 1699 70743 1733
rect 71045 1699 71079 1733
rect 71381 1699 71415 1733
rect 71717 1699 71751 1733
rect 72053 1699 72087 1733
rect 72389 1699 72423 1733
rect 72725 1699 72759 1733
rect 73061 1699 73095 1733
rect 73397 1699 73431 1733
rect 73733 1699 73767 1733
rect 74069 1699 74103 1733
rect 74405 1699 74439 1733
rect 74741 1699 74775 1733
rect 75077 1699 75111 1733
rect 75413 1699 75447 1733
rect 75749 1699 75783 1733
rect 76085 1699 76119 1733
rect 76421 1699 76455 1733
rect 76757 1699 76791 1733
rect 77093 1699 77127 1733
rect 77429 1699 77463 1733
rect 77765 1699 77799 1733
rect 78101 1699 78135 1733
rect 78437 1699 78471 1733
rect 78773 1699 78807 1733
rect 79109 1699 79143 1733
rect 79445 1699 79479 1733
rect 79781 1699 79815 1733
rect 80117 1699 80151 1733
rect 80453 1699 80487 1733
rect 80789 1699 80823 1733
rect 81125 1699 81159 1733
rect 81461 1699 81495 1733
rect 81797 1699 81831 1733
rect 82133 1699 82167 1733
rect 82469 1699 82503 1733
rect 82805 1699 82839 1733
rect 83141 1699 83175 1733
rect 83477 1699 83511 1733
rect 83813 1699 83847 1733
rect 84149 1699 84183 1733
rect 84485 1699 84519 1733
rect 84821 1699 84855 1733
rect 85157 1699 85191 1733
rect 85493 1699 85527 1733
rect 85829 1699 85863 1733
rect 86165 1699 86199 1733
rect 86501 1699 86535 1733
rect 86837 1699 86871 1733
rect 87173 1699 87207 1733
rect 87509 1699 87543 1733
rect 87845 1699 87879 1733
rect 88181 1699 88215 1733
rect 88517 1699 88551 1733
rect 88853 1699 88887 1733
rect 89189 1699 89223 1733
rect 89525 1699 89559 1733
rect 89861 1699 89895 1733
rect 90197 1699 90231 1733
rect 90533 1699 90567 1733
rect 90869 1699 90903 1733
rect 91205 1699 91239 1733
rect 91541 1699 91575 1733
rect 91877 1699 91911 1733
rect 92213 1699 92247 1733
rect 92549 1699 92583 1733
rect 92885 1699 92919 1733
rect 93221 1699 93255 1733
rect 93557 1699 93591 1733
<< metal1 >>
rect 1734 77806 94316 77892
rect 1734 77754 2156 77806
rect 2208 77797 3836 77806
rect 3888 77797 5516 77806
rect 5568 77797 7196 77806
rect 7248 77797 8876 77806
rect 8928 77797 10556 77806
rect 10608 77797 12236 77806
rect 12288 77797 13916 77806
rect 13968 77797 15596 77806
rect 15648 77797 17276 77806
rect 17328 77797 18956 77806
rect 19008 77797 20636 77806
rect 20688 77797 22316 77806
rect 22368 77797 23996 77806
rect 24048 77797 25676 77806
rect 25728 77797 27356 77806
rect 27408 77797 29036 77806
rect 29088 77797 30716 77806
rect 30768 77797 32396 77806
rect 32448 77797 34076 77806
rect 34128 77797 35756 77806
rect 35808 77797 37436 77806
rect 37488 77797 39116 77806
rect 39168 77797 40796 77806
rect 40848 77797 42476 77806
rect 42528 77797 44156 77806
rect 44208 77797 45836 77806
rect 45888 77797 47516 77806
rect 47568 77797 49196 77806
rect 49248 77797 50876 77806
rect 50928 77797 52556 77806
rect 52608 77797 54236 77806
rect 54288 77797 55916 77806
rect 55968 77797 57596 77806
rect 57648 77797 59276 77806
rect 59328 77797 60956 77806
rect 61008 77797 62636 77806
rect 62688 77797 64316 77806
rect 64368 77797 65996 77806
rect 66048 77797 67676 77806
rect 67728 77797 69356 77806
rect 69408 77797 71036 77806
rect 71088 77797 72716 77806
rect 72768 77797 74396 77806
rect 74448 77797 76076 77806
rect 76128 77797 77756 77806
rect 77808 77797 79436 77806
rect 79488 77797 81116 77806
rect 81168 77797 82796 77806
rect 82848 77797 84476 77806
rect 84528 77797 86156 77806
rect 86208 77797 87836 77806
rect 87888 77797 89516 77806
rect 89568 77797 91196 77806
rect 91248 77797 92876 77806
rect 92928 77797 94316 77806
rect 2208 77763 2501 77797
rect 2535 77763 2837 77797
rect 2871 77763 3173 77797
rect 3207 77763 3509 77797
rect 3543 77763 3836 77797
rect 3888 77763 4181 77797
rect 4215 77763 4517 77797
rect 4551 77763 4853 77797
rect 4887 77763 5189 77797
rect 5223 77763 5516 77797
rect 5568 77763 5861 77797
rect 5895 77763 6197 77797
rect 6231 77763 6533 77797
rect 6567 77763 6869 77797
rect 6903 77763 7196 77797
rect 7248 77763 7541 77797
rect 7575 77763 7877 77797
rect 7911 77763 8213 77797
rect 8247 77763 8549 77797
rect 8583 77763 8876 77797
rect 8928 77763 9221 77797
rect 9255 77763 9557 77797
rect 9591 77763 9893 77797
rect 9927 77763 10229 77797
rect 10263 77763 10556 77797
rect 10608 77763 10901 77797
rect 10935 77763 11237 77797
rect 11271 77763 11573 77797
rect 11607 77763 11909 77797
rect 11943 77763 12236 77797
rect 12288 77763 12581 77797
rect 12615 77763 12917 77797
rect 12951 77763 13253 77797
rect 13287 77763 13589 77797
rect 13623 77763 13916 77797
rect 13968 77763 14261 77797
rect 14295 77763 14597 77797
rect 14631 77763 14933 77797
rect 14967 77763 15269 77797
rect 15303 77763 15596 77797
rect 15648 77763 15941 77797
rect 15975 77763 16277 77797
rect 16311 77763 16613 77797
rect 16647 77763 16949 77797
rect 16983 77763 17276 77797
rect 17328 77763 17621 77797
rect 17655 77763 17957 77797
rect 17991 77763 18293 77797
rect 18327 77763 18629 77797
rect 18663 77763 18956 77797
rect 19008 77763 19301 77797
rect 19335 77763 19637 77797
rect 19671 77763 19973 77797
rect 20007 77763 20309 77797
rect 20343 77763 20636 77797
rect 20688 77763 20981 77797
rect 21015 77763 21317 77797
rect 21351 77763 21653 77797
rect 21687 77763 21989 77797
rect 22023 77763 22316 77797
rect 22368 77763 22661 77797
rect 22695 77763 22997 77797
rect 23031 77763 23333 77797
rect 23367 77763 23669 77797
rect 23703 77763 23996 77797
rect 24048 77763 24341 77797
rect 24375 77763 24677 77797
rect 24711 77763 25013 77797
rect 25047 77763 25349 77797
rect 25383 77763 25676 77797
rect 25728 77763 26021 77797
rect 26055 77763 26357 77797
rect 26391 77763 26693 77797
rect 26727 77763 27029 77797
rect 27063 77763 27356 77797
rect 27408 77763 27701 77797
rect 27735 77763 28037 77797
rect 28071 77763 28373 77797
rect 28407 77763 28709 77797
rect 28743 77763 29036 77797
rect 29088 77763 29381 77797
rect 29415 77763 29717 77797
rect 29751 77763 30053 77797
rect 30087 77763 30389 77797
rect 30423 77763 30716 77797
rect 30768 77763 31061 77797
rect 31095 77763 31397 77797
rect 31431 77763 31733 77797
rect 31767 77763 32069 77797
rect 32103 77763 32396 77797
rect 32448 77763 32741 77797
rect 32775 77763 33077 77797
rect 33111 77763 33413 77797
rect 33447 77763 33749 77797
rect 33783 77763 34076 77797
rect 34128 77763 34421 77797
rect 34455 77763 34757 77797
rect 34791 77763 35093 77797
rect 35127 77763 35429 77797
rect 35463 77763 35756 77797
rect 35808 77763 36101 77797
rect 36135 77763 36437 77797
rect 36471 77763 36773 77797
rect 36807 77763 37109 77797
rect 37143 77763 37436 77797
rect 37488 77763 37781 77797
rect 37815 77763 38117 77797
rect 38151 77763 38453 77797
rect 38487 77763 38789 77797
rect 38823 77763 39116 77797
rect 39168 77763 39461 77797
rect 39495 77763 39797 77797
rect 39831 77763 40133 77797
rect 40167 77763 40469 77797
rect 40503 77763 40796 77797
rect 40848 77763 41141 77797
rect 41175 77763 41477 77797
rect 41511 77763 41813 77797
rect 41847 77763 42149 77797
rect 42183 77763 42476 77797
rect 42528 77763 42821 77797
rect 42855 77763 43157 77797
rect 43191 77763 43493 77797
rect 43527 77763 43829 77797
rect 43863 77763 44156 77797
rect 44208 77763 44501 77797
rect 44535 77763 44837 77797
rect 44871 77763 45173 77797
rect 45207 77763 45509 77797
rect 45543 77763 45836 77797
rect 45888 77763 46181 77797
rect 46215 77763 46517 77797
rect 46551 77763 46853 77797
rect 46887 77763 47189 77797
rect 47223 77763 47516 77797
rect 47568 77763 47861 77797
rect 47895 77763 48197 77797
rect 48231 77763 48533 77797
rect 48567 77763 48869 77797
rect 48903 77763 49196 77797
rect 49248 77763 49541 77797
rect 49575 77763 49877 77797
rect 49911 77763 50213 77797
rect 50247 77763 50549 77797
rect 50583 77763 50876 77797
rect 50928 77763 51221 77797
rect 51255 77763 51557 77797
rect 51591 77763 51893 77797
rect 51927 77763 52229 77797
rect 52263 77763 52556 77797
rect 52608 77763 52901 77797
rect 52935 77763 53237 77797
rect 53271 77763 53573 77797
rect 53607 77763 53909 77797
rect 53943 77763 54236 77797
rect 54288 77763 54581 77797
rect 54615 77763 54917 77797
rect 54951 77763 55253 77797
rect 55287 77763 55589 77797
rect 55623 77763 55916 77797
rect 55968 77763 56261 77797
rect 56295 77763 56597 77797
rect 56631 77763 56933 77797
rect 56967 77763 57269 77797
rect 57303 77763 57596 77797
rect 57648 77763 57941 77797
rect 57975 77763 58277 77797
rect 58311 77763 58613 77797
rect 58647 77763 58949 77797
rect 58983 77763 59276 77797
rect 59328 77763 59621 77797
rect 59655 77763 59957 77797
rect 59991 77763 60293 77797
rect 60327 77763 60629 77797
rect 60663 77763 60956 77797
rect 61008 77763 61301 77797
rect 61335 77763 61637 77797
rect 61671 77763 61973 77797
rect 62007 77763 62309 77797
rect 62343 77763 62636 77797
rect 62688 77763 62981 77797
rect 63015 77763 63317 77797
rect 63351 77763 63653 77797
rect 63687 77763 63989 77797
rect 64023 77763 64316 77797
rect 64368 77763 64661 77797
rect 64695 77763 64997 77797
rect 65031 77763 65333 77797
rect 65367 77763 65669 77797
rect 65703 77763 65996 77797
rect 66048 77763 66341 77797
rect 66375 77763 66677 77797
rect 66711 77763 67013 77797
rect 67047 77763 67349 77797
rect 67383 77763 67676 77797
rect 67728 77763 68021 77797
rect 68055 77763 68357 77797
rect 68391 77763 68693 77797
rect 68727 77763 69029 77797
rect 69063 77763 69356 77797
rect 69408 77763 69701 77797
rect 69735 77763 70037 77797
rect 70071 77763 70373 77797
rect 70407 77763 70709 77797
rect 70743 77763 71036 77797
rect 71088 77763 71381 77797
rect 71415 77763 71717 77797
rect 71751 77763 72053 77797
rect 72087 77763 72389 77797
rect 72423 77763 72716 77797
rect 72768 77763 73061 77797
rect 73095 77763 73397 77797
rect 73431 77763 73733 77797
rect 73767 77763 74069 77797
rect 74103 77763 74396 77797
rect 74448 77763 74741 77797
rect 74775 77763 75077 77797
rect 75111 77763 75413 77797
rect 75447 77763 75749 77797
rect 75783 77763 76076 77797
rect 76128 77763 76421 77797
rect 76455 77763 76757 77797
rect 76791 77763 77093 77797
rect 77127 77763 77429 77797
rect 77463 77763 77756 77797
rect 77808 77763 78101 77797
rect 78135 77763 78437 77797
rect 78471 77763 78773 77797
rect 78807 77763 79109 77797
rect 79143 77763 79436 77797
rect 79488 77763 79781 77797
rect 79815 77763 80117 77797
rect 80151 77763 80453 77797
rect 80487 77763 80789 77797
rect 80823 77763 81116 77797
rect 81168 77763 81461 77797
rect 81495 77763 81797 77797
rect 81831 77763 82133 77797
rect 82167 77763 82469 77797
rect 82503 77763 82796 77797
rect 82848 77763 83141 77797
rect 83175 77763 83477 77797
rect 83511 77763 83813 77797
rect 83847 77763 84149 77797
rect 84183 77763 84476 77797
rect 84528 77763 84821 77797
rect 84855 77763 85157 77797
rect 85191 77763 85493 77797
rect 85527 77763 85829 77797
rect 85863 77763 86156 77797
rect 86208 77763 86501 77797
rect 86535 77763 86837 77797
rect 86871 77763 87173 77797
rect 87207 77763 87509 77797
rect 87543 77763 87836 77797
rect 87888 77763 88181 77797
rect 88215 77763 88517 77797
rect 88551 77763 88853 77797
rect 88887 77763 89189 77797
rect 89223 77763 89516 77797
rect 89568 77763 89861 77797
rect 89895 77763 90197 77797
rect 90231 77763 90533 77797
rect 90567 77763 90869 77797
rect 90903 77763 91196 77797
rect 91248 77763 91541 77797
rect 91575 77763 91877 77797
rect 91911 77763 92213 77797
rect 92247 77763 92549 77797
rect 92583 77763 92876 77797
rect 92928 77763 93221 77797
rect 93255 77763 93557 77797
rect 93591 77763 94316 77797
rect 2208 77754 3836 77763
rect 3888 77754 5516 77763
rect 5568 77754 7196 77763
rect 7248 77754 8876 77763
rect 8928 77754 10556 77763
rect 10608 77754 12236 77763
rect 12288 77754 13916 77763
rect 13968 77754 15596 77763
rect 15648 77754 17276 77763
rect 17328 77754 18956 77763
rect 19008 77754 20636 77763
rect 20688 77754 22316 77763
rect 22368 77754 23996 77763
rect 24048 77754 25676 77763
rect 25728 77754 27356 77763
rect 27408 77754 29036 77763
rect 29088 77754 30716 77763
rect 30768 77754 32396 77763
rect 32448 77754 34076 77763
rect 34128 77754 35756 77763
rect 35808 77754 37436 77763
rect 37488 77754 39116 77763
rect 39168 77754 40796 77763
rect 40848 77754 42476 77763
rect 42528 77754 44156 77763
rect 44208 77754 45836 77763
rect 45888 77754 47516 77763
rect 47568 77754 49196 77763
rect 49248 77754 50876 77763
rect 50928 77754 52556 77763
rect 52608 77754 54236 77763
rect 54288 77754 55916 77763
rect 55968 77754 57596 77763
rect 57648 77754 59276 77763
rect 59328 77754 60956 77763
rect 61008 77754 62636 77763
rect 62688 77754 64316 77763
rect 64368 77754 65996 77763
rect 66048 77754 67676 77763
rect 67728 77754 69356 77763
rect 69408 77754 71036 77763
rect 71088 77754 72716 77763
rect 72768 77754 74396 77763
rect 74448 77754 76076 77763
rect 76128 77754 77756 77763
rect 77808 77754 79436 77763
rect 79488 77754 81116 77763
rect 81168 77754 82796 77763
rect 82848 77754 84476 77763
rect 84528 77754 86156 77763
rect 86208 77754 87836 77763
rect 87888 77754 89516 77763
rect 89568 77754 91196 77763
rect 91248 77754 92876 77763
rect 92928 77754 94316 77763
rect 1734 77668 94316 77754
rect 1814 77290 1820 77342
rect 1872 77290 1878 77342
rect 94172 77290 94178 77342
rect 94230 77290 94236 77342
rect 1814 76954 1820 77006
rect 1872 76954 1878 77006
rect 94172 76954 94178 77006
rect 94230 76954 94236 77006
rect 1814 76618 1820 76670
rect 1872 76618 1878 76670
rect 94172 76618 94178 76670
rect 94230 76618 94236 76670
rect 1814 76282 1820 76334
rect 1872 76282 1878 76334
rect 94172 76282 94178 76334
rect 94230 76282 94236 76334
rect 1814 75946 1820 75998
rect 1872 75946 1878 75998
rect 94172 75946 94178 75998
rect 94230 75946 94236 75998
rect 1814 75610 1820 75662
rect 1872 75610 1878 75662
rect 94172 75610 94178 75662
rect 94230 75610 94236 75662
rect 1814 75274 1820 75326
rect 1872 75274 1878 75326
rect 94172 75274 94178 75326
rect 94230 75274 94236 75326
rect 1814 74938 1820 74990
rect 1872 74938 1878 74990
rect 94172 74938 94178 74990
rect 94230 74938 94236 74990
rect 1814 74602 1820 74654
rect 1872 74602 1878 74654
rect 94172 74602 94178 74654
rect 94230 74602 94236 74654
rect 1814 74266 1820 74318
rect 1872 74266 1878 74318
rect 94172 74266 94178 74318
rect 94230 74266 94236 74318
rect 28206 74049 28212 74101
rect 28264 74049 28270 74101
rect 29454 74049 29460 74101
rect 29512 74049 29518 74101
rect 30702 74049 30708 74101
rect 30760 74049 30766 74101
rect 31950 74049 31956 74101
rect 32008 74049 32014 74101
rect 33198 74049 33204 74101
rect 33256 74049 33262 74101
rect 34446 74049 34452 74101
rect 34504 74049 34510 74101
rect 35694 74049 35700 74101
rect 35752 74049 35758 74101
rect 36942 74049 36948 74101
rect 37000 74049 37006 74101
rect 38190 74049 38196 74101
rect 38248 74049 38254 74101
rect 39438 74049 39444 74101
rect 39496 74049 39502 74101
rect 40686 74049 40692 74101
rect 40744 74049 40750 74101
rect 41934 74049 41940 74101
rect 41992 74049 41998 74101
rect 43182 74049 43188 74101
rect 43240 74049 43246 74101
rect 44430 74049 44436 74101
rect 44488 74049 44494 74101
rect 45678 74049 45684 74101
rect 45736 74049 45742 74101
rect 46926 74049 46932 74101
rect 46984 74049 46990 74101
rect 48174 74049 48180 74101
rect 48232 74049 48238 74101
rect 49422 74049 49428 74101
rect 49480 74049 49486 74101
rect 50670 74049 50676 74101
rect 50728 74049 50734 74101
rect 51918 74049 51924 74101
rect 51976 74049 51982 74101
rect 53166 74049 53172 74101
rect 53224 74049 53230 74101
rect 54414 74049 54420 74101
rect 54472 74049 54478 74101
rect 55662 74049 55668 74101
rect 55720 74049 55726 74101
rect 56910 74049 56916 74101
rect 56968 74049 56974 74101
rect 58158 74049 58164 74101
rect 58216 74049 58222 74101
rect 59406 74049 59412 74101
rect 59464 74049 59470 74101
rect 60654 74049 60660 74101
rect 60712 74049 60718 74101
rect 61902 74049 61908 74101
rect 61960 74049 61966 74101
rect 63150 74049 63156 74101
rect 63208 74049 63214 74101
rect 64398 74049 64404 74101
rect 64456 74049 64462 74101
rect 65646 74049 65652 74101
rect 65704 74049 65710 74101
rect 66894 74049 66900 74101
rect 66952 74049 66958 74101
rect 1814 73930 1820 73982
rect 1872 73930 1878 73982
rect 94172 73930 94178 73982
rect 94230 73930 94236 73982
rect 1814 73594 1820 73646
rect 1872 73594 1878 73646
rect 94172 73594 94178 73646
rect 94230 73594 94236 73646
rect 1814 73258 1820 73310
rect 1872 73258 1878 73310
rect 94172 73258 94178 73310
rect 94230 73258 94236 73310
rect 1814 72922 1820 72974
rect 1872 72922 1878 72974
rect 94172 72922 94178 72974
rect 94230 72922 94236 72974
rect 1814 72586 1820 72638
rect 1872 72586 1878 72638
rect 94172 72586 94178 72638
rect 94230 72586 94236 72638
rect 1814 72250 1820 72302
rect 1872 72250 1878 72302
rect 94172 72250 94178 72302
rect 94230 72250 94236 72302
rect 1814 71914 1820 71966
rect 1872 71914 1878 71966
rect 94172 71914 94178 71966
rect 94230 71914 94236 71966
rect 1814 71578 1820 71630
rect 1872 71578 1878 71630
rect 94172 71578 94178 71630
rect 94230 71578 94236 71630
rect 1814 71242 1820 71294
rect 1872 71242 1878 71294
rect 94172 71242 94178 71294
rect 94230 71242 94236 71294
rect 1814 70906 1820 70958
rect 1872 70906 1878 70958
rect 94172 70906 94178 70958
rect 94230 70906 94236 70958
rect 1814 70570 1820 70622
rect 1872 70570 1878 70622
rect 94172 70570 94178 70622
rect 94230 70570 94236 70622
rect 1814 70234 1820 70286
rect 1872 70234 1878 70286
rect 94172 70234 94178 70286
rect 94230 70234 94236 70286
rect 1814 69898 1820 69950
rect 1872 69898 1878 69950
rect 94172 69898 94178 69950
rect 94230 69898 94236 69950
rect 1814 69562 1820 69614
rect 1872 69562 1878 69614
rect 94172 69562 94178 69614
rect 94230 69562 94236 69614
rect 1814 69226 1820 69278
rect 1872 69226 1878 69278
rect 94172 69226 94178 69278
rect 94230 69226 94236 69278
rect 1814 68890 1820 68942
rect 1872 68890 1878 68942
rect 94172 68890 94178 68942
rect 94230 68890 94236 68942
rect 1814 68554 1820 68606
rect 1872 68554 1878 68606
rect 94172 68554 94178 68606
rect 94230 68554 94236 68606
rect 1814 68218 1820 68270
rect 1872 68218 1878 68270
rect 94172 68218 94178 68270
rect 94230 68218 94236 68270
rect 1814 67882 1820 67934
rect 1872 67882 1878 67934
rect 94172 67882 94178 67934
rect 94230 67882 94236 67934
rect 1814 67546 1820 67598
rect 1872 67546 1878 67598
rect 94172 67546 94178 67598
rect 94230 67546 94236 67598
rect 1814 67210 1820 67262
rect 1872 67210 1878 67262
rect 94172 67210 94178 67262
rect 94230 67210 94236 67262
rect 1814 66874 1820 66926
rect 1872 66874 1878 66926
rect 94172 66874 94178 66926
rect 94230 66874 94236 66926
rect 1814 66538 1820 66590
rect 1872 66538 1878 66590
rect 94172 66538 94178 66590
rect 94230 66538 94236 66590
rect 1814 66202 1820 66254
rect 1872 66202 1878 66254
rect 94172 66202 94178 66254
rect 94230 66202 94236 66254
rect 1814 65866 1820 65918
rect 1872 65866 1878 65918
rect 94172 65866 94178 65918
rect 94230 65866 94236 65918
rect 1814 65530 1820 65582
rect 1872 65530 1878 65582
rect 94172 65530 94178 65582
rect 94230 65530 94236 65582
rect 1814 65194 1820 65246
rect 1872 65194 1878 65246
rect 94172 65194 94178 65246
rect 94230 65194 94236 65246
rect 1814 64858 1820 64910
rect 1872 64858 1878 64910
rect 94172 64858 94178 64910
rect 94230 64858 94236 64910
rect 1814 64522 1820 64574
rect 1872 64522 1878 64574
rect 94172 64522 94178 64574
rect 94230 64522 94236 64574
rect 1814 64186 1820 64238
rect 1872 64186 1878 64238
rect 94172 64186 94178 64238
rect 94230 64186 94236 64238
rect 1814 63850 1820 63902
rect 1872 63850 1878 63902
rect 94172 63850 94178 63902
rect 94230 63850 94236 63902
rect 1814 63514 1820 63566
rect 1872 63514 1878 63566
rect 94172 63514 94178 63566
rect 94230 63514 94236 63566
rect 1814 63178 1820 63230
rect 1872 63178 1878 63230
rect 94172 63178 94178 63230
rect 94230 63178 94236 63230
rect 1814 62842 1820 62894
rect 1872 62842 1878 62894
rect 94172 62842 94178 62894
rect 94230 62842 94236 62894
rect 1814 62506 1820 62558
rect 1872 62506 1878 62558
rect 94172 62506 94178 62558
rect 94230 62506 94236 62558
rect 1814 62170 1820 62222
rect 1872 62170 1878 62222
rect 94172 62170 94178 62222
rect 94230 62170 94236 62222
rect 1814 61834 1820 61886
rect 1872 61834 1878 61886
rect 94172 61834 94178 61886
rect 94230 61834 94236 61886
rect 1814 61498 1820 61550
rect 1872 61498 1878 61550
rect 94172 61498 94178 61550
rect 94230 61498 94236 61550
rect 1814 61162 1820 61214
rect 1872 61162 1878 61214
rect 94172 61162 94178 61214
rect 94230 61162 94236 61214
rect 1814 60826 1820 60878
rect 1872 60826 1878 60878
rect 94172 60826 94178 60878
rect 94230 60826 94236 60878
rect 1814 60490 1820 60542
rect 1872 60490 1878 60542
rect 94172 60490 94178 60542
rect 94230 60490 94236 60542
rect 1814 60154 1820 60206
rect 1872 60154 1878 60206
rect 94172 60154 94178 60206
rect 94230 60154 94236 60206
rect 1814 59818 1820 59870
rect 1872 59818 1878 59870
rect 94172 59818 94178 59870
rect 94230 59818 94236 59870
rect 1814 59482 1820 59534
rect 1872 59482 1878 59534
rect 94172 59482 94178 59534
rect 94230 59482 94236 59534
rect 1814 59146 1820 59198
rect 1872 59146 1878 59198
rect 94172 59146 94178 59198
rect 94230 59146 94236 59198
rect 1814 58810 1820 58862
rect 1872 58810 1878 58862
rect 94172 58810 94178 58862
rect 94230 58810 94236 58862
rect 1814 58474 1820 58526
rect 1872 58474 1878 58526
rect 94172 58474 94178 58526
rect 94230 58474 94236 58526
rect 1814 58138 1820 58190
rect 1872 58138 1878 58190
rect 94172 58138 94178 58190
rect 94230 58138 94236 58190
rect 1814 57802 1820 57854
rect 1872 57802 1878 57854
rect 94172 57802 94178 57854
rect 94230 57802 94236 57854
rect 1814 57466 1820 57518
rect 1872 57466 1878 57518
rect 94172 57466 94178 57518
rect 94230 57466 94236 57518
rect 1814 57130 1820 57182
rect 1872 57130 1878 57182
rect 94172 57130 94178 57182
rect 94230 57130 94236 57182
rect 1814 56794 1820 56846
rect 1872 56794 1878 56846
rect 94172 56794 94178 56846
rect 94230 56794 94236 56846
rect 1814 56458 1820 56510
rect 1872 56458 1878 56510
rect 94172 56458 94178 56510
rect 94230 56458 94236 56510
rect 1814 56122 1820 56174
rect 1872 56122 1878 56174
rect 94172 56122 94178 56174
rect 94230 56122 94236 56174
rect 1814 55786 1820 55838
rect 1872 55786 1878 55838
rect 94172 55786 94178 55838
rect 94230 55786 94236 55838
rect 1814 55450 1820 55502
rect 1872 55450 1878 55502
rect 94172 55450 94178 55502
rect 94230 55450 94236 55502
rect 1814 55114 1820 55166
rect 1872 55114 1878 55166
rect 94172 55114 94178 55166
rect 94230 55114 94236 55166
rect 1814 54778 1820 54830
rect 1872 54778 1878 54830
rect 94172 54778 94178 54830
rect 94230 54778 94236 54830
rect 1814 54442 1820 54494
rect 1872 54442 1878 54494
rect 94172 54442 94178 54494
rect 94230 54442 94236 54494
rect 1814 54106 1820 54158
rect 1872 54106 1878 54158
rect 94172 54106 94178 54158
rect 94230 54106 94236 54158
rect 1814 53770 1820 53822
rect 1872 53770 1878 53822
rect 94172 53770 94178 53822
rect 94230 53770 94236 53822
rect 1814 53434 1820 53486
rect 1872 53434 1878 53486
rect 94172 53434 94178 53486
rect 94230 53434 94236 53486
rect 1814 53098 1820 53150
rect 1872 53098 1878 53150
rect 94172 53098 94178 53150
rect 94230 53098 94236 53150
rect 1814 52762 1820 52814
rect 1872 52762 1878 52814
rect 94172 52762 94178 52814
rect 94230 52762 94236 52814
rect 1814 52426 1820 52478
rect 1872 52426 1878 52478
rect 94172 52426 94178 52478
rect 94230 52426 94236 52478
rect 1814 52090 1820 52142
rect 1872 52090 1878 52142
rect 94172 52090 94178 52142
rect 94230 52090 94236 52142
rect 1814 51754 1820 51806
rect 1872 51754 1878 51806
rect 94172 51754 94178 51806
rect 94230 51754 94236 51806
rect 1814 51418 1820 51470
rect 1872 51418 1878 51470
rect 94172 51418 94178 51470
rect 94230 51418 94236 51470
rect 1814 51082 1820 51134
rect 1872 51082 1878 51134
rect 94172 51082 94178 51134
rect 94230 51082 94236 51134
rect 1814 50746 1820 50798
rect 1872 50746 1878 50798
rect 94172 50746 94178 50798
rect 94230 50746 94236 50798
rect 1814 50410 1820 50462
rect 1872 50410 1878 50462
rect 94172 50410 94178 50462
rect 94230 50410 94236 50462
rect 1814 50074 1820 50126
rect 1872 50074 1878 50126
rect 94172 50074 94178 50126
rect 94230 50074 94236 50126
rect 1814 49738 1820 49790
rect 1872 49738 1878 49790
rect 94172 49738 94178 49790
rect 94230 49738 94236 49790
rect 1814 49402 1820 49454
rect 1872 49402 1878 49454
rect 94172 49402 94178 49454
rect 94230 49402 94236 49454
rect 1814 49066 1820 49118
rect 1872 49066 1878 49118
rect 94172 49066 94178 49118
rect 94230 49066 94236 49118
rect 1814 48730 1820 48782
rect 1872 48730 1878 48782
rect 94172 48730 94178 48782
rect 94230 48730 94236 48782
rect 1814 48394 1820 48446
rect 1872 48394 1878 48446
rect 94172 48394 94178 48446
rect 94230 48394 94236 48446
rect 1814 48058 1820 48110
rect 1872 48058 1878 48110
rect 94172 48058 94178 48110
rect 94230 48058 94236 48110
rect 1814 47722 1820 47774
rect 1872 47722 1878 47774
rect 94172 47722 94178 47774
rect 94230 47722 94236 47774
rect 1814 47386 1820 47438
rect 1872 47386 1878 47438
rect 94172 47386 94178 47438
rect 94230 47386 94236 47438
rect 1814 47050 1820 47102
rect 1872 47050 1878 47102
rect 94172 47050 94178 47102
rect 94230 47050 94236 47102
rect 1814 46714 1820 46766
rect 1872 46714 1878 46766
rect 94172 46714 94178 46766
rect 94230 46714 94236 46766
rect 1814 46378 1820 46430
rect 1872 46378 1878 46430
rect 94172 46378 94178 46430
rect 94230 46378 94236 46430
rect 1814 46042 1820 46094
rect 1872 46042 1878 46094
rect 94172 46042 94178 46094
rect 94230 46042 94236 46094
rect 1814 45706 1820 45758
rect 1872 45706 1878 45758
rect 94172 45706 94178 45758
rect 94230 45706 94236 45758
rect 1814 45370 1820 45422
rect 1872 45370 1878 45422
rect 94172 45370 94178 45422
rect 94230 45370 94236 45422
rect 1814 45034 1820 45086
rect 1872 45034 1878 45086
rect 94172 45034 94178 45086
rect 94230 45034 94236 45086
rect 1814 44698 1820 44750
rect 1872 44698 1878 44750
rect 94172 44698 94178 44750
rect 94230 44698 94236 44750
rect 1814 44362 1820 44414
rect 1872 44362 1878 44414
rect 94172 44362 94178 44414
rect 94230 44362 94236 44414
rect 1814 44026 1820 44078
rect 1872 44026 1878 44078
rect 94172 44026 94178 44078
rect 94230 44026 94236 44078
rect 1814 43690 1820 43742
rect 1872 43690 1878 43742
rect 94172 43690 94178 43742
rect 94230 43690 94236 43742
rect 1814 43354 1820 43406
rect 1872 43354 1878 43406
rect 94172 43354 94178 43406
rect 94230 43354 94236 43406
rect 1814 43018 1820 43070
rect 1872 43018 1878 43070
rect 94172 43018 94178 43070
rect 94230 43018 94236 43070
rect 1814 42682 1820 42734
rect 1872 42682 1878 42734
rect 94172 42682 94178 42734
rect 94230 42682 94236 42734
rect 1814 42346 1820 42398
rect 1872 42346 1878 42398
rect 94172 42346 94178 42398
rect 94230 42346 94236 42398
rect 1814 42010 1820 42062
rect 1872 42010 1878 42062
rect 94172 42010 94178 42062
rect 94230 42010 94236 42062
rect 1814 41674 1820 41726
rect 1872 41674 1878 41726
rect 94172 41674 94178 41726
rect 94230 41674 94236 41726
rect 1814 41338 1820 41390
rect 1872 41338 1878 41390
rect 94172 41338 94178 41390
rect 94230 41338 94236 41390
rect 1814 41002 1820 41054
rect 1872 41002 1878 41054
rect 94172 41002 94178 41054
rect 94230 41002 94236 41054
rect 1814 40666 1820 40718
rect 1872 40666 1878 40718
rect 94172 40666 94178 40718
rect 94230 40666 94236 40718
rect 1814 40330 1820 40382
rect 1872 40330 1878 40382
rect 94172 40330 94178 40382
rect 94230 40330 94236 40382
rect 1814 39994 1820 40046
rect 1872 39994 1878 40046
rect 94172 39994 94178 40046
rect 94230 39994 94236 40046
rect 1814 39658 1820 39710
rect 1872 39658 1878 39710
rect 94172 39658 94178 39710
rect 94230 39658 94236 39710
rect 1814 39322 1820 39374
rect 1872 39322 1878 39374
rect 94172 39322 94178 39374
rect 94230 39322 94236 39374
rect 1814 38986 1820 39038
rect 1872 38986 1878 39038
rect 94172 38986 94178 39038
rect 94230 38986 94236 39038
rect 1814 38650 1820 38702
rect 1872 38650 1878 38702
rect 94172 38650 94178 38702
rect 94230 38650 94236 38702
rect 1814 38314 1820 38366
rect 1872 38314 1878 38366
rect 94172 38314 94178 38366
rect 94230 38314 94236 38366
rect 1814 37978 1820 38030
rect 1872 37978 1878 38030
rect 94172 37978 94178 38030
rect 94230 37978 94236 38030
rect 1814 37642 1820 37694
rect 1872 37642 1878 37694
rect 94172 37642 94178 37694
rect 94230 37642 94236 37694
rect 1814 37306 1820 37358
rect 1872 37306 1878 37358
rect 94172 37306 94178 37358
rect 94230 37306 94236 37358
rect 1814 36970 1820 37022
rect 1872 36970 1878 37022
rect 94172 36970 94178 37022
rect 94230 36970 94236 37022
rect 1814 36634 1820 36686
rect 1872 36634 1878 36686
rect 94172 36634 94178 36686
rect 94230 36634 94236 36686
rect 1814 36298 1820 36350
rect 1872 36298 1878 36350
rect 94172 36298 94178 36350
rect 94230 36298 94236 36350
rect 1814 35962 1820 36014
rect 1872 35962 1878 36014
rect 94172 35962 94178 36014
rect 94230 35962 94236 36014
rect 1814 35626 1820 35678
rect 1872 35626 1878 35678
rect 94172 35626 94178 35678
rect 94230 35626 94236 35678
rect 1814 35290 1820 35342
rect 1872 35290 1878 35342
rect 94172 35290 94178 35342
rect 94230 35290 94236 35342
rect 1814 34954 1820 35006
rect 1872 34954 1878 35006
rect 94172 34954 94178 35006
rect 94230 34954 94236 35006
rect 1814 34618 1820 34670
rect 1872 34618 1878 34670
rect 94172 34618 94178 34670
rect 94230 34618 94236 34670
rect 1814 34282 1820 34334
rect 1872 34282 1878 34334
rect 94172 34282 94178 34334
rect 94230 34282 94236 34334
rect 14935 34143 14941 34195
rect 14993 34143 14999 34195
rect 1814 33946 1820 33998
rect 1872 33946 1878 33998
rect 1814 33610 1820 33662
rect 1872 33610 1878 33662
rect 1814 33274 1820 33326
rect 1872 33274 1878 33326
rect 1814 32938 1820 32990
rect 1872 32938 1878 32990
rect 14855 32873 14861 32925
rect 14913 32873 14919 32925
rect 1814 32602 1820 32654
rect 1872 32602 1878 32654
rect 1814 32266 1820 32318
rect 1872 32266 1878 32318
rect 1814 31930 1820 31982
rect 1872 31930 1878 31982
rect 1814 31594 1820 31646
rect 1872 31594 1878 31646
rect 14775 31315 14781 31367
rect 14833 31315 14839 31367
rect 1814 31258 1820 31310
rect 1872 31258 1878 31310
rect 1814 30922 1820 30974
rect 1872 30922 1878 30974
rect 1814 30586 1820 30638
rect 1872 30586 1878 30638
rect 1814 30250 1820 30302
rect 1872 30250 1878 30302
rect 14695 30045 14701 30097
rect 14753 30045 14759 30097
rect 1814 29914 1820 29966
rect 1872 29914 1878 29966
rect 1814 29578 1820 29630
rect 1872 29578 1878 29630
rect 1814 29242 1820 29294
rect 1872 29242 1878 29294
rect 1814 28906 1820 28958
rect 1872 28906 1878 28958
rect 1814 28570 1820 28622
rect 1872 28570 1878 28622
rect 14615 28487 14621 28539
rect 14673 28487 14679 28539
rect 1814 28234 1820 28286
rect 1872 28234 1878 28286
rect 1814 27898 1820 27950
rect 1872 27898 1878 27950
rect 1814 27562 1820 27614
rect 1872 27562 1878 27614
rect 1814 27226 1820 27278
rect 1872 27226 1878 27278
rect 14535 27217 14541 27269
rect 14593 27217 14599 27269
rect 1814 26890 1820 26942
rect 1872 26890 1878 26942
rect 1814 26554 1820 26606
rect 1872 26554 1878 26606
rect 1814 26218 1820 26270
rect 1872 26218 1878 26270
rect 1814 25882 1820 25934
rect 1872 25882 1878 25934
rect 14455 25659 14461 25711
rect 14513 25659 14519 25711
rect 1814 25546 1820 25598
rect 1872 25546 1878 25598
rect 1814 25210 1820 25262
rect 1872 25210 1878 25262
rect 1814 24874 1820 24926
rect 1872 24874 1878 24926
rect 1814 24538 1820 24590
rect 1872 24538 1878 24590
rect 1814 24202 1820 24254
rect 1872 24202 1878 24254
rect 1814 23866 1820 23918
rect 1872 23866 1878 23918
rect 1814 23530 1820 23582
rect 1872 23530 1878 23582
rect 1814 23194 1820 23246
rect 1872 23194 1878 23246
rect 1814 22858 1820 22910
rect 1872 22858 1878 22910
rect 1814 22522 1820 22574
rect 1872 22522 1878 22574
rect 1814 22186 1820 22238
rect 1872 22186 1878 22238
rect 1814 21850 1820 21902
rect 1872 21850 1878 21902
rect 1814 21514 1820 21566
rect 1872 21514 1878 21566
rect 1814 21178 1820 21230
rect 1872 21178 1878 21230
rect 14473 21100 14501 25659
rect 14553 21100 14581 27217
rect 14633 21100 14661 28487
rect 14713 21100 14741 30045
rect 14793 21100 14821 31315
rect 14873 21100 14901 32873
rect 14953 21100 14981 34143
rect 94172 33946 94178 33998
rect 94230 33946 94236 33998
rect 94172 33610 94178 33662
rect 94230 33610 94236 33662
rect 94172 33274 94178 33326
rect 94230 33274 94236 33326
rect 94172 32938 94178 32990
rect 94230 32938 94236 32990
rect 94172 32602 94178 32654
rect 94230 32602 94236 32654
rect 94172 32266 94178 32318
rect 94230 32266 94236 32318
rect 94172 31930 94178 31982
rect 94230 31930 94236 31982
rect 94172 31594 94178 31646
rect 94230 31594 94236 31646
rect 94172 31258 94178 31310
rect 94230 31258 94236 31310
rect 94172 30922 94178 30974
rect 94230 30922 94236 30974
rect 94172 30586 94178 30638
rect 94230 30586 94236 30638
rect 94172 30250 94178 30302
rect 94230 30250 94236 30302
rect 94172 29914 94178 29966
rect 94230 29914 94236 29966
rect 94172 29578 94178 29630
rect 94230 29578 94236 29630
rect 94172 29242 94178 29294
rect 94230 29242 94236 29294
rect 94172 28906 94178 28958
rect 94230 28906 94236 28958
rect 94172 28570 94178 28622
rect 94230 28570 94236 28622
rect 94172 28234 94178 28286
rect 94230 28234 94236 28286
rect 94172 27898 94178 27950
rect 94230 27898 94236 27950
rect 94172 27562 94178 27614
rect 94230 27562 94236 27614
rect 94172 27226 94178 27278
rect 94230 27226 94236 27278
rect 94172 26890 94178 26942
rect 94230 26890 94236 26942
rect 94172 26554 94178 26606
rect 94230 26554 94236 26606
rect 94172 26218 94178 26270
rect 94230 26218 94236 26270
rect 94172 25882 94178 25934
rect 94230 25882 94236 25934
rect 94172 25546 94178 25598
rect 94230 25546 94236 25598
rect 94172 25210 94178 25262
rect 94230 25210 94236 25262
rect 94172 24874 94178 24926
rect 94230 24874 94236 24926
rect 94172 24538 94178 24590
rect 94230 24538 94236 24590
rect 94172 24202 94178 24254
rect 94230 24202 94236 24254
rect 94172 23866 94178 23918
rect 94230 23866 94236 23918
rect 94172 23530 94178 23582
rect 94230 23530 94236 23582
rect 94172 23194 94178 23246
rect 94230 23194 94236 23246
rect 94172 22858 94178 22910
rect 94230 22858 94236 22910
rect 94172 22522 94178 22574
rect 94230 22522 94236 22574
rect 94172 22186 94178 22238
rect 94230 22186 94236 22238
rect 94172 21850 94178 21902
rect 94230 21850 94236 21902
rect 94172 21514 94178 21566
rect 94230 21514 94236 21566
rect 94172 21178 94178 21230
rect 94230 21178 94236 21230
rect 1814 20842 1820 20894
rect 1872 20842 1878 20894
rect 1814 20506 1820 20558
rect 1872 20506 1878 20558
rect 1814 20170 1820 20222
rect 1872 20170 1878 20222
rect 1814 19834 1820 19886
rect 1872 19834 1878 19886
rect 1814 19498 1820 19550
rect 1872 19498 1878 19550
rect 1814 19162 1820 19214
rect 1872 19162 1878 19214
rect 1814 18826 1820 18878
rect 1872 18826 1878 18878
rect 1814 18490 1820 18542
rect 1872 18490 1878 18542
rect 1814 18154 1820 18206
rect 1872 18154 1878 18206
rect 1814 17818 1820 17870
rect 1872 17818 1878 17870
rect 1814 17482 1820 17534
rect 1872 17482 1878 17534
rect 1814 17146 1820 17198
rect 1872 17146 1878 17198
rect 1814 16810 1820 16862
rect 1872 16810 1878 16862
rect 1814 16474 1820 16526
rect 1872 16474 1878 16526
rect 1814 16138 1820 16190
rect 1872 16138 1878 16190
rect 1814 15802 1820 15854
rect 1872 15802 1878 15854
rect 1814 15466 1820 15518
rect 1872 15466 1878 15518
rect 1814 15130 1820 15182
rect 1872 15130 1878 15182
rect 1814 14794 1820 14846
rect 1872 14794 1878 14846
rect 1814 14458 1820 14510
rect 1872 14458 1878 14510
rect 1814 14122 1820 14174
rect 1872 14122 1878 14174
rect 1814 13786 1820 13838
rect 1872 13786 1878 13838
rect 1814 13450 1820 13502
rect 1872 13450 1878 13502
rect 1814 13114 1820 13166
rect 1872 13114 1878 13166
rect 1814 12778 1820 12830
rect 1872 12778 1878 12830
rect 1814 12442 1820 12494
rect 1872 12442 1878 12494
rect 1814 12106 1820 12158
rect 1872 12106 1878 12158
rect 1814 11770 1820 11822
rect 1872 11770 1878 11822
rect 1814 11434 1820 11486
rect 1872 11434 1878 11486
rect 1814 11098 1820 11150
rect 1872 11098 1878 11150
rect 1814 10762 1820 10814
rect 1872 10762 1878 10814
rect 28206 10759 28212 10811
rect 28264 10759 28270 10811
rect 29454 10759 29460 10811
rect 29512 10759 29518 10811
rect 30702 10759 30708 10811
rect 30760 10759 30766 10811
rect 31950 10759 31956 10811
rect 32008 10759 32014 10811
rect 33198 10759 33204 10811
rect 33256 10759 33262 10811
rect 34446 10759 34452 10811
rect 34504 10759 34510 10811
rect 35694 10759 35700 10811
rect 35752 10759 35758 10811
rect 36942 10759 36948 10811
rect 37000 10759 37006 10811
rect 38190 10759 38196 10811
rect 38248 10759 38254 10811
rect 39438 10759 39444 10811
rect 39496 10759 39502 10811
rect 40686 10759 40692 10811
rect 40744 10759 40750 10811
rect 41934 10759 41940 10811
rect 41992 10759 41998 10811
rect 43182 10759 43188 10811
rect 43240 10759 43246 10811
rect 44430 10759 44436 10811
rect 44488 10759 44494 10811
rect 45678 10759 45684 10811
rect 45736 10759 45742 10811
rect 46926 10759 46932 10811
rect 46984 10759 46990 10811
rect 48174 10759 48180 10811
rect 48232 10759 48238 10811
rect 49422 10759 49428 10811
rect 49480 10759 49486 10811
rect 50670 10759 50676 10811
rect 50728 10759 50734 10811
rect 51918 10759 51924 10811
rect 51976 10759 51982 10811
rect 53166 10759 53172 10811
rect 53224 10759 53230 10811
rect 54414 10759 54420 10811
rect 54472 10759 54478 10811
rect 55662 10759 55668 10811
rect 55720 10759 55726 10811
rect 56910 10759 56916 10811
rect 56968 10759 56974 10811
rect 58158 10759 58164 10811
rect 58216 10759 58222 10811
rect 59406 10759 59412 10811
rect 59464 10759 59470 10811
rect 60654 10759 60660 10811
rect 60712 10759 60718 10811
rect 61902 10759 61908 10811
rect 61960 10759 61966 10811
rect 63150 10759 63156 10811
rect 63208 10759 63214 10811
rect 64398 10759 64404 10811
rect 64456 10759 64462 10811
rect 65646 10759 65652 10811
rect 65704 10759 65710 10811
rect 66894 10759 66900 10811
rect 66952 10759 66958 10811
rect 1814 10426 1820 10478
rect 1872 10426 1878 10478
rect 1814 10090 1820 10142
rect 1872 10090 1878 10142
rect 1814 9754 1820 9806
rect 1872 9754 1878 9806
rect 1814 9418 1820 9470
rect 1872 9418 1878 9470
rect 1814 9082 1820 9134
rect 1872 9082 1878 9134
rect 1814 8746 1820 8798
rect 1872 8746 1878 8798
rect 1814 8410 1820 8462
rect 1872 8410 1878 8462
rect 1814 8074 1820 8126
rect 1872 8074 1878 8126
rect 81177 8057 81205 21100
rect 81257 9327 81285 21100
rect 81337 10885 81365 21100
rect 81417 12155 81445 21100
rect 81497 13713 81525 21100
rect 81577 14983 81605 21100
rect 81657 16541 81685 21100
rect 94172 20842 94178 20894
rect 94230 20842 94236 20894
rect 94172 20506 94178 20558
rect 94230 20506 94236 20558
rect 94172 20170 94178 20222
rect 94230 20170 94236 20222
rect 94172 19834 94178 19886
rect 94230 19834 94236 19886
rect 94172 19498 94178 19550
rect 94230 19498 94236 19550
rect 94172 19162 94178 19214
rect 94230 19162 94236 19214
rect 94172 18826 94178 18878
rect 94230 18826 94236 18878
rect 94172 18490 94178 18542
rect 94230 18490 94236 18542
rect 94172 18154 94178 18206
rect 94230 18154 94236 18206
rect 94172 17818 94178 17870
rect 94230 17818 94236 17870
rect 94172 17482 94178 17534
rect 94230 17482 94236 17534
rect 94172 17146 94178 17198
rect 94230 17146 94236 17198
rect 94172 16810 94178 16862
rect 94230 16810 94236 16862
rect 81639 16489 81645 16541
rect 81697 16489 81703 16541
rect 94172 16474 94178 16526
rect 94230 16474 94236 16526
rect 94172 16138 94178 16190
rect 94230 16138 94236 16190
rect 94172 15802 94178 15854
rect 94230 15802 94236 15854
rect 94172 15466 94178 15518
rect 94230 15466 94236 15518
rect 94172 15130 94178 15182
rect 94230 15130 94236 15182
rect 81559 14931 81565 14983
rect 81617 14931 81623 14983
rect 94172 14794 94178 14846
rect 94230 14794 94236 14846
rect 94172 14458 94178 14510
rect 94230 14458 94236 14510
rect 94172 14122 94178 14174
rect 94230 14122 94236 14174
rect 94172 13786 94178 13838
rect 94230 13786 94236 13838
rect 81479 13661 81485 13713
rect 81537 13661 81543 13713
rect 94172 13450 94178 13502
rect 94230 13450 94236 13502
rect 94172 13114 94178 13166
rect 94230 13114 94236 13166
rect 94172 12778 94178 12830
rect 94230 12778 94236 12830
rect 94172 12442 94178 12494
rect 94230 12442 94236 12494
rect 81399 12103 81405 12155
rect 81457 12103 81463 12155
rect 94172 12106 94178 12158
rect 94230 12106 94236 12158
rect 94172 11770 94178 11822
rect 94230 11770 94236 11822
rect 94172 11434 94178 11486
rect 94230 11434 94236 11486
rect 94172 11098 94178 11150
rect 94230 11098 94236 11150
rect 81319 10833 81325 10885
rect 81377 10833 81383 10885
rect 94172 10762 94178 10814
rect 94230 10762 94236 10814
rect 94172 10426 94178 10478
rect 94230 10426 94236 10478
rect 94172 10090 94178 10142
rect 94230 10090 94236 10142
rect 94172 9754 94178 9806
rect 94230 9754 94236 9806
rect 94172 9418 94178 9470
rect 94230 9418 94236 9470
rect 81239 9275 81245 9327
rect 81297 9275 81303 9327
rect 94172 9082 94178 9134
rect 94230 9082 94236 9134
rect 94172 8746 94178 8798
rect 94230 8746 94236 8798
rect 94172 8410 94178 8462
rect 94230 8410 94236 8462
rect 94172 8074 94178 8126
rect 94230 8074 94236 8126
rect 81159 8005 81165 8057
rect 81217 8005 81223 8057
rect 1814 7738 1820 7790
rect 1872 7738 1878 7790
rect 94172 7738 94178 7790
rect 94230 7738 94236 7790
rect 1814 7402 1820 7454
rect 1872 7402 1878 7454
rect 94172 7402 94178 7454
rect 94230 7402 94236 7454
rect 1814 7066 1820 7118
rect 1872 7066 1878 7118
rect 94172 7066 94178 7118
rect 94230 7066 94236 7118
rect 1814 6730 1820 6782
rect 1872 6730 1878 6782
rect 94172 6730 94178 6782
rect 94230 6730 94236 6782
rect 1814 6394 1820 6446
rect 1872 6394 1878 6446
rect 94172 6394 94178 6446
rect 94230 6394 94236 6446
rect 1814 6058 1820 6110
rect 1872 6058 1878 6110
rect 94172 6058 94178 6110
rect 94230 6058 94236 6110
rect 1814 5722 1820 5774
rect 1872 5722 1878 5774
rect 94172 5722 94178 5774
rect 94230 5722 94236 5774
rect 1814 5386 1820 5438
rect 1872 5386 1878 5438
rect 94172 5386 94178 5438
rect 94230 5386 94236 5438
rect 1814 5050 1820 5102
rect 1872 5050 1878 5102
rect 94172 5050 94178 5102
rect 94230 5050 94236 5102
rect 1814 4714 1820 4766
rect 1872 4714 1878 4766
rect 94172 4714 94178 4766
rect 94230 4714 94236 4766
rect 1814 4378 1820 4430
rect 1872 4378 1878 4430
rect 94172 4378 94178 4430
rect 94230 4378 94236 4430
rect 1814 4042 1820 4094
rect 1872 4042 1878 4094
rect 94172 4042 94178 4094
rect 94230 4042 94236 4094
rect 1814 3706 1820 3758
rect 1872 3706 1878 3758
rect 94172 3706 94178 3758
rect 94230 3706 94236 3758
rect 1814 3370 1820 3422
rect 1872 3370 1878 3422
rect 94172 3370 94178 3422
rect 94230 3370 94236 3422
rect 1814 3034 1820 3086
rect 1872 3034 1878 3086
rect 94172 3034 94178 3086
rect 94230 3034 94236 3086
rect 1814 2698 1820 2750
rect 1872 2698 1878 2750
rect 94172 2698 94178 2750
rect 94230 2698 94236 2750
rect 1814 2362 1820 2414
rect 1872 2362 1878 2414
rect 94172 2362 94178 2414
rect 94230 2362 94236 2414
rect 1814 2026 1820 2078
rect 1872 2026 1878 2078
rect 94172 2026 94178 2078
rect 94230 2026 94236 2078
rect 1734 1742 94316 1828
rect 1734 1690 2156 1742
rect 2208 1733 3836 1742
rect 3888 1733 5516 1742
rect 5568 1733 7196 1742
rect 7248 1733 8876 1742
rect 8928 1733 10556 1742
rect 10608 1733 12236 1742
rect 12288 1733 13916 1742
rect 13968 1733 15596 1742
rect 15648 1733 17276 1742
rect 17328 1733 18956 1742
rect 19008 1733 20636 1742
rect 20688 1733 22316 1742
rect 22368 1733 23996 1742
rect 24048 1733 25676 1742
rect 25728 1733 27356 1742
rect 27408 1733 29036 1742
rect 29088 1733 30716 1742
rect 30768 1733 32396 1742
rect 32448 1733 34076 1742
rect 34128 1733 35756 1742
rect 35808 1733 37436 1742
rect 37488 1733 39116 1742
rect 39168 1733 40796 1742
rect 40848 1733 42476 1742
rect 42528 1733 44156 1742
rect 44208 1733 45836 1742
rect 45888 1733 47516 1742
rect 47568 1733 49196 1742
rect 49248 1733 50876 1742
rect 50928 1733 52556 1742
rect 52608 1733 54236 1742
rect 54288 1733 55916 1742
rect 55968 1733 57596 1742
rect 57648 1733 59276 1742
rect 59328 1733 60956 1742
rect 61008 1733 62636 1742
rect 62688 1733 64316 1742
rect 64368 1733 65996 1742
rect 66048 1733 67676 1742
rect 67728 1733 69356 1742
rect 69408 1733 71036 1742
rect 71088 1733 72716 1742
rect 72768 1733 74396 1742
rect 74448 1733 76076 1742
rect 76128 1733 77756 1742
rect 77808 1733 79436 1742
rect 79488 1733 81116 1742
rect 81168 1733 82796 1742
rect 82848 1733 84476 1742
rect 84528 1733 86156 1742
rect 86208 1733 87836 1742
rect 87888 1733 89516 1742
rect 89568 1733 91196 1742
rect 91248 1733 92876 1742
rect 92928 1733 94316 1742
rect 2208 1699 2501 1733
rect 2535 1699 2837 1733
rect 2871 1699 3173 1733
rect 3207 1699 3509 1733
rect 3543 1699 3836 1733
rect 3888 1699 4181 1733
rect 4215 1699 4517 1733
rect 4551 1699 4853 1733
rect 4887 1699 5189 1733
rect 5223 1699 5516 1733
rect 5568 1699 5861 1733
rect 5895 1699 6197 1733
rect 6231 1699 6533 1733
rect 6567 1699 6869 1733
rect 6903 1699 7196 1733
rect 7248 1699 7541 1733
rect 7575 1699 7877 1733
rect 7911 1699 8213 1733
rect 8247 1699 8549 1733
rect 8583 1699 8876 1733
rect 8928 1699 9221 1733
rect 9255 1699 9557 1733
rect 9591 1699 9893 1733
rect 9927 1699 10229 1733
rect 10263 1699 10556 1733
rect 10608 1699 10901 1733
rect 10935 1699 11237 1733
rect 11271 1699 11573 1733
rect 11607 1699 11909 1733
rect 11943 1699 12236 1733
rect 12288 1699 12581 1733
rect 12615 1699 12917 1733
rect 12951 1699 13253 1733
rect 13287 1699 13589 1733
rect 13623 1699 13916 1733
rect 13968 1699 14261 1733
rect 14295 1699 14597 1733
rect 14631 1699 14933 1733
rect 14967 1699 15269 1733
rect 15303 1699 15596 1733
rect 15648 1699 15941 1733
rect 15975 1699 16277 1733
rect 16311 1699 16613 1733
rect 16647 1699 16949 1733
rect 16983 1699 17276 1733
rect 17328 1699 17621 1733
rect 17655 1699 17957 1733
rect 17991 1699 18293 1733
rect 18327 1699 18629 1733
rect 18663 1699 18956 1733
rect 19008 1699 19301 1733
rect 19335 1699 19637 1733
rect 19671 1699 19973 1733
rect 20007 1699 20309 1733
rect 20343 1699 20636 1733
rect 20688 1699 20981 1733
rect 21015 1699 21317 1733
rect 21351 1699 21653 1733
rect 21687 1699 21989 1733
rect 22023 1699 22316 1733
rect 22368 1699 22661 1733
rect 22695 1699 22997 1733
rect 23031 1699 23333 1733
rect 23367 1699 23669 1733
rect 23703 1699 23996 1733
rect 24048 1699 24341 1733
rect 24375 1699 24677 1733
rect 24711 1699 25013 1733
rect 25047 1699 25349 1733
rect 25383 1699 25676 1733
rect 25728 1699 26021 1733
rect 26055 1699 26357 1733
rect 26391 1699 26693 1733
rect 26727 1699 27029 1733
rect 27063 1699 27356 1733
rect 27408 1699 27701 1733
rect 27735 1699 28037 1733
rect 28071 1699 28373 1733
rect 28407 1699 28709 1733
rect 28743 1699 29036 1733
rect 29088 1699 29381 1733
rect 29415 1699 29717 1733
rect 29751 1699 30053 1733
rect 30087 1699 30389 1733
rect 30423 1699 30716 1733
rect 30768 1699 31061 1733
rect 31095 1699 31397 1733
rect 31431 1699 31733 1733
rect 31767 1699 32069 1733
rect 32103 1699 32396 1733
rect 32448 1699 32741 1733
rect 32775 1699 33077 1733
rect 33111 1699 33413 1733
rect 33447 1699 33749 1733
rect 33783 1699 34076 1733
rect 34128 1699 34421 1733
rect 34455 1699 34757 1733
rect 34791 1699 35093 1733
rect 35127 1699 35429 1733
rect 35463 1699 35756 1733
rect 35808 1699 36101 1733
rect 36135 1699 36437 1733
rect 36471 1699 36773 1733
rect 36807 1699 37109 1733
rect 37143 1699 37436 1733
rect 37488 1699 37781 1733
rect 37815 1699 38117 1733
rect 38151 1699 38453 1733
rect 38487 1699 38789 1733
rect 38823 1699 39116 1733
rect 39168 1699 39461 1733
rect 39495 1699 39797 1733
rect 39831 1699 40133 1733
rect 40167 1699 40469 1733
rect 40503 1699 40796 1733
rect 40848 1699 41141 1733
rect 41175 1699 41477 1733
rect 41511 1699 41813 1733
rect 41847 1699 42149 1733
rect 42183 1699 42476 1733
rect 42528 1699 42821 1733
rect 42855 1699 43157 1733
rect 43191 1699 43493 1733
rect 43527 1699 43829 1733
rect 43863 1699 44156 1733
rect 44208 1699 44501 1733
rect 44535 1699 44837 1733
rect 44871 1699 45173 1733
rect 45207 1699 45509 1733
rect 45543 1699 45836 1733
rect 45888 1699 46181 1733
rect 46215 1699 46517 1733
rect 46551 1699 46853 1733
rect 46887 1699 47189 1733
rect 47223 1699 47516 1733
rect 47568 1699 47861 1733
rect 47895 1699 48197 1733
rect 48231 1699 48533 1733
rect 48567 1699 48869 1733
rect 48903 1699 49196 1733
rect 49248 1699 49541 1733
rect 49575 1699 49877 1733
rect 49911 1699 50213 1733
rect 50247 1699 50549 1733
rect 50583 1699 50876 1733
rect 50928 1699 51221 1733
rect 51255 1699 51557 1733
rect 51591 1699 51893 1733
rect 51927 1699 52229 1733
rect 52263 1699 52556 1733
rect 52608 1699 52901 1733
rect 52935 1699 53237 1733
rect 53271 1699 53573 1733
rect 53607 1699 53909 1733
rect 53943 1699 54236 1733
rect 54288 1699 54581 1733
rect 54615 1699 54917 1733
rect 54951 1699 55253 1733
rect 55287 1699 55589 1733
rect 55623 1699 55916 1733
rect 55968 1699 56261 1733
rect 56295 1699 56597 1733
rect 56631 1699 56933 1733
rect 56967 1699 57269 1733
rect 57303 1699 57596 1733
rect 57648 1699 57941 1733
rect 57975 1699 58277 1733
rect 58311 1699 58613 1733
rect 58647 1699 58949 1733
rect 58983 1699 59276 1733
rect 59328 1699 59621 1733
rect 59655 1699 59957 1733
rect 59991 1699 60293 1733
rect 60327 1699 60629 1733
rect 60663 1699 60956 1733
rect 61008 1699 61301 1733
rect 61335 1699 61637 1733
rect 61671 1699 61973 1733
rect 62007 1699 62309 1733
rect 62343 1699 62636 1733
rect 62688 1699 62981 1733
rect 63015 1699 63317 1733
rect 63351 1699 63653 1733
rect 63687 1699 63989 1733
rect 64023 1699 64316 1733
rect 64368 1699 64661 1733
rect 64695 1699 64997 1733
rect 65031 1699 65333 1733
rect 65367 1699 65669 1733
rect 65703 1699 65996 1733
rect 66048 1699 66341 1733
rect 66375 1699 66677 1733
rect 66711 1699 67013 1733
rect 67047 1699 67349 1733
rect 67383 1699 67676 1733
rect 67728 1699 68021 1733
rect 68055 1699 68357 1733
rect 68391 1699 68693 1733
rect 68727 1699 69029 1733
rect 69063 1699 69356 1733
rect 69408 1699 69701 1733
rect 69735 1699 70037 1733
rect 70071 1699 70373 1733
rect 70407 1699 70709 1733
rect 70743 1699 71036 1733
rect 71088 1699 71381 1733
rect 71415 1699 71717 1733
rect 71751 1699 72053 1733
rect 72087 1699 72389 1733
rect 72423 1699 72716 1733
rect 72768 1699 73061 1733
rect 73095 1699 73397 1733
rect 73431 1699 73733 1733
rect 73767 1699 74069 1733
rect 74103 1699 74396 1733
rect 74448 1699 74741 1733
rect 74775 1699 75077 1733
rect 75111 1699 75413 1733
rect 75447 1699 75749 1733
rect 75783 1699 76076 1733
rect 76128 1699 76421 1733
rect 76455 1699 76757 1733
rect 76791 1699 77093 1733
rect 77127 1699 77429 1733
rect 77463 1699 77756 1733
rect 77808 1699 78101 1733
rect 78135 1699 78437 1733
rect 78471 1699 78773 1733
rect 78807 1699 79109 1733
rect 79143 1699 79436 1733
rect 79488 1699 79781 1733
rect 79815 1699 80117 1733
rect 80151 1699 80453 1733
rect 80487 1699 80789 1733
rect 80823 1699 81116 1733
rect 81168 1699 81461 1733
rect 81495 1699 81797 1733
rect 81831 1699 82133 1733
rect 82167 1699 82469 1733
rect 82503 1699 82796 1733
rect 82848 1699 83141 1733
rect 83175 1699 83477 1733
rect 83511 1699 83813 1733
rect 83847 1699 84149 1733
rect 84183 1699 84476 1733
rect 84528 1699 84821 1733
rect 84855 1699 85157 1733
rect 85191 1699 85493 1733
rect 85527 1699 85829 1733
rect 85863 1699 86156 1733
rect 86208 1699 86501 1733
rect 86535 1699 86837 1733
rect 86871 1699 87173 1733
rect 87207 1699 87509 1733
rect 87543 1699 87836 1733
rect 87888 1699 88181 1733
rect 88215 1699 88517 1733
rect 88551 1699 88853 1733
rect 88887 1699 89189 1733
rect 89223 1699 89516 1733
rect 89568 1699 89861 1733
rect 89895 1699 90197 1733
rect 90231 1699 90533 1733
rect 90567 1699 90869 1733
rect 90903 1699 91196 1733
rect 91248 1699 91541 1733
rect 91575 1699 91877 1733
rect 91911 1699 92213 1733
rect 92247 1699 92549 1733
rect 92583 1699 92876 1733
rect 92928 1699 93221 1733
rect 93255 1699 93557 1733
rect 93591 1699 94316 1733
rect 2208 1690 3836 1699
rect 3888 1690 5516 1699
rect 5568 1690 7196 1699
rect 7248 1690 8876 1699
rect 8928 1690 10556 1699
rect 10608 1690 12236 1699
rect 12288 1690 13916 1699
rect 13968 1690 15596 1699
rect 15648 1690 17276 1699
rect 17328 1690 18956 1699
rect 19008 1690 20636 1699
rect 20688 1690 22316 1699
rect 22368 1690 23996 1699
rect 24048 1690 25676 1699
rect 25728 1690 27356 1699
rect 27408 1690 29036 1699
rect 29088 1690 30716 1699
rect 30768 1690 32396 1699
rect 32448 1690 34076 1699
rect 34128 1690 35756 1699
rect 35808 1690 37436 1699
rect 37488 1690 39116 1699
rect 39168 1690 40796 1699
rect 40848 1690 42476 1699
rect 42528 1690 44156 1699
rect 44208 1690 45836 1699
rect 45888 1690 47516 1699
rect 47568 1690 49196 1699
rect 49248 1690 50876 1699
rect 50928 1690 52556 1699
rect 52608 1690 54236 1699
rect 54288 1690 55916 1699
rect 55968 1690 57596 1699
rect 57648 1690 59276 1699
rect 59328 1690 60956 1699
rect 61008 1690 62636 1699
rect 62688 1690 64316 1699
rect 64368 1690 65996 1699
rect 66048 1690 67676 1699
rect 67728 1690 69356 1699
rect 69408 1690 71036 1699
rect 71088 1690 72716 1699
rect 72768 1690 74396 1699
rect 74448 1690 76076 1699
rect 76128 1690 77756 1699
rect 77808 1690 79436 1699
rect 79488 1690 81116 1699
rect 81168 1690 82796 1699
rect 82848 1690 84476 1699
rect 84528 1690 86156 1699
rect 86208 1690 87836 1699
rect 87888 1690 89516 1699
rect 89568 1690 91196 1699
rect 91248 1690 92876 1699
rect 92928 1690 94316 1699
rect 1734 1604 94316 1690
<< via1 >>
rect 2156 77797 2208 77806
rect 3836 77797 3888 77806
rect 5516 77797 5568 77806
rect 7196 77797 7248 77806
rect 8876 77797 8928 77806
rect 10556 77797 10608 77806
rect 12236 77797 12288 77806
rect 13916 77797 13968 77806
rect 15596 77797 15648 77806
rect 17276 77797 17328 77806
rect 18956 77797 19008 77806
rect 20636 77797 20688 77806
rect 22316 77797 22368 77806
rect 23996 77797 24048 77806
rect 25676 77797 25728 77806
rect 27356 77797 27408 77806
rect 29036 77797 29088 77806
rect 30716 77797 30768 77806
rect 32396 77797 32448 77806
rect 34076 77797 34128 77806
rect 35756 77797 35808 77806
rect 37436 77797 37488 77806
rect 39116 77797 39168 77806
rect 40796 77797 40848 77806
rect 42476 77797 42528 77806
rect 44156 77797 44208 77806
rect 45836 77797 45888 77806
rect 47516 77797 47568 77806
rect 49196 77797 49248 77806
rect 50876 77797 50928 77806
rect 52556 77797 52608 77806
rect 54236 77797 54288 77806
rect 55916 77797 55968 77806
rect 57596 77797 57648 77806
rect 59276 77797 59328 77806
rect 60956 77797 61008 77806
rect 62636 77797 62688 77806
rect 64316 77797 64368 77806
rect 65996 77797 66048 77806
rect 67676 77797 67728 77806
rect 69356 77797 69408 77806
rect 71036 77797 71088 77806
rect 72716 77797 72768 77806
rect 74396 77797 74448 77806
rect 76076 77797 76128 77806
rect 77756 77797 77808 77806
rect 79436 77797 79488 77806
rect 81116 77797 81168 77806
rect 82796 77797 82848 77806
rect 84476 77797 84528 77806
rect 86156 77797 86208 77806
rect 87836 77797 87888 77806
rect 89516 77797 89568 77806
rect 91196 77797 91248 77806
rect 92876 77797 92928 77806
rect 2156 77763 2165 77797
rect 2165 77763 2199 77797
rect 2199 77763 2208 77797
rect 3836 77763 3845 77797
rect 3845 77763 3879 77797
rect 3879 77763 3888 77797
rect 5516 77763 5525 77797
rect 5525 77763 5559 77797
rect 5559 77763 5568 77797
rect 7196 77763 7205 77797
rect 7205 77763 7239 77797
rect 7239 77763 7248 77797
rect 8876 77763 8885 77797
rect 8885 77763 8919 77797
rect 8919 77763 8928 77797
rect 10556 77763 10565 77797
rect 10565 77763 10599 77797
rect 10599 77763 10608 77797
rect 12236 77763 12245 77797
rect 12245 77763 12279 77797
rect 12279 77763 12288 77797
rect 13916 77763 13925 77797
rect 13925 77763 13959 77797
rect 13959 77763 13968 77797
rect 15596 77763 15605 77797
rect 15605 77763 15639 77797
rect 15639 77763 15648 77797
rect 17276 77763 17285 77797
rect 17285 77763 17319 77797
rect 17319 77763 17328 77797
rect 18956 77763 18965 77797
rect 18965 77763 18999 77797
rect 18999 77763 19008 77797
rect 20636 77763 20645 77797
rect 20645 77763 20679 77797
rect 20679 77763 20688 77797
rect 22316 77763 22325 77797
rect 22325 77763 22359 77797
rect 22359 77763 22368 77797
rect 23996 77763 24005 77797
rect 24005 77763 24039 77797
rect 24039 77763 24048 77797
rect 25676 77763 25685 77797
rect 25685 77763 25719 77797
rect 25719 77763 25728 77797
rect 27356 77763 27365 77797
rect 27365 77763 27399 77797
rect 27399 77763 27408 77797
rect 29036 77763 29045 77797
rect 29045 77763 29079 77797
rect 29079 77763 29088 77797
rect 30716 77763 30725 77797
rect 30725 77763 30759 77797
rect 30759 77763 30768 77797
rect 32396 77763 32405 77797
rect 32405 77763 32439 77797
rect 32439 77763 32448 77797
rect 34076 77763 34085 77797
rect 34085 77763 34119 77797
rect 34119 77763 34128 77797
rect 35756 77763 35765 77797
rect 35765 77763 35799 77797
rect 35799 77763 35808 77797
rect 37436 77763 37445 77797
rect 37445 77763 37479 77797
rect 37479 77763 37488 77797
rect 39116 77763 39125 77797
rect 39125 77763 39159 77797
rect 39159 77763 39168 77797
rect 40796 77763 40805 77797
rect 40805 77763 40839 77797
rect 40839 77763 40848 77797
rect 42476 77763 42485 77797
rect 42485 77763 42519 77797
rect 42519 77763 42528 77797
rect 44156 77763 44165 77797
rect 44165 77763 44199 77797
rect 44199 77763 44208 77797
rect 45836 77763 45845 77797
rect 45845 77763 45879 77797
rect 45879 77763 45888 77797
rect 47516 77763 47525 77797
rect 47525 77763 47559 77797
rect 47559 77763 47568 77797
rect 49196 77763 49205 77797
rect 49205 77763 49239 77797
rect 49239 77763 49248 77797
rect 50876 77763 50885 77797
rect 50885 77763 50919 77797
rect 50919 77763 50928 77797
rect 52556 77763 52565 77797
rect 52565 77763 52599 77797
rect 52599 77763 52608 77797
rect 54236 77763 54245 77797
rect 54245 77763 54279 77797
rect 54279 77763 54288 77797
rect 55916 77763 55925 77797
rect 55925 77763 55959 77797
rect 55959 77763 55968 77797
rect 57596 77763 57605 77797
rect 57605 77763 57639 77797
rect 57639 77763 57648 77797
rect 59276 77763 59285 77797
rect 59285 77763 59319 77797
rect 59319 77763 59328 77797
rect 60956 77763 60965 77797
rect 60965 77763 60999 77797
rect 60999 77763 61008 77797
rect 62636 77763 62645 77797
rect 62645 77763 62679 77797
rect 62679 77763 62688 77797
rect 64316 77763 64325 77797
rect 64325 77763 64359 77797
rect 64359 77763 64368 77797
rect 65996 77763 66005 77797
rect 66005 77763 66039 77797
rect 66039 77763 66048 77797
rect 67676 77763 67685 77797
rect 67685 77763 67719 77797
rect 67719 77763 67728 77797
rect 69356 77763 69365 77797
rect 69365 77763 69399 77797
rect 69399 77763 69408 77797
rect 71036 77763 71045 77797
rect 71045 77763 71079 77797
rect 71079 77763 71088 77797
rect 72716 77763 72725 77797
rect 72725 77763 72759 77797
rect 72759 77763 72768 77797
rect 74396 77763 74405 77797
rect 74405 77763 74439 77797
rect 74439 77763 74448 77797
rect 76076 77763 76085 77797
rect 76085 77763 76119 77797
rect 76119 77763 76128 77797
rect 77756 77763 77765 77797
rect 77765 77763 77799 77797
rect 77799 77763 77808 77797
rect 79436 77763 79445 77797
rect 79445 77763 79479 77797
rect 79479 77763 79488 77797
rect 81116 77763 81125 77797
rect 81125 77763 81159 77797
rect 81159 77763 81168 77797
rect 82796 77763 82805 77797
rect 82805 77763 82839 77797
rect 82839 77763 82848 77797
rect 84476 77763 84485 77797
rect 84485 77763 84519 77797
rect 84519 77763 84528 77797
rect 86156 77763 86165 77797
rect 86165 77763 86199 77797
rect 86199 77763 86208 77797
rect 87836 77763 87845 77797
rect 87845 77763 87879 77797
rect 87879 77763 87888 77797
rect 89516 77763 89525 77797
rect 89525 77763 89559 77797
rect 89559 77763 89568 77797
rect 91196 77763 91205 77797
rect 91205 77763 91239 77797
rect 91239 77763 91248 77797
rect 92876 77763 92885 77797
rect 92885 77763 92919 77797
rect 92919 77763 92928 77797
rect 2156 77754 2208 77763
rect 3836 77754 3888 77763
rect 5516 77754 5568 77763
rect 7196 77754 7248 77763
rect 8876 77754 8928 77763
rect 10556 77754 10608 77763
rect 12236 77754 12288 77763
rect 13916 77754 13968 77763
rect 15596 77754 15648 77763
rect 17276 77754 17328 77763
rect 18956 77754 19008 77763
rect 20636 77754 20688 77763
rect 22316 77754 22368 77763
rect 23996 77754 24048 77763
rect 25676 77754 25728 77763
rect 27356 77754 27408 77763
rect 29036 77754 29088 77763
rect 30716 77754 30768 77763
rect 32396 77754 32448 77763
rect 34076 77754 34128 77763
rect 35756 77754 35808 77763
rect 37436 77754 37488 77763
rect 39116 77754 39168 77763
rect 40796 77754 40848 77763
rect 42476 77754 42528 77763
rect 44156 77754 44208 77763
rect 45836 77754 45888 77763
rect 47516 77754 47568 77763
rect 49196 77754 49248 77763
rect 50876 77754 50928 77763
rect 52556 77754 52608 77763
rect 54236 77754 54288 77763
rect 55916 77754 55968 77763
rect 57596 77754 57648 77763
rect 59276 77754 59328 77763
rect 60956 77754 61008 77763
rect 62636 77754 62688 77763
rect 64316 77754 64368 77763
rect 65996 77754 66048 77763
rect 67676 77754 67728 77763
rect 69356 77754 69408 77763
rect 71036 77754 71088 77763
rect 72716 77754 72768 77763
rect 74396 77754 74448 77763
rect 76076 77754 76128 77763
rect 77756 77754 77808 77763
rect 79436 77754 79488 77763
rect 81116 77754 81168 77763
rect 82796 77754 82848 77763
rect 84476 77754 84528 77763
rect 86156 77754 86208 77763
rect 87836 77754 87888 77763
rect 89516 77754 89568 77763
rect 91196 77754 91248 77763
rect 92876 77754 92928 77763
rect 1820 77333 1872 77342
rect 1820 77299 1829 77333
rect 1829 77299 1863 77333
rect 1863 77299 1872 77333
rect 1820 77290 1872 77299
rect 94178 77333 94230 77342
rect 94178 77299 94187 77333
rect 94187 77299 94221 77333
rect 94221 77299 94230 77333
rect 94178 77290 94230 77299
rect 1820 76997 1872 77006
rect 1820 76963 1829 76997
rect 1829 76963 1863 76997
rect 1863 76963 1872 76997
rect 1820 76954 1872 76963
rect 94178 76997 94230 77006
rect 94178 76963 94187 76997
rect 94187 76963 94221 76997
rect 94221 76963 94230 76997
rect 94178 76954 94230 76963
rect 1820 76661 1872 76670
rect 1820 76627 1829 76661
rect 1829 76627 1863 76661
rect 1863 76627 1872 76661
rect 1820 76618 1872 76627
rect 94178 76661 94230 76670
rect 94178 76627 94187 76661
rect 94187 76627 94221 76661
rect 94221 76627 94230 76661
rect 94178 76618 94230 76627
rect 1820 76325 1872 76334
rect 1820 76291 1829 76325
rect 1829 76291 1863 76325
rect 1863 76291 1872 76325
rect 1820 76282 1872 76291
rect 94178 76325 94230 76334
rect 94178 76291 94187 76325
rect 94187 76291 94221 76325
rect 94221 76291 94230 76325
rect 94178 76282 94230 76291
rect 1820 75989 1872 75998
rect 1820 75955 1829 75989
rect 1829 75955 1863 75989
rect 1863 75955 1872 75989
rect 1820 75946 1872 75955
rect 94178 75989 94230 75998
rect 94178 75955 94187 75989
rect 94187 75955 94221 75989
rect 94221 75955 94230 75989
rect 94178 75946 94230 75955
rect 1820 75653 1872 75662
rect 1820 75619 1829 75653
rect 1829 75619 1863 75653
rect 1863 75619 1872 75653
rect 1820 75610 1872 75619
rect 94178 75653 94230 75662
rect 94178 75619 94187 75653
rect 94187 75619 94221 75653
rect 94221 75619 94230 75653
rect 94178 75610 94230 75619
rect 1820 75317 1872 75326
rect 1820 75283 1829 75317
rect 1829 75283 1863 75317
rect 1863 75283 1872 75317
rect 1820 75274 1872 75283
rect 94178 75317 94230 75326
rect 94178 75283 94187 75317
rect 94187 75283 94221 75317
rect 94221 75283 94230 75317
rect 94178 75274 94230 75283
rect 1820 74981 1872 74990
rect 1820 74947 1829 74981
rect 1829 74947 1863 74981
rect 1863 74947 1872 74981
rect 1820 74938 1872 74947
rect 94178 74981 94230 74990
rect 94178 74947 94187 74981
rect 94187 74947 94221 74981
rect 94221 74947 94230 74981
rect 94178 74938 94230 74947
rect 1820 74645 1872 74654
rect 1820 74611 1829 74645
rect 1829 74611 1863 74645
rect 1863 74611 1872 74645
rect 1820 74602 1872 74611
rect 94178 74645 94230 74654
rect 94178 74611 94187 74645
rect 94187 74611 94221 74645
rect 94221 74611 94230 74645
rect 94178 74602 94230 74611
rect 1820 74309 1872 74318
rect 1820 74275 1829 74309
rect 1829 74275 1863 74309
rect 1863 74275 1872 74309
rect 1820 74266 1872 74275
rect 94178 74309 94230 74318
rect 94178 74275 94187 74309
rect 94187 74275 94221 74309
rect 94221 74275 94230 74309
rect 94178 74266 94230 74275
rect 28212 74049 28264 74101
rect 29460 74049 29512 74101
rect 30708 74049 30760 74101
rect 31956 74049 32008 74101
rect 33204 74049 33256 74101
rect 34452 74049 34504 74101
rect 35700 74049 35752 74101
rect 36948 74049 37000 74101
rect 38196 74049 38248 74101
rect 39444 74049 39496 74101
rect 40692 74049 40744 74101
rect 41940 74049 41992 74101
rect 43188 74049 43240 74101
rect 44436 74049 44488 74101
rect 45684 74049 45736 74101
rect 46932 74049 46984 74101
rect 48180 74049 48232 74101
rect 49428 74049 49480 74101
rect 50676 74049 50728 74101
rect 51924 74049 51976 74101
rect 53172 74049 53224 74101
rect 54420 74049 54472 74101
rect 55668 74049 55720 74101
rect 56916 74049 56968 74101
rect 58164 74049 58216 74101
rect 59412 74049 59464 74101
rect 60660 74049 60712 74101
rect 61908 74049 61960 74101
rect 63156 74049 63208 74101
rect 64404 74049 64456 74101
rect 65652 74049 65704 74101
rect 66900 74049 66952 74101
rect 1820 73973 1872 73982
rect 1820 73939 1829 73973
rect 1829 73939 1863 73973
rect 1863 73939 1872 73973
rect 1820 73930 1872 73939
rect 94178 73973 94230 73982
rect 94178 73939 94187 73973
rect 94187 73939 94221 73973
rect 94221 73939 94230 73973
rect 94178 73930 94230 73939
rect 1820 73637 1872 73646
rect 1820 73603 1829 73637
rect 1829 73603 1863 73637
rect 1863 73603 1872 73637
rect 1820 73594 1872 73603
rect 94178 73637 94230 73646
rect 94178 73603 94187 73637
rect 94187 73603 94221 73637
rect 94221 73603 94230 73637
rect 94178 73594 94230 73603
rect 1820 73301 1872 73310
rect 1820 73267 1829 73301
rect 1829 73267 1863 73301
rect 1863 73267 1872 73301
rect 1820 73258 1872 73267
rect 94178 73301 94230 73310
rect 94178 73267 94187 73301
rect 94187 73267 94221 73301
rect 94221 73267 94230 73301
rect 94178 73258 94230 73267
rect 1820 72965 1872 72974
rect 1820 72931 1829 72965
rect 1829 72931 1863 72965
rect 1863 72931 1872 72965
rect 1820 72922 1872 72931
rect 94178 72965 94230 72974
rect 94178 72931 94187 72965
rect 94187 72931 94221 72965
rect 94221 72931 94230 72965
rect 94178 72922 94230 72931
rect 1820 72629 1872 72638
rect 1820 72595 1829 72629
rect 1829 72595 1863 72629
rect 1863 72595 1872 72629
rect 1820 72586 1872 72595
rect 94178 72629 94230 72638
rect 94178 72595 94187 72629
rect 94187 72595 94221 72629
rect 94221 72595 94230 72629
rect 94178 72586 94230 72595
rect 1820 72293 1872 72302
rect 1820 72259 1829 72293
rect 1829 72259 1863 72293
rect 1863 72259 1872 72293
rect 1820 72250 1872 72259
rect 94178 72293 94230 72302
rect 94178 72259 94187 72293
rect 94187 72259 94221 72293
rect 94221 72259 94230 72293
rect 94178 72250 94230 72259
rect 1820 71957 1872 71966
rect 1820 71923 1829 71957
rect 1829 71923 1863 71957
rect 1863 71923 1872 71957
rect 1820 71914 1872 71923
rect 94178 71957 94230 71966
rect 94178 71923 94187 71957
rect 94187 71923 94221 71957
rect 94221 71923 94230 71957
rect 94178 71914 94230 71923
rect 1820 71621 1872 71630
rect 1820 71587 1829 71621
rect 1829 71587 1863 71621
rect 1863 71587 1872 71621
rect 1820 71578 1872 71587
rect 94178 71621 94230 71630
rect 94178 71587 94187 71621
rect 94187 71587 94221 71621
rect 94221 71587 94230 71621
rect 94178 71578 94230 71587
rect 1820 71285 1872 71294
rect 1820 71251 1829 71285
rect 1829 71251 1863 71285
rect 1863 71251 1872 71285
rect 1820 71242 1872 71251
rect 94178 71285 94230 71294
rect 94178 71251 94187 71285
rect 94187 71251 94221 71285
rect 94221 71251 94230 71285
rect 94178 71242 94230 71251
rect 1820 70949 1872 70958
rect 1820 70915 1829 70949
rect 1829 70915 1863 70949
rect 1863 70915 1872 70949
rect 1820 70906 1872 70915
rect 94178 70949 94230 70958
rect 94178 70915 94187 70949
rect 94187 70915 94221 70949
rect 94221 70915 94230 70949
rect 94178 70906 94230 70915
rect 1820 70613 1872 70622
rect 1820 70579 1829 70613
rect 1829 70579 1863 70613
rect 1863 70579 1872 70613
rect 1820 70570 1872 70579
rect 94178 70613 94230 70622
rect 94178 70579 94187 70613
rect 94187 70579 94221 70613
rect 94221 70579 94230 70613
rect 94178 70570 94230 70579
rect 1820 70277 1872 70286
rect 1820 70243 1829 70277
rect 1829 70243 1863 70277
rect 1863 70243 1872 70277
rect 1820 70234 1872 70243
rect 94178 70277 94230 70286
rect 94178 70243 94187 70277
rect 94187 70243 94221 70277
rect 94221 70243 94230 70277
rect 94178 70234 94230 70243
rect 1820 69941 1872 69950
rect 1820 69907 1829 69941
rect 1829 69907 1863 69941
rect 1863 69907 1872 69941
rect 1820 69898 1872 69907
rect 94178 69941 94230 69950
rect 94178 69907 94187 69941
rect 94187 69907 94221 69941
rect 94221 69907 94230 69941
rect 94178 69898 94230 69907
rect 1820 69605 1872 69614
rect 1820 69571 1829 69605
rect 1829 69571 1863 69605
rect 1863 69571 1872 69605
rect 1820 69562 1872 69571
rect 94178 69605 94230 69614
rect 94178 69571 94187 69605
rect 94187 69571 94221 69605
rect 94221 69571 94230 69605
rect 94178 69562 94230 69571
rect 1820 69269 1872 69278
rect 1820 69235 1829 69269
rect 1829 69235 1863 69269
rect 1863 69235 1872 69269
rect 1820 69226 1872 69235
rect 94178 69269 94230 69278
rect 94178 69235 94187 69269
rect 94187 69235 94221 69269
rect 94221 69235 94230 69269
rect 94178 69226 94230 69235
rect 1820 68933 1872 68942
rect 1820 68899 1829 68933
rect 1829 68899 1863 68933
rect 1863 68899 1872 68933
rect 1820 68890 1872 68899
rect 94178 68933 94230 68942
rect 94178 68899 94187 68933
rect 94187 68899 94221 68933
rect 94221 68899 94230 68933
rect 94178 68890 94230 68899
rect 1820 68597 1872 68606
rect 1820 68563 1829 68597
rect 1829 68563 1863 68597
rect 1863 68563 1872 68597
rect 1820 68554 1872 68563
rect 94178 68597 94230 68606
rect 94178 68563 94187 68597
rect 94187 68563 94221 68597
rect 94221 68563 94230 68597
rect 94178 68554 94230 68563
rect 1820 68261 1872 68270
rect 1820 68227 1829 68261
rect 1829 68227 1863 68261
rect 1863 68227 1872 68261
rect 1820 68218 1872 68227
rect 94178 68261 94230 68270
rect 94178 68227 94187 68261
rect 94187 68227 94221 68261
rect 94221 68227 94230 68261
rect 94178 68218 94230 68227
rect 1820 67925 1872 67934
rect 1820 67891 1829 67925
rect 1829 67891 1863 67925
rect 1863 67891 1872 67925
rect 1820 67882 1872 67891
rect 94178 67925 94230 67934
rect 94178 67891 94187 67925
rect 94187 67891 94221 67925
rect 94221 67891 94230 67925
rect 94178 67882 94230 67891
rect 1820 67589 1872 67598
rect 1820 67555 1829 67589
rect 1829 67555 1863 67589
rect 1863 67555 1872 67589
rect 1820 67546 1872 67555
rect 94178 67589 94230 67598
rect 94178 67555 94187 67589
rect 94187 67555 94221 67589
rect 94221 67555 94230 67589
rect 94178 67546 94230 67555
rect 1820 67253 1872 67262
rect 1820 67219 1829 67253
rect 1829 67219 1863 67253
rect 1863 67219 1872 67253
rect 1820 67210 1872 67219
rect 94178 67253 94230 67262
rect 94178 67219 94187 67253
rect 94187 67219 94221 67253
rect 94221 67219 94230 67253
rect 94178 67210 94230 67219
rect 1820 66917 1872 66926
rect 1820 66883 1829 66917
rect 1829 66883 1863 66917
rect 1863 66883 1872 66917
rect 1820 66874 1872 66883
rect 94178 66917 94230 66926
rect 94178 66883 94187 66917
rect 94187 66883 94221 66917
rect 94221 66883 94230 66917
rect 94178 66874 94230 66883
rect 1820 66581 1872 66590
rect 1820 66547 1829 66581
rect 1829 66547 1863 66581
rect 1863 66547 1872 66581
rect 1820 66538 1872 66547
rect 94178 66581 94230 66590
rect 94178 66547 94187 66581
rect 94187 66547 94221 66581
rect 94221 66547 94230 66581
rect 94178 66538 94230 66547
rect 1820 66245 1872 66254
rect 1820 66211 1829 66245
rect 1829 66211 1863 66245
rect 1863 66211 1872 66245
rect 1820 66202 1872 66211
rect 94178 66245 94230 66254
rect 94178 66211 94187 66245
rect 94187 66211 94221 66245
rect 94221 66211 94230 66245
rect 94178 66202 94230 66211
rect 1820 65909 1872 65918
rect 1820 65875 1829 65909
rect 1829 65875 1863 65909
rect 1863 65875 1872 65909
rect 1820 65866 1872 65875
rect 94178 65909 94230 65918
rect 94178 65875 94187 65909
rect 94187 65875 94221 65909
rect 94221 65875 94230 65909
rect 94178 65866 94230 65875
rect 1820 65573 1872 65582
rect 1820 65539 1829 65573
rect 1829 65539 1863 65573
rect 1863 65539 1872 65573
rect 1820 65530 1872 65539
rect 94178 65573 94230 65582
rect 94178 65539 94187 65573
rect 94187 65539 94221 65573
rect 94221 65539 94230 65573
rect 94178 65530 94230 65539
rect 1820 65237 1872 65246
rect 1820 65203 1829 65237
rect 1829 65203 1863 65237
rect 1863 65203 1872 65237
rect 1820 65194 1872 65203
rect 94178 65237 94230 65246
rect 94178 65203 94187 65237
rect 94187 65203 94221 65237
rect 94221 65203 94230 65237
rect 94178 65194 94230 65203
rect 1820 64901 1872 64910
rect 1820 64867 1829 64901
rect 1829 64867 1863 64901
rect 1863 64867 1872 64901
rect 1820 64858 1872 64867
rect 94178 64901 94230 64910
rect 94178 64867 94187 64901
rect 94187 64867 94221 64901
rect 94221 64867 94230 64901
rect 94178 64858 94230 64867
rect 1820 64565 1872 64574
rect 1820 64531 1829 64565
rect 1829 64531 1863 64565
rect 1863 64531 1872 64565
rect 1820 64522 1872 64531
rect 94178 64565 94230 64574
rect 94178 64531 94187 64565
rect 94187 64531 94221 64565
rect 94221 64531 94230 64565
rect 94178 64522 94230 64531
rect 1820 64229 1872 64238
rect 1820 64195 1829 64229
rect 1829 64195 1863 64229
rect 1863 64195 1872 64229
rect 1820 64186 1872 64195
rect 94178 64229 94230 64238
rect 94178 64195 94187 64229
rect 94187 64195 94221 64229
rect 94221 64195 94230 64229
rect 94178 64186 94230 64195
rect 1820 63893 1872 63902
rect 1820 63859 1829 63893
rect 1829 63859 1863 63893
rect 1863 63859 1872 63893
rect 1820 63850 1872 63859
rect 94178 63893 94230 63902
rect 94178 63859 94187 63893
rect 94187 63859 94221 63893
rect 94221 63859 94230 63893
rect 94178 63850 94230 63859
rect 1820 63557 1872 63566
rect 1820 63523 1829 63557
rect 1829 63523 1863 63557
rect 1863 63523 1872 63557
rect 1820 63514 1872 63523
rect 94178 63557 94230 63566
rect 94178 63523 94187 63557
rect 94187 63523 94221 63557
rect 94221 63523 94230 63557
rect 94178 63514 94230 63523
rect 1820 63221 1872 63230
rect 1820 63187 1829 63221
rect 1829 63187 1863 63221
rect 1863 63187 1872 63221
rect 1820 63178 1872 63187
rect 94178 63221 94230 63230
rect 94178 63187 94187 63221
rect 94187 63187 94221 63221
rect 94221 63187 94230 63221
rect 94178 63178 94230 63187
rect 1820 62885 1872 62894
rect 1820 62851 1829 62885
rect 1829 62851 1863 62885
rect 1863 62851 1872 62885
rect 1820 62842 1872 62851
rect 94178 62885 94230 62894
rect 94178 62851 94187 62885
rect 94187 62851 94221 62885
rect 94221 62851 94230 62885
rect 94178 62842 94230 62851
rect 1820 62549 1872 62558
rect 1820 62515 1829 62549
rect 1829 62515 1863 62549
rect 1863 62515 1872 62549
rect 1820 62506 1872 62515
rect 94178 62549 94230 62558
rect 94178 62515 94187 62549
rect 94187 62515 94221 62549
rect 94221 62515 94230 62549
rect 94178 62506 94230 62515
rect 1820 62213 1872 62222
rect 1820 62179 1829 62213
rect 1829 62179 1863 62213
rect 1863 62179 1872 62213
rect 1820 62170 1872 62179
rect 94178 62213 94230 62222
rect 94178 62179 94187 62213
rect 94187 62179 94221 62213
rect 94221 62179 94230 62213
rect 94178 62170 94230 62179
rect 1820 61877 1872 61886
rect 1820 61843 1829 61877
rect 1829 61843 1863 61877
rect 1863 61843 1872 61877
rect 1820 61834 1872 61843
rect 94178 61877 94230 61886
rect 94178 61843 94187 61877
rect 94187 61843 94221 61877
rect 94221 61843 94230 61877
rect 94178 61834 94230 61843
rect 1820 61541 1872 61550
rect 1820 61507 1829 61541
rect 1829 61507 1863 61541
rect 1863 61507 1872 61541
rect 1820 61498 1872 61507
rect 94178 61541 94230 61550
rect 94178 61507 94187 61541
rect 94187 61507 94221 61541
rect 94221 61507 94230 61541
rect 94178 61498 94230 61507
rect 1820 61205 1872 61214
rect 1820 61171 1829 61205
rect 1829 61171 1863 61205
rect 1863 61171 1872 61205
rect 1820 61162 1872 61171
rect 94178 61205 94230 61214
rect 94178 61171 94187 61205
rect 94187 61171 94221 61205
rect 94221 61171 94230 61205
rect 94178 61162 94230 61171
rect 1820 60869 1872 60878
rect 1820 60835 1829 60869
rect 1829 60835 1863 60869
rect 1863 60835 1872 60869
rect 1820 60826 1872 60835
rect 94178 60869 94230 60878
rect 94178 60835 94187 60869
rect 94187 60835 94221 60869
rect 94221 60835 94230 60869
rect 94178 60826 94230 60835
rect 1820 60533 1872 60542
rect 1820 60499 1829 60533
rect 1829 60499 1863 60533
rect 1863 60499 1872 60533
rect 1820 60490 1872 60499
rect 94178 60533 94230 60542
rect 94178 60499 94187 60533
rect 94187 60499 94221 60533
rect 94221 60499 94230 60533
rect 94178 60490 94230 60499
rect 1820 60197 1872 60206
rect 1820 60163 1829 60197
rect 1829 60163 1863 60197
rect 1863 60163 1872 60197
rect 1820 60154 1872 60163
rect 94178 60197 94230 60206
rect 94178 60163 94187 60197
rect 94187 60163 94221 60197
rect 94221 60163 94230 60197
rect 94178 60154 94230 60163
rect 1820 59861 1872 59870
rect 1820 59827 1829 59861
rect 1829 59827 1863 59861
rect 1863 59827 1872 59861
rect 1820 59818 1872 59827
rect 94178 59861 94230 59870
rect 94178 59827 94187 59861
rect 94187 59827 94221 59861
rect 94221 59827 94230 59861
rect 94178 59818 94230 59827
rect 1820 59525 1872 59534
rect 1820 59491 1829 59525
rect 1829 59491 1863 59525
rect 1863 59491 1872 59525
rect 1820 59482 1872 59491
rect 94178 59525 94230 59534
rect 94178 59491 94187 59525
rect 94187 59491 94221 59525
rect 94221 59491 94230 59525
rect 94178 59482 94230 59491
rect 1820 59189 1872 59198
rect 1820 59155 1829 59189
rect 1829 59155 1863 59189
rect 1863 59155 1872 59189
rect 1820 59146 1872 59155
rect 94178 59189 94230 59198
rect 94178 59155 94187 59189
rect 94187 59155 94221 59189
rect 94221 59155 94230 59189
rect 94178 59146 94230 59155
rect 1820 58853 1872 58862
rect 1820 58819 1829 58853
rect 1829 58819 1863 58853
rect 1863 58819 1872 58853
rect 1820 58810 1872 58819
rect 94178 58853 94230 58862
rect 94178 58819 94187 58853
rect 94187 58819 94221 58853
rect 94221 58819 94230 58853
rect 94178 58810 94230 58819
rect 1820 58517 1872 58526
rect 1820 58483 1829 58517
rect 1829 58483 1863 58517
rect 1863 58483 1872 58517
rect 1820 58474 1872 58483
rect 94178 58517 94230 58526
rect 94178 58483 94187 58517
rect 94187 58483 94221 58517
rect 94221 58483 94230 58517
rect 94178 58474 94230 58483
rect 1820 58181 1872 58190
rect 1820 58147 1829 58181
rect 1829 58147 1863 58181
rect 1863 58147 1872 58181
rect 1820 58138 1872 58147
rect 94178 58181 94230 58190
rect 94178 58147 94187 58181
rect 94187 58147 94221 58181
rect 94221 58147 94230 58181
rect 94178 58138 94230 58147
rect 1820 57845 1872 57854
rect 1820 57811 1829 57845
rect 1829 57811 1863 57845
rect 1863 57811 1872 57845
rect 1820 57802 1872 57811
rect 94178 57845 94230 57854
rect 94178 57811 94187 57845
rect 94187 57811 94221 57845
rect 94221 57811 94230 57845
rect 94178 57802 94230 57811
rect 1820 57509 1872 57518
rect 1820 57475 1829 57509
rect 1829 57475 1863 57509
rect 1863 57475 1872 57509
rect 1820 57466 1872 57475
rect 94178 57509 94230 57518
rect 94178 57475 94187 57509
rect 94187 57475 94221 57509
rect 94221 57475 94230 57509
rect 94178 57466 94230 57475
rect 1820 57173 1872 57182
rect 1820 57139 1829 57173
rect 1829 57139 1863 57173
rect 1863 57139 1872 57173
rect 1820 57130 1872 57139
rect 94178 57173 94230 57182
rect 94178 57139 94187 57173
rect 94187 57139 94221 57173
rect 94221 57139 94230 57173
rect 94178 57130 94230 57139
rect 1820 56837 1872 56846
rect 1820 56803 1829 56837
rect 1829 56803 1863 56837
rect 1863 56803 1872 56837
rect 1820 56794 1872 56803
rect 94178 56837 94230 56846
rect 94178 56803 94187 56837
rect 94187 56803 94221 56837
rect 94221 56803 94230 56837
rect 94178 56794 94230 56803
rect 1820 56501 1872 56510
rect 1820 56467 1829 56501
rect 1829 56467 1863 56501
rect 1863 56467 1872 56501
rect 1820 56458 1872 56467
rect 94178 56501 94230 56510
rect 94178 56467 94187 56501
rect 94187 56467 94221 56501
rect 94221 56467 94230 56501
rect 94178 56458 94230 56467
rect 1820 56165 1872 56174
rect 1820 56131 1829 56165
rect 1829 56131 1863 56165
rect 1863 56131 1872 56165
rect 1820 56122 1872 56131
rect 94178 56165 94230 56174
rect 94178 56131 94187 56165
rect 94187 56131 94221 56165
rect 94221 56131 94230 56165
rect 94178 56122 94230 56131
rect 1820 55829 1872 55838
rect 1820 55795 1829 55829
rect 1829 55795 1863 55829
rect 1863 55795 1872 55829
rect 1820 55786 1872 55795
rect 94178 55829 94230 55838
rect 94178 55795 94187 55829
rect 94187 55795 94221 55829
rect 94221 55795 94230 55829
rect 94178 55786 94230 55795
rect 1820 55493 1872 55502
rect 1820 55459 1829 55493
rect 1829 55459 1863 55493
rect 1863 55459 1872 55493
rect 1820 55450 1872 55459
rect 94178 55493 94230 55502
rect 94178 55459 94187 55493
rect 94187 55459 94221 55493
rect 94221 55459 94230 55493
rect 94178 55450 94230 55459
rect 1820 55157 1872 55166
rect 1820 55123 1829 55157
rect 1829 55123 1863 55157
rect 1863 55123 1872 55157
rect 1820 55114 1872 55123
rect 94178 55157 94230 55166
rect 94178 55123 94187 55157
rect 94187 55123 94221 55157
rect 94221 55123 94230 55157
rect 94178 55114 94230 55123
rect 1820 54821 1872 54830
rect 1820 54787 1829 54821
rect 1829 54787 1863 54821
rect 1863 54787 1872 54821
rect 1820 54778 1872 54787
rect 94178 54821 94230 54830
rect 94178 54787 94187 54821
rect 94187 54787 94221 54821
rect 94221 54787 94230 54821
rect 94178 54778 94230 54787
rect 1820 54485 1872 54494
rect 1820 54451 1829 54485
rect 1829 54451 1863 54485
rect 1863 54451 1872 54485
rect 1820 54442 1872 54451
rect 94178 54485 94230 54494
rect 94178 54451 94187 54485
rect 94187 54451 94221 54485
rect 94221 54451 94230 54485
rect 94178 54442 94230 54451
rect 1820 54149 1872 54158
rect 1820 54115 1829 54149
rect 1829 54115 1863 54149
rect 1863 54115 1872 54149
rect 1820 54106 1872 54115
rect 94178 54149 94230 54158
rect 94178 54115 94187 54149
rect 94187 54115 94221 54149
rect 94221 54115 94230 54149
rect 94178 54106 94230 54115
rect 1820 53813 1872 53822
rect 1820 53779 1829 53813
rect 1829 53779 1863 53813
rect 1863 53779 1872 53813
rect 1820 53770 1872 53779
rect 94178 53813 94230 53822
rect 94178 53779 94187 53813
rect 94187 53779 94221 53813
rect 94221 53779 94230 53813
rect 94178 53770 94230 53779
rect 1820 53477 1872 53486
rect 1820 53443 1829 53477
rect 1829 53443 1863 53477
rect 1863 53443 1872 53477
rect 1820 53434 1872 53443
rect 94178 53477 94230 53486
rect 94178 53443 94187 53477
rect 94187 53443 94221 53477
rect 94221 53443 94230 53477
rect 94178 53434 94230 53443
rect 1820 53141 1872 53150
rect 1820 53107 1829 53141
rect 1829 53107 1863 53141
rect 1863 53107 1872 53141
rect 1820 53098 1872 53107
rect 94178 53141 94230 53150
rect 94178 53107 94187 53141
rect 94187 53107 94221 53141
rect 94221 53107 94230 53141
rect 94178 53098 94230 53107
rect 1820 52805 1872 52814
rect 1820 52771 1829 52805
rect 1829 52771 1863 52805
rect 1863 52771 1872 52805
rect 1820 52762 1872 52771
rect 94178 52805 94230 52814
rect 94178 52771 94187 52805
rect 94187 52771 94221 52805
rect 94221 52771 94230 52805
rect 94178 52762 94230 52771
rect 1820 52469 1872 52478
rect 1820 52435 1829 52469
rect 1829 52435 1863 52469
rect 1863 52435 1872 52469
rect 1820 52426 1872 52435
rect 94178 52469 94230 52478
rect 94178 52435 94187 52469
rect 94187 52435 94221 52469
rect 94221 52435 94230 52469
rect 94178 52426 94230 52435
rect 1820 52133 1872 52142
rect 1820 52099 1829 52133
rect 1829 52099 1863 52133
rect 1863 52099 1872 52133
rect 1820 52090 1872 52099
rect 94178 52133 94230 52142
rect 94178 52099 94187 52133
rect 94187 52099 94221 52133
rect 94221 52099 94230 52133
rect 94178 52090 94230 52099
rect 1820 51797 1872 51806
rect 1820 51763 1829 51797
rect 1829 51763 1863 51797
rect 1863 51763 1872 51797
rect 1820 51754 1872 51763
rect 94178 51797 94230 51806
rect 94178 51763 94187 51797
rect 94187 51763 94221 51797
rect 94221 51763 94230 51797
rect 94178 51754 94230 51763
rect 1820 51461 1872 51470
rect 1820 51427 1829 51461
rect 1829 51427 1863 51461
rect 1863 51427 1872 51461
rect 1820 51418 1872 51427
rect 94178 51461 94230 51470
rect 94178 51427 94187 51461
rect 94187 51427 94221 51461
rect 94221 51427 94230 51461
rect 94178 51418 94230 51427
rect 1820 51125 1872 51134
rect 1820 51091 1829 51125
rect 1829 51091 1863 51125
rect 1863 51091 1872 51125
rect 1820 51082 1872 51091
rect 94178 51125 94230 51134
rect 94178 51091 94187 51125
rect 94187 51091 94221 51125
rect 94221 51091 94230 51125
rect 94178 51082 94230 51091
rect 1820 50789 1872 50798
rect 1820 50755 1829 50789
rect 1829 50755 1863 50789
rect 1863 50755 1872 50789
rect 1820 50746 1872 50755
rect 94178 50789 94230 50798
rect 94178 50755 94187 50789
rect 94187 50755 94221 50789
rect 94221 50755 94230 50789
rect 94178 50746 94230 50755
rect 1820 50453 1872 50462
rect 1820 50419 1829 50453
rect 1829 50419 1863 50453
rect 1863 50419 1872 50453
rect 1820 50410 1872 50419
rect 94178 50453 94230 50462
rect 94178 50419 94187 50453
rect 94187 50419 94221 50453
rect 94221 50419 94230 50453
rect 94178 50410 94230 50419
rect 1820 50117 1872 50126
rect 1820 50083 1829 50117
rect 1829 50083 1863 50117
rect 1863 50083 1872 50117
rect 1820 50074 1872 50083
rect 94178 50117 94230 50126
rect 94178 50083 94187 50117
rect 94187 50083 94221 50117
rect 94221 50083 94230 50117
rect 94178 50074 94230 50083
rect 1820 49781 1872 49790
rect 1820 49747 1829 49781
rect 1829 49747 1863 49781
rect 1863 49747 1872 49781
rect 1820 49738 1872 49747
rect 94178 49781 94230 49790
rect 94178 49747 94187 49781
rect 94187 49747 94221 49781
rect 94221 49747 94230 49781
rect 94178 49738 94230 49747
rect 1820 49445 1872 49454
rect 1820 49411 1829 49445
rect 1829 49411 1863 49445
rect 1863 49411 1872 49445
rect 1820 49402 1872 49411
rect 94178 49445 94230 49454
rect 94178 49411 94187 49445
rect 94187 49411 94221 49445
rect 94221 49411 94230 49445
rect 94178 49402 94230 49411
rect 1820 49109 1872 49118
rect 1820 49075 1829 49109
rect 1829 49075 1863 49109
rect 1863 49075 1872 49109
rect 1820 49066 1872 49075
rect 94178 49109 94230 49118
rect 94178 49075 94187 49109
rect 94187 49075 94221 49109
rect 94221 49075 94230 49109
rect 94178 49066 94230 49075
rect 1820 48773 1872 48782
rect 1820 48739 1829 48773
rect 1829 48739 1863 48773
rect 1863 48739 1872 48773
rect 1820 48730 1872 48739
rect 94178 48773 94230 48782
rect 94178 48739 94187 48773
rect 94187 48739 94221 48773
rect 94221 48739 94230 48773
rect 94178 48730 94230 48739
rect 1820 48437 1872 48446
rect 1820 48403 1829 48437
rect 1829 48403 1863 48437
rect 1863 48403 1872 48437
rect 1820 48394 1872 48403
rect 94178 48437 94230 48446
rect 94178 48403 94187 48437
rect 94187 48403 94221 48437
rect 94221 48403 94230 48437
rect 94178 48394 94230 48403
rect 1820 48101 1872 48110
rect 1820 48067 1829 48101
rect 1829 48067 1863 48101
rect 1863 48067 1872 48101
rect 1820 48058 1872 48067
rect 94178 48101 94230 48110
rect 94178 48067 94187 48101
rect 94187 48067 94221 48101
rect 94221 48067 94230 48101
rect 94178 48058 94230 48067
rect 1820 47765 1872 47774
rect 1820 47731 1829 47765
rect 1829 47731 1863 47765
rect 1863 47731 1872 47765
rect 1820 47722 1872 47731
rect 94178 47765 94230 47774
rect 94178 47731 94187 47765
rect 94187 47731 94221 47765
rect 94221 47731 94230 47765
rect 94178 47722 94230 47731
rect 1820 47429 1872 47438
rect 1820 47395 1829 47429
rect 1829 47395 1863 47429
rect 1863 47395 1872 47429
rect 1820 47386 1872 47395
rect 94178 47429 94230 47438
rect 94178 47395 94187 47429
rect 94187 47395 94221 47429
rect 94221 47395 94230 47429
rect 94178 47386 94230 47395
rect 1820 47093 1872 47102
rect 1820 47059 1829 47093
rect 1829 47059 1863 47093
rect 1863 47059 1872 47093
rect 1820 47050 1872 47059
rect 94178 47093 94230 47102
rect 94178 47059 94187 47093
rect 94187 47059 94221 47093
rect 94221 47059 94230 47093
rect 94178 47050 94230 47059
rect 1820 46757 1872 46766
rect 1820 46723 1829 46757
rect 1829 46723 1863 46757
rect 1863 46723 1872 46757
rect 1820 46714 1872 46723
rect 94178 46757 94230 46766
rect 94178 46723 94187 46757
rect 94187 46723 94221 46757
rect 94221 46723 94230 46757
rect 94178 46714 94230 46723
rect 1820 46421 1872 46430
rect 1820 46387 1829 46421
rect 1829 46387 1863 46421
rect 1863 46387 1872 46421
rect 1820 46378 1872 46387
rect 94178 46421 94230 46430
rect 94178 46387 94187 46421
rect 94187 46387 94221 46421
rect 94221 46387 94230 46421
rect 94178 46378 94230 46387
rect 1820 46085 1872 46094
rect 1820 46051 1829 46085
rect 1829 46051 1863 46085
rect 1863 46051 1872 46085
rect 1820 46042 1872 46051
rect 94178 46085 94230 46094
rect 94178 46051 94187 46085
rect 94187 46051 94221 46085
rect 94221 46051 94230 46085
rect 94178 46042 94230 46051
rect 1820 45749 1872 45758
rect 1820 45715 1829 45749
rect 1829 45715 1863 45749
rect 1863 45715 1872 45749
rect 1820 45706 1872 45715
rect 94178 45749 94230 45758
rect 94178 45715 94187 45749
rect 94187 45715 94221 45749
rect 94221 45715 94230 45749
rect 94178 45706 94230 45715
rect 1820 45413 1872 45422
rect 1820 45379 1829 45413
rect 1829 45379 1863 45413
rect 1863 45379 1872 45413
rect 1820 45370 1872 45379
rect 94178 45413 94230 45422
rect 94178 45379 94187 45413
rect 94187 45379 94221 45413
rect 94221 45379 94230 45413
rect 94178 45370 94230 45379
rect 1820 45077 1872 45086
rect 1820 45043 1829 45077
rect 1829 45043 1863 45077
rect 1863 45043 1872 45077
rect 1820 45034 1872 45043
rect 94178 45077 94230 45086
rect 94178 45043 94187 45077
rect 94187 45043 94221 45077
rect 94221 45043 94230 45077
rect 94178 45034 94230 45043
rect 1820 44741 1872 44750
rect 1820 44707 1829 44741
rect 1829 44707 1863 44741
rect 1863 44707 1872 44741
rect 1820 44698 1872 44707
rect 94178 44741 94230 44750
rect 94178 44707 94187 44741
rect 94187 44707 94221 44741
rect 94221 44707 94230 44741
rect 94178 44698 94230 44707
rect 1820 44405 1872 44414
rect 1820 44371 1829 44405
rect 1829 44371 1863 44405
rect 1863 44371 1872 44405
rect 1820 44362 1872 44371
rect 94178 44405 94230 44414
rect 94178 44371 94187 44405
rect 94187 44371 94221 44405
rect 94221 44371 94230 44405
rect 94178 44362 94230 44371
rect 1820 44069 1872 44078
rect 1820 44035 1829 44069
rect 1829 44035 1863 44069
rect 1863 44035 1872 44069
rect 1820 44026 1872 44035
rect 94178 44069 94230 44078
rect 94178 44035 94187 44069
rect 94187 44035 94221 44069
rect 94221 44035 94230 44069
rect 94178 44026 94230 44035
rect 1820 43733 1872 43742
rect 1820 43699 1829 43733
rect 1829 43699 1863 43733
rect 1863 43699 1872 43733
rect 1820 43690 1872 43699
rect 94178 43733 94230 43742
rect 94178 43699 94187 43733
rect 94187 43699 94221 43733
rect 94221 43699 94230 43733
rect 94178 43690 94230 43699
rect 1820 43397 1872 43406
rect 1820 43363 1829 43397
rect 1829 43363 1863 43397
rect 1863 43363 1872 43397
rect 1820 43354 1872 43363
rect 94178 43397 94230 43406
rect 94178 43363 94187 43397
rect 94187 43363 94221 43397
rect 94221 43363 94230 43397
rect 94178 43354 94230 43363
rect 1820 43061 1872 43070
rect 1820 43027 1829 43061
rect 1829 43027 1863 43061
rect 1863 43027 1872 43061
rect 1820 43018 1872 43027
rect 94178 43061 94230 43070
rect 94178 43027 94187 43061
rect 94187 43027 94221 43061
rect 94221 43027 94230 43061
rect 94178 43018 94230 43027
rect 1820 42725 1872 42734
rect 1820 42691 1829 42725
rect 1829 42691 1863 42725
rect 1863 42691 1872 42725
rect 1820 42682 1872 42691
rect 94178 42725 94230 42734
rect 94178 42691 94187 42725
rect 94187 42691 94221 42725
rect 94221 42691 94230 42725
rect 94178 42682 94230 42691
rect 1820 42389 1872 42398
rect 1820 42355 1829 42389
rect 1829 42355 1863 42389
rect 1863 42355 1872 42389
rect 1820 42346 1872 42355
rect 94178 42389 94230 42398
rect 94178 42355 94187 42389
rect 94187 42355 94221 42389
rect 94221 42355 94230 42389
rect 94178 42346 94230 42355
rect 1820 42053 1872 42062
rect 1820 42019 1829 42053
rect 1829 42019 1863 42053
rect 1863 42019 1872 42053
rect 1820 42010 1872 42019
rect 94178 42053 94230 42062
rect 94178 42019 94187 42053
rect 94187 42019 94221 42053
rect 94221 42019 94230 42053
rect 94178 42010 94230 42019
rect 1820 41717 1872 41726
rect 1820 41683 1829 41717
rect 1829 41683 1863 41717
rect 1863 41683 1872 41717
rect 1820 41674 1872 41683
rect 94178 41717 94230 41726
rect 94178 41683 94187 41717
rect 94187 41683 94221 41717
rect 94221 41683 94230 41717
rect 94178 41674 94230 41683
rect 1820 41381 1872 41390
rect 1820 41347 1829 41381
rect 1829 41347 1863 41381
rect 1863 41347 1872 41381
rect 1820 41338 1872 41347
rect 94178 41381 94230 41390
rect 94178 41347 94187 41381
rect 94187 41347 94221 41381
rect 94221 41347 94230 41381
rect 94178 41338 94230 41347
rect 1820 41045 1872 41054
rect 1820 41011 1829 41045
rect 1829 41011 1863 41045
rect 1863 41011 1872 41045
rect 1820 41002 1872 41011
rect 94178 41045 94230 41054
rect 94178 41011 94187 41045
rect 94187 41011 94221 41045
rect 94221 41011 94230 41045
rect 94178 41002 94230 41011
rect 1820 40709 1872 40718
rect 1820 40675 1829 40709
rect 1829 40675 1863 40709
rect 1863 40675 1872 40709
rect 1820 40666 1872 40675
rect 94178 40709 94230 40718
rect 94178 40675 94187 40709
rect 94187 40675 94221 40709
rect 94221 40675 94230 40709
rect 94178 40666 94230 40675
rect 1820 40373 1872 40382
rect 1820 40339 1829 40373
rect 1829 40339 1863 40373
rect 1863 40339 1872 40373
rect 1820 40330 1872 40339
rect 94178 40373 94230 40382
rect 94178 40339 94187 40373
rect 94187 40339 94221 40373
rect 94221 40339 94230 40373
rect 94178 40330 94230 40339
rect 1820 40037 1872 40046
rect 1820 40003 1829 40037
rect 1829 40003 1863 40037
rect 1863 40003 1872 40037
rect 1820 39994 1872 40003
rect 94178 40037 94230 40046
rect 94178 40003 94187 40037
rect 94187 40003 94221 40037
rect 94221 40003 94230 40037
rect 94178 39994 94230 40003
rect 1820 39701 1872 39710
rect 1820 39667 1829 39701
rect 1829 39667 1863 39701
rect 1863 39667 1872 39701
rect 1820 39658 1872 39667
rect 94178 39701 94230 39710
rect 94178 39667 94187 39701
rect 94187 39667 94221 39701
rect 94221 39667 94230 39701
rect 94178 39658 94230 39667
rect 1820 39365 1872 39374
rect 1820 39331 1829 39365
rect 1829 39331 1863 39365
rect 1863 39331 1872 39365
rect 1820 39322 1872 39331
rect 94178 39365 94230 39374
rect 94178 39331 94187 39365
rect 94187 39331 94221 39365
rect 94221 39331 94230 39365
rect 94178 39322 94230 39331
rect 1820 39029 1872 39038
rect 1820 38995 1829 39029
rect 1829 38995 1863 39029
rect 1863 38995 1872 39029
rect 1820 38986 1872 38995
rect 94178 39029 94230 39038
rect 94178 38995 94187 39029
rect 94187 38995 94221 39029
rect 94221 38995 94230 39029
rect 94178 38986 94230 38995
rect 1820 38693 1872 38702
rect 1820 38659 1829 38693
rect 1829 38659 1863 38693
rect 1863 38659 1872 38693
rect 1820 38650 1872 38659
rect 94178 38693 94230 38702
rect 94178 38659 94187 38693
rect 94187 38659 94221 38693
rect 94221 38659 94230 38693
rect 94178 38650 94230 38659
rect 1820 38357 1872 38366
rect 1820 38323 1829 38357
rect 1829 38323 1863 38357
rect 1863 38323 1872 38357
rect 1820 38314 1872 38323
rect 94178 38357 94230 38366
rect 94178 38323 94187 38357
rect 94187 38323 94221 38357
rect 94221 38323 94230 38357
rect 94178 38314 94230 38323
rect 1820 38021 1872 38030
rect 1820 37987 1829 38021
rect 1829 37987 1863 38021
rect 1863 37987 1872 38021
rect 1820 37978 1872 37987
rect 94178 38021 94230 38030
rect 94178 37987 94187 38021
rect 94187 37987 94221 38021
rect 94221 37987 94230 38021
rect 94178 37978 94230 37987
rect 1820 37685 1872 37694
rect 1820 37651 1829 37685
rect 1829 37651 1863 37685
rect 1863 37651 1872 37685
rect 1820 37642 1872 37651
rect 94178 37685 94230 37694
rect 94178 37651 94187 37685
rect 94187 37651 94221 37685
rect 94221 37651 94230 37685
rect 94178 37642 94230 37651
rect 1820 37349 1872 37358
rect 1820 37315 1829 37349
rect 1829 37315 1863 37349
rect 1863 37315 1872 37349
rect 1820 37306 1872 37315
rect 94178 37349 94230 37358
rect 94178 37315 94187 37349
rect 94187 37315 94221 37349
rect 94221 37315 94230 37349
rect 94178 37306 94230 37315
rect 1820 37013 1872 37022
rect 1820 36979 1829 37013
rect 1829 36979 1863 37013
rect 1863 36979 1872 37013
rect 1820 36970 1872 36979
rect 94178 37013 94230 37022
rect 94178 36979 94187 37013
rect 94187 36979 94221 37013
rect 94221 36979 94230 37013
rect 94178 36970 94230 36979
rect 1820 36677 1872 36686
rect 1820 36643 1829 36677
rect 1829 36643 1863 36677
rect 1863 36643 1872 36677
rect 1820 36634 1872 36643
rect 94178 36677 94230 36686
rect 94178 36643 94187 36677
rect 94187 36643 94221 36677
rect 94221 36643 94230 36677
rect 94178 36634 94230 36643
rect 1820 36341 1872 36350
rect 1820 36307 1829 36341
rect 1829 36307 1863 36341
rect 1863 36307 1872 36341
rect 1820 36298 1872 36307
rect 94178 36341 94230 36350
rect 94178 36307 94187 36341
rect 94187 36307 94221 36341
rect 94221 36307 94230 36341
rect 94178 36298 94230 36307
rect 1820 36005 1872 36014
rect 1820 35971 1829 36005
rect 1829 35971 1863 36005
rect 1863 35971 1872 36005
rect 1820 35962 1872 35971
rect 94178 36005 94230 36014
rect 94178 35971 94187 36005
rect 94187 35971 94221 36005
rect 94221 35971 94230 36005
rect 94178 35962 94230 35971
rect 1820 35669 1872 35678
rect 1820 35635 1829 35669
rect 1829 35635 1863 35669
rect 1863 35635 1872 35669
rect 1820 35626 1872 35635
rect 94178 35669 94230 35678
rect 94178 35635 94187 35669
rect 94187 35635 94221 35669
rect 94221 35635 94230 35669
rect 94178 35626 94230 35635
rect 1820 35333 1872 35342
rect 1820 35299 1829 35333
rect 1829 35299 1863 35333
rect 1863 35299 1872 35333
rect 1820 35290 1872 35299
rect 94178 35333 94230 35342
rect 94178 35299 94187 35333
rect 94187 35299 94221 35333
rect 94221 35299 94230 35333
rect 94178 35290 94230 35299
rect 1820 34997 1872 35006
rect 1820 34963 1829 34997
rect 1829 34963 1863 34997
rect 1863 34963 1872 34997
rect 1820 34954 1872 34963
rect 94178 34997 94230 35006
rect 94178 34963 94187 34997
rect 94187 34963 94221 34997
rect 94221 34963 94230 34997
rect 94178 34954 94230 34963
rect 1820 34661 1872 34670
rect 1820 34627 1829 34661
rect 1829 34627 1863 34661
rect 1863 34627 1872 34661
rect 1820 34618 1872 34627
rect 94178 34661 94230 34670
rect 94178 34627 94187 34661
rect 94187 34627 94221 34661
rect 94221 34627 94230 34661
rect 94178 34618 94230 34627
rect 1820 34325 1872 34334
rect 1820 34291 1829 34325
rect 1829 34291 1863 34325
rect 1863 34291 1872 34325
rect 1820 34282 1872 34291
rect 94178 34325 94230 34334
rect 94178 34291 94187 34325
rect 94187 34291 94221 34325
rect 94221 34291 94230 34325
rect 94178 34282 94230 34291
rect 14941 34143 14993 34195
rect 1820 33989 1872 33998
rect 1820 33955 1829 33989
rect 1829 33955 1863 33989
rect 1863 33955 1872 33989
rect 1820 33946 1872 33955
rect 1820 33653 1872 33662
rect 1820 33619 1829 33653
rect 1829 33619 1863 33653
rect 1863 33619 1872 33653
rect 1820 33610 1872 33619
rect 1820 33317 1872 33326
rect 1820 33283 1829 33317
rect 1829 33283 1863 33317
rect 1863 33283 1872 33317
rect 1820 33274 1872 33283
rect 1820 32981 1872 32990
rect 1820 32947 1829 32981
rect 1829 32947 1863 32981
rect 1863 32947 1872 32981
rect 1820 32938 1872 32947
rect 14861 32873 14913 32925
rect 1820 32645 1872 32654
rect 1820 32611 1829 32645
rect 1829 32611 1863 32645
rect 1863 32611 1872 32645
rect 1820 32602 1872 32611
rect 1820 32309 1872 32318
rect 1820 32275 1829 32309
rect 1829 32275 1863 32309
rect 1863 32275 1872 32309
rect 1820 32266 1872 32275
rect 1820 31973 1872 31982
rect 1820 31939 1829 31973
rect 1829 31939 1863 31973
rect 1863 31939 1872 31973
rect 1820 31930 1872 31939
rect 1820 31637 1872 31646
rect 1820 31603 1829 31637
rect 1829 31603 1863 31637
rect 1863 31603 1872 31637
rect 1820 31594 1872 31603
rect 14781 31315 14833 31367
rect 1820 31301 1872 31310
rect 1820 31267 1829 31301
rect 1829 31267 1863 31301
rect 1863 31267 1872 31301
rect 1820 31258 1872 31267
rect 1820 30965 1872 30974
rect 1820 30931 1829 30965
rect 1829 30931 1863 30965
rect 1863 30931 1872 30965
rect 1820 30922 1872 30931
rect 1820 30629 1872 30638
rect 1820 30595 1829 30629
rect 1829 30595 1863 30629
rect 1863 30595 1872 30629
rect 1820 30586 1872 30595
rect 1820 30293 1872 30302
rect 1820 30259 1829 30293
rect 1829 30259 1863 30293
rect 1863 30259 1872 30293
rect 1820 30250 1872 30259
rect 14701 30045 14753 30097
rect 1820 29957 1872 29966
rect 1820 29923 1829 29957
rect 1829 29923 1863 29957
rect 1863 29923 1872 29957
rect 1820 29914 1872 29923
rect 1820 29621 1872 29630
rect 1820 29587 1829 29621
rect 1829 29587 1863 29621
rect 1863 29587 1872 29621
rect 1820 29578 1872 29587
rect 1820 29285 1872 29294
rect 1820 29251 1829 29285
rect 1829 29251 1863 29285
rect 1863 29251 1872 29285
rect 1820 29242 1872 29251
rect 1820 28949 1872 28958
rect 1820 28915 1829 28949
rect 1829 28915 1863 28949
rect 1863 28915 1872 28949
rect 1820 28906 1872 28915
rect 1820 28613 1872 28622
rect 1820 28579 1829 28613
rect 1829 28579 1863 28613
rect 1863 28579 1872 28613
rect 1820 28570 1872 28579
rect 14621 28487 14673 28539
rect 1820 28277 1872 28286
rect 1820 28243 1829 28277
rect 1829 28243 1863 28277
rect 1863 28243 1872 28277
rect 1820 28234 1872 28243
rect 1820 27941 1872 27950
rect 1820 27907 1829 27941
rect 1829 27907 1863 27941
rect 1863 27907 1872 27941
rect 1820 27898 1872 27907
rect 1820 27605 1872 27614
rect 1820 27571 1829 27605
rect 1829 27571 1863 27605
rect 1863 27571 1872 27605
rect 1820 27562 1872 27571
rect 1820 27269 1872 27278
rect 1820 27235 1829 27269
rect 1829 27235 1863 27269
rect 1863 27235 1872 27269
rect 1820 27226 1872 27235
rect 14541 27217 14593 27269
rect 1820 26933 1872 26942
rect 1820 26899 1829 26933
rect 1829 26899 1863 26933
rect 1863 26899 1872 26933
rect 1820 26890 1872 26899
rect 1820 26597 1872 26606
rect 1820 26563 1829 26597
rect 1829 26563 1863 26597
rect 1863 26563 1872 26597
rect 1820 26554 1872 26563
rect 1820 26261 1872 26270
rect 1820 26227 1829 26261
rect 1829 26227 1863 26261
rect 1863 26227 1872 26261
rect 1820 26218 1872 26227
rect 1820 25925 1872 25934
rect 1820 25891 1829 25925
rect 1829 25891 1863 25925
rect 1863 25891 1872 25925
rect 1820 25882 1872 25891
rect 14461 25659 14513 25711
rect 1820 25589 1872 25598
rect 1820 25555 1829 25589
rect 1829 25555 1863 25589
rect 1863 25555 1872 25589
rect 1820 25546 1872 25555
rect 1820 25253 1872 25262
rect 1820 25219 1829 25253
rect 1829 25219 1863 25253
rect 1863 25219 1872 25253
rect 1820 25210 1872 25219
rect 1820 24917 1872 24926
rect 1820 24883 1829 24917
rect 1829 24883 1863 24917
rect 1863 24883 1872 24917
rect 1820 24874 1872 24883
rect 1820 24581 1872 24590
rect 1820 24547 1829 24581
rect 1829 24547 1863 24581
rect 1863 24547 1872 24581
rect 1820 24538 1872 24547
rect 1820 24245 1872 24254
rect 1820 24211 1829 24245
rect 1829 24211 1863 24245
rect 1863 24211 1872 24245
rect 1820 24202 1872 24211
rect 1820 23909 1872 23918
rect 1820 23875 1829 23909
rect 1829 23875 1863 23909
rect 1863 23875 1872 23909
rect 1820 23866 1872 23875
rect 1820 23573 1872 23582
rect 1820 23539 1829 23573
rect 1829 23539 1863 23573
rect 1863 23539 1872 23573
rect 1820 23530 1872 23539
rect 1820 23237 1872 23246
rect 1820 23203 1829 23237
rect 1829 23203 1863 23237
rect 1863 23203 1872 23237
rect 1820 23194 1872 23203
rect 1820 22901 1872 22910
rect 1820 22867 1829 22901
rect 1829 22867 1863 22901
rect 1863 22867 1872 22901
rect 1820 22858 1872 22867
rect 1820 22565 1872 22574
rect 1820 22531 1829 22565
rect 1829 22531 1863 22565
rect 1863 22531 1872 22565
rect 1820 22522 1872 22531
rect 1820 22229 1872 22238
rect 1820 22195 1829 22229
rect 1829 22195 1863 22229
rect 1863 22195 1872 22229
rect 1820 22186 1872 22195
rect 1820 21893 1872 21902
rect 1820 21859 1829 21893
rect 1829 21859 1863 21893
rect 1863 21859 1872 21893
rect 1820 21850 1872 21859
rect 1820 21557 1872 21566
rect 1820 21523 1829 21557
rect 1829 21523 1863 21557
rect 1863 21523 1872 21557
rect 1820 21514 1872 21523
rect 1820 21221 1872 21230
rect 1820 21187 1829 21221
rect 1829 21187 1863 21221
rect 1863 21187 1872 21221
rect 1820 21178 1872 21187
rect 94178 33989 94230 33998
rect 94178 33955 94187 33989
rect 94187 33955 94221 33989
rect 94221 33955 94230 33989
rect 94178 33946 94230 33955
rect 94178 33653 94230 33662
rect 94178 33619 94187 33653
rect 94187 33619 94221 33653
rect 94221 33619 94230 33653
rect 94178 33610 94230 33619
rect 94178 33317 94230 33326
rect 94178 33283 94187 33317
rect 94187 33283 94221 33317
rect 94221 33283 94230 33317
rect 94178 33274 94230 33283
rect 94178 32981 94230 32990
rect 94178 32947 94187 32981
rect 94187 32947 94221 32981
rect 94221 32947 94230 32981
rect 94178 32938 94230 32947
rect 94178 32645 94230 32654
rect 94178 32611 94187 32645
rect 94187 32611 94221 32645
rect 94221 32611 94230 32645
rect 94178 32602 94230 32611
rect 94178 32309 94230 32318
rect 94178 32275 94187 32309
rect 94187 32275 94221 32309
rect 94221 32275 94230 32309
rect 94178 32266 94230 32275
rect 94178 31973 94230 31982
rect 94178 31939 94187 31973
rect 94187 31939 94221 31973
rect 94221 31939 94230 31973
rect 94178 31930 94230 31939
rect 94178 31637 94230 31646
rect 94178 31603 94187 31637
rect 94187 31603 94221 31637
rect 94221 31603 94230 31637
rect 94178 31594 94230 31603
rect 94178 31301 94230 31310
rect 94178 31267 94187 31301
rect 94187 31267 94221 31301
rect 94221 31267 94230 31301
rect 94178 31258 94230 31267
rect 94178 30965 94230 30974
rect 94178 30931 94187 30965
rect 94187 30931 94221 30965
rect 94221 30931 94230 30965
rect 94178 30922 94230 30931
rect 94178 30629 94230 30638
rect 94178 30595 94187 30629
rect 94187 30595 94221 30629
rect 94221 30595 94230 30629
rect 94178 30586 94230 30595
rect 94178 30293 94230 30302
rect 94178 30259 94187 30293
rect 94187 30259 94221 30293
rect 94221 30259 94230 30293
rect 94178 30250 94230 30259
rect 94178 29957 94230 29966
rect 94178 29923 94187 29957
rect 94187 29923 94221 29957
rect 94221 29923 94230 29957
rect 94178 29914 94230 29923
rect 94178 29621 94230 29630
rect 94178 29587 94187 29621
rect 94187 29587 94221 29621
rect 94221 29587 94230 29621
rect 94178 29578 94230 29587
rect 94178 29285 94230 29294
rect 94178 29251 94187 29285
rect 94187 29251 94221 29285
rect 94221 29251 94230 29285
rect 94178 29242 94230 29251
rect 94178 28949 94230 28958
rect 94178 28915 94187 28949
rect 94187 28915 94221 28949
rect 94221 28915 94230 28949
rect 94178 28906 94230 28915
rect 94178 28613 94230 28622
rect 94178 28579 94187 28613
rect 94187 28579 94221 28613
rect 94221 28579 94230 28613
rect 94178 28570 94230 28579
rect 94178 28277 94230 28286
rect 94178 28243 94187 28277
rect 94187 28243 94221 28277
rect 94221 28243 94230 28277
rect 94178 28234 94230 28243
rect 94178 27941 94230 27950
rect 94178 27907 94187 27941
rect 94187 27907 94221 27941
rect 94221 27907 94230 27941
rect 94178 27898 94230 27907
rect 94178 27605 94230 27614
rect 94178 27571 94187 27605
rect 94187 27571 94221 27605
rect 94221 27571 94230 27605
rect 94178 27562 94230 27571
rect 94178 27269 94230 27278
rect 94178 27235 94187 27269
rect 94187 27235 94221 27269
rect 94221 27235 94230 27269
rect 94178 27226 94230 27235
rect 94178 26933 94230 26942
rect 94178 26899 94187 26933
rect 94187 26899 94221 26933
rect 94221 26899 94230 26933
rect 94178 26890 94230 26899
rect 94178 26597 94230 26606
rect 94178 26563 94187 26597
rect 94187 26563 94221 26597
rect 94221 26563 94230 26597
rect 94178 26554 94230 26563
rect 94178 26261 94230 26270
rect 94178 26227 94187 26261
rect 94187 26227 94221 26261
rect 94221 26227 94230 26261
rect 94178 26218 94230 26227
rect 94178 25925 94230 25934
rect 94178 25891 94187 25925
rect 94187 25891 94221 25925
rect 94221 25891 94230 25925
rect 94178 25882 94230 25891
rect 94178 25589 94230 25598
rect 94178 25555 94187 25589
rect 94187 25555 94221 25589
rect 94221 25555 94230 25589
rect 94178 25546 94230 25555
rect 94178 25253 94230 25262
rect 94178 25219 94187 25253
rect 94187 25219 94221 25253
rect 94221 25219 94230 25253
rect 94178 25210 94230 25219
rect 94178 24917 94230 24926
rect 94178 24883 94187 24917
rect 94187 24883 94221 24917
rect 94221 24883 94230 24917
rect 94178 24874 94230 24883
rect 94178 24581 94230 24590
rect 94178 24547 94187 24581
rect 94187 24547 94221 24581
rect 94221 24547 94230 24581
rect 94178 24538 94230 24547
rect 94178 24245 94230 24254
rect 94178 24211 94187 24245
rect 94187 24211 94221 24245
rect 94221 24211 94230 24245
rect 94178 24202 94230 24211
rect 94178 23909 94230 23918
rect 94178 23875 94187 23909
rect 94187 23875 94221 23909
rect 94221 23875 94230 23909
rect 94178 23866 94230 23875
rect 94178 23573 94230 23582
rect 94178 23539 94187 23573
rect 94187 23539 94221 23573
rect 94221 23539 94230 23573
rect 94178 23530 94230 23539
rect 94178 23237 94230 23246
rect 94178 23203 94187 23237
rect 94187 23203 94221 23237
rect 94221 23203 94230 23237
rect 94178 23194 94230 23203
rect 94178 22901 94230 22910
rect 94178 22867 94187 22901
rect 94187 22867 94221 22901
rect 94221 22867 94230 22901
rect 94178 22858 94230 22867
rect 94178 22565 94230 22574
rect 94178 22531 94187 22565
rect 94187 22531 94221 22565
rect 94221 22531 94230 22565
rect 94178 22522 94230 22531
rect 94178 22229 94230 22238
rect 94178 22195 94187 22229
rect 94187 22195 94221 22229
rect 94221 22195 94230 22229
rect 94178 22186 94230 22195
rect 94178 21893 94230 21902
rect 94178 21859 94187 21893
rect 94187 21859 94221 21893
rect 94221 21859 94230 21893
rect 94178 21850 94230 21859
rect 94178 21557 94230 21566
rect 94178 21523 94187 21557
rect 94187 21523 94221 21557
rect 94221 21523 94230 21557
rect 94178 21514 94230 21523
rect 94178 21221 94230 21230
rect 94178 21187 94187 21221
rect 94187 21187 94221 21221
rect 94221 21187 94230 21221
rect 94178 21178 94230 21187
rect 1820 20885 1872 20894
rect 1820 20851 1829 20885
rect 1829 20851 1863 20885
rect 1863 20851 1872 20885
rect 1820 20842 1872 20851
rect 1820 20549 1872 20558
rect 1820 20515 1829 20549
rect 1829 20515 1863 20549
rect 1863 20515 1872 20549
rect 1820 20506 1872 20515
rect 1820 20213 1872 20222
rect 1820 20179 1829 20213
rect 1829 20179 1863 20213
rect 1863 20179 1872 20213
rect 1820 20170 1872 20179
rect 1820 19877 1872 19886
rect 1820 19843 1829 19877
rect 1829 19843 1863 19877
rect 1863 19843 1872 19877
rect 1820 19834 1872 19843
rect 1820 19541 1872 19550
rect 1820 19507 1829 19541
rect 1829 19507 1863 19541
rect 1863 19507 1872 19541
rect 1820 19498 1872 19507
rect 1820 19205 1872 19214
rect 1820 19171 1829 19205
rect 1829 19171 1863 19205
rect 1863 19171 1872 19205
rect 1820 19162 1872 19171
rect 1820 18869 1872 18878
rect 1820 18835 1829 18869
rect 1829 18835 1863 18869
rect 1863 18835 1872 18869
rect 1820 18826 1872 18835
rect 1820 18533 1872 18542
rect 1820 18499 1829 18533
rect 1829 18499 1863 18533
rect 1863 18499 1872 18533
rect 1820 18490 1872 18499
rect 1820 18197 1872 18206
rect 1820 18163 1829 18197
rect 1829 18163 1863 18197
rect 1863 18163 1872 18197
rect 1820 18154 1872 18163
rect 1820 17861 1872 17870
rect 1820 17827 1829 17861
rect 1829 17827 1863 17861
rect 1863 17827 1872 17861
rect 1820 17818 1872 17827
rect 1820 17525 1872 17534
rect 1820 17491 1829 17525
rect 1829 17491 1863 17525
rect 1863 17491 1872 17525
rect 1820 17482 1872 17491
rect 1820 17189 1872 17198
rect 1820 17155 1829 17189
rect 1829 17155 1863 17189
rect 1863 17155 1872 17189
rect 1820 17146 1872 17155
rect 1820 16853 1872 16862
rect 1820 16819 1829 16853
rect 1829 16819 1863 16853
rect 1863 16819 1872 16853
rect 1820 16810 1872 16819
rect 1820 16517 1872 16526
rect 1820 16483 1829 16517
rect 1829 16483 1863 16517
rect 1863 16483 1872 16517
rect 1820 16474 1872 16483
rect 1820 16181 1872 16190
rect 1820 16147 1829 16181
rect 1829 16147 1863 16181
rect 1863 16147 1872 16181
rect 1820 16138 1872 16147
rect 1820 15845 1872 15854
rect 1820 15811 1829 15845
rect 1829 15811 1863 15845
rect 1863 15811 1872 15845
rect 1820 15802 1872 15811
rect 1820 15509 1872 15518
rect 1820 15475 1829 15509
rect 1829 15475 1863 15509
rect 1863 15475 1872 15509
rect 1820 15466 1872 15475
rect 1820 15173 1872 15182
rect 1820 15139 1829 15173
rect 1829 15139 1863 15173
rect 1863 15139 1872 15173
rect 1820 15130 1872 15139
rect 1820 14837 1872 14846
rect 1820 14803 1829 14837
rect 1829 14803 1863 14837
rect 1863 14803 1872 14837
rect 1820 14794 1872 14803
rect 1820 14501 1872 14510
rect 1820 14467 1829 14501
rect 1829 14467 1863 14501
rect 1863 14467 1872 14501
rect 1820 14458 1872 14467
rect 1820 14165 1872 14174
rect 1820 14131 1829 14165
rect 1829 14131 1863 14165
rect 1863 14131 1872 14165
rect 1820 14122 1872 14131
rect 1820 13829 1872 13838
rect 1820 13795 1829 13829
rect 1829 13795 1863 13829
rect 1863 13795 1872 13829
rect 1820 13786 1872 13795
rect 1820 13493 1872 13502
rect 1820 13459 1829 13493
rect 1829 13459 1863 13493
rect 1863 13459 1872 13493
rect 1820 13450 1872 13459
rect 1820 13157 1872 13166
rect 1820 13123 1829 13157
rect 1829 13123 1863 13157
rect 1863 13123 1872 13157
rect 1820 13114 1872 13123
rect 1820 12821 1872 12830
rect 1820 12787 1829 12821
rect 1829 12787 1863 12821
rect 1863 12787 1872 12821
rect 1820 12778 1872 12787
rect 1820 12485 1872 12494
rect 1820 12451 1829 12485
rect 1829 12451 1863 12485
rect 1863 12451 1872 12485
rect 1820 12442 1872 12451
rect 1820 12149 1872 12158
rect 1820 12115 1829 12149
rect 1829 12115 1863 12149
rect 1863 12115 1872 12149
rect 1820 12106 1872 12115
rect 1820 11813 1872 11822
rect 1820 11779 1829 11813
rect 1829 11779 1863 11813
rect 1863 11779 1872 11813
rect 1820 11770 1872 11779
rect 1820 11477 1872 11486
rect 1820 11443 1829 11477
rect 1829 11443 1863 11477
rect 1863 11443 1872 11477
rect 1820 11434 1872 11443
rect 1820 11141 1872 11150
rect 1820 11107 1829 11141
rect 1829 11107 1863 11141
rect 1863 11107 1872 11141
rect 1820 11098 1872 11107
rect 1820 10805 1872 10814
rect 1820 10771 1829 10805
rect 1829 10771 1863 10805
rect 1863 10771 1872 10805
rect 1820 10762 1872 10771
rect 28212 10759 28264 10811
rect 29460 10759 29512 10811
rect 30708 10759 30760 10811
rect 31956 10759 32008 10811
rect 33204 10759 33256 10811
rect 34452 10759 34504 10811
rect 35700 10759 35752 10811
rect 36948 10759 37000 10811
rect 38196 10759 38248 10811
rect 39444 10759 39496 10811
rect 40692 10759 40744 10811
rect 41940 10759 41992 10811
rect 43188 10759 43240 10811
rect 44436 10759 44488 10811
rect 45684 10759 45736 10811
rect 46932 10759 46984 10811
rect 48180 10759 48232 10811
rect 49428 10759 49480 10811
rect 50676 10759 50728 10811
rect 51924 10759 51976 10811
rect 53172 10759 53224 10811
rect 54420 10759 54472 10811
rect 55668 10759 55720 10811
rect 56916 10759 56968 10811
rect 58164 10759 58216 10811
rect 59412 10759 59464 10811
rect 60660 10759 60712 10811
rect 61908 10759 61960 10811
rect 63156 10759 63208 10811
rect 64404 10759 64456 10811
rect 65652 10759 65704 10811
rect 66900 10759 66952 10811
rect 1820 10469 1872 10478
rect 1820 10435 1829 10469
rect 1829 10435 1863 10469
rect 1863 10435 1872 10469
rect 1820 10426 1872 10435
rect 1820 10133 1872 10142
rect 1820 10099 1829 10133
rect 1829 10099 1863 10133
rect 1863 10099 1872 10133
rect 1820 10090 1872 10099
rect 1820 9797 1872 9806
rect 1820 9763 1829 9797
rect 1829 9763 1863 9797
rect 1863 9763 1872 9797
rect 1820 9754 1872 9763
rect 1820 9461 1872 9470
rect 1820 9427 1829 9461
rect 1829 9427 1863 9461
rect 1863 9427 1872 9461
rect 1820 9418 1872 9427
rect 1820 9125 1872 9134
rect 1820 9091 1829 9125
rect 1829 9091 1863 9125
rect 1863 9091 1872 9125
rect 1820 9082 1872 9091
rect 1820 8789 1872 8798
rect 1820 8755 1829 8789
rect 1829 8755 1863 8789
rect 1863 8755 1872 8789
rect 1820 8746 1872 8755
rect 1820 8453 1872 8462
rect 1820 8419 1829 8453
rect 1829 8419 1863 8453
rect 1863 8419 1872 8453
rect 1820 8410 1872 8419
rect 1820 8117 1872 8126
rect 1820 8083 1829 8117
rect 1829 8083 1863 8117
rect 1863 8083 1872 8117
rect 1820 8074 1872 8083
rect 94178 20885 94230 20894
rect 94178 20851 94187 20885
rect 94187 20851 94221 20885
rect 94221 20851 94230 20885
rect 94178 20842 94230 20851
rect 94178 20549 94230 20558
rect 94178 20515 94187 20549
rect 94187 20515 94221 20549
rect 94221 20515 94230 20549
rect 94178 20506 94230 20515
rect 94178 20213 94230 20222
rect 94178 20179 94187 20213
rect 94187 20179 94221 20213
rect 94221 20179 94230 20213
rect 94178 20170 94230 20179
rect 94178 19877 94230 19886
rect 94178 19843 94187 19877
rect 94187 19843 94221 19877
rect 94221 19843 94230 19877
rect 94178 19834 94230 19843
rect 94178 19541 94230 19550
rect 94178 19507 94187 19541
rect 94187 19507 94221 19541
rect 94221 19507 94230 19541
rect 94178 19498 94230 19507
rect 94178 19205 94230 19214
rect 94178 19171 94187 19205
rect 94187 19171 94221 19205
rect 94221 19171 94230 19205
rect 94178 19162 94230 19171
rect 94178 18869 94230 18878
rect 94178 18835 94187 18869
rect 94187 18835 94221 18869
rect 94221 18835 94230 18869
rect 94178 18826 94230 18835
rect 94178 18533 94230 18542
rect 94178 18499 94187 18533
rect 94187 18499 94221 18533
rect 94221 18499 94230 18533
rect 94178 18490 94230 18499
rect 94178 18197 94230 18206
rect 94178 18163 94187 18197
rect 94187 18163 94221 18197
rect 94221 18163 94230 18197
rect 94178 18154 94230 18163
rect 94178 17861 94230 17870
rect 94178 17827 94187 17861
rect 94187 17827 94221 17861
rect 94221 17827 94230 17861
rect 94178 17818 94230 17827
rect 94178 17525 94230 17534
rect 94178 17491 94187 17525
rect 94187 17491 94221 17525
rect 94221 17491 94230 17525
rect 94178 17482 94230 17491
rect 94178 17189 94230 17198
rect 94178 17155 94187 17189
rect 94187 17155 94221 17189
rect 94221 17155 94230 17189
rect 94178 17146 94230 17155
rect 94178 16853 94230 16862
rect 94178 16819 94187 16853
rect 94187 16819 94221 16853
rect 94221 16819 94230 16853
rect 94178 16810 94230 16819
rect 81645 16489 81697 16541
rect 94178 16517 94230 16526
rect 94178 16483 94187 16517
rect 94187 16483 94221 16517
rect 94221 16483 94230 16517
rect 94178 16474 94230 16483
rect 94178 16181 94230 16190
rect 94178 16147 94187 16181
rect 94187 16147 94221 16181
rect 94221 16147 94230 16181
rect 94178 16138 94230 16147
rect 94178 15845 94230 15854
rect 94178 15811 94187 15845
rect 94187 15811 94221 15845
rect 94221 15811 94230 15845
rect 94178 15802 94230 15811
rect 94178 15509 94230 15518
rect 94178 15475 94187 15509
rect 94187 15475 94221 15509
rect 94221 15475 94230 15509
rect 94178 15466 94230 15475
rect 94178 15173 94230 15182
rect 94178 15139 94187 15173
rect 94187 15139 94221 15173
rect 94221 15139 94230 15173
rect 94178 15130 94230 15139
rect 81565 14931 81617 14983
rect 94178 14837 94230 14846
rect 94178 14803 94187 14837
rect 94187 14803 94221 14837
rect 94221 14803 94230 14837
rect 94178 14794 94230 14803
rect 94178 14501 94230 14510
rect 94178 14467 94187 14501
rect 94187 14467 94221 14501
rect 94221 14467 94230 14501
rect 94178 14458 94230 14467
rect 94178 14165 94230 14174
rect 94178 14131 94187 14165
rect 94187 14131 94221 14165
rect 94221 14131 94230 14165
rect 94178 14122 94230 14131
rect 94178 13829 94230 13838
rect 94178 13795 94187 13829
rect 94187 13795 94221 13829
rect 94221 13795 94230 13829
rect 94178 13786 94230 13795
rect 81485 13661 81537 13713
rect 94178 13493 94230 13502
rect 94178 13459 94187 13493
rect 94187 13459 94221 13493
rect 94221 13459 94230 13493
rect 94178 13450 94230 13459
rect 94178 13157 94230 13166
rect 94178 13123 94187 13157
rect 94187 13123 94221 13157
rect 94221 13123 94230 13157
rect 94178 13114 94230 13123
rect 94178 12821 94230 12830
rect 94178 12787 94187 12821
rect 94187 12787 94221 12821
rect 94221 12787 94230 12821
rect 94178 12778 94230 12787
rect 94178 12485 94230 12494
rect 94178 12451 94187 12485
rect 94187 12451 94221 12485
rect 94221 12451 94230 12485
rect 94178 12442 94230 12451
rect 81405 12103 81457 12155
rect 94178 12149 94230 12158
rect 94178 12115 94187 12149
rect 94187 12115 94221 12149
rect 94221 12115 94230 12149
rect 94178 12106 94230 12115
rect 94178 11813 94230 11822
rect 94178 11779 94187 11813
rect 94187 11779 94221 11813
rect 94221 11779 94230 11813
rect 94178 11770 94230 11779
rect 94178 11477 94230 11486
rect 94178 11443 94187 11477
rect 94187 11443 94221 11477
rect 94221 11443 94230 11477
rect 94178 11434 94230 11443
rect 94178 11141 94230 11150
rect 94178 11107 94187 11141
rect 94187 11107 94221 11141
rect 94221 11107 94230 11141
rect 94178 11098 94230 11107
rect 81325 10833 81377 10885
rect 94178 10805 94230 10814
rect 94178 10771 94187 10805
rect 94187 10771 94221 10805
rect 94221 10771 94230 10805
rect 94178 10762 94230 10771
rect 94178 10469 94230 10478
rect 94178 10435 94187 10469
rect 94187 10435 94221 10469
rect 94221 10435 94230 10469
rect 94178 10426 94230 10435
rect 94178 10133 94230 10142
rect 94178 10099 94187 10133
rect 94187 10099 94221 10133
rect 94221 10099 94230 10133
rect 94178 10090 94230 10099
rect 94178 9797 94230 9806
rect 94178 9763 94187 9797
rect 94187 9763 94221 9797
rect 94221 9763 94230 9797
rect 94178 9754 94230 9763
rect 94178 9461 94230 9470
rect 94178 9427 94187 9461
rect 94187 9427 94221 9461
rect 94221 9427 94230 9461
rect 94178 9418 94230 9427
rect 81245 9275 81297 9327
rect 94178 9125 94230 9134
rect 94178 9091 94187 9125
rect 94187 9091 94221 9125
rect 94221 9091 94230 9125
rect 94178 9082 94230 9091
rect 94178 8789 94230 8798
rect 94178 8755 94187 8789
rect 94187 8755 94221 8789
rect 94221 8755 94230 8789
rect 94178 8746 94230 8755
rect 94178 8453 94230 8462
rect 94178 8419 94187 8453
rect 94187 8419 94221 8453
rect 94221 8419 94230 8453
rect 94178 8410 94230 8419
rect 94178 8117 94230 8126
rect 94178 8083 94187 8117
rect 94187 8083 94221 8117
rect 94221 8083 94230 8117
rect 94178 8074 94230 8083
rect 81165 8005 81217 8057
rect 1820 7781 1872 7790
rect 1820 7747 1829 7781
rect 1829 7747 1863 7781
rect 1863 7747 1872 7781
rect 1820 7738 1872 7747
rect 94178 7781 94230 7790
rect 94178 7747 94187 7781
rect 94187 7747 94221 7781
rect 94221 7747 94230 7781
rect 94178 7738 94230 7747
rect 1820 7445 1872 7454
rect 1820 7411 1829 7445
rect 1829 7411 1863 7445
rect 1863 7411 1872 7445
rect 1820 7402 1872 7411
rect 94178 7445 94230 7454
rect 94178 7411 94187 7445
rect 94187 7411 94221 7445
rect 94221 7411 94230 7445
rect 94178 7402 94230 7411
rect 1820 7109 1872 7118
rect 1820 7075 1829 7109
rect 1829 7075 1863 7109
rect 1863 7075 1872 7109
rect 1820 7066 1872 7075
rect 94178 7109 94230 7118
rect 94178 7075 94187 7109
rect 94187 7075 94221 7109
rect 94221 7075 94230 7109
rect 94178 7066 94230 7075
rect 1820 6773 1872 6782
rect 1820 6739 1829 6773
rect 1829 6739 1863 6773
rect 1863 6739 1872 6773
rect 1820 6730 1872 6739
rect 94178 6773 94230 6782
rect 94178 6739 94187 6773
rect 94187 6739 94221 6773
rect 94221 6739 94230 6773
rect 94178 6730 94230 6739
rect 1820 6437 1872 6446
rect 1820 6403 1829 6437
rect 1829 6403 1863 6437
rect 1863 6403 1872 6437
rect 1820 6394 1872 6403
rect 94178 6437 94230 6446
rect 94178 6403 94187 6437
rect 94187 6403 94221 6437
rect 94221 6403 94230 6437
rect 94178 6394 94230 6403
rect 1820 6101 1872 6110
rect 1820 6067 1829 6101
rect 1829 6067 1863 6101
rect 1863 6067 1872 6101
rect 1820 6058 1872 6067
rect 94178 6101 94230 6110
rect 94178 6067 94187 6101
rect 94187 6067 94221 6101
rect 94221 6067 94230 6101
rect 94178 6058 94230 6067
rect 1820 5765 1872 5774
rect 1820 5731 1829 5765
rect 1829 5731 1863 5765
rect 1863 5731 1872 5765
rect 1820 5722 1872 5731
rect 94178 5765 94230 5774
rect 94178 5731 94187 5765
rect 94187 5731 94221 5765
rect 94221 5731 94230 5765
rect 94178 5722 94230 5731
rect 1820 5429 1872 5438
rect 1820 5395 1829 5429
rect 1829 5395 1863 5429
rect 1863 5395 1872 5429
rect 1820 5386 1872 5395
rect 94178 5429 94230 5438
rect 94178 5395 94187 5429
rect 94187 5395 94221 5429
rect 94221 5395 94230 5429
rect 94178 5386 94230 5395
rect 1820 5093 1872 5102
rect 1820 5059 1829 5093
rect 1829 5059 1863 5093
rect 1863 5059 1872 5093
rect 1820 5050 1872 5059
rect 94178 5093 94230 5102
rect 94178 5059 94187 5093
rect 94187 5059 94221 5093
rect 94221 5059 94230 5093
rect 94178 5050 94230 5059
rect 1820 4757 1872 4766
rect 1820 4723 1829 4757
rect 1829 4723 1863 4757
rect 1863 4723 1872 4757
rect 1820 4714 1872 4723
rect 94178 4757 94230 4766
rect 94178 4723 94187 4757
rect 94187 4723 94221 4757
rect 94221 4723 94230 4757
rect 94178 4714 94230 4723
rect 1820 4421 1872 4430
rect 1820 4387 1829 4421
rect 1829 4387 1863 4421
rect 1863 4387 1872 4421
rect 1820 4378 1872 4387
rect 94178 4421 94230 4430
rect 94178 4387 94187 4421
rect 94187 4387 94221 4421
rect 94221 4387 94230 4421
rect 94178 4378 94230 4387
rect 1820 4085 1872 4094
rect 1820 4051 1829 4085
rect 1829 4051 1863 4085
rect 1863 4051 1872 4085
rect 1820 4042 1872 4051
rect 94178 4085 94230 4094
rect 94178 4051 94187 4085
rect 94187 4051 94221 4085
rect 94221 4051 94230 4085
rect 94178 4042 94230 4051
rect 1820 3749 1872 3758
rect 1820 3715 1829 3749
rect 1829 3715 1863 3749
rect 1863 3715 1872 3749
rect 1820 3706 1872 3715
rect 94178 3749 94230 3758
rect 94178 3715 94187 3749
rect 94187 3715 94221 3749
rect 94221 3715 94230 3749
rect 94178 3706 94230 3715
rect 1820 3413 1872 3422
rect 1820 3379 1829 3413
rect 1829 3379 1863 3413
rect 1863 3379 1872 3413
rect 1820 3370 1872 3379
rect 94178 3413 94230 3422
rect 94178 3379 94187 3413
rect 94187 3379 94221 3413
rect 94221 3379 94230 3413
rect 94178 3370 94230 3379
rect 1820 3077 1872 3086
rect 1820 3043 1829 3077
rect 1829 3043 1863 3077
rect 1863 3043 1872 3077
rect 1820 3034 1872 3043
rect 94178 3077 94230 3086
rect 94178 3043 94187 3077
rect 94187 3043 94221 3077
rect 94221 3043 94230 3077
rect 94178 3034 94230 3043
rect 1820 2741 1872 2750
rect 1820 2707 1829 2741
rect 1829 2707 1863 2741
rect 1863 2707 1872 2741
rect 1820 2698 1872 2707
rect 94178 2741 94230 2750
rect 94178 2707 94187 2741
rect 94187 2707 94221 2741
rect 94221 2707 94230 2741
rect 94178 2698 94230 2707
rect 1820 2405 1872 2414
rect 1820 2371 1829 2405
rect 1829 2371 1863 2405
rect 1863 2371 1872 2405
rect 1820 2362 1872 2371
rect 94178 2405 94230 2414
rect 94178 2371 94187 2405
rect 94187 2371 94221 2405
rect 94221 2371 94230 2405
rect 94178 2362 94230 2371
rect 1820 2069 1872 2078
rect 1820 2035 1829 2069
rect 1829 2035 1863 2069
rect 1863 2035 1872 2069
rect 1820 2026 1872 2035
rect 94178 2069 94230 2078
rect 94178 2035 94187 2069
rect 94187 2035 94221 2069
rect 94221 2035 94230 2069
rect 94178 2026 94230 2035
rect 2156 1733 2208 1742
rect 3836 1733 3888 1742
rect 5516 1733 5568 1742
rect 7196 1733 7248 1742
rect 8876 1733 8928 1742
rect 10556 1733 10608 1742
rect 12236 1733 12288 1742
rect 13916 1733 13968 1742
rect 15596 1733 15648 1742
rect 17276 1733 17328 1742
rect 18956 1733 19008 1742
rect 20636 1733 20688 1742
rect 22316 1733 22368 1742
rect 23996 1733 24048 1742
rect 25676 1733 25728 1742
rect 27356 1733 27408 1742
rect 29036 1733 29088 1742
rect 30716 1733 30768 1742
rect 32396 1733 32448 1742
rect 34076 1733 34128 1742
rect 35756 1733 35808 1742
rect 37436 1733 37488 1742
rect 39116 1733 39168 1742
rect 40796 1733 40848 1742
rect 42476 1733 42528 1742
rect 44156 1733 44208 1742
rect 45836 1733 45888 1742
rect 47516 1733 47568 1742
rect 49196 1733 49248 1742
rect 50876 1733 50928 1742
rect 52556 1733 52608 1742
rect 54236 1733 54288 1742
rect 55916 1733 55968 1742
rect 57596 1733 57648 1742
rect 59276 1733 59328 1742
rect 60956 1733 61008 1742
rect 62636 1733 62688 1742
rect 64316 1733 64368 1742
rect 65996 1733 66048 1742
rect 67676 1733 67728 1742
rect 69356 1733 69408 1742
rect 71036 1733 71088 1742
rect 72716 1733 72768 1742
rect 74396 1733 74448 1742
rect 76076 1733 76128 1742
rect 77756 1733 77808 1742
rect 79436 1733 79488 1742
rect 81116 1733 81168 1742
rect 82796 1733 82848 1742
rect 84476 1733 84528 1742
rect 86156 1733 86208 1742
rect 87836 1733 87888 1742
rect 89516 1733 89568 1742
rect 91196 1733 91248 1742
rect 92876 1733 92928 1742
rect 2156 1699 2165 1733
rect 2165 1699 2199 1733
rect 2199 1699 2208 1733
rect 3836 1699 3845 1733
rect 3845 1699 3879 1733
rect 3879 1699 3888 1733
rect 5516 1699 5525 1733
rect 5525 1699 5559 1733
rect 5559 1699 5568 1733
rect 7196 1699 7205 1733
rect 7205 1699 7239 1733
rect 7239 1699 7248 1733
rect 8876 1699 8885 1733
rect 8885 1699 8919 1733
rect 8919 1699 8928 1733
rect 10556 1699 10565 1733
rect 10565 1699 10599 1733
rect 10599 1699 10608 1733
rect 12236 1699 12245 1733
rect 12245 1699 12279 1733
rect 12279 1699 12288 1733
rect 13916 1699 13925 1733
rect 13925 1699 13959 1733
rect 13959 1699 13968 1733
rect 15596 1699 15605 1733
rect 15605 1699 15639 1733
rect 15639 1699 15648 1733
rect 17276 1699 17285 1733
rect 17285 1699 17319 1733
rect 17319 1699 17328 1733
rect 18956 1699 18965 1733
rect 18965 1699 18999 1733
rect 18999 1699 19008 1733
rect 20636 1699 20645 1733
rect 20645 1699 20679 1733
rect 20679 1699 20688 1733
rect 22316 1699 22325 1733
rect 22325 1699 22359 1733
rect 22359 1699 22368 1733
rect 23996 1699 24005 1733
rect 24005 1699 24039 1733
rect 24039 1699 24048 1733
rect 25676 1699 25685 1733
rect 25685 1699 25719 1733
rect 25719 1699 25728 1733
rect 27356 1699 27365 1733
rect 27365 1699 27399 1733
rect 27399 1699 27408 1733
rect 29036 1699 29045 1733
rect 29045 1699 29079 1733
rect 29079 1699 29088 1733
rect 30716 1699 30725 1733
rect 30725 1699 30759 1733
rect 30759 1699 30768 1733
rect 32396 1699 32405 1733
rect 32405 1699 32439 1733
rect 32439 1699 32448 1733
rect 34076 1699 34085 1733
rect 34085 1699 34119 1733
rect 34119 1699 34128 1733
rect 35756 1699 35765 1733
rect 35765 1699 35799 1733
rect 35799 1699 35808 1733
rect 37436 1699 37445 1733
rect 37445 1699 37479 1733
rect 37479 1699 37488 1733
rect 39116 1699 39125 1733
rect 39125 1699 39159 1733
rect 39159 1699 39168 1733
rect 40796 1699 40805 1733
rect 40805 1699 40839 1733
rect 40839 1699 40848 1733
rect 42476 1699 42485 1733
rect 42485 1699 42519 1733
rect 42519 1699 42528 1733
rect 44156 1699 44165 1733
rect 44165 1699 44199 1733
rect 44199 1699 44208 1733
rect 45836 1699 45845 1733
rect 45845 1699 45879 1733
rect 45879 1699 45888 1733
rect 47516 1699 47525 1733
rect 47525 1699 47559 1733
rect 47559 1699 47568 1733
rect 49196 1699 49205 1733
rect 49205 1699 49239 1733
rect 49239 1699 49248 1733
rect 50876 1699 50885 1733
rect 50885 1699 50919 1733
rect 50919 1699 50928 1733
rect 52556 1699 52565 1733
rect 52565 1699 52599 1733
rect 52599 1699 52608 1733
rect 54236 1699 54245 1733
rect 54245 1699 54279 1733
rect 54279 1699 54288 1733
rect 55916 1699 55925 1733
rect 55925 1699 55959 1733
rect 55959 1699 55968 1733
rect 57596 1699 57605 1733
rect 57605 1699 57639 1733
rect 57639 1699 57648 1733
rect 59276 1699 59285 1733
rect 59285 1699 59319 1733
rect 59319 1699 59328 1733
rect 60956 1699 60965 1733
rect 60965 1699 60999 1733
rect 60999 1699 61008 1733
rect 62636 1699 62645 1733
rect 62645 1699 62679 1733
rect 62679 1699 62688 1733
rect 64316 1699 64325 1733
rect 64325 1699 64359 1733
rect 64359 1699 64368 1733
rect 65996 1699 66005 1733
rect 66005 1699 66039 1733
rect 66039 1699 66048 1733
rect 67676 1699 67685 1733
rect 67685 1699 67719 1733
rect 67719 1699 67728 1733
rect 69356 1699 69365 1733
rect 69365 1699 69399 1733
rect 69399 1699 69408 1733
rect 71036 1699 71045 1733
rect 71045 1699 71079 1733
rect 71079 1699 71088 1733
rect 72716 1699 72725 1733
rect 72725 1699 72759 1733
rect 72759 1699 72768 1733
rect 74396 1699 74405 1733
rect 74405 1699 74439 1733
rect 74439 1699 74448 1733
rect 76076 1699 76085 1733
rect 76085 1699 76119 1733
rect 76119 1699 76128 1733
rect 77756 1699 77765 1733
rect 77765 1699 77799 1733
rect 77799 1699 77808 1733
rect 79436 1699 79445 1733
rect 79445 1699 79479 1733
rect 79479 1699 79488 1733
rect 81116 1699 81125 1733
rect 81125 1699 81159 1733
rect 81159 1699 81168 1733
rect 82796 1699 82805 1733
rect 82805 1699 82839 1733
rect 82839 1699 82848 1733
rect 84476 1699 84485 1733
rect 84485 1699 84519 1733
rect 84519 1699 84528 1733
rect 86156 1699 86165 1733
rect 86165 1699 86199 1733
rect 86199 1699 86208 1733
rect 87836 1699 87845 1733
rect 87845 1699 87879 1733
rect 87879 1699 87888 1733
rect 89516 1699 89525 1733
rect 89525 1699 89559 1733
rect 89559 1699 89568 1733
rect 91196 1699 91205 1733
rect 91205 1699 91239 1733
rect 91239 1699 91248 1733
rect 92876 1699 92885 1733
rect 92885 1699 92919 1733
rect 92919 1699 92928 1733
rect 2156 1690 2208 1699
rect 3836 1690 3888 1699
rect 5516 1690 5568 1699
rect 7196 1690 7248 1699
rect 8876 1690 8928 1699
rect 10556 1690 10608 1699
rect 12236 1690 12288 1699
rect 13916 1690 13968 1699
rect 15596 1690 15648 1699
rect 17276 1690 17328 1699
rect 18956 1690 19008 1699
rect 20636 1690 20688 1699
rect 22316 1690 22368 1699
rect 23996 1690 24048 1699
rect 25676 1690 25728 1699
rect 27356 1690 27408 1699
rect 29036 1690 29088 1699
rect 30716 1690 30768 1699
rect 32396 1690 32448 1699
rect 34076 1690 34128 1699
rect 35756 1690 35808 1699
rect 37436 1690 37488 1699
rect 39116 1690 39168 1699
rect 40796 1690 40848 1699
rect 42476 1690 42528 1699
rect 44156 1690 44208 1699
rect 45836 1690 45888 1699
rect 47516 1690 47568 1699
rect 49196 1690 49248 1699
rect 50876 1690 50928 1699
rect 52556 1690 52608 1699
rect 54236 1690 54288 1699
rect 55916 1690 55968 1699
rect 57596 1690 57648 1699
rect 59276 1690 59328 1699
rect 60956 1690 61008 1699
rect 62636 1690 62688 1699
rect 64316 1690 64368 1699
rect 65996 1690 66048 1699
rect 67676 1690 67728 1699
rect 69356 1690 69408 1699
rect 71036 1690 71088 1699
rect 72716 1690 72768 1699
rect 74396 1690 74448 1699
rect 76076 1690 76128 1699
rect 77756 1690 77808 1699
rect 79436 1690 79488 1699
rect 81116 1690 81168 1699
rect 82796 1690 82848 1699
rect 84476 1690 84528 1699
rect 86156 1690 86208 1699
rect 87836 1690 87888 1699
rect 89516 1690 89568 1699
rect 91196 1690 91248 1699
rect 92876 1690 92928 1699
<< metal2 >>
rect 1734 77342 1958 77892
rect 2154 77808 2210 77817
rect 2154 77743 2210 77752
rect 3834 77808 3890 77817
rect 3834 77743 3890 77752
rect 5514 77808 5570 77817
rect 5514 77743 5570 77752
rect 7194 77808 7250 77817
rect 7194 77743 7250 77752
rect 8874 77808 8930 77817
rect 8874 77743 8930 77752
rect 10554 77808 10610 77817
rect 10554 77743 10610 77752
rect 12234 77808 12290 77817
rect 12234 77743 12290 77752
rect 13914 77808 13970 77817
rect 13914 77743 13970 77752
rect 15594 77808 15650 77817
rect 15594 77743 15650 77752
rect 17274 77808 17330 77817
rect 17274 77743 17330 77752
rect 18954 77808 19010 77817
rect 18954 77743 19010 77752
rect 20634 77808 20690 77817
rect 20634 77743 20690 77752
rect 22314 77808 22370 77817
rect 22314 77743 22370 77752
rect 23994 77808 24050 77817
rect 23994 77743 24050 77752
rect 25674 77808 25730 77817
rect 25674 77743 25730 77752
rect 27354 77808 27410 77817
rect 27354 77743 27410 77752
rect 29034 77808 29090 77817
rect 29034 77743 29090 77752
rect 30714 77808 30770 77817
rect 30714 77743 30770 77752
rect 32394 77808 32450 77817
rect 32394 77743 32450 77752
rect 34074 77808 34130 77817
rect 34074 77743 34130 77752
rect 35754 77808 35810 77817
rect 35754 77743 35810 77752
rect 37434 77808 37490 77817
rect 37434 77743 37490 77752
rect 39114 77808 39170 77817
rect 39114 77743 39170 77752
rect 40794 77808 40850 77817
rect 40794 77743 40850 77752
rect 42474 77808 42530 77817
rect 42474 77743 42530 77752
rect 44154 77808 44210 77817
rect 44154 77743 44210 77752
rect 45834 77808 45890 77817
rect 45834 77743 45890 77752
rect 47514 77808 47570 77817
rect 47514 77743 47570 77752
rect 49194 77808 49250 77817
rect 49194 77743 49250 77752
rect 50874 77808 50930 77817
rect 50874 77743 50930 77752
rect 52554 77808 52610 77817
rect 52554 77743 52610 77752
rect 54234 77808 54290 77817
rect 54234 77743 54290 77752
rect 55914 77808 55970 77817
rect 55914 77743 55970 77752
rect 57594 77808 57650 77817
rect 57594 77743 57650 77752
rect 59274 77808 59330 77817
rect 59274 77743 59330 77752
rect 60954 77808 61010 77817
rect 60954 77743 61010 77752
rect 62634 77808 62690 77817
rect 62634 77743 62690 77752
rect 64314 77808 64370 77817
rect 64314 77743 64370 77752
rect 65994 77808 66050 77817
rect 65994 77743 66050 77752
rect 67674 77808 67730 77817
rect 67674 77743 67730 77752
rect 69354 77808 69410 77817
rect 69354 77743 69410 77752
rect 71034 77808 71090 77817
rect 71034 77743 71090 77752
rect 72714 77808 72770 77817
rect 72714 77743 72770 77752
rect 74394 77808 74450 77817
rect 74394 77743 74450 77752
rect 76074 77808 76130 77817
rect 76074 77743 76130 77752
rect 77754 77808 77810 77817
rect 77754 77743 77810 77752
rect 79434 77808 79490 77817
rect 79434 77743 79490 77752
rect 81114 77808 81170 77817
rect 81114 77743 81170 77752
rect 82794 77808 82850 77817
rect 82794 77743 82850 77752
rect 84474 77808 84530 77817
rect 84474 77743 84530 77752
rect 86154 77808 86210 77817
rect 86154 77743 86210 77752
rect 87834 77808 87890 77817
rect 87834 77743 87890 77752
rect 89514 77808 89570 77817
rect 89514 77743 89570 77752
rect 91194 77808 91250 77817
rect 91194 77743 91250 77752
rect 92874 77808 92930 77817
rect 92874 77743 92930 77752
rect 1734 77290 1820 77342
rect 1872 77290 1958 77342
rect 1734 77006 1958 77290
rect 1734 76954 1820 77006
rect 1872 76954 1958 77006
rect 1734 76670 1958 76954
rect 1734 76618 1820 76670
rect 1872 76618 1958 76670
rect 1734 76334 1958 76618
rect 94092 77342 94316 77892
rect 94092 77290 94178 77342
rect 94230 77290 94316 77342
rect 94092 77006 94316 77290
rect 94092 76954 94178 77006
rect 94230 76954 94316 77006
rect 94092 76670 94316 76954
rect 94092 76618 94178 76670
rect 94230 76618 94316 76670
rect 93216 76572 93272 76581
rect 93216 76507 93272 76516
rect 90079 76467 90135 76476
rect 1734 76282 1820 76334
rect 1872 76282 1958 76334
rect 1734 76000 1958 76282
rect 81858 76387 81956 76415
rect 90079 76402 90135 76411
rect 81858 76112 81886 76387
rect 94092 76334 94316 76618
rect 94092 76282 94178 76334
rect 94230 76282 94316 76334
rect 81844 76103 81900 76112
rect 81844 76038 81900 76047
rect 1734 75944 1818 76000
rect 1874 75944 1958 76000
rect 1734 75662 1958 75944
rect 79422 75847 79478 75856
rect 79422 75782 79478 75791
rect 1734 75610 1820 75662
rect 1872 75610 1958 75662
rect 1734 75326 1958 75610
rect 1734 75274 1820 75326
rect 1872 75274 1958 75326
rect 1734 74990 1958 75274
rect 1734 74938 1820 74990
rect 1872 74938 1958 74990
rect 1734 74654 1958 74938
rect 1734 74602 1820 74654
rect 1872 74602 1958 74654
rect 1734 74320 1958 74602
rect 1734 74264 1818 74320
rect 1874 74264 1958 74320
rect 1734 73982 1958 74264
rect 28210 74103 28266 74112
rect 28210 74038 28266 74047
rect 29458 74103 29514 74112
rect 29458 74038 29514 74047
rect 30706 74103 30762 74112
rect 30706 74038 30762 74047
rect 31954 74103 32010 74112
rect 31954 74038 32010 74047
rect 33202 74103 33258 74112
rect 33202 74038 33258 74047
rect 34450 74103 34506 74112
rect 34450 74038 34506 74047
rect 35698 74103 35754 74112
rect 35698 74038 35754 74047
rect 36946 74103 37002 74112
rect 36946 74038 37002 74047
rect 38194 74103 38250 74112
rect 38194 74038 38250 74047
rect 39442 74103 39498 74112
rect 39442 74038 39498 74047
rect 40690 74103 40746 74112
rect 40690 74038 40746 74047
rect 41938 74103 41994 74112
rect 41938 74038 41994 74047
rect 43186 74103 43242 74112
rect 43186 74038 43242 74047
rect 44434 74103 44490 74112
rect 44434 74038 44490 74047
rect 45682 74103 45738 74112
rect 45682 74038 45738 74047
rect 46930 74103 46986 74112
rect 46930 74038 46986 74047
rect 48178 74103 48234 74112
rect 48178 74038 48234 74047
rect 49426 74103 49482 74112
rect 49426 74038 49482 74047
rect 50674 74103 50730 74112
rect 50674 74038 50730 74047
rect 51922 74103 51978 74112
rect 51922 74038 51978 74047
rect 53170 74103 53226 74112
rect 53170 74038 53226 74047
rect 54418 74103 54474 74112
rect 54418 74038 54474 74047
rect 55666 74103 55722 74112
rect 55666 74038 55722 74047
rect 56914 74103 56970 74112
rect 56914 74038 56970 74047
rect 58162 74103 58218 74112
rect 58162 74038 58218 74047
rect 59410 74103 59466 74112
rect 59410 74038 59466 74047
rect 60658 74103 60714 74112
rect 60658 74038 60714 74047
rect 61906 74103 61962 74112
rect 61906 74038 61962 74047
rect 63154 74103 63210 74112
rect 63154 74038 63210 74047
rect 64402 74103 64458 74112
rect 64402 74038 64458 74047
rect 65650 74103 65706 74112
rect 65650 74038 65706 74047
rect 66898 74103 66954 74112
rect 66898 74038 66954 74047
rect 1734 73930 1820 73982
rect 1872 73930 1958 73982
rect 1734 73646 1958 73930
rect 1734 73594 1820 73646
rect 1872 73594 1958 73646
rect 1734 73310 1958 73594
rect 1734 73258 1820 73310
rect 1872 73258 1958 73310
rect 1734 72974 1958 73258
rect 1734 72922 1820 72974
rect 1872 72922 1958 72974
rect 1734 72640 1958 72922
rect 1734 72584 1818 72640
rect 1874 72584 1958 72640
rect 1734 72302 1958 72584
rect 1734 72250 1820 72302
rect 1872 72250 1958 72302
rect 1734 71966 1958 72250
rect 69731 72196 69759 74300
rect 69717 72187 69773 72196
rect 69717 72122 69773 72131
rect 1734 71914 1820 71966
rect 1872 71914 1958 71966
rect 1734 71630 1958 71914
rect 1734 71578 1820 71630
rect 1872 71578 1958 71630
rect 1734 71294 1958 71578
rect 1734 71242 1820 71294
rect 1872 71242 1958 71294
rect 1734 70960 1958 71242
rect 1734 70904 1818 70960
rect 1874 70904 1958 70960
rect 1734 70622 1958 70904
rect 69841 70773 69897 70782
rect 69841 70708 69897 70717
rect 1734 70570 1820 70622
rect 1872 70570 1958 70622
rect 1734 70286 1958 70570
rect 1734 70234 1820 70286
rect 1872 70234 1958 70286
rect 1734 69950 1958 70234
rect 1734 69898 1820 69950
rect 1872 69898 1958 69950
rect 1734 69614 1958 69898
rect 1734 69562 1820 69614
rect 1872 69562 1958 69614
rect 1734 69280 1958 69562
rect 1734 69224 1818 69280
rect 1874 69224 1958 69280
rect 1734 68942 1958 69224
rect 1734 68890 1820 68942
rect 1872 68890 1958 68942
rect 1734 68606 1958 68890
rect 1734 68554 1820 68606
rect 1872 68554 1958 68606
rect 1734 68270 1958 68554
rect 69855 68486 69883 70708
rect 73702 69359 73758 69368
rect 73702 69294 73758 69303
rect 1734 68218 1820 68270
rect 1872 68218 1958 68270
rect 1734 67934 1958 68218
rect 73716 68009 73744 69294
rect 1734 67882 1820 67934
rect 1872 67882 1958 67934
rect 1734 67600 1958 67882
rect 1734 67544 1818 67600
rect 1874 67544 1958 67600
rect 1734 67262 1958 67544
rect 1734 67210 1820 67262
rect 1872 67210 1958 67262
rect 1734 66926 1958 67210
rect 1734 66874 1820 66926
rect 1872 66874 1958 66926
rect 1734 66590 1958 66874
rect 1734 66538 1820 66590
rect 1872 66538 1958 66590
rect 1734 66254 1958 66538
rect 1734 66202 1820 66254
rect 1872 66202 1958 66254
rect 1734 65920 1958 66202
rect 1734 65864 1818 65920
rect 1874 65864 1958 65920
rect 1734 65582 1958 65864
rect 1734 65530 1820 65582
rect 1872 65530 1958 65582
rect 1734 65246 1958 65530
rect 1734 65194 1820 65246
rect 1872 65194 1958 65246
rect 1734 64910 1958 65194
rect 1734 64858 1820 64910
rect 1872 64858 1958 64910
rect 1734 64574 1958 64858
rect 1734 64522 1820 64574
rect 1872 64522 1958 64574
rect 1734 64240 1958 64522
rect 1734 64184 1818 64240
rect 1874 64184 1958 64240
rect 1734 63902 1958 64184
rect 1734 63850 1820 63902
rect 1872 63850 1958 63902
rect 1734 63566 1958 63850
rect 1734 63514 1820 63566
rect 1872 63514 1958 63566
rect 1734 63230 1958 63514
rect 1734 63178 1820 63230
rect 1872 63178 1958 63230
rect 1734 62894 1958 63178
rect 1734 62842 1820 62894
rect 1872 62842 1958 62894
rect 1734 62560 1958 62842
rect 1734 62504 1818 62560
rect 1874 62504 1958 62560
rect 1734 62222 1958 62504
rect 1734 62170 1820 62222
rect 1872 62170 1958 62222
rect 1734 61886 1958 62170
rect 1734 61834 1820 61886
rect 1872 61834 1958 61886
rect 1734 61550 1958 61834
rect 1734 61498 1820 61550
rect 1872 61498 1958 61550
rect 1734 61214 1958 61498
rect 1734 61162 1820 61214
rect 1872 61162 1958 61214
rect 1734 60880 1958 61162
rect 1734 60824 1818 60880
rect 1874 60824 1958 60880
rect 1734 60542 1958 60824
rect 1734 60490 1820 60542
rect 1872 60490 1958 60542
rect 1734 60206 1958 60490
rect 1734 60154 1820 60206
rect 1872 60154 1958 60206
rect 1734 59870 1958 60154
rect 1734 59818 1820 59870
rect 1872 59818 1958 59870
rect 1734 59534 1958 59818
rect 1734 59482 1820 59534
rect 1872 59482 1958 59534
rect 1734 59200 1958 59482
rect 1734 59144 1818 59200
rect 1874 59144 1958 59200
rect 1734 58862 1958 59144
rect 1734 58810 1820 58862
rect 1872 58810 1958 58862
rect 1734 58526 1958 58810
rect 1734 58474 1820 58526
rect 1872 58474 1958 58526
rect 1734 58190 1958 58474
rect 1734 58138 1820 58190
rect 1872 58138 1958 58190
rect 1734 57854 1958 58138
rect 1734 57802 1820 57854
rect 1872 57802 1958 57854
rect 1734 57520 1958 57802
rect 1734 57464 1818 57520
rect 1874 57464 1958 57520
rect 1734 57182 1958 57464
rect 1734 57130 1820 57182
rect 1872 57130 1958 57182
rect 1734 56846 1958 57130
rect 1734 56794 1820 56846
rect 1872 56794 1958 56846
rect 1734 56510 1958 56794
rect 1734 56458 1820 56510
rect 1872 56458 1958 56510
rect 1734 56174 1958 56458
rect 1734 56122 1820 56174
rect 1872 56122 1958 56174
rect 1734 55840 1958 56122
rect 1734 55784 1818 55840
rect 1874 55784 1958 55840
rect 1734 55502 1958 55784
rect 1734 55450 1820 55502
rect 1872 55450 1958 55502
rect 1734 55166 1958 55450
rect 1734 55114 1820 55166
rect 1872 55114 1958 55166
rect 1734 54830 1958 55114
rect 1734 54778 1820 54830
rect 1872 54778 1958 54830
rect 1734 54494 1958 54778
rect 1734 54442 1820 54494
rect 1872 54442 1958 54494
rect 1734 54160 1958 54442
rect 1734 54104 1818 54160
rect 1874 54104 1958 54160
rect 1734 53822 1958 54104
rect 1734 53770 1820 53822
rect 1872 53770 1958 53822
rect 1734 53486 1958 53770
rect 1734 53434 1820 53486
rect 1872 53434 1958 53486
rect 1734 53150 1958 53434
rect 1734 53098 1820 53150
rect 1872 53098 1958 53150
rect 1734 52814 1958 53098
rect 1734 52762 1820 52814
rect 1872 52762 1958 52814
rect 1734 52480 1958 52762
rect 1734 52424 1818 52480
rect 1874 52424 1958 52480
rect 1734 52142 1958 52424
rect 1734 52090 1820 52142
rect 1872 52090 1958 52142
rect 1734 51806 1958 52090
rect 1734 51754 1820 51806
rect 1872 51754 1958 51806
rect 1734 51470 1958 51754
rect 1734 51418 1820 51470
rect 1872 51418 1958 51470
rect 1734 51134 1958 51418
rect 1734 51082 1820 51134
rect 1872 51082 1958 51134
rect 1734 50800 1958 51082
rect 1734 50744 1818 50800
rect 1874 50744 1958 50800
rect 1734 50462 1958 50744
rect 1734 50410 1820 50462
rect 1872 50410 1958 50462
rect 1734 50126 1958 50410
rect 1734 50074 1820 50126
rect 1872 50074 1958 50126
rect 1734 49790 1958 50074
rect 1734 49738 1820 49790
rect 1872 49738 1958 49790
rect 1734 49454 1958 49738
rect 1734 49402 1820 49454
rect 1872 49402 1958 49454
rect 1734 49120 1958 49402
rect 1734 49064 1818 49120
rect 1874 49064 1958 49120
rect 1734 48782 1958 49064
rect 1734 48730 1820 48782
rect 1872 48730 1958 48782
rect 1734 48446 1958 48730
rect 1734 48394 1820 48446
rect 1872 48394 1958 48446
rect 1734 48110 1958 48394
rect 1734 48058 1820 48110
rect 1872 48058 1958 48110
rect 1734 47774 1958 48058
rect 1734 47722 1820 47774
rect 1872 47722 1958 47774
rect 1734 47440 1958 47722
rect 1734 47384 1818 47440
rect 1874 47384 1958 47440
rect 1734 47102 1958 47384
rect 1734 47050 1820 47102
rect 1872 47050 1958 47102
rect 1734 46766 1958 47050
rect 1734 46714 1820 46766
rect 1872 46714 1958 46766
rect 1734 46430 1958 46714
rect 1734 46378 1820 46430
rect 1872 46378 1958 46430
rect 1734 46094 1958 46378
rect 1734 46042 1820 46094
rect 1872 46042 1958 46094
rect 1734 45760 1958 46042
rect 1734 45704 1818 45760
rect 1874 45704 1958 45760
rect 1734 45422 1958 45704
rect 1734 45370 1820 45422
rect 1872 45370 1958 45422
rect 1734 45086 1958 45370
rect 1734 45034 1820 45086
rect 1872 45034 1958 45086
rect 1734 44750 1958 45034
rect 1734 44698 1820 44750
rect 1872 44698 1958 44750
rect 1734 44414 1958 44698
rect 1734 44362 1820 44414
rect 1872 44362 1958 44414
rect 1734 44080 1958 44362
rect 1734 44024 1818 44080
rect 1874 44024 1958 44080
rect 1734 43742 1958 44024
rect 1734 43690 1820 43742
rect 1872 43690 1958 43742
rect 1734 43406 1958 43690
rect 1734 43354 1820 43406
rect 1872 43354 1958 43406
rect 1734 43070 1958 43354
rect 1734 43018 1820 43070
rect 1872 43018 1958 43070
rect 1734 42734 1958 43018
rect 1734 42682 1820 42734
rect 1872 42682 1958 42734
rect 1734 42400 1958 42682
rect 1734 42344 1818 42400
rect 1874 42344 1958 42400
rect 1734 42062 1958 42344
rect 1734 42010 1820 42062
rect 1872 42010 1958 42062
rect 1734 41726 1958 42010
rect 1734 41674 1820 41726
rect 1872 41674 1958 41726
rect 1734 41390 1958 41674
rect 1734 41338 1820 41390
rect 1872 41338 1958 41390
rect 1734 41054 1958 41338
rect 1734 41002 1820 41054
rect 1872 41002 1958 41054
rect 1734 40720 1958 41002
rect 1734 40664 1818 40720
rect 1874 40664 1958 40720
rect 1734 40382 1958 40664
rect 1734 40330 1820 40382
rect 1872 40330 1958 40382
rect 1734 40046 1958 40330
rect 1734 39994 1820 40046
rect 1872 39994 1958 40046
rect 1734 39710 1958 39994
rect 1734 39658 1820 39710
rect 1872 39658 1958 39710
rect 1734 39374 1958 39658
rect 1734 39322 1820 39374
rect 1872 39322 1958 39374
rect 1734 39040 1958 39322
rect 1734 38984 1818 39040
rect 1874 38984 1958 39040
rect 1734 38702 1958 38984
rect 1734 38650 1820 38702
rect 1872 38650 1958 38702
rect 1734 38366 1958 38650
rect 1734 38314 1820 38366
rect 1872 38314 1958 38366
rect 1734 38030 1958 38314
rect 1734 37978 1820 38030
rect 1872 37978 1958 38030
rect 1734 37694 1958 37978
rect 1734 37642 1820 37694
rect 1872 37642 1958 37694
rect 1734 37360 1958 37642
rect 1734 37304 1818 37360
rect 1874 37304 1958 37360
rect 1734 37022 1958 37304
rect 1734 36970 1820 37022
rect 1872 36970 1958 37022
rect 1734 36686 1958 36970
rect 1734 36634 1820 36686
rect 1872 36634 1958 36686
rect 1734 36350 1958 36634
rect 1734 36298 1820 36350
rect 1872 36298 1958 36350
rect 1734 36014 1958 36298
rect 1734 35962 1820 36014
rect 1872 35962 1958 36014
rect 1734 35680 1958 35962
rect 1734 35624 1818 35680
rect 1874 35624 1958 35680
rect 1734 35342 1958 35624
rect 1734 35290 1820 35342
rect 1872 35290 1958 35342
rect 1734 35006 1958 35290
rect 1734 34954 1820 35006
rect 1872 34954 1958 35006
rect 1734 34670 1958 34954
rect 1734 34618 1820 34670
rect 1872 34618 1958 34670
rect 1734 34334 1958 34618
rect 1734 34282 1820 34334
rect 1872 34282 1958 34334
rect 1734 34000 1958 34282
rect 14205 34197 14261 34206
rect 13260 34126 13316 34135
rect 14205 34132 14261 34141
rect 14939 34197 14995 34206
rect 14939 34132 14995 34141
rect 13260 34061 13316 34070
rect 1734 33944 1818 34000
rect 1874 33944 1958 34000
rect 1734 33662 1958 33944
rect 1734 33610 1820 33662
rect 1872 33610 1958 33662
rect 1734 33326 1958 33610
rect 1734 33274 1820 33326
rect 1872 33274 1958 33326
rect 1734 32990 1958 33274
rect 1734 32938 1820 32990
rect 1872 32938 1958 32990
rect 1734 32654 1958 32938
rect 13260 32998 13316 33007
rect 13260 32933 13316 32942
rect 14205 32927 14261 32936
rect 14205 32862 14261 32871
rect 14859 32927 14915 32936
rect 14859 32862 14915 32871
rect 1734 32602 1820 32654
rect 1872 32602 1958 32654
rect 1734 32320 1958 32602
rect 1734 32264 1818 32320
rect 1874 32264 1958 32320
rect 1734 31982 1958 32264
rect 1734 31930 1820 31982
rect 1872 31930 1958 31982
rect 1734 31646 1958 31930
rect 1734 31594 1820 31646
rect 1872 31594 1958 31646
rect 1734 31310 1958 31594
rect 1734 31258 1820 31310
rect 1872 31258 1958 31310
rect 14205 31369 14261 31378
rect 1734 30974 1958 31258
rect 13260 31298 13316 31307
rect 14205 31304 14261 31313
rect 14779 31369 14835 31378
rect 14779 31304 14835 31313
rect 13260 31233 13316 31242
rect 1734 30922 1820 30974
rect 1872 30922 1958 30974
rect 1734 30640 1958 30922
rect 1734 30584 1818 30640
rect 1874 30584 1958 30640
rect 1734 30302 1958 30584
rect 1734 30250 1820 30302
rect 1872 30250 1958 30302
rect 1734 29966 1958 30250
rect 13260 30170 13316 30179
rect 13260 30105 13316 30114
rect 14205 30099 14261 30108
rect 14205 30034 14261 30043
rect 14699 30099 14755 30108
rect 14699 30034 14755 30043
rect 1734 29914 1820 29966
rect 1872 29914 1958 29966
rect 1734 29630 1958 29914
rect 1734 29578 1820 29630
rect 1872 29578 1958 29630
rect 1734 29294 1958 29578
rect 1734 29242 1820 29294
rect 1872 29242 1958 29294
rect 1734 28960 1958 29242
rect 1734 28904 1818 28960
rect 1874 28904 1958 28960
rect 1734 28622 1958 28904
rect 1734 28570 1820 28622
rect 1872 28570 1958 28622
rect 1734 28286 1958 28570
rect 14205 28541 14261 28550
rect 13260 28470 13316 28479
rect 14205 28476 14261 28485
rect 14619 28541 14675 28550
rect 14619 28476 14675 28485
rect 13260 28405 13316 28414
rect 1734 28234 1820 28286
rect 1872 28234 1958 28286
rect 1734 27950 1958 28234
rect 1734 27898 1820 27950
rect 1872 27898 1958 27950
rect 1734 27614 1958 27898
rect 1734 27562 1820 27614
rect 1872 27562 1958 27614
rect 1734 27280 1958 27562
rect 1734 27224 1818 27280
rect 1874 27224 1958 27280
rect 13260 27342 13316 27351
rect 13260 27277 13316 27286
rect 1734 26942 1958 27224
rect 14205 27271 14261 27280
rect 14205 27206 14261 27215
rect 14539 27271 14595 27280
rect 14539 27206 14595 27215
rect 1734 26890 1820 26942
rect 1872 26890 1958 26942
rect 1734 26606 1958 26890
rect 1734 26554 1820 26606
rect 1872 26554 1958 26606
rect 1734 26270 1958 26554
rect 1734 26218 1820 26270
rect 1872 26218 1958 26270
rect 1734 25934 1958 26218
rect 1734 25882 1820 25934
rect 1872 25882 1958 25934
rect 1734 25600 1958 25882
rect 14205 25713 14261 25722
rect 1734 25544 1818 25600
rect 1874 25544 1958 25600
rect 13260 25642 13316 25651
rect 14205 25648 14261 25657
rect 14459 25713 14515 25722
rect 14459 25648 14515 25657
rect 13260 25577 13316 25586
rect 1734 25262 1958 25544
rect 14342 25386 14398 25395
rect 14342 25321 14398 25330
rect 1734 25210 1820 25262
rect 1872 25210 1958 25262
rect 1734 24926 1958 25210
rect 1734 24874 1820 24926
rect 1872 24874 1958 24926
rect 1734 24590 1958 24874
rect 1734 24538 1820 24590
rect 1872 24538 1958 24590
rect 1734 24254 1958 24538
rect 1734 24202 1820 24254
rect 1872 24202 1958 24254
rect 1734 23920 1958 24202
rect 1734 23864 1818 23920
rect 1874 23864 1958 23920
rect 1734 23582 1958 23864
rect 1734 23530 1820 23582
rect 1872 23530 1958 23582
rect 1734 23246 1958 23530
rect 1734 23194 1820 23246
rect 1872 23194 1958 23246
rect 1734 22910 1958 23194
rect 1734 22858 1820 22910
rect 1872 22858 1958 22910
rect 1734 22574 1958 22858
rect 2565 22665 2621 22674
rect 2565 22600 2621 22609
rect 1734 22522 1820 22574
rect 1872 22522 1958 22574
rect 1734 22240 1958 22522
rect 1734 22184 1818 22240
rect 1874 22184 1958 22240
rect 1734 21902 1958 22184
rect 1734 21850 1820 21902
rect 1872 21850 1958 21902
rect 1734 21566 1958 21850
rect 1734 21514 1820 21566
rect 1872 21514 1958 21566
rect 1734 21230 1958 21514
rect 1734 21178 1820 21230
rect 1872 21178 1958 21230
rect 1734 20894 1958 21178
rect 1734 20842 1820 20894
rect 1872 20842 1958 20894
rect 1734 20560 1958 20842
rect 1734 20504 1818 20560
rect 1874 20504 1958 20560
rect 1734 20222 1958 20504
rect 1734 20170 1820 20222
rect 1872 20170 1958 20222
rect 1734 19886 1958 20170
rect 1734 19834 1820 19886
rect 1872 19834 1958 19886
rect 1734 19550 1958 19834
rect 1734 19498 1820 19550
rect 1872 19498 1958 19550
rect 1734 19214 1958 19498
rect 1734 19162 1820 19214
rect 1872 19162 1958 19214
rect 1734 18880 1958 19162
rect 1734 18824 1818 18880
rect 1874 18824 1958 18880
rect 1734 18542 1958 18824
rect 1734 18490 1820 18542
rect 1872 18490 1958 18542
rect 1734 18206 1958 18490
rect 1734 18154 1820 18206
rect 1872 18154 1958 18206
rect 1734 17870 1958 18154
rect 1734 17818 1820 17870
rect 1872 17818 1958 17870
rect 1734 17534 1958 17818
rect 1734 17482 1820 17534
rect 1872 17482 1958 17534
rect 1734 17200 1958 17482
rect 1734 17144 1818 17200
rect 1874 17144 1958 17200
rect 1734 16862 1958 17144
rect 1734 16810 1820 16862
rect 1872 16810 1958 16862
rect 1734 16526 1958 16810
rect 1734 16474 1820 16526
rect 1872 16474 1958 16526
rect 1734 16190 1958 16474
rect 1734 16138 1820 16190
rect 1872 16138 1958 16190
rect 1734 15854 1958 16138
rect 1734 15802 1820 15854
rect 1872 15802 1958 15854
rect 1734 15520 1958 15802
rect 1734 15464 1818 15520
rect 1874 15464 1958 15520
rect 14258 15557 14314 15566
rect 14258 15492 14314 15501
rect 1734 15182 1958 15464
rect 1734 15130 1820 15182
rect 1872 15130 1958 15182
rect 1734 14846 1958 15130
rect 1734 14794 1820 14846
rect 1872 14794 1958 14846
rect 1734 14510 1958 14794
rect 1734 14458 1820 14510
rect 1872 14458 1958 14510
rect 1734 14174 1958 14458
rect 1734 14122 1820 14174
rect 1872 14122 1958 14174
rect 1734 13840 1958 14122
rect 1734 13784 1818 13840
rect 1874 13784 1958 13840
rect 1734 13502 1958 13784
rect 1734 13450 1820 13502
rect 1872 13450 1958 13502
rect 1734 13166 1958 13450
rect 1734 13114 1820 13166
rect 1872 13114 1958 13166
rect 1734 12830 1958 13114
rect 1734 12778 1820 12830
rect 1872 12778 1958 12830
rect 1734 12494 1958 12778
rect 14258 12729 14314 12738
rect 14258 12664 14314 12673
rect 1734 12442 1820 12494
rect 1872 12442 1958 12494
rect 1734 12160 1958 12442
rect 1734 12104 1818 12160
rect 1874 12104 1958 12160
rect 1734 11822 1958 12104
rect 1734 11770 1820 11822
rect 1872 11770 1958 11822
rect 1734 11486 1958 11770
rect 1734 11434 1820 11486
rect 1872 11434 1958 11486
rect 1734 11150 1958 11434
rect 14258 11315 14314 11324
rect 14258 11250 14314 11259
rect 1734 11098 1820 11150
rect 1872 11098 1958 11150
rect 1734 10814 1958 11098
rect 1734 10762 1820 10814
rect 1872 10762 1958 10814
rect 1734 10480 1958 10762
rect 1734 10424 1818 10480
rect 1874 10424 1958 10480
rect 1734 10142 1958 10424
rect 1734 10090 1820 10142
rect 1872 10090 1958 10142
rect 1734 9806 1958 10090
rect 14258 9901 14314 9910
rect 14258 9836 14314 9845
rect 1734 9754 1820 9806
rect 1872 9754 1958 9806
rect 1734 9470 1958 9754
rect 1734 9418 1820 9470
rect 1872 9418 1958 9470
rect 1734 9134 1958 9418
rect 1734 9082 1820 9134
rect 1872 9082 1958 9134
rect 1734 8800 1958 9082
rect 1734 8744 1818 8800
rect 1874 8744 1958 8800
rect 1734 8462 1958 8744
rect 1734 8410 1820 8462
rect 1872 8410 1958 8462
rect 1734 8126 1958 8410
rect 1734 8074 1820 8126
rect 1872 8074 1958 8126
rect 1734 7790 1958 8074
rect 1734 7738 1820 7790
rect 1872 7738 1958 7790
rect 1734 7454 1958 7738
rect 1734 7402 1820 7454
rect 1872 7402 1958 7454
rect 1734 7120 1958 7402
rect 2778 7216 2834 7225
rect 2778 7151 2834 7160
rect 1734 7064 1818 7120
rect 1874 7064 1958 7120
rect 1734 6782 1958 7064
rect 1734 6730 1820 6782
rect 1872 6730 1958 6782
rect 1734 6446 1958 6730
rect 1734 6394 1820 6446
rect 1872 6394 1958 6446
rect 1734 6110 1958 6394
rect 1734 6058 1820 6110
rect 1872 6058 1958 6110
rect 1734 5774 1958 6058
rect 1734 5722 1820 5774
rect 1872 5722 1958 5774
rect 1734 5440 1958 5722
rect 14356 5645 14384 25321
rect 81858 16879 81886 76038
rect 94092 76000 94316 76282
rect 94092 75944 94176 76000
rect 94232 75944 94316 76000
rect 94092 75662 94316 75944
rect 94092 75610 94178 75662
rect 94230 75610 94316 75662
rect 94092 75326 94316 75610
rect 94092 75274 94178 75326
rect 94230 75274 94316 75326
rect 94092 74990 94316 75274
rect 94092 74938 94178 74990
rect 94230 74938 94316 74990
rect 94092 74654 94316 74938
rect 94092 74602 94178 74654
rect 94230 74602 94316 74654
rect 94092 74320 94316 74602
rect 94092 74264 94176 74320
rect 94232 74264 94316 74320
rect 94092 73982 94316 74264
rect 94092 73930 94178 73982
rect 94230 73930 94316 73982
rect 94092 73646 94316 73930
rect 94092 73594 94178 73646
rect 94230 73594 94316 73646
rect 94092 73310 94316 73594
rect 94092 73258 94178 73310
rect 94230 73258 94316 73310
rect 94092 72974 94316 73258
rect 94092 72922 94178 72974
rect 94230 72922 94316 72974
rect 94092 72640 94316 72922
rect 94092 72584 94176 72640
rect 94232 72584 94316 72640
rect 94092 72302 94316 72584
rect 94092 72250 94178 72302
rect 94230 72250 94316 72302
rect 81928 72187 81984 72196
rect 81928 72122 81984 72131
rect 94092 71966 94316 72250
rect 94092 71914 94178 71966
rect 94230 71914 94316 71966
rect 94092 71630 94316 71914
rect 94092 71578 94178 71630
rect 94230 71578 94316 71630
rect 94092 71294 94316 71578
rect 94092 71242 94178 71294
rect 94230 71242 94316 71294
rect 94092 70960 94316 71242
rect 94092 70904 94176 70960
rect 94232 70904 94316 70960
rect 81928 70773 81984 70782
rect 81928 70708 81984 70717
rect 94092 70622 94316 70904
rect 94092 70570 94178 70622
rect 94230 70570 94316 70622
rect 94092 70286 94316 70570
rect 94092 70234 94178 70286
rect 94230 70234 94316 70286
rect 94092 69950 94316 70234
rect 94092 69898 94178 69950
rect 94230 69898 94316 69950
rect 94092 69614 94316 69898
rect 94092 69562 94178 69614
rect 94230 69562 94316 69614
rect 81928 69359 81984 69368
rect 81928 69294 81984 69303
rect 94092 69280 94316 69562
rect 94092 69224 94176 69280
rect 94232 69224 94316 69280
rect 94092 68942 94316 69224
rect 94092 68890 94178 68942
rect 94230 68890 94316 68942
rect 94092 68606 94316 68890
rect 94092 68554 94178 68606
rect 94230 68554 94316 68606
rect 94092 68270 94316 68554
rect 94092 68218 94178 68270
rect 94230 68218 94316 68270
rect 94092 67934 94316 68218
rect 94092 67882 94178 67934
rect 94230 67882 94316 67934
rect 94092 67600 94316 67882
rect 94092 67544 94176 67600
rect 94232 67544 94316 67600
rect 94092 67262 94316 67544
rect 94092 67210 94178 67262
rect 94230 67210 94316 67262
rect 94092 66926 94316 67210
rect 94092 66874 94178 66926
rect 94230 66874 94316 66926
rect 94092 66590 94316 66874
rect 94092 66538 94178 66590
rect 94230 66538 94316 66590
rect 94092 66254 94316 66538
rect 94092 66202 94178 66254
rect 94230 66202 94316 66254
rect 94092 65920 94316 66202
rect 94092 65864 94176 65920
rect 94232 65864 94316 65920
rect 94092 65582 94316 65864
rect 94092 65530 94178 65582
rect 94230 65530 94316 65582
rect 94092 65246 94316 65530
rect 94092 65194 94178 65246
rect 94230 65194 94316 65246
rect 94092 64910 94316 65194
rect 94092 64858 94178 64910
rect 94230 64858 94316 64910
rect 94092 64574 94316 64858
rect 94092 64522 94178 64574
rect 94230 64522 94316 64574
rect 94092 64240 94316 64522
rect 94092 64184 94176 64240
rect 94232 64184 94316 64240
rect 94092 63902 94316 64184
rect 94092 63850 94178 63902
rect 94230 63850 94316 63902
rect 94092 63566 94316 63850
rect 94092 63514 94178 63566
rect 94230 63514 94316 63566
rect 94092 63230 94316 63514
rect 94092 63178 94178 63230
rect 94230 63178 94316 63230
rect 94092 62894 94316 63178
rect 94092 62842 94178 62894
rect 94230 62842 94316 62894
rect 94092 62560 94316 62842
rect 94092 62504 94176 62560
rect 94232 62504 94316 62560
rect 94092 62222 94316 62504
rect 94092 62170 94178 62222
rect 94230 62170 94316 62222
rect 94092 61886 94316 62170
rect 94092 61834 94178 61886
rect 94230 61834 94316 61886
rect 94092 61550 94316 61834
rect 94092 61498 94178 61550
rect 94230 61498 94316 61550
rect 94092 61214 94316 61498
rect 94092 61162 94178 61214
rect 94230 61162 94316 61214
rect 94092 60880 94316 61162
rect 94092 60824 94176 60880
rect 94232 60824 94316 60880
rect 94092 60542 94316 60824
rect 94092 60490 94178 60542
rect 94230 60490 94316 60542
rect 94092 60206 94316 60490
rect 94092 60154 94178 60206
rect 94230 60154 94316 60206
rect 94092 59870 94316 60154
rect 94092 59818 94178 59870
rect 94230 59818 94316 59870
rect 94092 59534 94316 59818
rect 94092 59482 94178 59534
rect 94230 59482 94316 59534
rect 93429 59423 93485 59432
rect 93429 59358 93485 59367
rect 94092 59200 94316 59482
rect 94092 59144 94176 59200
rect 94232 59144 94316 59200
rect 94092 58862 94316 59144
rect 94092 58810 94178 58862
rect 94230 58810 94316 58862
rect 94092 58526 94316 58810
rect 94092 58474 94178 58526
rect 94230 58474 94316 58526
rect 94092 58190 94316 58474
rect 94092 58138 94178 58190
rect 94230 58138 94316 58190
rect 94092 57854 94316 58138
rect 94092 57802 94178 57854
rect 94230 57802 94316 57854
rect 94092 57520 94316 57802
rect 94092 57464 94176 57520
rect 94232 57464 94316 57520
rect 94092 57182 94316 57464
rect 94092 57130 94178 57182
rect 94230 57130 94316 57182
rect 94092 56846 94316 57130
rect 94092 56794 94178 56846
rect 94230 56794 94316 56846
rect 94092 56510 94316 56794
rect 94092 56458 94178 56510
rect 94230 56458 94316 56510
rect 94092 56174 94316 56458
rect 94092 56122 94178 56174
rect 94230 56122 94316 56174
rect 94092 55840 94316 56122
rect 94092 55784 94176 55840
rect 94232 55784 94316 55840
rect 94092 55502 94316 55784
rect 94092 55450 94178 55502
rect 94230 55450 94316 55502
rect 94092 55166 94316 55450
rect 94092 55114 94178 55166
rect 94230 55114 94316 55166
rect 94092 54830 94316 55114
rect 94092 54778 94178 54830
rect 94230 54778 94316 54830
rect 94092 54494 94316 54778
rect 94092 54442 94178 54494
rect 94230 54442 94316 54494
rect 94092 54160 94316 54442
rect 94092 54104 94176 54160
rect 94232 54104 94316 54160
rect 94092 53822 94316 54104
rect 94092 53770 94178 53822
rect 94230 53770 94316 53822
rect 94092 53486 94316 53770
rect 94092 53434 94178 53486
rect 94230 53434 94316 53486
rect 94092 53150 94316 53434
rect 94092 53098 94178 53150
rect 94230 53098 94316 53150
rect 94092 52814 94316 53098
rect 94092 52762 94178 52814
rect 94230 52762 94316 52814
rect 94092 52480 94316 52762
rect 94092 52424 94176 52480
rect 94232 52424 94316 52480
rect 94092 52142 94316 52424
rect 94092 52090 94178 52142
rect 94230 52090 94316 52142
rect 94092 51806 94316 52090
rect 94092 51754 94178 51806
rect 94230 51754 94316 51806
rect 94092 51470 94316 51754
rect 94092 51418 94178 51470
rect 94230 51418 94316 51470
rect 94092 51134 94316 51418
rect 94092 51082 94178 51134
rect 94230 51082 94316 51134
rect 94092 50800 94316 51082
rect 94092 50744 94176 50800
rect 94232 50744 94316 50800
rect 94092 50462 94316 50744
rect 94092 50410 94178 50462
rect 94230 50410 94316 50462
rect 94092 50126 94316 50410
rect 94092 50074 94178 50126
rect 94230 50074 94316 50126
rect 94092 49790 94316 50074
rect 94092 49738 94178 49790
rect 94230 49738 94316 49790
rect 94092 49454 94316 49738
rect 94092 49402 94178 49454
rect 94230 49402 94316 49454
rect 94092 49120 94316 49402
rect 94092 49064 94176 49120
rect 94232 49064 94316 49120
rect 94092 48782 94316 49064
rect 94092 48730 94178 48782
rect 94230 48730 94316 48782
rect 94092 48446 94316 48730
rect 94092 48394 94178 48446
rect 94230 48394 94316 48446
rect 94092 48110 94316 48394
rect 94092 48058 94178 48110
rect 94230 48058 94316 48110
rect 94092 47774 94316 48058
rect 94092 47722 94178 47774
rect 94230 47722 94316 47774
rect 94092 47440 94316 47722
rect 94092 47384 94176 47440
rect 94232 47384 94316 47440
rect 94092 47102 94316 47384
rect 94092 47050 94178 47102
rect 94230 47050 94316 47102
rect 94092 46766 94316 47050
rect 94092 46714 94178 46766
rect 94230 46714 94316 46766
rect 94092 46430 94316 46714
rect 94092 46378 94178 46430
rect 94230 46378 94316 46430
rect 94092 46094 94316 46378
rect 94092 46042 94178 46094
rect 94230 46042 94316 46094
rect 94092 45760 94316 46042
rect 94092 45704 94176 45760
rect 94232 45704 94316 45760
rect 94092 45422 94316 45704
rect 94092 45370 94178 45422
rect 94230 45370 94316 45422
rect 94092 45086 94316 45370
rect 94092 45034 94178 45086
rect 94230 45034 94316 45086
rect 94092 44750 94316 45034
rect 94092 44698 94178 44750
rect 94230 44698 94316 44750
rect 94092 44414 94316 44698
rect 94092 44362 94178 44414
rect 94230 44362 94316 44414
rect 94092 44080 94316 44362
rect 94092 44024 94176 44080
rect 94232 44024 94316 44080
rect 94092 43742 94316 44024
rect 94092 43690 94178 43742
rect 94230 43690 94316 43742
rect 94092 43406 94316 43690
rect 94092 43354 94178 43406
rect 94230 43354 94316 43406
rect 94092 43070 94316 43354
rect 94092 43018 94178 43070
rect 94230 43018 94316 43070
rect 94092 42734 94316 43018
rect 94092 42682 94178 42734
rect 94230 42682 94316 42734
rect 94092 42400 94316 42682
rect 94092 42344 94176 42400
rect 94232 42344 94316 42400
rect 94092 42062 94316 42344
rect 94092 42010 94178 42062
rect 94230 42010 94316 42062
rect 94092 41726 94316 42010
rect 94092 41674 94178 41726
rect 94230 41674 94316 41726
rect 94092 41390 94316 41674
rect 94092 41338 94178 41390
rect 94230 41338 94316 41390
rect 94092 41054 94316 41338
rect 94092 41002 94178 41054
rect 94230 41002 94316 41054
rect 94092 40720 94316 41002
rect 94092 40664 94176 40720
rect 94232 40664 94316 40720
rect 94092 40382 94316 40664
rect 94092 40330 94178 40382
rect 94230 40330 94316 40382
rect 94092 40046 94316 40330
rect 94092 39994 94178 40046
rect 94230 39994 94316 40046
rect 94092 39710 94316 39994
rect 94092 39658 94178 39710
rect 94230 39658 94316 39710
rect 94092 39374 94316 39658
rect 94092 39322 94178 39374
rect 94230 39322 94316 39374
rect 94092 39040 94316 39322
rect 94092 38984 94176 39040
rect 94232 38984 94316 39040
rect 94092 38702 94316 38984
rect 94092 38650 94178 38702
rect 94230 38650 94316 38702
rect 94092 38366 94316 38650
rect 94092 38314 94178 38366
rect 94230 38314 94316 38366
rect 94092 38030 94316 38314
rect 94092 37978 94178 38030
rect 94230 37978 94316 38030
rect 94092 37694 94316 37978
rect 94092 37642 94178 37694
rect 94230 37642 94316 37694
rect 94092 37360 94316 37642
rect 94092 37304 94176 37360
rect 94232 37304 94316 37360
rect 94092 37022 94316 37304
rect 94092 36970 94178 37022
rect 94230 36970 94316 37022
rect 94092 36686 94316 36970
rect 94092 36634 94178 36686
rect 94230 36634 94316 36686
rect 94092 36350 94316 36634
rect 94092 36298 94178 36350
rect 94230 36298 94316 36350
rect 94092 36014 94316 36298
rect 94092 35962 94178 36014
rect 94230 35962 94316 36014
rect 94092 35680 94316 35962
rect 94092 35624 94176 35680
rect 94232 35624 94316 35680
rect 94092 35342 94316 35624
rect 94092 35290 94178 35342
rect 94230 35290 94316 35342
rect 94092 35006 94316 35290
rect 94092 34954 94178 35006
rect 94230 34954 94316 35006
rect 94092 34670 94316 34954
rect 94092 34618 94178 34670
rect 94230 34618 94316 34670
rect 94092 34334 94316 34618
rect 94092 34282 94178 34334
rect 94230 34282 94316 34334
rect 94092 34000 94316 34282
rect 94092 33944 94176 34000
rect 94232 33944 94316 34000
rect 94092 33662 94316 33944
rect 94092 33610 94178 33662
rect 94230 33610 94316 33662
rect 94092 33326 94316 33610
rect 94092 33274 94178 33326
rect 94230 33274 94316 33326
rect 94092 32990 94316 33274
rect 94092 32938 94178 32990
rect 94230 32938 94316 32990
rect 94092 32654 94316 32938
rect 94092 32602 94178 32654
rect 94230 32602 94316 32654
rect 94092 32320 94316 32602
rect 94092 32264 94176 32320
rect 94232 32264 94316 32320
rect 94092 31982 94316 32264
rect 94092 31930 94178 31982
rect 94230 31930 94316 31982
rect 94092 31646 94316 31930
rect 94092 31594 94178 31646
rect 94230 31594 94316 31646
rect 94092 31310 94316 31594
rect 94092 31258 94178 31310
rect 94230 31258 94316 31310
rect 94092 30974 94316 31258
rect 94092 30922 94178 30974
rect 94230 30922 94316 30974
rect 94092 30640 94316 30922
rect 94092 30584 94176 30640
rect 94232 30584 94316 30640
rect 94092 30302 94316 30584
rect 94092 30250 94178 30302
rect 94230 30250 94316 30302
rect 94092 29966 94316 30250
rect 94092 29914 94178 29966
rect 94230 29914 94316 29966
rect 94092 29630 94316 29914
rect 94092 29578 94178 29630
rect 94230 29578 94316 29630
rect 94092 29294 94316 29578
rect 94092 29242 94178 29294
rect 94230 29242 94316 29294
rect 94092 28960 94316 29242
rect 94092 28904 94176 28960
rect 94232 28904 94316 28960
rect 94092 28622 94316 28904
rect 94092 28570 94178 28622
rect 94230 28570 94316 28622
rect 94092 28286 94316 28570
rect 94092 28234 94178 28286
rect 94230 28234 94316 28286
rect 94092 27950 94316 28234
rect 94092 27898 94178 27950
rect 94230 27898 94316 27950
rect 94092 27614 94316 27898
rect 94092 27562 94178 27614
rect 94230 27562 94316 27614
rect 94092 27280 94316 27562
rect 94092 27224 94176 27280
rect 94232 27224 94316 27280
rect 94092 26942 94316 27224
rect 94092 26890 94178 26942
rect 94230 26890 94316 26942
rect 94092 26606 94316 26890
rect 94092 26554 94178 26606
rect 94230 26554 94316 26606
rect 94092 26270 94316 26554
rect 94092 26218 94178 26270
rect 94230 26218 94316 26270
rect 94092 25934 94316 26218
rect 94092 25882 94178 25934
rect 94230 25882 94316 25934
rect 94092 25600 94316 25882
rect 94092 25544 94176 25600
rect 94232 25544 94316 25600
rect 94092 25262 94316 25544
rect 94092 25210 94178 25262
rect 94230 25210 94316 25262
rect 94092 24926 94316 25210
rect 94092 24874 94178 24926
rect 94230 24874 94316 24926
rect 94092 24590 94316 24874
rect 94092 24538 94178 24590
rect 94230 24538 94316 24590
rect 94092 24254 94316 24538
rect 94092 24202 94178 24254
rect 94230 24202 94316 24254
rect 94092 23920 94316 24202
rect 94092 23864 94176 23920
rect 94232 23864 94316 23920
rect 94092 23582 94316 23864
rect 94092 23530 94178 23582
rect 94230 23530 94316 23582
rect 94092 23246 94316 23530
rect 94092 23194 94178 23246
rect 94230 23194 94316 23246
rect 94092 22910 94316 23194
rect 94092 22858 94178 22910
rect 94230 22858 94316 22910
rect 94092 22574 94316 22858
rect 94092 22522 94178 22574
rect 94230 22522 94316 22574
rect 94092 22240 94316 22522
rect 94092 22184 94176 22240
rect 94232 22184 94316 22240
rect 94092 21902 94316 22184
rect 94092 21850 94178 21902
rect 94230 21850 94316 21902
rect 94092 21566 94316 21850
rect 94092 21514 94178 21566
rect 94230 21514 94316 21566
rect 94092 21230 94316 21514
rect 94092 21178 94178 21230
rect 94230 21178 94316 21230
rect 94092 20894 94316 21178
rect 94092 20842 94178 20894
rect 94230 20842 94316 20894
rect 94092 20560 94316 20842
rect 94092 20504 94176 20560
rect 94232 20504 94316 20560
rect 94092 20222 94316 20504
rect 94092 20170 94178 20222
rect 94230 20170 94316 20222
rect 94092 19886 94316 20170
rect 94092 19834 94178 19886
rect 94230 19834 94316 19886
rect 94092 19550 94316 19834
rect 94092 19498 94178 19550
rect 94230 19498 94316 19550
rect 94092 19214 94316 19498
rect 94092 19162 94178 19214
rect 94230 19162 94316 19214
rect 94092 18880 94316 19162
rect 94092 18824 94176 18880
rect 94232 18824 94316 18880
rect 94092 18542 94316 18824
rect 94092 18490 94178 18542
rect 94230 18490 94316 18542
rect 94092 18206 94316 18490
rect 94092 18154 94178 18206
rect 94230 18154 94316 18206
rect 94092 17870 94316 18154
rect 94092 17818 94178 17870
rect 94230 17818 94316 17870
rect 94092 17534 94316 17818
rect 94092 17482 94178 17534
rect 94230 17482 94316 17534
rect 94092 17200 94316 17482
rect 94092 17144 94176 17200
rect 94232 17144 94316 17200
rect 81844 16870 81900 16879
rect 22414 15566 22442 16851
rect 81844 16805 81900 16814
rect 94092 16862 94316 17144
rect 94092 16810 94178 16862
rect 94230 16810 94316 16862
rect 82926 16614 82982 16623
rect 81643 16543 81699 16552
rect 81643 16478 81699 16487
rect 81981 16543 82037 16552
rect 82926 16549 82982 16558
rect 81981 16478 82037 16487
rect 94092 16526 94316 16810
rect 94092 16474 94178 16526
rect 94230 16474 94316 16526
rect 22400 15557 22456 15566
rect 22400 15492 22456 15501
rect 26117 12738 26145 16374
rect 94092 16190 94316 16474
rect 94092 16138 94178 16190
rect 94230 16138 94316 16190
rect 94092 15854 94316 16138
rect 94092 15802 94178 15854
rect 94230 15802 94316 15854
rect 94092 15520 94316 15802
rect 94092 15464 94176 15520
rect 94232 15464 94316 15520
rect 94092 15182 94316 15464
rect 94092 15130 94178 15182
rect 94230 15130 94316 15182
rect 81563 14985 81619 14994
rect 81563 14920 81619 14929
rect 81981 14985 82037 14994
rect 81981 14920 82037 14929
rect 82926 14914 82982 14923
rect 82926 14849 82982 14858
rect 94092 14846 94316 15130
rect 94092 14794 94178 14846
rect 94230 14794 94316 14846
rect 94092 14510 94316 14794
rect 94092 14458 94178 14510
rect 94230 14458 94316 14510
rect 94092 14174 94316 14458
rect 94092 14122 94178 14174
rect 94230 14122 94316 14174
rect 94092 13840 94316 14122
rect 82926 13786 82982 13795
rect 81483 13715 81539 13724
rect 81483 13650 81539 13659
rect 81981 13715 82037 13724
rect 82926 13721 82982 13730
rect 94092 13784 94176 13840
rect 94232 13784 94316 13840
rect 81981 13650 82037 13659
rect 94092 13502 94316 13784
rect 94092 13450 94178 13502
rect 94230 13450 94316 13502
rect 94092 13166 94316 13450
rect 94092 13114 94178 13166
rect 94230 13114 94316 13166
rect 94092 12830 94316 13114
rect 94092 12778 94178 12830
rect 94230 12778 94316 12830
rect 26103 12729 26159 12738
rect 26103 12664 26159 12673
rect 94092 12494 94316 12778
rect 94092 12442 94178 12494
rect 94230 12442 94316 12494
rect 81403 12157 81459 12166
rect 81403 12092 81459 12101
rect 81981 12157 82037 12166
rect 81981 12092 82037 12101
rect 94092 12160 94316 12442
rect 94092 12104 94176 12160
rect 94232 12104 94316 12160
rect 82926 12086 82982 12095
rect 82926 12021 82982 12030
rect 94092 11822 94316 12104
rect 94092 11770 94178 11822
rect 94230 11770 94316 11822
rect 94092 11486 94316 11770
rect 94092 11434 94178 11486
rect 94230 11434 94316 11486
rect 26351 11315 26407 11324
rect 26351 11250 26407 11259
rect 26227 9901 26283 9910
rect 26227 9836 26283 9845
rect 26241 7009 26269 9836
rect 26365 7009 26393 11250
rect 94092 11150 94316 11434
rect 94092 11098 94178 11150
rect 94230 11098 94316 11150
rect 82926 10958 82982 10967
rect 81323 10887 81379 10896
rect 81323 10822 81379 10831
rect 81981 10887 82037 10896
rect 82926 10893 82982 10902
rect 81981 10822 82037 10831
rect 28210 10813 28266 10822
rect 28210 10748 28266 10757
rect 29458 10813 29514 10822
rect 29458 10748 29514 10757
rect 30706 10813 30762 10822
rect 30706 10748 30762 10757
rect 31954 10813 32010 10822
rect 31954 10748 32010 10757
rect 33202 10813 33258 10822
rect 33202 10748 33258 10757
rect 34450 10813 34506 10822
rect 34450 10748 34506 10757
rect 35698 10813 35754 10822
rect 35698 10748 35754 10757
rect 36946 10813 37002 10822
rect 36946 10748 37002 10757
rect 38194 10813 38250 10822
rect 38194 10748 38250 10757
rect 39442 10813 39498 10822
rect 39442 10748 39498 10757
rect 40690 10813 40746 10822
rect 40690 10748 40746 10757
rect 41938 10813 41994 10822
rect 41938 10748 41994 10757
rect 43186 10813 43242 10822
rect 43186 10748 43242 10757
rect 44434 10813 44490 10822
rect 44434 10748 44490 10757
rect 45682 10813 45738 10822
rect 45682 10748 45738 10757
rect 46930 10813 46986 10822
rect 46930 10748 46986 10757
rect 48178 10813 48234 10822
rect 48178 10748 48234 10757
rect 49426 10813 49482 10822
rect 49426 10748 49482 10757
rect 50674 10813 50730 10822
rect 50674 10748 50730 10757
rect 51922 10813 51978 10822
rect 51922 10748 51978 10757
rect 53170 10813 53226 10822
rect 53170 10748 53226 10757
rect 54418 10813 54474 10822
rect 54418 10748 54474 10757
rect 55666 10813 55722 10822
rect 55666 10748 55722 10757
rect 56914 10813 56970 10822
rect 56914 10748 56970 10757
rect 58162 10813 58218 10822
rect 58162 10748 58218 10757
rect 59410 10813 59466 10822
rect 59410 10748 59466 10757
rect 60658 10813 60714 10822
rect 60658 10748 60714 10757
rect 61906 10813 61962 10822
rect 61906 10748 61962 10757
rect 63154 10813 63210 10822
rect 63154 10748 63210 10757
rect 64402 10813 64458 10822
rect 64402 10748 64458 10757
rect 65650 10813 65706 10822
rect 65650 10748 65706 10757
rect 66898 10813 66954 10822
rect 66898 10748 66954 10757
rect 94092 10814 94316 11098
rect 94092 10762 94178 10814
rect 94230 10762 94316 10814
rect 94092 10480 94316 10762
rect 94092 10424 94176 10480
rect 94232 10424 94316 10480
rect 94092 10142 94316 10424
rect 94092 10090 94178 10142
rect 94230 10090 94316 10142
rect 94092 9806 94316 10090
rect 94092 9754 94178 9806
rect 94230 9754 94316 9806
rect 94092 9470 94316 9754
rect 94092 9418 94178 9470
rect 94230 9418 94316 9470
rect 81243 9329 81299 9338
rect 81243 9264 81299 9273
rect 81981 9329 82037 9338
rect 81981 9264 82037 9273
rect 82926 9258 82982 9267
rect 82926 9193 82982 9202
rect 94092 9134 94316 9418
rect 94092 9082 94178 9134
rect 94230 9082 94316 9134
rect 94092 8800 94316 9082
rect 94092 8744 94176 8800
rect 94232 8744 94316 8800
rect 94092 8462 94316 8744
rect 94092 8410 94178 8462
rect 94230 8410 94316 8462
rect 82926 8130 82982 8139
rect 81163 8059 81219 8068
rect 81163 7994 81219 8003
rect 81981 8059 82037 8068
rect 82926 8065 82982 8074
rect 94092 8126 94316 8410
rect 94092 8074 94178 8126
rect 94230 8074 94316 8126
rect 81981 7994 82037 8003
rect 94092 7790 94316 8074
rect 94092 7738 94178 7790
rect 94230 7738 94316 7790
rect 94092 7454 94316 7738
rect 94092 7402 94178 7454
rect 94230 7402 94316 7454
rect 94092 7120 94316 7402
rect 94092 7064 94176 7120
rect 94232 7064 94316 7120
rect 5999 5621 6055 5630
rect 14286 5617 14384 5645
rect 5999 5556 6055 5565
rect 2778 5516 2834 5525
rect 2778 5451 2834 5460
rect 1734 5384 1818 5440
rect 1874 5384 1958 5440
rect 1734 5102 1958 5384
rect 1734 5050 1820 5102
rect 1872 5050 1958 5102
rect 1734 4766 1958 5050
rect 1734 4714 1820 4766
rect 1872 4714 1958 4766
rect 1734 4430 1958 4714
rect 1734 4378 1820 4430
rect 1872 4378 1958 4430
rect 1734 4094 1958 4378
rect 1734 4042 1820 4094
rect 1872 4042 1958 4094
rect 1734 3760 1958 4042
rect 1734 3704 1818 3760
rect 1874 3704 1958 3760
rect 1734 3422 1958 3704
rect 1734 3370 1820 3422
rect 1872 3370 1958 3422
rect 1734 3086 1958 3370
rect 1734 3034 1820 3086
rect 1872 3034 1958 3086
rect 1734 2750 1958 3034
rect 1734 2698 1820 2750
rect 1872 2698 1958 2750
rect 14356 2733 14384 5617
rect 94092 6782 94316 7064
rect 94092 6730 94178 6782
rect 94230 6730 94316 6782
rect 94092 6446 94316 6730
rect 94092 6394 94178 6446
rect 94230 6394 94316 6446
rect 94092 6110 94316 6394
rect 94092 6058 94178 6110
rect 94230 6058 94316 6110
rect 94092 5774 94316 6058
rect 94092 5722 94178 5774
rect 94230 5722 94316 5774
rect 94092 5440 94316 5722
rect 94092 5384 94176 5440
rect 94232 5384 94316 5440
rect 94092 5102 94316 5384
rect 94092 5050 94178 5102
rect 94230 5050 94316 5102
rect 94092 4766 94316 5050
rect 94092 4714 94178 4766
rect 94230 4714 94316 4766
rect 94092 4430 94316 4714
rect 94092 4378 94178 4430
rect 94230 4378 94316 4430
rect 94092 4094 94316 4378
rect 94092 4042 94178 4094
rect 94230 4042 94316 4094
rect 94092 3760 94316 4042
rect 94092 3704 94176 3760
rect 94232 3704 94316 3760
rect 94092 3422 94316 3704
rect 94092 3370 94178 3422
rect 94230 3370 94316 3422
rect 94092 3086 94316 3370
rect 94092 3034 94178 3086
rect 94230 3034 94316 3086
rect 15596 2980 15652 2989
rect 15596 2915 15652 2924
rect 16764 2980 16820 2989
rect 16764 2915 16820 2924
rect 17932 2980 17988 2989
rect 17932 2915 17988 2924
rect 19100 2980 19156 2989
rect 19100 2915 19156 2924
rect 20268 2980 20324 2989
rect 20268 2915 20324 2924
rect 21436 2980 21492 2989
rect 21436 2915 21492 2924
rect 22604 2980 22660 2989
rect 22604 2915 22660 2924
rect 23772 2980 23828 2989
rect 23772 2915 23828 2924
rect 24940 2980 24996 2989
rect 24940 2915 24996 2924
rect 26108 2980 26164 2989
rect 26108 2915 26164 2924
rect 27276 2980 27332 2989
rect 27276 2915 27332 2924
rect 28444 2980 28500 2989
rect 28444 2915 28500 2924
rect 29612 2980 29668 2989
rect 29612 2915 29668 2924
rect 30780 2980 30836 2989
rect 30780 2915 30836 2924
rect 31948 2980 32004 2989
rect 31948 2915 32004 2924
rect 33116 2980 33172 2989
rect 33116 2915 33172 2924
rect 34284 2980 34340 2989
rect 34284 2915 34340 2924
rect 35452 2980 35508 2989
rect 35452 2915 35508 2924
rect 36620 2980 36676 2989
rect 36620 2915 36676 2924
rect 37788 2980 37844 2989
rect 37788 2915 37844 2924
rect 38956 2980 39012 2989
rect 38956 2915 39012 2924
rect 40124 2980 40180 2989
rect 40124 2915 40180 2924
rect 41292 2980 41348 2989
rect 41292 2915 41348 2924
rect 42460 2980 42516 2989
rect 42460 2915 42516 2924
rect 43628 2980 43684 2989
rect 43628 2915 43684 2924
rect 44796 2980 44852 2989
rect 44796 2915 44852 2924
rect 45964 2980 46020 2989
rect 45964 2915 46020 2924
rect 47132 2980 47188 2989
rect 47132 2915 47188 2924
rect 48300 2980 48356 2989
rect 48300 2915 48356 2924
rect 49468 2980 49524 2989
rect 49468 2915 49524 2924
rect 50636 2980 50692 2989
rect 50636 2915 50692 2924
rect 51804 2980 51860 2989
rect 51804 2915 51860 2924
rect 52972 2980 53028 2989
rect 52972 2915 53028 2924
rect 54140 2980 54196 2989
rect 54140 2915 54196 2924
rect 55308 2980 55364 2989
rect 55308 2915 55364 2924
rect 56476 2980 56532 2989
rect 56476 2915 56532 2924
rect 57644 2980 57700 2989
rect 57644 2915 57700 2924
rect 94092 2750 94316 3034
rect 1734 2414 1958 2698
rect 14342 2724 14398 2733
rect 14342 2659 14398 2668
rect 94092 2698 94178 2750
rect 94230 2698 94316 2750
rect 1734 2362 1820 2414
rect 1872 2362 1958 2414
rect 1734 2080 1958 2362
rect 1734 2024 1818 2080
rect 1874 2024 1958 2080
rect 1734 1604 1958 2024
rect 94092 2414 94316 2698
rect 94092 2362 94178 2414
rect 94230 2362 94316 2414
rect 94092 2080 94316 2362
rect 94092 2024 94176 2080
rect 94232 2024 94316 2080
rect 2154 1744 2210 1753
rect 2154 1679 2210 1688
rect 3834 1744 3890 1753
rect 3834 1679 3890 1688
rect 5514 1744 5570 1753
rect 5514 1679 5570 1688
rect 7194 1744 7250 1753
rect 7194 1679 7250 1688
rect 8874 1744 8930 1753
rect 8874 1679 8930 1688
rect 10554 1744 10610 1753
rect 10554 1679 10610 1688
rect 12234 1744 12290 1753
rect 12234 1679 12290 1688
rect 13914 1744 13970 1753
rect 13914 1679 13970 1688
rect 15594 1744 15650 1753
rect 15594 1679 15650 1688
rect 17274 1744 17330 1753
rect 17274 1679 17330 1688
rect 18954 1744 19010 1753
rect 18954 1679 19010 1688
rect 20634 1744 20690 1753
rect 20634 1679 20690 1688
rect 22314 1744 22370 1753
rect 22314 1679 22370 1688
rect 23994 1744 24050 1753
rect 23994 1679 24050 1688
rect 25674 1744 25730 1753
rect 25674 1679 25730 1688
rect 27354 1744 27410 1753
rect 27354 1679 27410 1688
rect 29034 1744 29090 1753
rect 29034 1679 29090 1688
rect 30714 1744 30770 1753
rect 30714 1679 30770 1688
rect 32394 1744 32450 1753
rect 32394 1679 32450 1688
rect 34074 1744 34130 1753
rect 34074 1679 34130 1688
rect 35754 1744 35810 1753
rect 35754 1679 35810 1688
rect 37434 1744 37490 1753
rect 37434 1679 37490 1688
rect 39114 1744 39170 1753
rect 39114 1679 39170 1688
rect 40794 1744 40850 1753
rect 40794 1679 40850 1688
rect 42474 1744 42530 1753
rect 42474 1679 42530 1688
rect 44154 1744 44210 1753
rect 44154 1679 44210 1688
rect 45834 1744 45890 1753
rect 45834 1679 45890 1688
rect 47514 1744 47570 1753
rect 47514 1679 47570 1688
rect 49194 1744 49250 1753
rect 49194 1679 49250 1688
rect 50874 1744 50930 1753
rect 50874 1679 50930 1688
rect 52554 1744 52610 1753
rect 52554 1679 52610 1688
rect 54234 1744 54290 1753
rect 54234 1679 54290 1688
rect 55914 1744 55970 1753
rect 55914 1679 55970 1688
rect 57594 1744 57650 1753
rect 57594 1679 57650 1688
rect 59274 1744 59330 1753
rect 59274 1679 59330 1688
rect 60954 1744 61010 1753
rect 60954 1679 61010 1688
rect 62634 1744 62690 1753
rect 62634 1679 62690 1688
rect 64314 1744 64370 1753
rect 64314 1679 64370 1688
rect 65994 1744 66050 1753
rect 65994 1679 66050 1688
rect 67674 1744 67730 1753
rect 67674 1679 67730 1688
rect 69354 1744 69410 1753
rect 69354 1679 69410 1688
rect 71034 1744 71090 1753
rect 71034 1679 71090 1688
rect 72714 1744 72770 1753
rect 72714 1679 72770 1688
rect 74394 1744 74450 1753
rect 74394 1679 74450 1688
rect 76074 1744 76130 1753
rect 76074 1679 76130 1688
rect 77754 1744 77810 1753
rect 77754 1679 77810 1688
rect 79434 1744 79490 1753
rect 79434 1679 79490 1688
rect 81114 1744 81170 1753
rect 81114 1679 81170 1688
rect 82794 1744 82850 1753
rect 82794 1679 82850 1688
rect 84474 1744 84530 1753
rect 84474 1679 84530 1688
rect 86154 1744 86210 1753
rect 86154 1679 86210 1688
rect 87834 1744 87890 1753
rect 87834 1679 87890 1688
rect 89514 1744 89570 1753
rect 89514 1679 89570 1688
rect 91194 1744 91250 1753
rect 91194 1679 91250 1688
rect 92874 1744 92930 1753
rect 92874 1679 92930 1688
rect 94092 1604 94316 2024
<< via2 >>
rect 2154 77806 2210 77808
rect 2154 77754 2156 77806
rect 2156 77754 2208 77806
rect 2208 77754 2210 77806
rect 2154 77752 2210 77754
rect 3834 77806 3890 77808
rect 3834 77754 3836 77806
rect 3836 77754 3888 77806
rect 3888 77754 3890 77806
rect 3834 77752 3890 77754
rect 5514 77806 5570 77808
rect 5514 77754 5516 77806
rect 5516 77754 5568 77806
rect 5568 77754 5570 77806
rect 5514 77752 5570 77754
rect 7194 77806 7250 77808
rect 7194 77754 7196 77806
rect 7196 77754 7248 77806
rect 7248 77754 7250 77806
rect 7194 77752 7250 77754
rect 8874 77806 8930 77808
rect 8874 77754 8876 77806
rect 8876 77754 8928 77806
rect 8928 77754 8930 77806
rect 8874 77752 8930 77754
rect 10554 77806 10610 77808
rect 10554 77754 10556 77806
rect 10556 77754 10608 77806
rect 10608 77754 10610 77806
rect 10554 77752 10610 77754
rect 12234 77806 12290 77808
rect 12234 77754 12236 77806
rect 12236 77754 12288 77806
rect 12288 77754 12290 77806
rect 12234 77752 12290 77754
rect 13914 77806 13970 77808
rect 13914 77754 13916 77806
rect 13916 77754 13968 77806
rect 13968 77754 13970 77806
rect 13914 77752 13970 77754
rect 15594 77806 15650 77808
rect 15594 77754 15596 77806
rect 15596 77754 15648 77806
rect 15648 77754 15650 77806
rect 15594 77752 15650 77754
rect 17274 77806 17330 77808
rect 17274 77754 17276 77806
rect 17276 77754 17328 77806
rect 17328 77754 17330 77806
rect 17274 77752 17330 77754
rect 18954 77806 19010 77808
rect 18954 77754 18956 77806
rect 18956 77754 19008 77806
rect 19008 77754 19010 77806
rect 18954 77752 19010 77754
rect 20634 77806 20690 77808
rect 20634 77754 20636 77806
rect 20636 77754 20688 77806
rect 20688 77754 20690 77806
rect 20634 77752 20690 77754
rect 22314 77806 22370 77808
rect 22314 77754 22316 77806
rect 22316 77754 22368 77806
rect 22368 77754 22370 77806
rect 22314 77752 22370 77754
rect 23994 77806 24050 77808
rect 23994 77754 23996 77806
rect 23996 77754 24048 77806
rect 24048 77754 24050 77806
rect 23994 77752 24050 77754
rect 25674 77806 25730 77808
rect 25674 77754 25676 77806
rect 25676 77754 25728 77806
rect 25728 77754 25730 77806
rect 25674 77752 25730 77754
rect 27354 77806 27410 77808
rect 27354 77754 27356 77806
rect 27356 77754 27408 77806
rect 27408 77754 27410 77806
rect 27354 77752 27410 77754
rect 29034 77806 29090 77808
rect 29034 77754 29036 77806
rect 29036 77754 29088 77806
rect 29088 77754 29090 77806
rect 29034 77752 29090 77754
rect 30714 77806 30770 77808
rect 30714 77754 30716 77806
rect 30716 77754 30768 77806
rect 30768 77754 30770 77806
rect 30714 77752 30770 77754
rect 32394 77806 32450 77808
rect 32394 77754 32396 77806
rect 32396 77754 32448 77806
rect 32448 77754 32450 77806
rect 32394 77752 32450 77754
rect 34074 77806 34130 77808
rect 34074 77754 34076 77806
rect 34076 77754 34128 77806
rect 34128 77754 34130 77806
rect 34074 77752 34130 77754
rect 35754 77806 35810 77808
rect 35754 77754 35756 77806
rect 35756 77754 35808 77806
rect 35808 77754 35810 77806
rect 35754 77752 35810 77754
rect 37434 77806 37490 77808
rect 37434 77754 37436 77806
rect 37436 77754 37488 77806
rect 37488 77754 37490 77806
rect 37434 77752 37490 77754
rect 39114 77806 39170 77808
rect 39114 77754 39116 77806
rect 39116 77754 39168 77806
rect 39168 77754 39170 77806
rect 39114 77752 39170 77754
rect 40794 77806 40850 77808
rect 40794 77754 40796 77806
rect 40796 77754 40848 77806
rect 40848 77754 40850 77806
rect 40794 77752 40850 77754
rect 42474 77806 42530 77808
rect 42474 77754 42476 77806
rect 42476 77754 42528 77806
rect 42528 77754 42530 77806
rect 42474 77752 42530 77754
rect 44154 77806 44210 77808
rect 44154 77754 44156 77806
rect 44156 77754 44208 77806
rect 44208 77754 44210 77806
rect 44154 77752 44210 77754
rect 45834 77806 45890 77808
rect 45834 77754 45836 77806
rect 45836 77754 45888 77806
rect 45888 77754 45890 77806
rect 45834 77752 45890 77754
rect 47514 77806 47570 77808
rect 47514 77754 47516 77806
rect 47516 77754 47568 77806
rect 47568 77754 47570 77806
rect 47514 77752 47570 77754
rect 49194 77806 49250 77808
rect 49194 77754 49196 77806
rect 49196 77754 49248 77806
rect 49248 77754 49250 77806
rect 49194 77752 49250 77754
rect 50874 77806 50930 77808
rect 50874 77754 50876 77806
rect 50876 77754 50928 77806
rect 50928 77754 50930 77806
rect 50874 77752 50930 77754
rect 52554 77806 52610 77808
rect 52554 77754 52556 77806
rect 52556 77754 52608 77806
rect 52608 77754 52610 77806
rect 52554 77752 52610 77754
rect 54234 77806 54290 77808
rect 54234 77754 54236 77806
rect 54236 77754 54288 77806
rect 54288 77754 54290 77806
rect 54234 77752 54290 77754
rect 55914 77806 55970 77808
rect 55914 77754 55916 77806
rect 55916 77754 55968 77806
rect 55968 77754 55970 77806
rect 55914 77752 55970 77754
rect 57594 77806 57650 77808
rect 57594 77754 57596 77806
rect 57596 77754 57648 77806
rect 57648 77754 57650 77806
rect 57594 77752 57650 77754
rect 59274 77806 59330 77808
rect 59274 77754 59276 77806
rect 59276 77754 59328 77806
rect 59328 77754 59330 77806
rect 59274 77752 59330 77754
rect 60954 77806 61010 77808
rect 60954 77754 60956 77806
rect 60956 77754 61008 77806
rect 61008 77754 61010 77806
rect 60954 77752 61010 77754
rect 62634 77806 62690 77808
rect 62634 77754 62636 77806
rect 62636 77754 62688 77806
rect 62688 77754 62690 77806
rect 62634 77752 62690 77754
rect 64314 77806 64370 77808
rect 64314 77754 64316 77806
rect 64316 77754 64368 77806
rect 64368 77754 64370 77806
rect 64314 77752 64370 77754
rect 65994 77806 66050 77808
rect 65994 77754 65996 77806
rect 65996 77754 66048 77806
rect 66048 77754 66050 77806
rect 65994 77752 66050 77754
rect 67674 77806 67730 77808
rect 67674 77754 67676 77806
rect 67676 77754 67728 77806
rect 67728 77754 67730 77806
rect 67674 77752 67730 77754
rect 69354 77806 69410 77808
rect 69354 77754 69356 77806
rect 69356 77754 69408 77806
rect 69408 77754 69410 77806
rect 69354 77752 69410 77754
rect 71034 77806 71090 77808
rect 71034 77754 71036 77806
rect 71036 77754 71088 77806
rect 71088 77754 71090 77806
rect 71034 77752 71090 77754
rect 72714 77806 72770 77808
rect 72714 77754 72716 77806
rect 72716 77754 72768 77806
rect 72768 77754 72770 77806
rect 72714 77752 72770 77754
rect 74394 77806 74450 77808
rect 74394 77754 74396 77806
rect 74396 77754 74448 77806
rect 74448 77754 74450 77806
rect 74394 77752 74450 77754
rect 76074 77806 76130 77808
rect 76074 77754 76076 77806
rect 76076 77754 76128 77806
rect 76128 77754 76130 77806
rect 76074 77752 76130 77754
rect 77754 77806 77810 77808
rect 77754 77754 77756 77806
rect 77756 77754 77808 77806
rect 77808 77754 77810 77806
rect 77754 77752 77810 77754
rect 79434 77806 79490 77808
rect 79434 77754 79436 77806
rect 79436 77754 79488 77806
rect 79488 77754 79490 77806
rect 79434 77752 79490 77754
rect 81114 77806 81170 77808
rect 81114 77754 81116 77806
rect 81116 77754 81168 77806
rect 81168 77754 81170 77806
rect 81114 77752 81170 77754
rect 82794 77806 82850 77808
rect 82794 77754 82796 77806
rect 82796 77754 82848 77806
rect 82848 77754 82850 77806
rect 82794 77752 82850 77754
rect 84474 77806 84530 77808
rect 84474 77754 84476 77806
rect 84476 77754 84528 77806
rect 84528 77754 84530 77806
rect 84474 77752 84530 77754
rect 86154 77806 86210 77808
rect 86154 77754 86156 77806
rect 86156 77754 86208 77806
rect 86208 77754 86210 77806
rect 86154 77752 86210 77754
rect 87834 77806 87890 77808
rect 87834 77754 87836 77806
rect 87836 77754 87888 77806
rect 87888 77754 87890 77806
rect 87834 77752 87890 77754
rect 89514 77806 89570 77808
rect 89514 77754 89516 77806
rect 89516 77754 89568 77806
rect 89568 77754 89570 77806
rect 89514 77752 89570 77754
rect 91194 77806 91250 77808
rect 91194 77754 91196 77806
rect 91196 77754 91248 77806
rect 91248 77754 91250 77806
rect 91194 77752 91250 77754
rect 92874 77806 92930 77808
rect 92874 77754 92876 77806
rect 92876 77754 92928 77806
rect 92928 77754 92930 77806
rect 92874 77752 92930 77754
rect 93216 76516 93272 76572
rect 90079 76411 90135 76467
rect 81844 76047 81900 76103
rect 1818 75998 1874 76000
rect 1818 75946 1820 75998
rect 1820 75946 1872 75998
rect 1872 75946 1874 75998
rect 1818 75944 1874 75946
rect 79422 75791 79478 75847
rect 1818 74318 1874 74320
rect 1818 74266 1820 74318
rect 1820 74266 1872 74318
rect 1872 74266 1874 74318
rect 1818 74264 1874 74266
rect 28210 74101 28266 74103
rect 28210 74049 28212 74101
rect 28212 74049 28264 74101
rect 28264 74049 28266 74101
rect 28210 74047 28266 74049
rect 29458 74101 29514 74103
rect 29458 74049 29460 74101
rect 29460 74049 29512 74101
rect 29512 74049 29514 74101
rect 29458 74047 29514 74049
rect 30706 74101 30762 74103
rect 30706 74049 30708 74101
rect 30708 74049 30760 74101
rect 30760 74049 30762 74101
rect 30706 74047 30762 74049
rect 31954 74101 32010 74103
rect 31954 74049 31956 74101
rect 31956 74049 32008 74101
rect 32008 74049 32010 74101
rect 31954 74047 32010 74049
rect 33202 74101 33258 74103
rect 33202 74049 33204 74101
rect 33204 74049 33256 74101
rect 33256 74049 33258 74101
rect 33202 74047 33258 74049
rect 34450 74101 34506 74103
rect 34450 74049 34452 74101
rect 34452 74049 34504 74101
rect 34504 74049 34506 74101
rect 34450 74047 34506 74049
rect 35698 74101 35754 74103
rect 35698 74049 35700 74101
rect 35700 74049 35752 74101
rect 35752 74049 35754 74101
rect 35698 74047 35754 74049
rect 36946 74101 37002 74103
rect 36946 74049 36948 74101
rect 36948 74049 37000 74101
rect 37000 74049 37002 74101
rect 36946 74047 37002 74049
rect 38194 74101 38250 74103
rect 38194 74049 38196 74101
rect 38196 74049 38248 74101
rect 38248 74049 38250 74101
rect 38194 74047 38250 74049
rect 39442 74101 39498 74103
rect 39442 74049 39444 74101
rect 39444 74049 39496 74101
rect 39496 74049 39498 74101
rect 39442 74047 39498 74049
rect 40690 74101 40746 74103
rect 40690 74049 40692 74101
rect 40692 74049 40744 74101
rect 40744 74049 40746 74101
rect 40690 74047 40746 74049
rect 41938 74101 41994 74103
rect 41938 74049 41940 74101
rect 41940 74049 41992 74101
rect 41992 74049 41994 74101
rect 41938 74047 41994 74049
rect 43186 74101 43242 74103
rect 43186 74049 43188 74101
rect 43188 74049 43240 74101
rect 43240 74049 43242 74101
rect 43186 74047 43242 74049
rect 44434 74101 44490 74103
rect 44434 74049 44436 74101
rect 44436 74049 44488 74101
rect 44488 74049 44490 74101
rect 44434 74047 44490 74049
rect 45682 74101 45738 74103
rect 45682 74049 45684 74101
rect 45684 74049 45736 74101
rect 45736 74049 45738 74101
rect 45682 74047 45738 74049
rect 46930 74101 46986 74103
rect 46930 74049 46932 74101
rect 46932 74049 46984 74101
rect 46984 74049 46986 74101
rect 46930 74047 46986 74049
rect 48178 74101 48234 74103
rect 48178 74049 48180 74101
rect 48180 74049 48232 74101
rect 48232 74049 48234 74101
rect 48178 74047 48234 74049
rect 49426 74101 49482 74103
rect 49426 74049 49428 74101
rect 49428 74049 49480 74101
rect 49480 74049 49482 74101
rect 49426 74047 49482 74049
rect 50674 74101 50730 74103
rect 50674 74049 50676 74101
rect 50676 74049 50728 74101
rect 50728 74049 50730 74101
rect 50674 74047 50730 74049
rect 51922 74101 51978 74103
rect 51922 74049 51924 74101
rect 51924 74049 51976 74101
rect 51976 74049 51978 74101
rect 51922 74047 51978 74049
rect 53170 74101 53226 74103
rect 53170 74049 53172 74101
rect 53172 74049 53224 74101
rect 53224 74049 53226 74101
rect 53170 74047 53226 74049
rect 54418 74101 54474 74103
rect 54418 74049 54420 74101
rect 54420 74049 54472 74101
rect 54472 74049 54474 74101
rect 54418 74047 54474 74049
rect 55666 74101 55722 74103
rect 55666 74049 55668 74101
rect 55668 74049 55720 74101
rect 55720 74049 55722 74101
rect 55666 74047 55722 74049
rect 56914 74101 56970 74103
rect 56914 74049 56916 74101
rect 56916 74049 56968 74101
rect 56968 74049 56970 74101
rect 56914 74047 56970 74049
rect 58162 74101 58218 74103
rect 58162 74049 58164 74101
rect 58164 74049 58216 74101
rect 58216 74049 58218 74101
rect 58162 74047 58218 74049
rect 59410 74101 59466 74103
rect 59410 74049 59412 74101
rect 59412 74049 59464 74101
rect 59464 74049 59466 74101
rect 59410 74047 59466 74049
rect 60658 74101 60714 74103
rect 60658 74049 60660 74101
rect 60660 74049 60712 74101
rect 60712 74049 60714 74101
rect 60658 74047 60714 74049
rect 61906 74101 61962 74103
rect 61906 74049 61908 74101
rect 61908 74049 61960 74101
rect 61960 74049 61962 74101
rect 61906 74047 61962 74049
rect 63154 74101 63210 74103
rect 63154 74049 63156 74101
rect 63156 74049 63208 74101
rect 63208 74049 63210 74101
rect 63154 74047 63210 74049
rect 64402 74101 64458 74103
rect 64402 74049 64404 74101
rect 64404 74049 64456 74101
rect 64456 74049 64458 74101
rect 64402 74047 64458 74049
rect 65650 74101 65706 74103
rect 65650 74049 65652 74101
rect 65652 74049 65704 74101
rect 65704 74049 65706 74101
rect 65650 74047 65706 74049
rect 66898 74101 66954 74103
rect 66898 74049 66900 74101
rect 66900 74049 66952 74101
rect 66952 74049 66954 74101
rect 66898 74047 66954 74049
rect 1818 72638 1874 72640
rect 1818 72586 1820 72638
rect 1820 72586 1872 72638
rect 1872 72586 1874 72638
rect 1818 72584 1874 72586
rect 69717 72131 69773 72187
rect 1818 70958 1874 70960
rect 1818 70906 1820 70958
rect 1820 70906 1872 70958
rect 1872 70906 1874 70958
rect 1818 70904 1874 70906
rect 69841 70717 69897 70773
rect 1818 69278 1874 69280
rect 1818 69226 1820 69278
rect 1820 69226 1872 69278
rect 1872 69226 1874 69278
rect 1818 69224 1874 69226
rect 73702 69303 73758 69359
rect 1818 67598 1874 67600
rect 1818 67546 1820 67598
rect 1820 67546 1872 67598
rect 1872 67546 1874 67598
rect 1818 67544 1874 67546
rect 1818 65918 1874 65920
rect 1818 65866 1820 65918
rect 1820 65866 1872 65918
rect 1872 65866 1874 65918
rect 1818 65864 1874 65866
rect 1818 64238 1874 64240
rect 1818 64186 1820 64238
rect 1820 64186 1872 64238
rect 1872 64186 1874 64238
rect 1818 64184 1874 64186
rect 1818 62558 1874 62560
rect 1818 62506 1820 62558
rect 1820 62506 1872 62558
rect 1872 62506 1874 62558
rect 1818 62504 1874 62506
rect 1818 60878 1874 60880
rect 1818 60826 1820 60878
rect 1820 60826 1872 60878
rect 1872 60826 1874 60878
rect 1818 60824 1874 60826
rect 1818 59198 1874 59200
rect 1818 59146 1820 59198
rect 1820 59146 1872 59198
rect 1872 59146 1874 59198
rect 1818 59144 1874 59146
rect 1818 57518 1874 57520
rect 1818 57466 1820 57518
rect 1820 57466 1872 57518
rect 1872 57466 1874 57518
rect 1818 57464 1874 57466
rect 1818 55838 1874 55840
rect 1818 55786 1820 55838
rect 1820 55786 1872 55838
rect 1872 55786 1874 55838
rect 1818 55784 1874 55786
rect 1818 54158 1874 54160
rect 1818 54106 1820 54158
rect 1820 54106 1872 54158
rect 1872 54106 1874 54158
rect 1818 54104 1874 54106
rect 1818 52478 1874 52480
rect 1818 52426 1820 52478
rect 1820 52426 1872 52478
rect 1872 52426 1874 52478
rect 1818 52424 1874 52426
rect 1818 50798 1874 50800
rect 1818 50746 1820 50798
rect 1820 50746 1872 50798
rect 1872 50746 1874 50798
rect 1818 50744 1874 50746
rect 1818 49118 1874 49120
rect 1818 49066 1820 49118
rect 1820 49066 1872 49118
rect 1872 49066 1874 49118
rect 1818 49064 1874 49066
rect 1818 47438 1874 47440
rect 1818 47386 1820 47438
rect 1820 47386 1872 47438
rect 1872 47386 1874 47438
rect 1818 47384 1874 47386
rect 1818 45758 1874 45760
rect 1818 45706 1820 45758
rect 1820 45706 1872 45758
rect 1872 45706 1874 45758
rect 1818 45704 1874 45706
rect 1818 44078 1874 44080
rect 1818 44026 1820 44078
rect 1820 44026 1872 44078
rect 1872 44026 1874 44078
rect 1818 44024 1874 44026
rect 1818 42398 1874 42400
rect 1818 42346 1820 42398
rect 1820 42346 1872 42398
rect 1872 42346 1874 42398
rect 1818 42344 1874 42346
rect 1818 40718 1874 40720
rect 1818 40666 1820 40718
rect 1820 40666 1872 40718
rect 1872 40666 1874 40718
rect 1818 40664 1874 40666
rect 1818 39038 1874 39040
rect 1818 38986 1820 39038
rect 1820 38986 1872 39038
rect 1872 38986 1874 39038
rect 1818 38984 1874 38986
rect 1818 37358 1874 37360
rect 1818 37306 1820 37358
rect 1820 37306 1872 37358
rect 1872 37306 1874 37358
rect 1818 37304 1874 37306
rect 1818 35678 1874 35680
rect 1818 35626 1820 35678
rect 1820 35626 1872 35678
rect 1872 35626 1874 35678
rect 1818 35624 1874 35626
rect 14205 34141 14261 34197
rect 14939 34195 14995 34197
rect 14939 34143 14941 34195
rect 14941 34143 14993 34195
rect 14993 34143 14995 34195
rect 14939 34141 14995 34143
rect 13260 34070 13316 34126
rect 1818 33998 1874 34000
rect 1818 33946 1820 33998
rect 1820 33946 1872 33998
rect 1872 33946 1874 33998
rect 1818 33944 1874 33946
rect 13260 32942 13316 32998
rect 14205 32871 14261 32927
rect 14859 32925 14915 32927
rect 14859 32873 14861 32925
rect 14861 32873 14913 32925
rect 14913 32873 14915 32925
rect 14859 32871 14915 32873
rect 1818 32318 1874 32320
rect 1818 32266 1820 32318
rect 1820 32266 1872 32318
rect 1872 32266 1874 32318
rect 1818 32264 1874 32266
rect 14205 31313 14261 31369
rect 14779 31367 14835 31369
rect 14779 31315 14781 31367
rect 14781 31315 14833 31367
rect 14833 31315 14835 31367
rect 14779 31313 14835 31315
rect 13260 31242 13316 31298
rect 1818 30638 1874 30640
rect 1818 30586 1820 30638
rect 1820 30586 1872 30638
rect 1872 30586 1874 30638
rect 1818 30584 1874 30586
rect 13260 30114 13316 30170
rect 14205 30043 14261 30099
rect 14699 30097 14755 30099
rect 14699 30045 14701 30097
rect 14701 30045 14753 30097
rect 14753 30045 14755 30097
rect 14699 30043 14755 30045
rect 1818 28958 1874 28960
rect 1818 28906 1820 28958
rect 1820 28906 1872 28958
rect 1872 28906 1874 28958
rect 1818 28904 1874 28906
rect 14205 28485 14261 28541
rect 14619 28539 14675 28541
rect 14619 28487 14621 28539
rect 14621 28487 14673 28539
rect 14673 28487 14675 28539
rect 14619 28485 14675 28487
rect 13260 28414 13316 28470
rect 1818 27278 1874 27280
rect 1818 27226 1820 27278
rect 1820 27226 1872 27278
rect 1872 27226 1874 27278
rect 1818 27224 1874 27226
rect 13260 27286 13316 27342
rect 14205 27215 14261 27271
rect 14539 27269 14595 27271
rect 14539 27217 14541 27269
rect 14541 27217 14593 27269
rect 14593 27217 14595 27269
rect 14539 27215 14595 27217
rect 14205 25657 14261 25713
rect 1818 25598 1874 25600
rect 1818 25546 1820 25598
rect 1820 25546 1872 25598
rect 1872 25546 1874 25598
rect 1818 25544 1874 25546
rect 14459 25711 14515 25713
rect 14459 25659 14461 25711
rect 14461 25659 14513 25711
rect 14513 25659 14515 25711
rect 14459 25657 14515 25659
rect 13260 25586 13316 25642
rect 14342 25330 14398 25386
rect 1818 23918 1874 23920
rect 1818 23866 1820 23918
rect 1820 23866 1872 23918
rect 1872 23866 1874 23918
rect 1818 23864 1874 23866
rect 2565 22609 2621 22665
rect 1818 22238 1874 22240
rect 1818 22186 1820 22238
rect 1820 22186 1872 22238
rect 1872 22186 1874 22238
rect 1818 22184 1874 22186
rect 1818 20558 1874 20560
rect 1818 20506 1820 20558
rect 1820 20506 1872 20558
rect 1872 20506 1874 20558
rect 1818 20504 1874 20506
rect 1818 18878 1874 18880
rect 1818 18826 1820 18878
rect 1820 18826 1872 18878
rect 1872 18826 1874 18878
rect 1818 18824 1874 18826
rect 1818 17198 1874 17200
rect 1818 17146 1820 17198
rect 1820 17146 1872 17198
rect 1872 17146 1874 17198
rect 1818 17144 1874 17146
rect 1818 15518 1874 15520
rect 1818 15466 1820 15518
rect 1820 15466 1872 15518
rect 1872 15466 1874 15518
rect 1818 15464 1874 15466
rect 14258 15501 14314 15557
rect 1818 13838 1874 13840
rect 1818 13786 1820 13838
rect 1820 13786 1872 13838
rect 1872 13786 1874 13838
rect 1818 13784 1874 13786
rect 14258 12673 14314 12729
rect 1818 12158 1874 12160
rect 1818 12106 1820 12158
rect 1820 12106 1872 12158
rect 1872 12106 1874 12158
rect 1818 12104 1874 12106
rect 14258 11259 14314 11315
rect 1818 10478 1874 10480
rect 1818 10426 1820 10478
rect 1820 10426 1872 10478
rect 1872 10426 1874 10478
rect 1818 10424 1874 10426
rect 14258 9845 14314 9901
rect 1818 8798 1874 8800
rect 1818 8746 1820 8798
rect 1820 8746 1872 8798
rect 1872 8746 1874 8798
rect 1818 8744 1874 8746
rect 2778 7160 2834 7216
rect 1818 7118 1874 7120
rect 1818 7066 1820 7118
rect 1820 7066 1872 7118
rect 1872 7066 1874 7118
rect 1818 7064 1874 7066
rect 94176 75998 94232 76000
rect 94176 75946 94178 75998
rect 94178 75946 94230 75998
rect 94230 75946 94232 75998
rect 94176 75944 94232 75946
rect 94176 74318 94232 74320
rect 94176 74266 94178 74318
rect 94178 74266 94230 74318
rect 94230 74266 94232 74318
rect 94176 74264 94232 74266
rect 94176 72638 94232 72640
rect 94176 72586 94178 72638
rect 94178 72586 94230 72638
rect 94230 72586 94232 72638
rect 94176 72584 94232 72586
rect 81928 72131 81984 72187
rect 94176 70958 94232 70960
rect 94176 70906 94178 70958
rect 94178 70906 94230 70958
rect 94230 70906 94232 70958
rect 94176 70904 94232 70906
rect 81928 70717 81984 70773
rect 81928 69303 81984 69359
rect 94176 69278 94232 69280
rect 94176 69226 94178 69278
rect 94178 69226 94230 69278
rect 94230 69226 94232 69278
rect 94176 69224 94232 69226
rect 94176 67598 94232 67600
rect 94176 67546 94178 67598
rect 94178 67546 94230 67598
rect 94230 67546 94232 67598
rect 94176 67544 94232 67546
rect 94176 65918 94232 65920
rect 94176 65866 94178 65918
rect 94178 65866 94230 65918
rect 94230 65866 94232 65918
rect 94176 65864 94232 65866
rect 94176 64238 94232 64240
rect 94176 64186 94178 64238
rect 94178 64186 94230 64238
rect 94230 64186 94232 64238
rect 94176 64184 94232 64186
rect 94176 62558 94232 62560
rect 94176 62506 94178 62558
rect 94178 62506 94230 62558
rect 94230 62506 94232 62558
rect 94176 62504 94232 62506
rect 94176 60878 94232 60880
rect 94176 60826 94178 60878
rect 94178 60826 94230 60878
rect 94230 60826 94232 60878
rect 94176 60824 94232 60826
rect 93429 59367 93485 59423
rect 94176 59198 94232 59200
rect 94176 59146 94178 59198
rect 94178 59146 94230 59198
rect 94230 59146 94232 59198
rect 94176 59144 94232 59146
rect 94176 57518 94232 57520
rect 94176 57466 94178 57518
rect 94178 57466 94230 57518
rect 94230 57466 94232 57518
rect 94176 57464 94232 57466
rect 94176 55838 94232 55840
rect 94176 55786 94178 55838
rect 94178 55786 94230 55838
rect 94230 55786 94232 55838
rect 94176 55784 94232 55786
rect 94176 54158 94232 54160
rect 94176 54106 94178 54158
rect 94178 54106 94230 54158
rect 94230 54106 94232 54158
rect 94176 54104 94232 54106
rect 94176 52478 94232 52480
rect 94176 52426 94178 52478
rect 94178 52426 94230 52478
rect 94230 52426 94232 52478
rect 94176 52424 94232 52426
rect 94176 50798 94232 50800
rect 94176 50746 94178 50798
rect 94178 50746 94230 50798
rect 94230 50746 94232 50798
rect 94176 50744 94232 50746
rect 94176 49118 94232 49120
rect 94176 49066 94178 49118
rect 94178 49066 94230 49118
rect 94230 49066 94232 49118
rect 94176 49064 94232 49066
rect 94176 47438 94232 47440
rect 94176 47386 94178 47438
rect 94178 47386 94230 47438
rect 94230 47386 94232 47438
rect 94176 47384 94232 47386
rect 94176 45758 94232 45760
rect 94176 45706 94178 45758
rect 94178 45706 94230 45758
rect 94230 45706 94232 45758
rect 94176 45704 94232 45706
rect 94176 44078 94232 44080
rect 94176 44026 94178 44078
rect 94178 44026 94230 44078
rect 94230 44026 94232 44078
rect 94176 44024 94232 44026
rect 94176 42398 94232 42400
rect 94176 42346 94178 42398
rect 94178 42346 94230 42398
rect 94230 42346 94232 42398
rect 94176 42344 94232 42346
rect 94176 40718 94232 40720
rect 94176 40666 94178 40718
rect 94178 40666 94230 40718
rect 94230 40666 94232 40718
rect 94176 40664 94232 40666
rect 94176 39038 94232 39040
rect 94176 38986 94178 39038
rect 94178 38986 94230 39038
rect 94230 38986 94232 39038
rect 94176 38984 94232 38986
rect 94176 37358 94232 37360
rect 94176 37306 94178 37358
rect 94178 37306 94230 37358
rect 94230 37306 94232 37358
rect 94176 37304 94232 37306
rect 94176 35678 94232 35680
rect 94176 35626 94178 35678
rect 94178 35626 94230 35678
rect 94230 35626 94232 35678
rect 94176 35624 94232 35626
rect 94176 33998 94232 34000
rect 94176 33946 94178 33998
rect 94178 33946 94230 33998
rect 94230 33946 94232 33998
rect 94176 33944 94232 33946
rect 94176 32318 94232 32320
rect 94176 32266 94178 32318
rect 94178 32266 94230 32318
rect 94230 32266 94232 32318
rect 94176 32264 94232 32266
rect 94176 30638 94232 30640
rect 94176 30586 94178 30638
rect 94178 30586 94230 30638
rect 94230 30586 94232 30638
rect 94176 30584 94232 30586
rect 94176 28958 94232 28960
rect 94176 28906 94178 28958
rect 94178 28906 94230 28958
rect 94230 28906 94232 28958
rect 94176 28904 94232 28906
rect 94176 27278 94232 27280
rect 94176 27226 94178 27278
rect 94178 27226 94230 27278
rect 94230 27226 94232 27278
rect 94176 27224 94232 27226
rect 94176 25598 94232 25600
rect 94176 25546 94178 25598
rect 94178 25546 94230 25598
rect 94230 25546 94232 25598
rect 94176 25544 94232 25546
rect 94176 23918 94232 23920
rect 94176 23866 94178 23918
rect 94178 23866 94230 23918
rect 94230 23866 94232 23918
rect 94176 23864 94232 23866
rect 94176 22238 94232 22240
rect 94176 22186 94178 22238
rect 94178 22186 94230 22238
rect 94230 22186 94232 22238
rect 94176 22184 94232 22186
rect 94176 20558 94232 20560
rect 94176 20506 94178 20558
rect 94178 20506 94230 20558
rect 94230 20506 94232 20558
rect 94176 20504 94232 20506
rect 94176 18878 94232 18880
rect 94176 18826 94178 18878
rect 94178 18826 94230 18878
rect 94230 18826 94232 18878
rect 94176 18824 94232 18826
rect 94176 17198 94232 17200
rect 94176 17146 94178 17198
rect 94178 17146 94230 17198
rect 94230 17146 94232 17198
rect 94176 17144 94232 17146
rect 81844 16814 81900 16870
rect 82926 16558 82982 16614
rect 81643 16541 81699 16543
rect 81643 16489 81645 16541
rect 81645 16489 81697 16541
rect 81697 16489 81699 16541
rect 81643 16487 81699 16489
rect 81981 16487 82037 16543
rect 22400 15501 22456 15557
rect 94176 15518 94232 15520
rect 94176 15466 94178 15518
rect 94178 15466 94230 15518
rect 94230 15466 94232 15518
rect 94176 15464 94232 15466
rect 81563 14983 81619 14985
rect 81563 14931 81565 14983
rect 81565 14931 81617 14983
rect 81617 14931 81619 14983
rect 81563 14929 81619 14931
rect 81981 14929 82037 14985
rect 82926 14858 82982 14914
rect 82926 13730 82982 13786
rect 81483 13713 81539 13715
rect 81483 13661 81485 13713
rect 81485 13661 81537 13713
rect 81537 13661 81539 13713
rect 81483 13659 81539 13661
rect 94176 13838 94232 13840
rect 94176 13786 94178 13838
rect 94178 13786 94230 13838
rect 94230 13786 94232 13838
rect 94176 13784 94232 13786
rect 81981 13659 82037 13715
rect 26103 12673 26159 12729
rect 81403 12155 81459 12157
rect 81403 12103 81405 12155
rect 81405 12103 81457 12155
rect 81457 12103 81459 12155
rect 81403 12101 81459 12103
rect 81981 12101 82037 12157
rect 94176 12158 94232 12160
rect 94176 12106 94178 12158
rect 94178 12106 94230 12158
rect 94230 12106 94232 12158
rect 94176 12104 94232 12106
rect 82926 12030 82982 12086
rect 26351 11259 26407 11315
rect 26227 9845 26283 9901
rect 82926 10902 82982 10958
rect 81323 10885 81379 10887
rect 81323 10833 81325 10885
rect 81325 10833 81377 10885
rect 81377 10833 81379 10885
rect 81323 10831 81379 10833
rect 81981 10831 82037 10887
rect 28210 10811 28266 10813
rect 28210 10759 28212 10811
rect 28212 10759 28264 10811
rect 28264 10759 28266 10811
rect 28210 10757 28266 10759
rect 29458 10811 29514 10813
rect 29458 10759 29460 10811
rect 29460 10759 29512 10811
rect 29512 10759 29514 10811
rect 29458 10757 29514 10759
rect 30706 10811 30762 10813
rect 30706 10759 30708 10811
rect 30708 10759 30760 10811
rect 30760 10759 30762 10811
rect 30706 10757 30762 10759
rect 31954 10811 32010 10813
rect 31954 10759 31956 10811
rect 31956 10759 32008 10811
rect 32008 10759 32010 10811
rect 31954 10757 32010 10759
rect 33202 10811 33258 10813
rect 33202 10759 33204 10811
rect 33204 10759 33256 10811
rect 33256 10759 33258 10811
rect 33202 10757 33258 10759
rect 34450 10811 34506 10813
rect 34450 10759 34452 10811
rect 34452 10759 34504 10811
rect 34504 10759 34506 10811
rect 34450 10757 34506 10759
rect 35698 10811 35754 10813
rect 35698 10759 35700 10811
rect 35700 10759 35752 10811
rect 35752 10759 35754 10811
rect 35698 10757 35754 10759
rect 36946 10811 37002 10813
rect 36946 10759 36948 10811
rect 36948 10759 37000 10811
rect 37000 10759 37002 10811
rect 36946 10757 37002 10759
rect 38194 10811 38250 10813
rect 38194 10759 38196 10811
rect 38196 10759 38248 10811
rect 38248 10759 38250 10811
rect 38194 10757 38250 10759
rect 39442 10811 39498 10813
rect 39442 10759 39444 10811
rect 39444 10759 39496 10811
rect 39496 10759 39498 10811
rect 39442 10757 39498 10759
rect 40690 10811 40746 10813
rect 40690 10759 40692 10811
rect 40692 10759 40744 10811
rect 40744 10759 40746 10811
rect 40690 10757 40746 10759
rect 41938 10811 41994 10813
rect 41938 10759 41940 10811
rect 41940 10759 41992 10811
rect 41992 10759 41994 10811
rect 41938 10757 41994 10759
rect 43186 10811 43242 10813
rect 43186 10759 43188 10811
rect 43188 10759 43240 10811
rect 43240 10759 43242 10811
rect 43186 10757 43242 10759
rect 44434 10811 44490 10813
rect 44434 10759 44436 10811
rect 44436 10759 44488 10811
rect 44488 10759 44490 10811
rect 44434 10757 44490 10759
rect 45682 10811 45738 10813
rect 45682 10759 45684 10811
rect 45684 10759 45736 10811
rect 45736 10759 45738 10811
rect 45682 10757 45738 10759
rect 46930 10811 46986 10813
rect 46930 10759 46932 10811
rect 46932 10759 46984 10811
rect 46984 10759 46986 10811
rect 46930 10757 46986 10759
rect 48178 10811 48234 10813
rect 48178 10759 48180 10811
rect 48180 10759 48232 10811
rect 48232 10759 48234 10811
rect 48178 10757 48234 10759
rect 49426 10811 49482 10813
rect 49426 10759 49428 10811
rect 49428 10759 49480 10811
rect 49480 10759 49482 10811
rect 49426 10757 49482 10759
rect 50674 10811 50730 10813
rect 50674 10759 50676 10811
rect 50676 10759 50728 10811
rect 50728 10759 50730 10811
rect 50674 10757 50730 10759
rect 51922 10811 51978 10813
rect 51922 10759 51924 10811
rect 51924 10759 51976 10811
rect 51976 10759 51978 10811
rect 51922 10757 51978 10759
rect 53170 10811 53226 10813
rect 53170 10759 53172 10811
rect 53172 10759 53224 10811
rect 53224 10759 53226 10811
rect 53170 10757 53226 10759
rect 54418 10811 54474 10813
rect 54418 10759 54420 10811
rect 54420 10759 54472 10811
rect 54472 10759 54474 10811
rect 54418 10757 54474 10759
rect 55666 10811 55722 10813
rect 55666 10759 55668 10811
rect 55668 10759 55720 10811
rect 55720 10759 55722 10811
rect 55666 10757 55722 10759
rect 56914 10811 56970 10813
rect 56914 10759 56916 10811
rect 56916 10759 56968 10811
rect 56968 10759 56970 10811
rect 56914 10757 56970 10759
rect 58162 10811 58218 10813
rect 58162 10759 58164 10811
rect 58164 10759 58216 10811
rect 58216 10759 58218 10811
rect 58162 10757 58218 10759
rect 59410 10811 59466 10813
rect 59410 10759 59412 10811
rect 59412 10759 59464 10811
rect 59464 10759 59466 10811
rect 59410 10757 59466 10759
rect 60658 10811 60714 10813
rect 60658 10759 60660 10811
rect 60660 10759 60712 10811
rect 60712 10759 60714 10811
rect 60658 10757 60714 10759
rect 61906 10811 61962 10813
rect 61906 10759 61908 10811
rect 61908 10759 61960 10811
rect 61960 10759 61962 10811
rect 61906 10757 61962 10759
rect 63154 10811 63210 10813
rect 63154 10759 63156 10811
rect 63156 10759 63208 10811
rect 63208 10759 63210 10811
rect 63154 10757 63210 10759
rect 64402 10811 64458 10813
rect 64402 10759 64404 10811
rect 64404 10759 64456 10811
rect 64456 10759 64458 10811
rect 64402 10757 64458 10759
rect 65650 10811 65706 10813
rect 65650 10759 65652 10811
rect 65652 10759 65704 10811
rect 65704 10759 65706 10811
rect 65650 10757 65706 10759
rect 66898 10811 66954 10813
rect 66898 10759 66900 10811
rect 66900 10759 66952 10811
rect 66952 10759 66954 10811
rect 66898 10757 66954 10759
rect 94176 10478 94232 10480
rect 94176 10426 94178 10478
rect 94178 10426 94230 10478
rect 94230 10426 94232 10478
rect 94176 10424 94232 10426
rect 81243 9327 81299 9329
rect 81243 9275 81245 9327
rect 81245 9275 81297 9327
rect 81297 9275 81299 9327
rect 81243 9273 81299 9275
rect 81981 9273 82037 9329
rect 82926 9202 82982 9258
rect 94176 8798 94232 8800
rect 94176 8746 94178 8798
rect 94178 8746 94230 8798
rect 94230 8746 94232 8798
rect 94176 8744 94232 8746
rect 82926 8074 82982 8130
rect 81163 8057 81219 8059
rect 81163 8005 81165 8057
rect 81165 8005 81217 8057
rect 81217 8005 81219 8057
rect 81163 8003 81219 8005
rect 81981 8003 82037 8059
rect 94176 7118 94232 7120
rect 94176 7066 94178 7118
rect 94178 7066 94230 7118
rect 94230 7066 94232 7118
rect 94176 7064 94232 7066
rect 5999 5565 6055 5621
rect 2778 5460 2834 5516
rect 1818 5438 1874 5440
rect 1818 5386 1820 5438
rect 1820 5386 1872 5438
rect 1872 5386 1874 5438
rect 1818 5384 1874 5386
rect 1818 3758 1874 3760
rect 1818 3706 1820 3758
rect 1820 3706 1872 3758
rect 1872 3706 1874 3758
rect 1818 3704 1874 3706
rect 94176 5438 94232 5440
rect 94176 5386 94178 5438
rect 94178 5386 94230 5438
rect 94230 5386 94232 5438
rect 94176 5384 94232 5386
rect 94176 3758 94232 3760
rect 94176 3706 94178 3758
rect 94178 3706 94230 3758
rect 94230 3706 94232 3758
rect 94176 3704 94232 3706
rect 15596 2924 15652 2980
rect 16764 2924 16820 2980
rect 17932 2924 17988 2980
rect 19100 2924 19156 2980
rect 20268 2924 20324 2980
rect 21436 2924 21492 2980
rect 22604 2924 22660 2980
rect 23772 2924 23828 2980
rect 24940 2924 24996 2980
rect 26108 2924 26164 2980
rect 27276 2924 27332 2980
rect 28444 2924 28500 2980
rect 29612 2924 29668 2980
rect 30780 2924 30836 2980
rect 31948 2924 32004 2980
rect 33116 2924 33172 2980
rect 34284 2924 34340 2980
rect 35452 2924 35508 2980
rect 36620 2924 36676 2980
rect 37788 2924 37844 2980
rect 38956 2924 39012 2980
rect 40124 2924 40180 2980
rect 41292 2924 41348 2980
rect 42460 2924 42516 2980
rect 43628 2924 43684 2980
rect 44796 2924 44852 2980
rect 45964 2924 46020 2980
rect 47132 2924 47188 2980
rect 48300 2924 48356 2980
rect 49468 2924 49524 2980
rect 50636 2924 50692 2980
rect 51804 2924 51860 2980
rect 52972 2924 53028 2980
rect 54140 2924 54196 2980
rect 55308 2924 55364 2980
rect 56476 2924 56532 2980
rect 57644 2924 57700 2980
rect 14342 2668 14398 2724
rect 1818 2078 1874 2080
rect 1818 2026 1820 2078
rect 1820 2026 1872 2078
rect 1872 2026 1874 2078
rect 1818 2024 1874 2026
rect 94176 2078 94232 2080
rect 94176 2026 94178 2078
rect 94178 2026 94230 2078
rect 94230 2026 94232 2078
rect 94176 2024 94232 2026
rect 2154 1742 2210 1744
rect 2154 1690 2156 1742
rect 2156 1690 2208 1742
rect 2208 1690 2210 1742
rect 2154 1688 2210 1690
rect 3834 1742 3890 1744
rect 3834 1690 3836 1742
rect 3836 1690 3888 1742
rect 3888 1690 3890 1742
rect 3834 1688 3890 1690
rect 5514 1742 5570 1744
rect 5514 1690 5516 1742
rect 5516 1690 5568 1742
rect 5568 1690 5570 1742
rect 5514 1688 5570 1690
rect 7194 1742 7250 1744
rect 7194 1690 7196 1742
rect 7196 1690 7248 1742
rect 7248 1690 7250 1742
rect 7194 1688 7250 1690
rect 8874 1742 8930 1744
rect 8874 1690 8876 1742
rect 8876 1690 8928 1742
rect 8928 1690 8930 1742
rect 8874 1688 8930 1690
rect 10554 1742 10610 1744
rect 10554 1690 10556 1742
rect 10556 1690 10608 1742
rect 10608 1690 10610 1742
rect 10554 1688 10610 1690
rect 12234 1742 12290 1744
rect 12234 1690 12236 1742
rect 12236 1690 12288 1742
rect 12288 1690 12290 1742
rect 12234 1688 12290 1690
rect 13914 1742 13970 1744
rect 13914 1690 13916 1742
rect 13916 1690 13968 1742
rect 13968 1690 13970 1742
rect 13914 1688 13970 1690
rect 15594 1742 15650 1744
rect 15594 1690 15596 1742
rect 15596 1690 15648 1742
rect 15648 1690 15650 1742
rect 15594 1688 15650 1690
rect 17274 1742 17330 1744
rect 17274 1690 17276 1742
rect 17276 1690 17328 1742
rect 17328 1690 17330 1742
rect 17274 1688 17330 1690
rect 18954 1742 19010 1744
rect 18954 1690 18956 1742
rect 18956 1690 19008 1742
rect 19008 1690 19010 1742
rect 18954 1688 19010 1690
rect 20634 1742 20690 1744
rect 20634 1690 20636 1742
rect 20636 1690 20688 1742
rect 20688 1690 20690 1742
rect 20634 1688 20690 1690
rect 22314 1742 22370 1744
rect 22314 1690 22316 1742
rect 22316 1690 22368 1742
rect 22368 1690 22370 1742
rect 22314 1688 22370 1690
rect 23994 1742 24050 1744
rect 23994 1690 23996 1742
rect 23996 1690 24048 1742
rect 24048 1690 24050 1742
rect 23994 1688 24050 1690
rect 25674 1742 25730 1744
rect 25674 1690 25676 1742
rect 25676 1690 25728 1742
rect 25728 1690 25730 1742
rect 25674 1688 25730 1690
rect 27354 1742 27410 1744
rect 27354 1690 27356 1742
rect 27356 1690 27408 1742
rect 27408 1690 27410 1742
rect 27354 1688 27410 1690
rect 29034 1742 29090 1744
rect 29034 1690 29036 1742
rect 29036 1690 29088 1742
rect 29088 1690 29090 1742
rect 29034 1688 29090 1690
rect 30714 1742 30770 1744
rect 30714 1690 30716 1742
rect 30716 1690 30768 1742
rect 30768 1690 30770 1742
rect 30714 1688 30770 1690
rect 32394 1742 32450 1744
rect 32394 1690 32396 1742
rect 32396 1690 32448 1742
rect 32448 1690 32450 1742
rect 32394 1688 32450 1690
rect 34074 1742 34130 1744
rect 34074 1690 34076 1742
rect 34076 1690 34128 1742
rect 34128 1690 34130 1742
rect 34074 1688 34130 1690
rect 35754 1742 35810 1744
rect 35754 1690 35756 1742
rect 35756 1690 35808 1742
rect 35808 1690 35810 1742
rect 35754 1688 35810 1690
rect 37434 1742 37490 1744
rect 37434 1690 37436 1742
rect 37436 1690 37488 1742
rect 37488 1690 37490 1742
rect 37434 1688 37490 1690
rect 39114 1742 39170 1744
rect 39114 1690 39116 1742
rect 39116 1690 39168 1742
rect 39168 1690 39170 1742
rect 39114 1688 39170 1690
rect 40794 1742 40850 1744
rect 40794 1690 40796 1742
rect 40796 1690 40848 1742
rect 40848 1690 40850 1742
rect 40794 1688 40850 1690
rect 42474 1742 42530 1744
rect 42474 1690 42476 1742
rect 42476 1690 42528 1742
rect 42528 1690 42530 1742
rect 42474 1688 42530 1690
rect 44154 1742 44210 1744
rect 44154 1690 44156 1742
rect 44156 1690 44208 1742
rect 44208 1690 44210 1742
rect 44154 1688 44210 1690
rect 45834 1742 45890 1744
rect 45834 1690 45836 1742
rect 45836 1690 45888 1742
rect 45888 1690 45890 1742
rect 45834 1688 45890 1690
rect 47514 1742 47570 1744
rect 47514 1690 47516 1742
rect 47516 1690 47568 1742
rect 47568 1690 47570 1742
rect 47514 1688 47570 1690
rect 49194 1742 49250 1744
rect 49194 1690 49196 1742
rect 49196 1690 49248 1742
rect 49248 1690 49250 1742
rect 49194 1688 49250 1690
rect 50874 1742 50930 1744
rect 50874 1690 50876 1742
rect 50876 1690 50928 1742
rect 50928 1690 50930 1742
rect 50874 1688 50930 1690
rect 52554 1742 52610 1744
rect 52554 1690 52556 1742
rect 52556 1690 52608 1742
rect 52608 1690 52610 1742
rect 52554 1688 52610 1690
rect 54234 1742 54290 1744
rect 54234 1690 54236 1742
rect 54236 1690 54288 1742
rect 54288 1690 54290 1742
rect 54234 1688 54290 1690
rect 55914 1742 55970 1744
rect 55914 1690 55916 1742
rect 55916 1690 55968 1742
rect 55968 1690 55970 1742
rect 55914 1688 55970 1690
rect 57594 1742 57650 1744
rect 57594 1690 57596 1742
rect 57596 1690 57648 1742
rect 57648 1690 57650 1742
rect 57594 1688 57650 1690
rect 59274 1742 59330 1744
rect 59274 1690 59276 1742
rect 59276 1690 59328 1742
rect 59328 1690 59330 1742
rect 59274 1688 59330 1690
rect 60954 1742 61010 1744
rect 60954 1690 60956 1742
rect 60956 1690 61008 1742
rect 61008 1690 61010 1742
rect 60954 1688 61010 1690
rect 62634 1742 62690 1744
rect 62634 1690 62636 1742
rect 62636 1690 62688 1742
rect 62688 1690 62690 1742
rect 62634 1688 62690 1690
rect 64314 1742 64370 1744
rect 64314 1690 64316 1742
rect 64316 1690 64368 1742
rect 64368 1690 64370 1742
rect 64314 1688 64370 1690
rect 65994 1742 66050 1744
rect 65994 1690 65996 1742
rect 65996 1690 66048 1742
rect 66048 1690 66050 1742
rect 65994 1688 66050 1690
rect 67674 1742 67730 1744
rect 67674 1690 67676 1742
rect 67676 1690 67728 1742
rect 67728 1690 67730 1742
rect 67674 1688 67730 1690
rect 69354 1742 69410 1744
rect 69354 1690 69356 1742
rect 69356 1690 69408 1742
rect 69408 1690 69410 1742
rect 69354 1688 69410 1690
rect 71034 1742 71090 1744
rect 71034 1690 71036 1742
rect 71036 1690 71088 1742
rect 71088 1690 71090 1742
rect 71034 1688 71090 1690
rect 72714 1742 72770 1744
rect 72714 1690 72716 1742
rect 72716 1690 72768 1742
rect 72768 1690 72770 1742
rect 72714 1688 72770 1690
rect 74394 1742 74450 1744
rect 74394 1690 74396 1742
rect 74396 1690 74448 1742
rect 74448 1690 74450 1742
rect 74394 1688 74450 1690
rect 76074 1742 76130 1744
rect 76074 1690 76076 1742
rect 76076 1690 76128 1742
rect 76128 1690 76130 1742
rect 76074 1688 76130 1690
rect 77754 1742 77810 1744
rect 77754 1690 77756 1742
rect 77756 1690 77808 1742
rect 77808 1690 77810 1742
rect 77754 1688 77810 1690
rect 79434 1742 79490 1744
rect 79434 1690 79436 1742
rect 79436 1690 79488 1742
rect 79488 1690 79490 1742
rect 79434 1688 79490 1690
rect 81114 1742 81170 1744
rect 81114 1690 81116 1742
rect 81116 1690 81168 1742
rect 81168 1690 81170 1742
rect 81114 1688 81170 1690
rect 82794 1742 82850 1744
rect 82794 1690 82796 1742
rect 82796 1690 82848 1742
rect 82848 1690 82850 1742
rect 82794 1688 82850 1690
rect 84474 1742 84530 1744
rect 84474 1690 84476 1742
rect 84476 1690 84528 1742
rect 84528 1690 84530 1742
rect 84474 1688 84530 1690
rect 86154 1742 86210 1744
rect 86154 1690 86156 1742
rect 86156 1690 86208 1742
rect 86208 1690 86210 1742
rect 86154 1688 86210 1690
rect 87834 1742 87890 1744
rect 87834 1690 87836 1742
rect 87836 1690 87888 1742
rect 87888 1690 87890 1742
rect 87834 1688 87890 1690
rect 89514 1742 89570 1744
rect 89514 1690 89516 1742
rect 89516 1690 89568 1742
rect 89568 1690 89570 1742
rect 89514 1688 89570 1690
rect 91194 1742 91250 1744
rect 91194 1690 91196 1742
rect 91196 1690 91248 1742
rect 91248 1690 91250 1742
rect 91194 1688 91250 1690
rect 92874 1742 92930 1744
rect 92874 1690 92876 1742
rect 92876 1690 92928 1742
rect 92928 1690 92930 1742
rect 92874 1688 92930 1690
<< metal3 >>
rect 272 79222 95684 79228
rect 272 79158 278 79222
rect 342 79158 414 79222
rect 478 79158 550 79222
rect 614 79158 95342 79222
rect 95406 79158 95478 79222
rect 95542 79158 95614 79222
rect 95678 79158 95684 79222
rect 272 79086 95684 79158
rect 272 79022 278 79086
rect 342 79022 414 79086
rect 478 79022 550 79086
rect 614 79022 95342 79086
rect 95406 79022 95478 79086
rect 95542 79022 95614 79086
rect 95678 79022 95684 79086
rect 272 78950 95684 79022
rect 272 78886 278 78950
rect 342 78886 414 78950
rect 478 78886 550 78950
rect 614 78886 78886 78950
rect 78950 78886 82150 78950
rect 82214 78886 95342 78950
rect 95406 78886 95478 78950
rect 95542 78886 95614 78950
rect 95678 78886 95684 78950
rect 272 78880 95684 78886
rect 952 78542 95004 78548
rect 952 78478 958 78542
rect 1022 78478 1094 78542
rect 1158 78478 1230 78542
rect 1294 78478 94662 78542
rect 94726 78478 94798 78542
rect 94862 78478 94934 78542
rect 94998 78478 95004 78542
rect 952 78406 95004 78478
rect 952 78342 958 78406
rect 1022 78342 1094 78406
rect 1158 78342 1230 78406
rect 1294 78342 94662 78406
rect 94726 78342 94798 78406
rect 94862 78342 94934 78406
rect 94998 78342 95004 78406
rect 952 78270 95004 78342
rect 952 78206 958 78270
rect 1022 78206 1094 78270
rect 1158 78206 1230 78270
rect 1294 78206 2182 78270
rect 2246 78206 3950 78270
rect 4014 78206 5446 78270
rect 5510 78206 7214 78270
rect 7278 78206 8982 78270
rect 9046 78206 10478 78270
rect 10542 78206 12246 78270
rect 12310 78206 14014 78270
rect 14078 78206 15646 78270
rect 15710 78206 17414 78270
rect 17478 78206 18910 78270
rect 18974 78206 20678 78270
rect 20742 78206 22174 78270
rect 22238 78206 23942 78270
rect 24006 78206 25710 78270
rect 25774 78206 27478 78270
rect 27542 78206 28974 78270
rect 29038 78206 30878 78270
rect 30942 78206 32510 78270
rect 32574 78206 34142 78270
rect 34206 78206 35502 78270
rect 35566 78206 37406 78270
rect 37470 78206 39174 78270
rect 39238 78206 40534 78270
rect 40598 78206 42438 78270
rect 42502 78206 44206 78270
rect 44270 78206 45838 78270
rect 45902 78206 47470 78270
rect 47534 78206 49238 78270
rect 49302 78206 50734 78270
rect 50798 78206 52638 78270
rect 52702 78206 54134 78270
rect 54198 78206 55902 78270
rect 55966 78206 57670 78270
rect 57734 78206 59166 78270
rect 59230 78206 60934 78270
rect 60998 78206 62702 78270
rect 62766 78206 64062 78270
rect 64126 78206 65966 78270
rect 66030 78206 67734 78270
rect 67798 78206 69230 78270
rect 69294 78206 71134 78270
rect 71198 78206 72766 78270
rect 72830 78206 74398 78270
rect 74462 78206 76166 78270
rect 76230 78206 77662 78270
rect 77726 78206 79294 78270
rect 79358 78206 81198 78270
rect 81262 78206 82694 78270
rect 82758 78206 84462 78270
rect 84526 78206 86230 78270
rect 86294 78206 87726 78270
rect 87790 78206 89630 78270
rect 89694 78206 91262 78270
rect 91326 78206 92894 78270
rect 92958 78206 94662 78270
rect 94726 78206 94798 78270
rect 94862 78206 94934 78270
rect 94998 78206 95004 78270
rect 952 78200 95004 78206
rect 2040 77862 2252 77868
rect 2040 77808 2182 77862
rect 2040 77752 2154 77808
rect 2246 77798 2252 77862
rect 2210 77752 2252 77798
rect 2040 77656 2252 77752
rect 3808 77862 4020 77868
rect 3808 77808 3950 77862
rect 3808 77752 3834 77808
rect 3890 77798 3950 77808
rect 4014 77798 4020 77862
rect 3890 77752 4020 77798
rect 3808 77656 4020 77752
rect 5440 77862 5652 77868
rect 5440 77798 5446 77862
rect 5510 77808 5652 77862
rect 5510 77798 5514 77808
rect 5440 77752 5514 77798
rect 5570 77752 5652 77808
rect 5440 77656 5652 77752
rect 7072 77862 7284 77868
rect 7072 77808 7214 77862
rect 7072 77752 7194 77808
rect 7278 77798 7284 77862
rect 7250 77752 7284 77798
rect 7072 77656 7284 77752
rect 8840 77862 9052 77868
rect 8840 77808 8982 77862
rect 8840 77752 8874 77808
rect 8930 77798 8982 77808
rect 9046 77798 9052 77862
rect 8930 77752 9052 77798
rect 8840 77656 9052 77752
rect 10472 77862 10684 77868
rect 10472 77798 10478 77862
rect 10542 77808 10684 77862
rect 10542 77798 10554 77808
rect 10472 77752 10554 77798
rect 10610 77752 10684 77808
rect 10472 77656 10684 77752
rect 12104 77862 12316 77868
rect 12104 77808 12246 77862
rect 12104 77752 12234 77808
rect 12310 77798 12316 77862
rect 12290 77752 12316 77798
rect 12104 77656 12316 77752
rect 13872 77862 14084 77868
rect 13872 77808 14014 77862
rect 13872 77752 13914 77808
rect 13970 77798 14014 77808
rect 14078 77798 14084 77862
rect 13970 77752 14084 77798
rect 13872 77656 14084 77752
rect 15504 77862 15716 77868
rect 15504 77808 15646 77862
rect 15504 77752 15594 77808
rect 15710 77798 15716 77862
rect 15650 77752 15716 77798
rect 15504 77656 15716 77752
rect 17136 77862 17484 77868
rect 17136 77808 17414 77862
rect 17136 77752 17274 77808
rect 17330 77798 17414 77808
rect 17478 77798 17484 77862
rect 17330 77752 17484 77798
rect 17136 77656 17484 77752
rect 18904 77862 19116 77868
rect 18904 77798 18910 77862
rect 18974 77808 19116 77862
rect 18904 77752 18954 77798
rect 19010 77752 19116 77808
rect 18904 77656 19116 77752
rect 20536 77862 20748 77868
rect 20536 77808 20678 77862
rect 20536 77752 20634 77808
rect 20742 77798 20748 77862
rect 20690 77752 20748 77798
rect 20536 77656 20748 77752
rect 22168 77862 22516 77868
rect 22168 77798 22174 77862
rect 22238 77808 22516 77862
rect 22238 77798 22314 77808
rect 22168 77752 22314 77798
rect 22370 77752 22516 77808
rect 22168 77656 22516 77752
rect 23936 77862 24148 77868
rect 23936 77798 23942 77862
rect 24006 77808 24148 77862
rect 23936 77752 23994 77798
rect 24050 77752 24148 77808
rect 23936 77656 24148 77752
rect 25568 77862 25780 77868
rect 25568 77808 25710 77862
rect 25568 77752 25674 77808
rect 25774 77798 25780 77862
rect 25730 77752 25780 77798
rect 25568 77656 25780 77752
rect 27200 77862 27548 77868
rect 27200 77808 27478 77862
rect 27200 77752 27354 77808
rect 27410 77798 27478 77808
rect 27542 77798 27548 77862
rect 27410 77752 27548 77798
rect 27200 77656 27548 77752
rect 28968 77862 29180 77868
rect 28968 77798 28974 77862
rect 29038 77808 29180 77862
rect 28968 77752 29034 77798
rect 29090 77752 29180 77808
rect 28968 77732 29180 77752
rect 30600 77862 30948 77868
rect 30600 77808 30878 77862
rect 30600 77752 30714 77808
rect 30770 77798 30878 77808
rect 30942 77798 30948 77862
rect 30770 77792 30948 77798
rect 32368 77862 32580 77868
rect 32368 77808 32510 77862
rect 30770 77752 30812 77792
rect 28968 77726 29860 77732
rect 28968 77662 29790 77726
rect 29854 77662 29860 77726
rect 28968 77656 29860 77662
rect 30600 77656 30812 77752
rect 32368 77752 32394 77808
rect 32450 77798 32510 77808
rect 32574 77798 32580 77862
rect 32450 77752 32580 77798
rect 32368 77656 32580 77752
rect 34000 77862 34212 77868
rect 34000 77808 34142 77862
rect 34000 77752 34074 77808
rect 34130 77798 34142 77808
rect 34206 77798 34212 77862
rect 34130 77752 34212 77798
rect 35496 77862 35844 77868
rect 35496 77798 35502 77862
rect 35566 77808 35844 77862
rect 35566 77798 35754 77808
rect 35496 77792 35754 77798
rect 34000 77656 34212 77752
rect 35632 77752 35754 77792
rect 35810 77752 35844 77808
rect 35632 77656 35844 77752
rect 37400 77862 37612 77868
rect 37400 77798 37406 77862
rect 37470 77808 37612 77862
rect 37400 77752 37434 77798
rect 37490 77752 37612 77808
rect 37400 77656 37612 77752
rect 39032 77862 39244 77868
rect 39032 77808 39174 77862
rect 39032 77752 39114 77808
rect 39170 77798 39174 77808
rect 39238 77798 39244 77862
rect 39170 77752 39244 77798
rect 40528 77862 40876 77868
rect 40528 77798 40534 77862
rect 40598 77808 40876 77862
rect 40598 77798 40794 77808
rect 40528 77792 40794 77798
rect 39032 77656 39244 77752
rect 40664 77752 40794 77792
rect 40850 77752 40876 77808
rect 40664 77656 40876 77752
rect 42432 77862 42644 77868
rect 42432 77798 42438 77862
rect 42502 77808 42644 77862
rect 42432 77752 42474 77798
rect 42530 77752 42644 77808
rect 42432 77656 42644 77752
rect 44064 77862 44276 77868
rect 44064 77808 44206 77862
rect 44064 77752 44154 77808
rect 44270 77798 44276 77862
rect 44210 77752 44276 77798
rect 44064 77656 44276 77752
rect 45696 77862 46044 77868
rect 45696 77808 45838 77862
rect 45696 77752 45834 77808
rect 45902 77798 46044 77862
rect 45890 77752 46044 77798
rect 45696 77656 46044 77752
rect 47464 77862 47676 77868
rect 47464 77798 47470 77862
rect 47534 77808 47676 77862
rect 47464 77752 47514 77798
rect 47570 77752 47676 77808
rect 47464 77656 47676 77752
rect 49096 77862 49308 77868
rect 49096 77808 49238 77862
rect 49096 77752 49194 77808
rect 49302 77798 49308 77862
rect 49250 77752 49308 77798
rect 49096 77656 49308 77752
rect 50728 77862 51076 77868
rect 50728 77798 50734 77862
rect 50798 77808 51076 77862
rect 50798 77798 50874 77808
rect 50728 77752 50874 77798
rect 50930 77752 51076 77808
rect 50728 77656 51076 77752
rect 52496 77862 52708 77868
rect 52496 77808 52638 77862
rect 52496 77752 52554 77808
rect 52610 77798 52638 77808
rect 52702 77798 52708 77862
rect 52610 77752 52708 77798
rect 52496 77656 52708 77752
rect 54128 77862 54340 77868
rect 54128 77798 54134 77862
rect 54198 77808 54340 77862
rect 54198 77798 54234 77808
rect 54128 77752 54234 77798
rect 54290 77752 54340 77808
rect 54128 77656 54340 77752
rect 55760 77862 56108 77868
rect 55760 77798 55902 77862
rect 55966 77808 56108 77862
rect 55760 77752 55914 77798
rect 55970 77752 56108 77808
rect 55760 77656 56108 77752
rect 57528 77862 57740 77868
rect 57528 77808 57670 77862
rect 57528 77752 57594 77808
rect 57650 77798 57670 77808
rect 57734 77798 57740 77862
rect 57650 77752 57740 77798
rect 57528 77656 57740 77752
rect 59160 77862 59372 77868
rect 59160 77798 59166 77862
rect 59230 77808 59372 77862
rect 59230 77798 59274 77808
rect 59160 77752 59274 77798
rect 59330 77752 59372 77808
rect 59160 77656 59372 77752
rect 60928 77862 61140 77868
rect 60928 77798 60934 77862
rect 60998 77808 61140 77862
rect 60928 77752 60954 77798
rect 61010 77752 61140 77808
rect 60928 77656 61140 77752
rect 62560 77862 62772 77868
rect 62560 77808 62702 77862
rect 62560 77752 62634 77808
rect 62690 77798 62702 77808
rect 62766 77798 62772 77862
rect 62690 77752 62772 77798
rect 64056 77862 64404 77868
rect 64056 77798 64062 77862
rect 64126 77808 64404 77862
rect 64126 77798 64314 77808
rect 64056 77792 64314 77798
rect 62560 77656 62772 77752
rect 64192 77752 64314 77792
rect 64370 77752 64404 77808
rect 64192 77656 64404 77752
rect 65960 77862 66172 77868
rect 65960 77798 65966 77862
rect 66030 77808 66172 77862
rect 65960 77752 65994 77798
rect 66050 77752 66172 77808
rect 65960 77656 66172 77752
rect 67592 77862 67804 77868
rect 67592 77808 67734 77862
rect 67592 77752 67674 77808
rect 67730 77798 67734 77808
rect 67798 77798 67804 77862
rect 67730 77752 67804 77798
rect 67592 77656 67804 77752
rect 69224 77862 69436 77868
rect 69224 77798 69230 77862
rect 69294 77808 69436 77862
rect 69294 77798 69354 77808
rect 69224 77752 69354 77798
rect 69410 77752 69436 77808
rect 69224 77656 69436 77752
rect 70992 77862 71204 77868
rect 70992 77808 71134 77862
rect 70992 77752 71034 77808
rect 71090 77798 71134 77808
rect 71198 77798 71204 77862
rect 71090 77752 71204 77798
rect 70992 77656 71204 77752
rect 72624 77862 72836 77868
rect 72624 77808 72766 77862
rect 72624 77752 72714 77808
rect 72830 77798 72836 77862
rect 72770 77752 72836 77798
rect 72624 77656 72836 77752
rect 74256 77862 74604 77868
rect 74256 77808 74398 77862
rect 74256 77752 74394 77808
rect 74462 77798 74604 77862
rect 74450 77752 74604 77798
rect 74256 77656 74604 77752
rect 76024 77862 76236 77868
rect 76024 77808 76166 77862
rect 76024 77752 76074 77808
rect 76130 77798 76166 77808
rect 76230 77798 76236 77862
rect 76130 77752 76236 77798
rect 76024 77656 76236 77752
rect 77656 77862 77868 77868
rect 77656 77798 77662 77862
rect 77726 77808 77868 77862
rect 77726 77798 77754 77808
rect 77656 77752 77754 77798
rect 77810 77752 77868 77808
rect 77656 77656 77868 77752
rect 79288 77862 79636 77868
rect 79288 77798 79294 77862
rect 79358 77808 79636 77862
rect 79358 77798 79434 77808
rect 79288 77752 79434 77798
rect 79490 77752 79636 77808
rect 79288 77726 79636 77752
rect 79288 77662 79294 77726
rect 79358 77662 79636 77726
rect 79288 77656 79636 77662
rect 81056 77862 81268 77868
rect 81056 77808 81198 77862
rect 81056 77752 81114 77808
rect 81170 77798 81198 77808
rect 81262 77798 81268 77862
rect 81170 77752 81268 77798
rect 81056 77732 81268 77752
rect 82688 77862 82900 77868
rect 82688 77798 82694 77862
rect 82758 77808 82900 77862
rect 82758 77798 82794 77808
rect 82688 77752 82794 77798
rect 82850 77752 82900 77808
rect 81056 77726 81948 77732
rect 81056 77662 81878 77726
rect 81942 77662 81948 77726
rect 81056 77656 81948 77662
rect 82688 77656 82900 77752
rect 84320 77862 84668 77868
rect 84320 77798 84462 77862
rect 84526 77808 84668 77862
rect 84320 77752 84474 77798
rect 84530 77752 84668 77808
rect 84320 77656 84668 77752
rect 86088 77862 86300 77868
rect 86088 77808 86230 77862
rect 86088 77752 86154 77808
rect 86210 77798 86230 77808
rect 86294 77798 86300 77862
rect 86210 77752 86300 77798
rect 86088 77656 86300 77752
rect 87720 77862 87932 77868
rect 87720 77798 87726 77862
rect 87790 77808 87932 77862
rect 87790 77798 87834 77808
rect 87720 77752 87834 77798
rect 87890 77752 87932 77808
rect 87720 77656 87932 77752
rect 89488 77862 89700 77868
rect 89488 77808 89630 77862
rect 89488 77752 89514 77808
rect 89570 77798 89630 77808
rect 89694 77798 89700 77862
rect 89570 77752 89700 77798
rect 89488 77656 89700 77752
rect 91120 77862 91332 77868
rect 91120 77808 91262 77862
rect 91120 77752 91194 77808
rect 91250 77798 91262 77808
rect 91326 77798 91332 77862
rect 91250 77752 91332 77798
rect 91120 77656 91332 77752
rect 92752 77862 92964 77868
rect 92752 77808 92894 77862
rect 92752 77752 92874 77808
rect 92958 77798 92964 77862
rect 92930 77752 92964 77798
rect 92752 77656 92964 77752
rect 81872 77182 82220 77188
rect 81872 77118 82150 77182
rect 82214 77118 82220 77182
rect 81872 77046 82220 77118
rect 81872 76982 82014 77046
rect 82078 76982 82220 77046
rect 81872 76976 82220 76982
rect 93296 77182 95412 77188
rect 93296 77118 95342 77182
rect 95406 77118 95412 77182
rect 93296 77112 95412 77118
rect 93296 76976 93508 77112
rect 93160 76572 93372 76644
rect 93160 76516 93216 76572
rect 93272 76516 93372 76572
rect 93160 76508 93372 76516
rect 78880 76502 79092 76508
rect 78880 76438 78886 76502
rect 78950 76438 79092 76502
rect 78880 76296 79092 76438
rect 90032 76502 90244 76508
rect 90032 76438 90038 76502
rect 90102 76467 90244 76502
rect 90032 76411 90079 76438
rect 90135 76411 90244 76467
rect 93160 76432 95956 76508
rect 90032 76296 90244 76411
rect 81839 76105 81905 76108
rect 79036 76103 81905 76105
rect 1768 76000 1980 76100
rect 79036 76047 81844 76103
rect 81900 76047 81905 76103
rect 79036 76045 81905 76047
rect 81839 76042 81905 76045
rect 1768 75964 1818 76000
rect 1224 75958 1818 75964
rect 1224 75894 1230 75958
rect 1294 75944 1818 75958
rect 1874 75944 1980 76000
rect 94112 76000 94324 76100
rect 1294 75894 1980 75944
rect 1224 75888 1980 75894
rect 79288 75958 79500 75964
rect 79288 75894 79430 75958
rect 79494 75894 79500 75958
rect 79288 75847 79500 75894
rect 79288 75791 79422 75847
rect 79478 75791 79500 75847
rect 94112 75944 94176 76000
rect 94232 75964 94324 76000
rect 94232 75958 94732 75964
rect 94232 75944 94662 75958
rect 94112 75894 94662 75944
rect 94726 75894 94732 75958
rect 94112 75888 94732 75894
rect 94112 75828 94188 75888
rect 79288 75752 79500 75791
rect 81872 75822 82220 75828
rect 81872 75758 81878 75822
rect 81942 75758 82220 75822
rect 81872 75686 82220 75758
rect 81872 75622 81878 75686
rect 81942 75622 82220 75686
rect 81872 75616 82220 75622
rect 93296 75752 94188 75828
rect 93296 75616 93508 75752
rect 78880 75142 79364 75148
rect 78880 75078 79294 75142
rect 79358 75078 79364 75142
rect 78880 75072 79364 75078
rect 78880 74800 79092 75072
rect 1224 74462 1980 74468
rect 1224 74398 1230 74462
rect 1294 74398 1980 74462
rect 1224 74392 1980 74398
rect 1768 74320 1980 74392
rect 94112 74332 94324 74468
rect 1768 74264 1818 74320
rect 1874 74264 1980 74320
rect 1768 74120 1980 74264
rect 29240 74256 29860 74332
rect 29240 74196 29316 74256
rect 29784 74196 29860 74256
rect 30328 74256 30948 74332
rect 30328 74196 30404 74256
rect 30872 74196 30948 74256
rect 31688 74256 32308 74332
rect 31688 74196 31764 74256
rect 32232 74196 32308 74256
rect 32912 74256 33532 74332
rect 32912 74196 32988 74256
rect 33456 74196 33532 74256
rect 34272 74256 34892 74332
rect 34272 74196 34348 74256
rect 34816 74196 34892 74256
rect 35496 74256 36116 74332
rect 35496 74196 35572 74256
rect 36040 74196 36116 74256
rect 36584 74256 37204 74332
rect 36584 74196 36660 74256
rect 37128 74196 37204 74256
rect 37944 74256 38564 74332
rect 37944 74196 38020 74256
rect 38488 74196 38564 74256
rect 39168 74256 39788 74332
rect 39168 74196 39244 74256
rect 39712 74196 39788 74256
rect 40528 74256 41012 74332
rect 40528 74196 40604 74256
rect 40936 74196 41012 74256
rect 41752 74256 42372 74332
rect 41752 74196 41828 74256
rect 42296 74196 42372 74256
rect 42976 74256 43596 74332
rect 42976 74196 43052 74256
rect 43520 74196 43596 74256
rect 44200 74256 44820 74332
rect 44200 74196 44276 74256
rect 44744 74196 44820 74256
rect 45288 74256 46044 74332
rect 45288 74196 45364 74256
rect 45968 74196 46044 74256
rect 46648 74256 47268 74332
rect 46648 74196 46724 74256
rect 47192 74196 47268 74256
rect 48008 74256 48492 74332
rect 48008 74196 48084 74256
rect 48416 74196 48492 74256
rect 49232 74256 49716 74332
rect 49232 74196 49308 74256
rect 49640 74196 49716 74256
rect 50456 74256 51076 74332
rect 50456 74196 50532 74256
rect 51000 74196 51076 74256
rect 51544 74256 52300 74332
rect 51544 74196 51620 74256
rect 52224 74196 52300 74256
rect 52904 74256 53524 74332
rect 52904 74196 52980 74256
rect 53448 74196 53524 74256
rect 54128 74256 54748 74332
rect 54128 74196 54204 74256
rect 54672 74196 54748 74256
rect 55488 74256 55972 74332
rect 55488 74196 55564 74256
rect 55896 74196 55972 74256
rect 56712 74256 57332 74332
rect 56712 74196 56788 74256
rect 57256 74196 57332 74256
rect 57800 74256 58556 74332
rect 57800 74196 57876 74256
rect 58480 74196 58556 74256
rect 59160 74256 59780 74332
rect 59160 74196 59236 74256
rect 59704 74196 59780 74256
rect 60384 74256 61004 74332
rect 60384 74196 60460 74256
rect 60928 74196 61004 74256
rect 61744 74256 62228 74332
rect 61744 74196 61820 74256
rect 62152 74196 62228 74256
rect 62968 74256 63588 74332
rect 62968 74196 63044 74256
rect 63512 74196 63588 74256
rect 64056 74256 64812 74332
rect 64056 74196 64132 74256
rect 64736 74196 64812 74256
rect 65416 74256 66036 74332
rect 65416 74196 65492 74256
rect 65960 74196 66036 74256
rect 66504 74256 67124 74332
rect 66504 74196 66580 74256
rect 67048 74196 67124 74256
rect 81872 74326 82220 74332
rect 81872 74262 82014 74326
rect 82078 74262 82220 74326
rect 28152 74190 28364 74196
rect 28152 74126 28158 74190
rect 28222 74126 28364 74190
rect 28560 74143 29316 74196
rect 28152 74103 28364 74126
rect 28152 74047 28210 74103
rect 28266 74047 28364 74103
rect 28152 73984 28364 74047
rect 28443 74120 29316 74143
rect 29376 74190 29588 74196
rect 29376 74126 29518 74190
rect 29582 74126 29588 74190
rect 29784 74143 30404 74196
rect 28443 74045 28636 74120
rect 28560 73984 28636 74045
rect 29376 74103 29588 74126
rect 29376 74047 29458 74103
rect 29514 74047 29588 74103
rect 29376 73984 29588 74047
rect 29691 74120 30404 74143
rect 30600 74190 30812 74196
rect 30600 74126 30606 74190
rect 30670 74126 30812 74190
rect 29691 74045 29860 74120
rect 29784 73984 29860 74045
rect 30600 74103 30812 74126
rect 30600 74047 30706 74103
rect 30762 74047 30812 74103
rect 30600 73984 30812 74047
rect 30872 74120 31764 74196
rect 31824 74190 32036 74196
rect 31824 74126 31966 74190
rect 32030 74126 32036 74190
rect 32232 74143 32988 74196
rect 30872 74060 31084 74120
rect 31824 74103 32036 74126
rect 30872 74054 31220 74060
rect 30872 73990 31150 74054
rect 31214 73990 31220 74054
rect 30872 73984 31220 73990
rect 31824 74047 31954 74103
rect 32010 74047 32036 74103
rect 31824 73984 32036 74047
rect 32187 74120 32988 74143
rect 33048 74190 33260 74196
rect 33048 74126 33190 74190
rect 33254 74126 33260 74190
rect 33456 74143 34348 74196
rect 33048 74124 33260 74126
rect 32187 74045 32308 74120
rect 32232 73984 32308 74045
rect 33048 74103 33279 74124
rect 33048 74047 33202 74103
rect 33258 74047 33279 74103
rect 33048 74026 33279 74047
rect 33435 74120 34348 74143
rect 34408 74190 34620 74196
rect 34408 74126 34550 74190
rect 34614 74126 34620 74190
rect 34816 74143 35572 74196
rect 33435 74045 33668 74120
rect 33048 73984 33260 74026
rect 33456 73984 33668 74045
rect 34408 74103 34620 74126
rect 34408 74047 34450 74103
rect 34506 74047 34620 74103
rect 34408 73984 34620 74047
rect 34683 74120 35572 74143
rect 35632 74190 35844 74196
rect 35632 74126 35774 74190
rect 35838 74126 35844 74190
rect 36040 74143 36660 74196
rect 34683 74045 34892 74120
rect 34816 73984 34892 74045
rect 35632 74103 35844 74126
rect 35632 74047 35698 74103
rect 35754 74047 35844 74103
rect 35632 73984 35844 74047
rect 35931 74120 36660 74143
rect 36856 74190 37068 74196
rect 36856 74126 36862 74190
rect 36926 74126 37068 74190
rect 35931 74045 36116 74120
rect 36040 73984 36116 74045
rect 36856 74103 37068 74126
rect 36856 74047 36946 74103
rect 37002 74047 37068 74103
rect 36856 73984 37068 74047
rect 37128 74120 38020 74196
rect 38080 74190 38292 74196
rect 38080 74126 38222 74190
rect 38286 74126 38292 74190
rect 38488 74143 39244 74196
rect 37128 73984 37340 74120
rect 38080 74103 38292 74126
rect 38080 74047 38194 74103
rect 38250 74047 38292 74103
rect 38080 73984 38292 74047
rect 38427 74120 39244 74143
rect 39304 74190 39516 74196
rect 39304 74126 39310 74190
rect 39374 74126 39516 74190
rect 39712 74143 40604 74196
rect 39304 74124 39516 74126
rect 38427 74045 38564 74120
rect 38488 73984 38564 74045
rect 39304 74103 39519 74124
rect 39304 74047 39442 74103
rect 39498 74047 39519 74103
rect 39304 74026 39519 74047
rect 39675 74120 40604 74143
rect 40664 74190 40740 74196
rect 40664 74126 40670 74190
rect 40734 74126 40740 74190
rect 40936 74143 41828 74196
rect 40664 74124 40740 74126
rect 39675 74045 39788 74120
rect 39304 73984 39516 74026
rect 39712 73984 39788 74045
rect 40664 74103 40767 74124
rect 40664 74047 40690 74103
rect 40746 74047 40767 74103
rect 40664 74026 40767 74047
rect 40923 74120 41828 74143
rect 41888 74190 42100 74196
rect 41888 74126 41894 74190
rect 41958 74126 42100 74190
rect 42296 74143 43052 74196
rect 40923 74045 41148 74120
rect 40664 73984 40740 74026
rect 40936 73984 41148 74045
rect 41888 74103 42100 74126
rect 41888 74047 41938 74103
rect 41994 74047 42100 74103
rect 41888 73984 42100 74047
rect 42171 74120 43052 74143
rect 43112 74190 43324 74196
rect 43112 74126 43254 74190
rect 43318 74126 43324 74190
rect 43520 74143 44276 74196
rect 42171 74045 42372 74120
rect 42296 73984 42372 74045
rect 43112 74103 43324 74126
rect 43112 74047 43186 74103
rect 43242 74047 43324 74103
rect 43112 73984 43324 74047
rect 43419 74120 44276 74143
rect 44336 74190 44548 74196
rect 44336 74126 44342 74190
rect 44406 74126 44548 74190
rect 44744 74143 45364 74196
rect 43419 74045 43596 74120
rect 43520 73984 43596 74045
rect 44336 74103 44548 74126
rect 44336 74047 44434 74103
rect 44490 74047 44548 74103
rect 44336 73984 44548 74047
rect 44667 74120 45364 74143
rect 45560 74190 45772 74196
rect 45560 74126 45566 74190
rect 45630 74126 45772 74190
rect 45968 74143 46724 74196
rect 44667 74045 44820 74120
rect 44744 73984 44820 74045
rect 45560 74103 45772 74126
rect 45560 74047 45682 74103
rect 45738 74047 45772 74103
rect 45560 73984 45772 74047
rect 45915 74120 46724 74143
rect 46784 74190 46996 74196
rect 46784 74126 46926 74190
rect 46990 74126 46996 74190
rect 47192 74143 48084 74196
rect 46784 74124 46996 74126
rect 45915 74045 46044 74120
rect 45968 73984 46044 74045
rect 46784 74103 47007 74124
rect 46784 74047 46930 74103
rect 46986 74047 47007 74103
rect 46784 74026 47007 74047
rect 47163 74120 48084 74143
rect 48144 74190 48220 74196
rect 48144 74126 48150 74190
rect 48214 74126 48220 74190
rect 48416 74143 49308 74196
rect 48144 74124 48220 74126
rect 47163 74045 47268 74120
rect 46784 73984 46996 74026
rect 47192 73984 47268 74045
rect 48144 74103 48255 74124
rect 48144 74047 48178 74103
rect 48234 74047 48255 74103
rect 48144 74026 48255 74047
rect 48411 74120 49308 74143
rect 49368 74190 49580 74196
rect 49368 74126 49510 74190
rect 49574 74126 49580 74190
rect 48411 74045 48628 74120
rect 48144 73984 48220 74026
rect 48416 73984 48628 74045
rect 49368 74103 49580 74126
rect 49368 74047 49426 74103
rect 49482 74047 49580 74103
rect 49368 73984 49580 74047
rect 49640 74120 50532 74196
rect 50592 74190 50804 74196
rect 50592 74126 50598 74190
rect 50662 74126 50804 74190
rect 51000 74143 51620 74196
rect 49640 73984 49852 74120
rect 50592 74103 50804 74126
rect 50592 74047 50674 74103
rect 50730 74047 50804 74103
rect 50592 73984 50804 74047
rect 50907 74120 51620 74143
rect 51816 74190 52028 74196
rect 51816 74126 51958 74190
rect 52022 74126 52028 74190
rect 52224 74143 52980 74196
rect 50907 74045 51076 74120
rect 51000 73984 51076 74045
rect 51816 74103 52028 74126
rect 51816 74047 51922 74103
rect 51978 74047 52028 74103
rect 51816 73984 52028 74047
rect 52155 74120 52980 74143
rect 53040 74190 53252 74196
rect 53040 74126 53046 74190
rect 53110 74126 53252 74190
rect 53448 74143 54204 74196
rect 52155 74045 52300 74120
rect 52224 73984 52300 74045
rect 53040 74103 53252 74126
rect 53040 74047 53170 74103
rect 53226 74047 53252 74103
rect 53040 73984 53252 74047
rect 53403 74120 54204 74143
rect 54264 74190 54476 74196
rect 54264 74126 54270 74190
rect 54334 74126 54476 74190
rect 54672 74143 55564 74196
rect 54264 74124 54476 74126
rect 53403 74045 53524 74120
rect 53448 73984 53524 74045
rect 54264 74103 54495 74124
rect 54264 74047 54418 74103
rect 54474 74047 54495 74103
rect 54264 74026 54495 74047
rect 54651 74120 55564 74143
rect 55624 74190 55836 74196
rect 55624 74126 55630 74190
rect 55694 74126 55836 74190
rect 54651 74045 54884 74120
rect 54264 73984 54476 74026
rect 54672 73984 54884 74045
rect 55624 74103 55836 74126
rect 55624 74047 55666 74103
rect 55722 74047 55836 74103
rect 55624 73984 55836 74047
rect 55896 74120 56788 74196
rect 56848 74190 57060 74196
rect 56848 74126 56854 74190
rect 56918 74126 57060 74190
rect 57256 74143 57876 74196
rect 55896 73984 56108 74120
rect 56848 74103 57060 74126
rect 56848 74047 56914 74103
rect 56970 74047 57060 74103
rect 56848 73984 57060 74047
rect 57147 74120 57876 74143
rect 58072 74190 58284 74196
rect 58072 74126 58214 74190
rect 58278 74126 58284 74190
rect 58480 74143 59236 74196
rect 57147 74045 57332 74120
rect 57256 73984 57332 74045
rect 58072 74103 58284 74126
rect 58072 74047 58162 74103
rect 58218 74047 58284 74103
rect 58072 73984 58284 74047
rect 58395 74120 59236 74143
rect 59296 74190 59508 74196
rect 59296 74126 59302 74190
rect 59366 74126 59508 74190
rect 59704 74143 60460 74196
rect 58395 74045 58556 74120
rect 58480 73984 58556 74045
rect 59296 74103 59508 74126
rect 59296 74047 59410 74103
rect 59466 74047 59508 74103
rect 59296 73984 59508 74047
rect 59643 74120 60460 74143
rect 60520 74190 60732 74196
rect 60520 74126 60662 74190
rect 60726 74126 60732 74190
rect 60928 74143 61820 74196
rect 60520 74124 60732 74126
rect 59643 74045 59780 74120
rect 59704 73984 59780 74045
rect 60520 74103 60735 74124
rect 60520 74047 60658 74103
rect 60714 74047 60735 74103
rect 60520 74026 60735 74047
rect 60891 74120 61820 74143
rect 61880 74190 61956 74196
rect 61880 74126 61886 74190
rect 61950 74126 61956 74190
rect 62152 74143 63044 74196
rect 61880 74124 61956 74126
rect 60891 74045 61004 74120
rect 60520 73984 60732 74026
rect 60928 73984 61004 74045
rect 61880 74103 61983 74124
rect 61880 74047 61906 74103
rect 61962 74047 61983 74103
rect 61880 74026 61983 74047
rect 62139 74120 63044 74143
rect 63104 74190 63316 74196
rect 63104 74126 63246 74190
rect 63310 74126 63316 74190
rect 63512 74143 64132 74196
rect 62139 74045 62364 74120
rect 61880 73984 61956 74026
rect 62152 73984 62364 74045
rect 63104 74103 63316 74126
rect 63104 74047 63154 74103
rect 63210 74047 63316 74103
rect 63104 73984 63316 74047
rect 63387 74120 64132 74143
rect 64328 74190 64540 74196
rect 64328 74126 64334 74190
rect 64398 74126 64540 74190
rect 64736 74143 65492 74196
rect 63387 74045 63588 74120
rect 63512 73984 63588 74045
rect 64328 74103 64540 74126
rect 64328 74047 64402 74103
rect 64458 74047 64540 74103
rect 64328 73984 64540 74047
rect 64635 74120 65492 74143
rect 65552 74190 65764 74196
rect 65552 74126 65558 74190
rect 65622 74126 65764 74190
rect 65960 74143 66580 74196
rect 64635 74045 64812 74120
rect 64736 73984 64812 74045
rect 65552 74103 65764 74126
rect 65552 74047 65650 74103
rect 65706 74047 65764 74103
rect 65552 73984 65764 74047
rect 65883 74120 66580 74143
rect 66776 74190 66988 74196
rect 66776 74126 66918 74190
rect 66982 74126 66988 74190
rect 65883 74045 66036 74120
rect 65960 73984 66036 74045
rect 66776 74103 66988 74126
rect 66776 74047 66898 74103
rect 66954 74047 66988 74103
rect 66776 73984 66988 74047
rect 67048 73984 67260 74196
rect 81872 74190 82220 74262
rect 81872 74126 82014 74190
rect 82078 74126 82220 74190
rect 81872 74120 82220 74126
rect 94112 74326 94732 74332
rect 94112 74320 94662 74326
rect 94112 74264 94176 74320
rect 94232 74264 94662 74320
rect 94112 74262 94662 74264
rect 94726 74262 94732 74326
rect 94112 74256 94732 74262
rect 94112 74120 94324 74256
rect 28424 73788 28636 73924
rect 29648 73918 29860 73924
rect 29648 73854 29790 73918
rect 29854 73854 29860 73918
rect 29648 73788 29860 73854
rect 28424 73782 29860 73788
rect 28424 73718 28566 73782
rect 28630 73718 29790 73782
rect 29854 73718 29860 73782
rect 28424 73712 29860 73718
rect 30872 73848 32308 73924
rect 30872 73782 31084 73848
rect 30872 73718 31014 73782
rect 31078 73718 31084 73782
rect 30872 73712 31084 73718
rect 32096 73788 32308 73848
rect 33320 73848 34892 73924
rect 33320 73788 33668 73848
rect 32096 73782 33668 73788
rect 32096 73718 32102 73782
rect 32166 73718 33462 73782
rect 33526 73718 33668 73782
rect 32096 73712 33668 73718
rect 34680 73788 34892 73848
rect 35904 73848 37340 73924
rect 35904 73788 36116 73848
rect 34680 73782 36116 73788
rect 34680 73718 34686 73782
rect 34750 73718 36046 73782
rect 36110 73718 36116 73782
rect 34680 73712 36116 73718
rect 37128 73788 37340 73848
rect 38352 73788 38564 73924
rect 37128 73782 38564 73788
rect 37128 73718 37270 73782
rect 37334 73718 38494 73782
rect 38558 73718 38564 73782
rect 37128 73712 38564 73718
rect 39576 73848 41148 73924
rect 39576 73782 39788 73848
rect 39576 73718 39718 73782
rect 39782 73718 39788 73782
rect 39576 73712 39788 73718
rect 40800 73788 41148 73848
rect 42160 73848 43596 73924
rect 40800 73782 42100 73788
rect 40800 73718 40806 73782
rect 40870 73718 42030 73782
rect 42094 73718 42100 73782
rect 40800 73712 42100 73718
rect 42160 73782 42372 73848
rect 42160 73718 42302 73782
rect 42366 73718 42372 73782
rect 42160 73712 42372 73718
rect 43384 73788 43596 73848
rect 44608 73788 44820 73924
rect 43384 73782 44820 73788
rect 43384 73718 43390 73782
rect 43454 73718 44750 73782
rect 44814 73718 44820 73782
rect 43384 73712 44820 73718
rect 45832 73788 46044 73924
rect 47056 73788 47268 73924
rect 45832 73782 47268 73788
rect 45832 73718 45974 73782
rect 46038 73718 47198 73782
rect 47262 73718 47268 73782
rect 45832 73712 47268 73718
rect 48280 73782 48628 73924
rect 48280 73718 48558 73782
rect 48622 73718 48628 73782
rect 48280 73712 48628 73718
rect 49640 73782 49852 73924
rect 49640 73718 49782 73782
rect 49846 73718 49852 73782
rect 49640 73712 49852 73718
rect 50864 73782 51076 73924
rect 50864 73718 51006 73782
rect 51070 73718 51076 73782
rect 50864 73712 51076 73718
rect 52088 73782 52300 73924
rect 52088 73718 52094 73782
rect 52158 73718 52300 73782
rect 52088 73712 52300 73718
rect 53312 73848 54884 73924
rect 53312 73782 53524 73848
rect 53312 73718 53454 73782
rect 53518 73718 53524 73782
rect 53312 73712 53524 73718
rect 54536 73782 54884 73848
rect 54536 73718 54678 73782
rect 54742 73718 54884 73782
rect 54536 73712 54884 73718
rect 55896 73848 57332 73924
rect 55896 73782 56108 73848
rect 55896 73718 56038 73782
rect 56102 73718 56108 73782
rect 55896 73712 56108 73718
rect 57120 73788 57332 73848
rect 58344 73788 58556 73924
rect 57120 73782 58556 73788
rect 57120 73718 57262 73782
rect 57326 73718 58486 73782
rect 58550 73718 58556 73782
rect 57120 73712 58556 73718
rect 59568 73782 59780 73924
rect 59568 73718 59710 73782
rect 59774 73718 59780 73782
rect 59568 73712 59780 73718
rect 60792 73782 61004 73924
rect 60792 73718 60798 73782
rect 60862 73718 61004 73782
rect 60792 73712 61004 73718
rect 62016 73782 62364 73924
rect 62016 73718 62158 73782
rect 62222 73718 62364 73782
rect 62016 73712 62364 73718
rect 63376 73788 63588 73924
rect 64600 73788 64812 73924
rect 63376 73782 64812 73788
rect 63376 73718 63518 73782
rect 63582 73718 64742 73782
rect 64806 73718 64812 73782
rect 63376 73712 64812 73718
rect 65824 73788 66036 73924
rect 67048 73788 67260 73924
rect 65824 73782 67260 73788
rect 65824 73718 65966 73782
rect 66030 73718 67190 73782
rect 67254 73718 67260 73782
rect 65824 73712 67260 73718
rect 28424 73102 28636 73108
rect 28424 73038 28566 73102
rect 28630 73038 28636 73102
rect 28424 72760 28636 73038
rect 29648 73102 31084 73108
rect 29648 73038 29790 73102
rect 29854 73038 31014 73102
rect 31078 73038 31084 73102
rect 29648 73032 31084 73038
rect 29648 72760 29860 73032
rect 30872 72830 31084 73032
rect 30872 72766 30878 72830
rect 30942 72766 31084 72830
rect 30872 72760 31084 72766
rect 32096 73102 32308 73108
rect 32096 73038 32102 73102
rect 32166 73038 32308 73102
rect 32096 72760 32308 73038
rect 33320 73102 33532 73108
rect 33320 73038 33462 73102
rect 33526 73038 33532 73102
rect 33320 72760 33532 73038
rect 34544 73102 34892 73108
rect 34544 73038 34686 73102
rect 34750 73038 34892 73102
rect 34544 72760 34892 73038
rect 35904 73102 36116 73108
rect 35904 73038 36046 73102
rect 36110 73038 36116 73102
rect 35904 72760 36116 73038
rect 37128 73102 37340 73108
rect 37128 73038 37270 73102
rect 37334 73038 37340 73102
rect 37128 72760 37340 73038
rect 38352 73102 39788 73108
rect 38352 73038 38494 73102
rect 38558 73038 39718 73102
rect 39782 73038 39788 73102
rect 38352 73032 39788 73038
rect 38352 72760 38564 73032
rect 39576 72760 39788 73032
rect 40800 73102 41012 73108
rect 40800 73038 40806 73102
rect 40870 73038 41012 73102
rect 40800 72760 41012 73038
rect 42024 73102 42372 73108
rect 42024 73038 42030 73102
rect 42094 73038 42302 73102
rect 42366 73038 42372 73102
rect 42024 72760 42372 73038
rect 43384 73102 43596 73108
rect 43384 73038 43390 73102
rect 43454 73038 43596 73102
rect 43384 72760 43596 73038
rect 44608 73102 46044 73108
rect 44608 73038 44750 73102
rect 44814 73038 45974 73102
rect 46038 73038 46044 73102
rect 44608 73032 46044 73038
rect 44608 72760 44820 73032
rect 45832 72760 46044 73032
rect 47056 73102 49852 73108
rect 47056 73038 47198 73102
rect 47262 73038 48558 73102
rect 48622 73038 49782 73102
rect 49846 73038 49852 73102
rect 47056 73032 49852 73038
rect 47056 72760 47268 73032
rect 48280 72760 48628 73032
rect 49640 72836 49852 73032
rect 50864 73102 52300 73108
rect 50864 73038 51006 73102
rect 51070 73038 52094 73102
rect 52158 73038 52300 73102
rect 50864 73032 52300 73038
rect 50864 72836 51076 73032
rect 49640 72760 51076 72836
rect 52088 72972 52300 73032
rect 53312 73102 53524 73108
rect 53312 73038 53454 73102
rect 53518 73038 53524 73102
rect 53312 72972 53524 73038
rect 52088 72896 53524 72972
rect 52088 72760 52300 72896
rect 53312 72760 53524 72896
rect 54536 73102 54748 73108
rect 54536 73038 54678 73102
rect 54742 73038 54748 73102
rect 54536 72836 54748 73038
rect 55760 73102 56108 73108
rect 55760 73038 56038 73102
rect 56102 73038 56108 73102
rect 55760 72836 56108 73038
rect 54536 72760 56108 72836
rect 57120 73102 57332 73108
rect 57120 73038 57262 73102
rect 57326 73038 57332 73102
rect 57120 72760 57332 73038
rect 58344 73102 58556 73108
rect 58344 73038 58486 73102
rect 58550 73038 58556 73102
rect 58344 72836 58556 73038
rect 59568 73102 61004 73108
rect 59568 73038 59710 73102
rect 59774 73038 60798 73102
rect 60862 73038 61004 73102
rect 59568 73032 61004 73038
rect 59568 72836 59780 73032
rect 58344 72760 59780 72836
rect 60792 72972 61004 73032
rect 62016 73102 63588 73108
rect 62016 73038 62158 73102
rect 62222 73038 63518 73102
rect 63582 73038 63588 73102
rect 62016 73032 63588 73038
rect 62016 72972 62228 73032
rect 60792 72896 62228 72972
rect 60792 72760 61004 72896
rect 62016 72760 62228 72896
rect 63240 72760 63588 73032
rect 64600 73102 66036 73108
rect 64600 73038 64742 73102
rect 64806 73038 65966 73102
rect 66030 73038 66036 73102
rect 64600 73032 66036 73038
rect 64600 72760 64812 73032
rect 65824 72760 66036 73032
rect 67048 73102 67260 73108
rect 67048 73038 67190 73102
rect 67254 73038 67260 73102
rect 67048 72760 67260 73038
rect 74664 72966 74876 73244
rect 74664 72902 74806 72966
rect 74870 72902 74876 72966
rect 74664 72896 74876 72902
rect 81872 72966 82220 72972
rect 81872 72902 81878 72966
rect 81942 72902 82220 72966
rect 81872 72830 82220 72902
rect 81872 72766 82150 72830
rect 82214 72766 82220 72830
rect 81872 72760 82220 72766
rect 1768 72640 1980 72700
rect 1768 72584 1818 72640
rect 1874 72584 1980 72640
rect 1768 72564 1980 72584
rect 1224 72558 1980 72564
rect 1224 72494 1230 72558
rect 1294 72494 1980 72558
rect 1224 72488 1980 72494
rect 94112 72640 94324 72700
rect 94112 72584 94176 72640
rect 94232 72584 94324 72640
rect 94112 72564 94324 72584
rect 94112 72558 94732 72564
rect 94112 72494 94662 72558
rect 94726 72494 94732 72558
rect 94112 72488 94732 72494
rect 28424 72286 67396 72292
rect 28424 72222 28566 72286
rect 28630 72222 31150 72286
rect 31214 72222 67396 72286
rect 28424 72216 67396 72222
rect 28513 72111 28611 72216
rect 29761 72111 29859 72216
rect 31009 72111 31107 72216
rect 32257 72111 32355 72216
rect 33505 72111 33603 72216
rect 34753 72111 34851 72216
rect 36001 72111 36099 72216
rect 37249 72111 37347 72216
rect 38497 72111 38595 72216
rect 39745 72111 39843 72216
rect 40993 72111 41091 72216
rect 42241 72111 42339 72216
rect 43489 72111 43587 72216
rect 44737 72111 44835 72216
rect 45985 72111 46083 72216
rect 47233 72111 47331 72216
rect 48481 72111 48579 72216
rect 49729 72111 49827 72216
rect 50977 72111 51075 72216
rect 52225 72111 52323 72216
rect 53473 72111 53571 72216
rect 54721 72111 54819 72216
rect 55969 72111 56067 72216
rect 57217 72111 57315 72216
rect 58465 72111 58563 72216
rect 59713 72111 59811 72216
rect 60961 72111 61059 72216
rect 62209 72111 62307 72216
rect 63457 72111 63555 72216
rect 64705 72111 64803 72216
rect 65953 72111 66051 72216
rect 67201 72111 67299 72216
rect 69712 72189 69778 72192
rect 81923 72189 81989 72192
rect 69712 72187 81989 72189
rect 69712 72131 69717 72187
rect 69773 72131 81928 72187
rect 81984 72131 81989 72187
rect 69712 72129 81989 72131
rect 69712 72126 69778 72129
rect 81923 72126 81989 72129
rect 74664 71606 74876 71748
rect 74664 71542 74670 71606
rect 74734 71542 74876 71606
rect 74664 71536 74876 71542
rect 81872 71606 82220 71612
rect 81872 71542 82014 71606
rect 82078 71542 82220 71606
rect 81872 71470 82220 71542
rect 81872 71406 82014 71470
rect 82078 71406 82220 71470
rect 81872 71400 82220 71406
rect 91936 71476 92148 71612
rect 92616 71476 92828 71612
rect 91936 71470 94188 71476
rect 91936 71406 94118 71470
rect 94182 71406 94188 71470
rect 91936 71400 94188 71406
rect 1768 70960 1980 71068
rect 1768 70932 1818 70960
rect 1224 70926 1818 70932
rect 1224 70862 1230 70926
rect 1294 70904 1818 70926
rect 1874 70904 1980 70960
rect 1294 70862 1980 70904
rect 1224 70856 1980 70862
rect 94112 71062 94324 71068
rect 94112 70998 94118 71062
rect 94182 70998 94324 71062
rect 94112 70960 94324 70998
rect 94112 70904 94176 70960
rect 94232 70932 94324 70960
rect 94232 70926 94732 70932
rect 94232 70904 94662 70926
rect 94112 70862 94662 70904
rect 94726 70862 94732 70926
rect 94112 70856 94732 70862
rect 69836 70775 69902 70778
rect 81923 70775 81989 70778
rect 69836 70773 81989 70775
rect 69836 70717 69841 70773
rect 69897 70717 81928 70773
rect 81984 70717 81989 70773
rect 69836 70715 81989 70717
rect 69836 70712 69902 70715
rect 81923 70712 81989 70715
rect 28560 70518 28908 70524
rect 28560 70454 28566 70518
rect 28630 70454 28908 70518
rect 28560 70388 28908 70454
rect 29920 70388 30132 70524
rect 31144 70448 32580 70524
rect 31144 70388 31356 70448
rect 27646 70382 31356 70388
rect 27608 70318 27614 70382
rect 27678 70318 31356 70382
rect 27646 70312 31356 70318
rect 32368 70388 32580 70448
rect 33592 70448 35028 70524
rect 33592 70388 33804 70448
rect 32368 70312 33804 70388
rect 34816 70388 35028 70448
rect 36040 70448 38836 70524
rect 36040 70388 36388 70448
rect 34816 70312 36388 70388
rect 37400 70312 37612 70448
rect 38624 70388 38836 70448
rect 39848 70448 41284 70524
rect 39848 70388 40060 70448
rect 38624 70312 40060 70388
rect 41072 70388 41284 70448
rect 42296 70448 45092 70524
rect 42296 70388 42644 70448
rect 41072 70312 42644 70388
rect 43656 70312 43868 70448
rect 44880 70388 45092 70448
rect 46104 70448 47540 70524
rect 46104 70388 46316 70448
rect 44880 70312 46316 70388
rect 47328 70388 47540 70448
rect 48552 70448 50124 70524
rect 48552 70388 48764 70448
rect 47328 70312 48764 70388
rect 49776 70388 50124 70448
rect 51136 70388 51348 70524
rect 52360 70448 53796 70524
rect 52360 70388 52572 70448
rect 49776 70312 52572 70388
rect 53584 70388 53796 70448
rect 54808 70448 56244 70524
rect 54808 70388 55020 70448
rect 53584 70312 55020 70388
rect 56032 70388 56244 70448
rect 57256 70388 57604 70524
rect 58616 70448 60052 70524
rect 58616 70388 58828 70448
rect 56032 70312 58828 70388
rect 59840 70388 60052 70448
rect 61064 70448 62500 70524
rect 61064 70388 61276 70448
rect 59840 70312 61276 70388
rect 62288 70388 62500 70448
rect 63512 70448 66308 70524
rect 63512 70388 63860 70448
rect 62288 70312 63860 70388
rect 64872 70312 65084 70448
rect 66096 70388 66308 70448
rect 67320 70388 67532 70524
rect 66096 70382 69028 70388
rect 66096 70318 68958 70382
rect 69022 70318 69028 70382
rect 66096 70312 69028 70318
rect 74664 70382 74876 70388
rect 74664 70318 74806 70382
rect 74870 70318 74876 70382
rect 74664 70252 74876 70318
rect 74566 70246 74876 70252
rect 74528 70182 74534 70246
rect 74598 70182 74876 70246
rect 74566 70176 74876 70182
rect 81872 70110 82220 70116
rect 81872 70046 82150 70110
rect 82214 70046 82220 70110
rect 81872 69904 82220 70046
rect 91936 70040 92828 70116
rect 91936 69980 92148 70040
rect 91936 69974 92556 69980
rect 91936 69910 92486 69974
rect 92550 69910 92556 69974
rect 91936 69904 92556 69910
rect 92616 69904 92828 70040
rect 93419 69660 93425 69662
rect 74928 69600 74988 69660
rect 81788 69600 93425 69660
rect 93419 69598 93425 69600
rect 93489 69598 93495 69662
rect 1768 69280 1980 69436
rect 73697 69361 73763 69364
rect 81923 69361 81989 69364
rect 73697 69359 81989 69361
rect 73697 69303 73702 69359
rect 73758 69303 81928 69359
rect 81984 69303 81989 69359
rect 73697 69301 81989 69303
rect 73697 69298 73763 69301
rect 81923 69298 81989 69301
rect 94112 69300 94324 69436
rect 1768 69224 1818 69280
rect 1874 69224 1980 69280
rect 1768 69164 1980 69224
rect 1224 69158 1980 69164
rect 1224 69094 1230 69158
rect 1294 69094 1980 69158
rect 1224 69088 1980 69094
rect 94112 69294 94732 69300
rect 94112 69280 94662 69294
rect 94112 69224 94176 69280
rect 94232 69230 94662 69280
rect 94726 69230 94732 69294
rect 94232 69224 94732 69230
rect 94112 69158 94324 69224
rect 94112 69094 94118 69158
rect 94182 69094 94324 69158
rect 94112 69088 94324 69094
rect 28152 68750 28364 69028
rect 28152 68686 28294 68750
rect 28358 68686 28364 68750
rect 28152 68680 28364 68686
rect 29104 68892 29316 69028
rect 29376 68892 29724 69028
rect 29104 68816 29724 68892
rect 29104 68750 29316 68816
rect 29104 68686 29246 68750
rect 29310 68686 29316 68750
rect 29104 68680 29316 68686
rect 29376 68680 29724 68816
rect 30328 69022 30948 69028
rect 30328 68958 30878 69022
rect 30942 68958 30948 69022
rect 30328 68952 30948 68958
rect 30328 68756 30540 68952
rect 30328 68750 30676 68756
rect 30328 68686 30334 68750
rect 30398 68686 30606 68750
rect 30670 68686 30676 68750
rect 30328 68680 30676 68686
rect 30736 68680 30948 68952
rect 31552 68756 31764 69028
rect 31960 68756 32172 69028
rect 31552 68750 32172 68756
rect 31552 68686 31558 68750
rect 31622 68686 31694 68750
rect 31758 68686 32172 68750
rect 31552 68680 32172 68686
rect 32776 68952 33396 69028
rect 32776 68750 32988 68952
rect 32776 68686 32782 68750
rect 32846 68686 32988 68750
rect 32776 68680 32988 68686
rect 33184 68750 33396 68952
rect 33184 68686 33326 68750
rect 33390 68686 33396 68750
rect 33184 68680 33396 68686
rect 34000 68952 34620 69028
rect 34000 68750 34212 68952
rect 34000 68686 34142 68750
rect 34206 68686 34212 68750
rect 34000 68680 34212 68686
rect 34408 68756 34620 68952
rect 35224 68952 35844 69028
rect 35224 68756 35572 68952
rect 34408 68750 35572 68756
rect 34408 68686 35230 68750
rect 35294 68686 35572 68750
rect 34408 68680 35572 68686
rect 35632 68750 35844 68952
rect 35632 68686 35774 68750
rect 35838 68686 35844 68750
rect 35632 68680 35844 68686
rect 36584 68892 36796 69028
rect 36856 68892 37204 69028
rect 36584 68816 37204 68892
rect 36584 68750 36796 68816
rect 36584 68686 36590 68750
rect 36654 68686 36796 68750
rect 36584 68680 36796 68686
rect 36856 68680 37204 68816
rect 37808 68892 38020 69028
rect 38216 68892 38428 69028
rect 37808 68816 38428 68892
rect 37808 68750 38020 68816
rect 37808 68686 37814 68750
rect 37878 68686 38020 68750
rect 37808 68680 38020 68686
rect 38216 68750 38428 68816
rect 38216 68686 38358 68750
rect 38422 68686 38428 68750
rect 38216 68680 38428 68686
rect 39032 68952 39652 69028
rect 39032 68756 39244 68952
rect 39032 68750 39380 68756
rect 39032 68686 39038 68750
rect 39102 68686 39310 68750
rect 39374 68686 39380 68750
rect 39032 68680 39380 68686
rect 39440 68680 39652 68952
rect 40256 68756 40468 69028
rect 40664 68756 40876 69028
rect 40256 68750 40876 68756
rect 40256 68686 40262 68750
rect 40326 68686 40876 68750
rect 40256 68680 40876 68686
rect 41480 68892 41828 69028
rect 41888 68892 42100 69028
rect 41480 68816 42100 68892
rect 41480 68680 41828 68816
rect 41888 68750 42100 68816
rect 41888 68686 41894 68750
rect 41958 68686 42100 68750
rect 41888 68680 42100 68686
rect 42840 68756 43052 69028
rect 43112 68756 43460 69028
rect 44064 68952 44684 69028
rect 44064 68756 44276 68952
rect 42840 68750 44276 68756
rect 42840 68686 42846 68750
rect 42910 68686 43390 68750
rect 43454 68686 44070 68750
rect 44134 68686 44276 68750
rect 42840 68680 44276 68686
rect 44472 68680 44684 68952
rect 45288 68892 45500 69028
rect 45696 68892 45908 69028
rect 45288 68816 45908 68892
rect 45288 68680 45500 68816
rect 45696 68750 45908 68816
rect 45696 68686 45838 68750
rect 45902 68686 45908 68750
rect 45696 68680 45908 68686
rect 46512 68892 46724 69028
rect 46920 68892 47132 69028
rect 46512 68816 47132 68892
rect 46512 68750 46724 68816
rect 46512 68686 46518 68750
rect 46582 68686 46724 68750
rect 46512 68680 46724 68686
rect 46920 68750 47132 68816
rect 46920 68686 47062 68750
rect 47126 68686 47132 68750
rect 46920 68680 47132 68686
rect 47736 68952 48356 69028
rect 47736 68750 47948 68952
rect 47736 68686 47742 68750
rect 47806 68686 47948 68750
rect 47736 68680 47948 68686
rect 48144 68680 48356 68952
rect 48960 68892 49308 69028
rect 49368 68892 49580 69028
rect 48960 68816 49580 68892
rect 48960 68750 49308 68816
rect 48960 68686 48966 68750
rect 49030 68686 49308 68750
rect 48960 68680 49308 68686
rect 49368 68680 49580 68816
rect 50320 68892 50532 69028
rect 50592 68892 50940 69028
rect 50320 68816 50940 68892
rect 50320 68680 50532 68816
rect 50592 68750 50940 68816
rect 50592 68686 50598 68750
rect 50662 68686 50940 68750
rect 50592 68680 50940 68686
rect 51544 68756 51756 69028
rect 51952 68756 52164 69028
rect 51544 68750 52164 68756
rect 51544 68686 51550 68750
rect 51614 68686 52094 68750
rect 52158 68686 52164 68750
rect 51544 68680 52164 68686
rect 52768 68952 53388 69028
rect 52768 68756 52980 68952
rect 52768 68750 53116 68756
rect 52768 68686 52774 68750
rect 52838 68686 53046 68750
rect 53110 68686 53116 68750
rect 52768 68680 53116 68686
rect 53176 68680 53388 68952
rect 53992 68892 54204 69028
rect 54400 68892 54612 69028
rect 53992 68816 54612 68892
rect 53992 68750 54204 68816
rect 53992 68686 53998 68750
rect 54062 68686 54204 68750
rect 53992 68680 54204 68686
rect 54400 68680 54612 68816
rect 55216 68892 55428 69028
rect 55624 68892 55836 69028
rect 55216 68816 55836 68892
rect 55216 68750 55428 68816
rect 55216 68686 55222 68750
rect 55286 68686 55428 68750
rect 55216 68680 55428 68686
rect 55624 68750 55836 68816
rect 55624 68686 55766 68750
rect 55830 68686 55836 68750
rect 55624 68680 55836 68686
rect 56440 68892 56788 69028
rect 56848 68892 57060 69028
rect 56440 68816 57060 68892
rect 56440 68680 56788 68816
rect 56848 68750 57060 68816
rect 56848 68686 56854 68750
rect 56918 68686 57060 68750
rect 56848 68680 57060 68686
rect 57800 68892 58012 69028
rect 58072 68892 58420 69028
rect 57800 68816 58420 68892
rect 57800 68750 58012 68816
rect 57800 68686 57806 68750
rect 57870 68686 57942 68750
rect 58006 68686 58012 68750
rect 57800 68680 58012 68686
rect 58072 68680 58420 68816
rect 59024 68892 59236 69028
rect 59432 68892 59644 69028
rect 59024 68816 59644 68892
rect 59024 68750 59236 68816
rect 59024 68686 59030 68750
rect 59094 68686 59236 68750
rect 59024 68680 59236 68686
rect 59432 68750 59644 68816
rect 59432 68686 59574 68750
rect 59638 68686 59644 68750
rect 59432 68680 59644 68686
rect 60248 68756 60460 69028
rect 60656 68756 60868 69028
rect 60248 68750 60868 68756
rect 60248 68686 60254 68750
rect 60318 68686 60798 68750
rect 60862 68686 60868 68750
rect 60248 68680 60868 68686
rect 61472 68952 62092 69028
rect 61472 68750 61684 68952
rect 61472 68686 61478 68750
rect 61542 68686 61684 68750
rect 61472 68680 61684 68686
rect 61880 68756 62092 68952
rect 62696 68892 63044 69028
rect 63104 68892 63316 69028
rect 62696 68816 63316 68892
rect 62696 68756 63044 68816
rect 61880 68750 63044 68756
rect 61880 68686 62702 68750
rect 62766 68686 63044 68750
rect 61880 68680 63044 68686
rect 63104 68680 63316 68816
rect 64056 68952 64676 69028
rect 64056 68750 64268 68952
rect 64056 68686 64062 68750
rect 64126 68686 64268 68750
rect 64056 68680 64268 68686
rect 64328 68680 64676 68952
rect 65280 68892 65492 69028
rect 65688 68892 65900 69028
rect 65280 68816 65900 68892
rect 65280 68750 65492 68816
rect 65280 68686 65286 68750
rect 65350 68686 65492 68750
rect 65280 68680 65492 68686
rect 65688 68680 65900 68816
rect 66504 68892 66716 69028
rect 66912 68892 67124 69028
rect 66504 68816 67124 68892
rect 66504 68750 66716 68816
rect 66504 68686 66510 68750
rect 66574 68686 66716 68750
rect 66504 68680 66716 68686
rect 66912 68750 67124 68816
rect 66912 68686 67054 68750
rect 67118 68686 67124 68750
rect 66912 68680 67124 68686
rect 67728 68892 67940 69028
rect 68136 68892 68348 69028
rect 67728 68816 68348 68892
rect 67728 68750 67940 68816
rect 67728 68686 67734 68750
rect 67798 68686 67940 68750
rect 67728 68680 67940 68686
rect 68136 68750 68348 68816
rect 68136 68686 68278 68750
rect 68342 68686 68348 68750
rect 68136 68680 68348 68686
rect 81872 68750 82220 68756
rect 81872 68686 82014 68750
rect 82078 68686 82220 68750
rect 81872 68544 82220 68686
rect 91936 68750 94188 68756
rect 91936 68686 94118 68750
rect 94182 68686 94188 68750
rect 91936 68680 94188 68686
rect 91936 68544 92148 68680
rect 92616 68544 92828 68680
rect 27744 68212 27956 68348
rect 28288 68342 28500 68348
rect 28288 68278 28294 68342
rect 28358 68278 28500 68342
rect 28288 68212 28500 68278
rect 28968 68342 30404 68348
rect 30638 68342 31084 68348
rect 28968 68278 30334 68342
rect 30398 68278 30404 68342
rect 30600 68278 30606 68342
rect 30670 68278 31084 68342
rect 28968 68272 30404 68278
rect 30638 68272 31084 68278
rect 28968 68212 29180 68272
rect 29512 68212 29724 68272
rect 26656 68206 27684 68212
rect 26656 68142 27614 68206
rect 27678 68142 27684 68206
rect 26656 68136 27684 68142
rect 27744 68136 29180 68212
rect 29278 68206 29724 68212
rect 29240 68142 29246 68206
rect 29310 68142 29724 68206
rect 29278 68136 29724 68142
rect 30192 68136 30404 68272
rect 30736 68212 31084 68272
rect 31416 68342 31628 68348
rect 31726 68342 32308 68348
rect 31416 68278 31558 68342
rect 31622 68278 31628 68342
rect 31688 68278 31694 68342
rect 31758 68278 32308 68342
rect 31416 68212 31628 68278
rect 31726 68272 32308 68278
rect 30736 68136 31628 68212
rect 32096 68212 32308 68272
rect 32640 68342 32852 68348
rect 32640 68278 32782 68342
rect 32846 68278 32852 68342
rect 32640 68212 32852 68278
rect 32096 68136 32852 68212
rect 33320 68342 34756 68348
rect 33320 68278 33326 68342
rect 33390 68278 34142 68342
rect 34206 68278 34756 68342
rect 33320 68272 34756 68278
rect 33320 68136 33532 68272
rect 33864 68136 34212 68272
rect 34544 68136 34756 68272
rect 35224 68342 35436 68348
rect 35224 68278 35230 68342
rect 35294 68278 35436 68342
rect 35224 68136 35436 68278
rect 35768 68342 36660 68348
rect 35768 68278 35774 68342
rect 35838 68278 36590 68342
rect 36654 68278 36660 68342
rect 35768 68272 36660 68278
rect 35768 68136 35980 68272
rect 36448 68212 36660 68272
rect 36992 68342 37884 68348
rect 36992 68278 37814 68342
rect 37878 68278 37884 68342
rect 36992 68272 37884 68278
rect 36992 68212 37340 68272
rect 36448 68136 37340 68212
rect 37672 68136 37884 68272
rect 38352 68342 38564 68348
rect 38352 68278 38358 68342
rect 38422 68278 38564 68342
rect 38352 68212 38564 68278
rect 38896 68342 39108 68348
rect 39342 68342 41012 68348
rect 38896 68278 39038 68342
rect 39102 68278 39108 68342
rect 39304 68278 39310 68342
rect 39374 68278 40262 68342
rect 40326 68278 41012 68342
rect 38896 68212 39108 68278
rect 39342 68272 41012 68278
rect 38352 68136 39108 68212
rect 39576 68136 39788 68272
rect 40120 68136 40332 68272
rect 40800 68212 41012 68272
rect 41344 68342 41964 68348
rect 41344 68278 41894 68342
rect 41958 68278 41964 68342
rect 41344 68272 41964 68278
rect 42024 68342 42916 68348
rect 42024 68278 42846 68342
rect 42910 68278 42916 68342
rect 42024 68272 42916 68278
rect 41344 68212 41692 68272
rect 42024 68212 42236 68272
rect 40800 68136 42236 68212
rect 42704 68136 42916 68272
rect 43248 68342 43460 68348
rect 43248 68278 43390 68342
rect 43454 68278 43460 68342
rect 43248 68136 43460 68278
rect 43928 68342 45364 68348
rect 43928 68278 44070 68342
rect 44134 68278 45364 68342
rect 43928 68272 45364 68278
rect 43928 68136 44140 68272
rect 44472 68136 44820 68272
rect 45152 68212 45364 68272
rect 45832 68342 46588 68348
rect 45832 68278 45838 68342
rect 45902 68278 46518 68342
rect 46582 68278 46588 68342
rect 45832 68272 46588 68278
rect 45832 68212 46044 68272
rect 45152 68136 46044 68212
rect 46376 68136 46588 68272
rect 47056 68342 47268 68348
rect 47056 68278 47062 68342
rect 47126 68278 47268 68342
rect 47056 68212 47268 68278
rect 47600 68342 47948 68348
rect 47600 68278 47742 68342
rect 47806 68278 47948 68342
rect 47600 68212 47948 68278
rect 48280 68342 49172 68348
rect 48280 68278 48966 68342
rect 49030 68278 49172 68342
rect 48280 68272 49172 68278
rect 48280 68212 48492 68272
rect 47056 68136 48492 68212
rect 48960 68212 49172 68272
rect 49504 68212 49716 68348
rect 50184 68342 50668 68348
rect 50184 68278 50598 68342
rect 50662 68278 50668 68342
rect 50184 68272 50668 68278
rect 50728 68342 51620 68348
rect 50728 68278 51550 68342
rect 51614 68278 51620 68342
rect 50728 68272 51620 68278
rect 50184 68212 50396 68272
rect 50728 68212 50940 68272
rect 48960 68136 50940 68212
rect 51408 68136 51620 68272
rect 51952 68342 52300 68348
rect 51952 68278 52094 68342
rect 52158 68278 52300 68342
rect 51952 68212 52300 68278
rect 52632 68342 52844 68348
rect 53078 68342 53524 68348
rect 52632 68278 52774 68342
rect 52838 68278 52844 68342
rect 53040 68278 53046 68342
rect 53110 68278 53524 68342
rect 52632 68212 52844 68278
rect 53078 68272 53524 68278
rect 51952 68136 52844 68212
rect 53312 68212 53524 68272
rect 53856 68342 54068 68348
rect 53856 68278 53998 68342
rect 54062 68278 54068 68342
rect 53856 68212 54068 68278
rect 54536 68342 55428 68348
rect 54536 68278 55222 68342
rect 55286 68278 55428 68342
rect 54536 68272 55428 68278
rect 54536 68212 54748 68272
rect 53312 68136 54748 68212
rect 55080 68136 55428 68272
rect 55760 68342 55972 68348
rect 55760 68278 55766 68342
rect 55830 68278 55972 68342
rect 55760 68212 55972 68278
rect 56440 68342 56924 68348
rect 56440 68278 56854 68342
rect 56918 68278 56924 68342
rect 56440 68272 56924 68278
rect 56984 68342 57876 68348
rect 57974 68342 58556 68348
rect 56984 68278 57806 68342
rect 57870 68278 57876 68342
rect 57936 68278 57942 68342
rect 58006 68278 58556 68342
rect 56984 68272 57876 68278
rect 57974 68272 58556 68278
rect 56440 68212 56652 68272
rect 56984 68212 57196 68272
rect 55760 68136 57196 68212
rect 57664 68136 57876 68272
rect 58208 68212 58556 68272
rect 58888 68342 59100 68348
rect 58888 68278 59030 68342
rect 59094 68278 59100 68342
rect 58888 68212 59100 68278
rect 58208 68136 59100 68212
rect 59568 68342 59780 68348
rect 59568 68278 59574 68342
rect 59638 68278 59780 68342
rect 59568 68212 59780 68278
rect 60112 68342 60324 68348
rect 60112 68278 60254 68342
rect 60318 68278 60324 68342
rect 60112 68212 60324 68278
rect 59568 68136 60324 68212
rect 60792 68342 61548 68348
rect 60792 68278 60798 68342
rect 60862 68278 61478 68342
rect 61542 68278 61548 68342
rect 60792 68272 61548 68278
rect 60792 68136 61004 68272
rect 61336 68136 61548 68272
rect 62016 68212 62228 68348
rect 62560 68342 62908 68348
rect 62560 68278 62702 68342
rect 62766 68278 62908 68342
rect 62560 68212 62908 68278
rect 63240 68342 64132 68348
rect 63240 68278 64062 68342
rect 64126 68278 64132 68342
rect 63240 68272 64132 68278
rect 63240 68212 63452 68272
rect 62016 68136 63452 68212
rect 63920 68212 64132 68272
rect 64464 68212 64676 68348
rect 65144 68342 66580 68348
rect 65144 68278 65286 68342
rect 65350 68278 66510 68342
rect 66574 68278 66580 68342
rect 65144 68272 66580 68278
rect 65144 68212 65356 68272
rect 63920 68136 65356 68212
rect 65688 68136 66036 68272
rect 66368 68136 66580 68272
rect 67048 68342 67804 68348
rect 67048 68278 67054 68342
rect 67118 68278 67734 68342
rect 67798 68278 67804 68342
rect 67048 68272 67804 68278
rect 67048 68136 67260 68272
rect 67592 68136 67804 68272
rect 68272 68342 70388 68348
rect 68272 68278 68278 68342
rect 68342 68278 70318 68342
rect 70382 68278 70388 68342
rect 68272 68272 70388 68278
rect 68272 68136 68484 68272
rect 26656 68076 26868 68136
rect 26656 68070 27004 68076
rect 26656 68006 26934 68070
rect 26998 68006 27004 68070
rect 26656 68000 27004 68006
rect 69360 68070 69572 68212
rect 69360 68006 69366 68070
rect 69430 68006 69572 68070
rect 69360 68000 69572 68006
rect 70312 68070 70524 68076
rect 70312 68006 70318 68070
rect 70382 68006 70524 68070
rect 70312 67804 70524 68006
rect 73032 67940 73244 68076
rect 73848 68070 74740 68076
rect 73848 68006 74670 68070
rect 74734 68006 74740 68070
rect 73848 68000 74740 68006
rect 73848 67940 74060 68000
rect 73032 67864 74060 67940
rect 73032 67804 73244 67864
rect 26928 67798 27276 67804
rect 26928 67734 26934 67798
rect 26998 67734 27276 67798
rect 1224 67662 1980 67668
rect 1224 67598 1230 67662
rect 1294 67600 1980 67662
rect 1294 67598 1818 67600
rect 1224 67592 1818 67598
rect 1768 67544 1818 67592
rect 1874 67544 1980 67600
rect 26928 67592 27276 67734
rect 68952 67798 69436 67804
rect 68952 67734 68958 67798
rect 69022 67734 69366 67798
rect 69430 67734 69436 67798
rect 68952 67728 69436 67734
rect 70312 67728 73244 67804
rect 73848 67798 74060 67864
rect 73848 67734 73854 67798
rect 73918 67734 74060 67798
rect 73848 67728 74060 67734
rect 68952 67592 69164 67728
rect 1768 67456 1980 67544
rect 27200 67532 27276 67592
rect 69088 67532 69164 67592
rect 20400 67184 20612 67396
rect 20808 67254 21020 67396
rect 21216 67260 21564 67396
rect 21118 67254 21564 67260
rect 20808 67190 20950 67254
rect 21014 67190 21020 67254
rect 21080 67190 21086 67254
rect 21150 67190 21358 67254
rect 21422 67190 21564 67254
rect 20808 67184 21020 67190
rect 21118 67184 21564 67190
rect 21624 67254 21836 67396
rect 21624 67190 21766 67254
rect 21830 67190 21836 67254
rect 21624 67184 21836 67190
rect 22032 67254 22244 67396
rect 26928 67320 27276 67532
rect 68952 67320 69164 67532
rect 94112 67662 94732 67668
rect 94112 67600 94662 67662
rect 94112 67544 94176 67600
rect 94232 67598 94662 67600
rect 94726 67598 94732 67662
rect 94232 67592 94732 67598
rect 94232 67544 94324 67592
rect 94112 67456 94324 67544
rect 73848 67390 74060 67396
rect 73848 67326 73854 67390
rect 73918 67326 74060 67390
rect 27064 67260 27140 67320
rect 68952 67260 69028 67320
rect 22032 67190 22038 67254
rect 22102 67190 22244 67254
rect 22032 67184 22244 67190
rect 20400 67124 20476 67184
rect 20400 66982 20612 67124
rect 26928 67118 27276 67260
rect 26928 67054 27206 67118
rect 27270 67054 27276 67118
rect 26928 67048 27276 67054
rect 27200 66988 27276 67048
rect 20400 66918 20406 66982
rect 20470 66918 20612 66982
rect 20400 66912 20612 66918
rect 20808 66982 21156 66988
rect 20808 66918 20950 66982
rect 21014 66918 21086 66982
rect 21150 66918 21156 66982
rect 20808 66912 21156 66918
rect 21216 66982 21564 66988
rect 21216 66918 21358 66982
rect 21422 66918 21564 66982
rect 20808 66776 21020 66912
rect 21216 66776 21564 66918
rect 21624 66982 21836 66988
rect 21624 66918 21766 66982
rect 21830 66918 21836 66982
rect 21624 66846 21836 66918
rect 21624 66782 21630 66846
rect 21694 66782 21836 66846
rect 21624 66776 21836 66782
rect 22032 66982 22244 66988
rect 22032 66918 22038 66982
rect 22102 66918 22244 66982
rect 22032 66846 22244 66918
rect 22032 66782 22038 66846
rect 22102 66782 22244 66846
rect 22032 66776 22244 66782
rect 26928 66846 27276 66988
rect 26928 66782 27206 66846
rect 27270 66782 27276 66846
rect 20944 66716 21020 66776
rect 21488 66716 21564 66776
rect 20400 66710 20612 66716
rect 20400 66646 20406 66710
rect 20470 66646 20612 66710
rect 20400 66368 20612 66646
rect 20808 66368 21020 66716
rect 21216 66368 21564 66716
rect 21624 66574 21836 66580
rect 21624 66510 21630 66574
rect 21694 66510 21836 66574
rect 21624 66368 21836 66510
rect 22032 66574 22244 66580
rect 22032 66510 22038 66574
rect 22102 66510 22244 66574
rect 22032 66368 22244 66510
rect 20536 66308 20612 66368
rect 21216 66308 21292 66368
rect 20400 66166 20612 66308
rect 20944 66232 21292 66308
rect 21624 66308 21700 66368
rect 22168 66308 22244 66368
rect 20944 66172 21020 66232
rect 20400 66102 20542 66166
rect 20606 66102 20612 66166
rect 20400 66096 20612 66102
rect 20808 66096 21564 66172
rect 1224 66030 1980 66036
rect 1224 65966 1230 66030
rect 1294 65966 1980 66030
rect 1224 65960 1980 65966
rect 20808 65960 21020 66096
rect 21216 65960 21564 66096
rect 21624 65960 21836 66308
rect 1768 65920 1980 65960
rect 1768 65864 1818 65920
rect 1874 65864 1980 65920
rect 21352 65900 21428 65960
rect 21760 65900 21836 65960
rect 1768 65824 1980 65864
rect 20400 65894 20612 65900
rect 20400 65830 20542 65894
rect 20606 65830 20612 65894
rect 20400 65758 20612 65830
rect 20400 65694 20406 65758
rect 20470 65694 20612 65758
rect 20400 65688 20612 65694
rect 20808 65824 21564 65900
rect 20808 65758 21020 65824
rect 20808 65694 20814 65758
rect 20878 65694 21020 65758
rect 20808 65688 21020 65694
rect 21216 65688 21564 65824
rect 21624 65552 21836 65900
rect 22032 65960 22244 66308
rect 26928 66504 27276 66782
rect 68952 67118 69164 67260
rect 73848 67254 74060 67326
rect 73848 67190 73990 67254
rect 74054 67190 74060 67254
rect 73848 67184 74060 67190
rect 74256 67390 74604 67396
rect 74256 67326 74534 67390
rect 74598 67326 74604 67390
rect 74256 67320 74604 67326
rect 74664 67320 75284 67396
rect 74256 67254 74468 67320
rect 74256 67190 74398 67254
rect 74462 67190 74468 67254
rect 74256 67184 74468 67190
rect 74664 67254 74876 67320
rect 74664 67190 74670 67254
rect 74734 67190 74876 67254
rect 74664 67184 74876 67190
rect 75072 67184 75284 67320
rect 75480 67184 75692 67396
rect 68952 67054 69094 67118
rect 69158 67054 69164 67118
rect 68952 67048 69164 67054
rect 75480 67124 75556 67184
rect 91936 67124 92148 67260
rect 92518 67254 95412 67260
rect 92480 67190 92486 67254
rect 92550 67190 95342 67254
rect 95406 67190 95412 67254
rect 92518 67184 95412 67190
rect 92616 67124 92828 67184
rect 68952 66988 69028 67048
rect 68952 66846 69164 66988
rect 68952 66782 69094 66846
rect 69158 66782 69164 66846
rect 68952 66574 69164 66782
rect 73848 66982 74060 66988
rect 73848 66918 73990 66982
rect 74054 66918 74060 66982
rect 73848 66846 74060 66918
rect 73848 66782 73990 66846
rect 74054 66782 74060 66846
rect 73848 66776 74060 66782
rect 74256 66982 74468 66988
rect 74256 66918 74398 66982
rect 74462 66918 74468 66982
rect 74256 66846 74468 66918
rect 74256 66782 74262 66846
rect 74326 66782 74468 66846
rect 74256 66776 74468 66782
rect 74664 66982 74876 66988
rect 74664 66918 74670 66982
rect 74734 66918 74876 66982
rect 74664 66776 74876 66918
rect 75072 66852 75284 66988
rect 75480 66982 75692 67124
rect 91936 67118 92828 67124
rect 91936 67054 92622 67118
rect 92686 67054 92828 67118
rect 91936 67048 92828 67054
rect 75480 66918 75622 66982
rect 75686 66918 75692 66982
rect 75480 66912 75692 66918
rect 74936 66776 75284 66852
rect 74664 66716 74740 66776
rect 74936 66716 75012 66776
rect 74664 66640 75012 66716
rect 68952 66510 69094 66574
rect 69158 66510 69164 66574
rect 68952 66504 69164 66510
rect 73848 66574 74060 66580
rect 73848 66510 73990 66574
rect 74054 66510 74060 66574
rect 26928 66444 27004 66504
rect 22032 65900 22108 65960
rect 22032 65552 22244 65900
rect 26928 65894 27276 66444
rect 26928 65830 26934 65894
rect 26998 65830 27276 65894
rect 26928 65824 27276 65830
rect 68952 66302 69164 66444
rect 68952 66238 68958 66302
rect 69022 66238 69094 66302
rect 69158 66238 69164 66302
rect 68952 66030 69164 66238
rect 68952 65966 68958 66030
rect 69022 65966 69164 66030
rect 68952 65894 69164 65966
rect 68952 65830 68958 65894
rect 69022 65830 69164 65894
rect 68952 65824 69164 65830
rect 73848 66368 74060 66510
rect 74256 66574 74468 66580
rect 74256 66510 74262 66574
rect 74326 66510 74468 66574
rect 74256 66368 74468 66510
rect 74664 66444 74876 66640
rect 75072 66444 75284 66716
rect 74664 66438 75284 66444
rect 74664 66374 75078 66438
rect 75142 66374 75284 66438
rect 74664 66368 75284 66374
rect 75480 66710 75692 66716
rect 75480 66646 75622 66710
rect 75686 66646 75692 66710
rect 75480 66368 75692 66646
rect 73848 66308 73924 66368
rect 74392 66308 74468 66368
rect 73848 65960 74060 66308
rect 74256 65960 74468 66308
rect 75480 66308 75556 66368
rect 73848 65900 73924 65960
rect 74392 65900 74468 65960
rect 26928 65622 27276 65628
rect 26928 65558 26934 65622
rect 26998 65558 27276 65622
rect 21624 65492 21700 65552
rect 22032 65492 22108 65552
rect 20400 65486 20612 65492
rect 20400 65422 20406 65486
rect 20470 65422 20612 65486
rect 20400 65350 20612 65422
rect 20400 65286 20406 65350
rect 20470 65286 20612 65350
rect 20400 65280 20612 65286
rect 20808 65486 21020 65492
rect 20808 65422 20814 65486
rect 20878 65422 21020 65486
rect 20808 65144 21020 65422
rect 21216 65144 21564 65492
rect 21624 65350 21836 65492
rect 21624 65286 21766 65350
rect 21830 65286 21836 65350
rect 21624 65280 21836 65286
rect 22032 65350 22244 65492
rect 22032 65286 22038 65350
rect 22102 65286 22244 65350
rect 22032 65280 22244 65286
rect 26928 65486 27276 65558
rect 26928 65422 27206 65486
rect 27270 65422 27276 65486
rect 26928 65280 27276 65422
rect 68952 65622 69164 65628
rect 68952 65558 68958 65622
rect 69022 65558 69164 65622
rect 68952 65280 69164 65558
rect 73848 65552 74060 65900
rect 74256 65552 74468 65900
rect 74664 65960 74876 66172
rect 75072 66166 75284 66172
rect 75072 66102 75078 66166
rect 75142 66102 75284 66166
rect 75072 65960 75284 66102
rect 75480 66166 75692 66308
rect 75480 66102 75486 66166
rect 75550 66102 75692 66166
rect 75480 66096 75692 66102
rect 94112 66030 94732 66036
rect 94112 65966 94662 66030
rect 94726 65966 94732 66030
rect 94112 65960 94732 65966
rect 74664 65900 74740 65960
rect 75072 65900 75148 65960
rect 94112 65920 94324 65960
rect 94112 65900 94176 65920
rect 74664 65758 74876 65900
rect 75072 65764 75284 65900
rect 74974 65758 75284 65764
rect 74664 65694 74670 65758
rect 74734 65694 74876 65758
rect 74936 65694 74942 65758
rect 75006 65694 75284 65758
rect 74664 65688 74876 65694
rect 74974 65688 75284 65694
rect 75480 65894 75692 65900
rect 75480 65830 75486 65894
rect 75550 65830 75692 65894
rect 75480 65758 75692 65830
rect 75480 65694 75486 65758
rect 75550 65694 75692 65758
rect 75480 65688 75692 65694
rect 91936 65764 92148 65900
rect 92616 65864 94176 65900
rect 94232 65864 94324 65920
rect 92616 65824 94324 65864
rect 92616 65764 92828 65824
rect 91936 65688 92828 65764
rect 73848 65492 73924 65552
rect 74256 65492 74332 65552
rect 73848 65350 74060 65492
rect 73848 65286 73854 65350
rect 73918 65286 74060 65350
rect 73848 65280 74060 65286
rect 74256 65350 74468 65492
rect 74256 65286 74262 65350
rect 74326 65286 74468 65350
rect 74256 65280 74468 65286
rect 74664 65486 75012 65492
rect 74664 65422 74670 65486
rect 74734 65422 74942 65486
rect 75006 65422 75012 65486
rect 74664 65416 75012 65422
rect 74664 65356 74876 65416
rect 75072 65356 75284 65492
rect 74664 65280 75284 65356
rect 75480 65486 75692 65492
rect 75480 65422 75486 65486
rect 75550 65422 75692 65486
rect 75480 65350 75692 65422
rect 75480 65286 75622 65350
rect 75686 65286 75692 65350
rect 75480 65280 75692 65286
rect 27200 65220 27276 65280
rect 69088 65220 69164 65280
rect 20944 65084 21020 65144
rect 21488 65084 21564 65144
rect 26928 65214 27276 65220
rect 26928 65150 27206 65214
rect 27270 65150 27276 65214
rect 20400 65078 20612 65084
rect 20400 65014 20406 65078
rect 20470 65014 20612 65078
rect 20400 64942 20612 65014
rect 20400 64878 20406 64942
rect 20470 64878 20612 64942
rect 20400 64872 20612 64878
rect 20808 65008 21564 65084
rect 20808 64872 21020 65008
rect 21216 64942 21564 65008
rect 21216 64878 21494 64942
rect 21558 64878 21564 64942
rect 21216 64872 21564 64878
rect 21624 65078 21836 65084
rect 21624 65014 21766 65078
rect 21830 65014 21836 65078
rect 21624 64942 21836 65014
rect 21624 64878 21766 64942
rect 21830 64878 21836 64942
rect 21624 64872 21836 64878
rect 22032 65078 22244 65084
rect 22032 65014 22038 65078
rect 22102 65014 22244 65078
rect 22032 64942 22244 65014
rect 26928 65008 27276 65150
rect 27200 64948 27276 65008
rect 22032 64878 22038 64942
rect 22102 64878 22244 64942
rect 22032 64872 22244 64878
rect 26928 64736 27276 64948
rect 68952 65008 69164 65220
rect 74664 65220 74876 65280
rect 74664 65144 75012 65220
rect 75072 65144 75284 65280
rect 74800 65084 74876 65144
rect 73848 65078 74060 65084
rect 73848 65014 73854 65078
rect 73918 65014 74060 65078
rect 68952 64948 69028 65008
rect 68952 64736 69164 64948
rect 73848 64942 74060 65014
rect 73848 64878 73990 64942
rect 74054 64878 74060 64942
rect 73848 64872 74060 64878
rect 74256 65078 74468 65084
rect 74256 65014 74262 65078
rect 74326 65014 74468 65078
rect 74256 64942 74468 65014
rect 74256 64878 74262 64942
rect 74326 64878 74468 64942
rect 74256 64872 74468 64878
rect 74664 64872 74876 65084
rect 74936 65084 75012 65144
rect 74936 65008 75284 65084
rect 75072 64942 75284 65008
rect 75072 64878 75078 64942
rect 75142 64878 75284 64942
rect 75072 64872 75284 64878
rect 75480 65078 75692 65084
rect 75480 65014 75622 65078
rect 75686 65014 75692 65078
rect 75480 64942 75692 65014
rect 75480 64878 75486 64942
rect 75550 64878 75692 64942
rect 75480 64872 75692 64878
rect 27064 64676 27140 64736
rect 68952 64676 69028 64736
rect 20400 64670 20612 64676
rect 20400 64606 20406 64670
rect 20470 64606 20612 64670
rect 20400 64534 20612 64606
rect 20400 64470 20542 64534
rect 20606 64470 20612 64534
rect 20400 64464 20612 64470
rect 20808 64534 21020 64676
rect 20808 64470 20814 64534
rect 20878 64470 21020 64534
rect 20808 64464 21020 64470
rect 21216 64670 21564 64676
rect 21216 64606 21494 64670
rect 21558 64606 21564 64670
rect 21216 64534 21564 64606
rect 21216 64470 21494 64534
rect 21558 64470 21564 64534
rect 21216 64464 21564 64470
rect 21624 64670 21836 64676
rect 21624 64606 21766 64670
rect 21830 64606 21836 64670
rect 21624 64534 21836 64606
rect 21624 64470 21630 64534
rect 21694 64470 21836 64534
rect 21624 64464 21836 64470
rect 22032 64670 22244 64676
rect 22032 64606 22038 64670
rect 22102 64606 22244 64670
rect 22032 64534 22244 64606
rect 22032 64470 22038 64534
rect 22102 64470 22244 64534
rect 22032 64464 22244 64470
rect 26928 64464 27276 64676
rect 68952 64464 69164 64676
rect 73848 64670 74060 64676
rect 73848 64606 73990 64670
rect 74054 64606 74060 64670
rect 73848 64534 74060 64606
rect 73848 64470 73854 64534
rect 73918 64470 74060 64534
rect 73848 64464 74060 64470
rect 74256 64670 74468 64676
rect 74256 64606 74262 64670
rect 74326 64606 74468 64670
rect 74256 64534 74468 64606
rect 74256 64470 74398 64534
rect 74462 64470 74468 64534
rect 74256 64464 74468 64470
rect 74664 64540 74876 64676
rect 75072 64670 75284 64676
rect 75072 64606 75078 64670
rect 75142 64606 75284 64670
rect 75072 64540 75284 64606
rect 74664 64534 75284 64540
rect 74664 64470 74806 64534
rect 74870 64470 75284 64534
rect 74664 64464 75284 64470
rect 75480 64670 75692 64676
rect 75480 64606 75486 64670
rect 75550 64606 75692 64670
rect 75480 64534 75692 64606
rect 75480 64470 75622 64534
rect 75686 64470 75692 64534
rect 75480 64464 75692 64470
rect 91936 64534 92556 64540
rect 91936 64470 92486 64534
rect 92550 64470 92556 64534
rect 91936 64464 92556 64470
rect 26928 64404 27004 64464
rect 69088 64404 69164 64464
rect 1768 64240 1980 64268
rect 1768 64184 1818 64240
rect 1874 64184 1980 64240
rect 1768 64132 1980 64184
rect 1224 64126 1980 64132
rect 1224 64062 1230 64126
rect 1294 64062 1980 64126
rect 1224 64056 1980 64062
rect 20400 64262 20612 64268
rect 20400 64198 20542 64262
rect 20606 64198 20612 64262
rect 20400 64126 20612 64198
rect 20400 64062 20542 64126
rect 20606 64062 20612 64126
rect 20400 64056 20612 64062
rect 20808 64262 21020 64268
rect 20808 64198 20814 64262
rect 20878 64198 21020 64262
rect 20808 64126 21020 64198
rect 21216 64262 21564 64268
rect 21216 64198 21494 64262
rect 21558 64198 21564 64262
rect 21216 64132 21564 64198
rect 21118 64126 21564 64132
rect 20808 64062 20950 64126
rect 21014 64062 21020 64126
rect 21080 64062 21086 64126
rect 21150 64062 21222 64126
rect 21286 64062 21564 64126
rect 20808 64056 21020 64062
rect 21118 64056 21564 64062
rect 21624 64262 21836 64268
rect 21624 64198 21630 64262
rect 21694 64198 21836 64262
rect 21624 64126 21836 64198
rect 21624 64062 21766 64126
rect 21830 64062 21836 64126
rect 21624 64056 21836 64062
rect 22032 64262 22244 64268
rect 22032 64198 22038 64262
rect 22102 64198 22244 64262
rect 22032 64126 22244 64198
rect 26928 64192 27276 64404
rect 68952 64192 69164 64404
rect 74800 64404 74876 64464
rect 91936 64404 92148 64464
rect 92616 64404 92828 64540
rect 74800 64328 75148 64404
rect 91936 64328 92828 64404
rect 75072 64268 75148 64328
rect 27064 64132 27140 64192
rect 69088 64132 69164 64192
rect 22032 64062 22038 64126
rect 22102 64062 22244 64126
rect 22032 64056 22244 64062
rect 26928 63920 27276 64132
rect 27200 63860 27276 63920
rect 20400 63854 20612 63860
rect 20400 63790 20542 63854
rect 20606 63790 20612 63854
rect 20400 63718 20612 63790
rect 20400 63654 20542 63718
rect 20606 63654 20612 63718
rect 20400 63648 20612 63654
rect 20808 63854 21156 63860
rect 20808 63790 20950 63854
rect 21014 63790 21086 63854
rect 21150 63790 21156 63854
rect 20808 63784 21156 63790
rect 21216 63854 21564 63860
rect 21216 63790 21222 63854
rect 21286 63790 21564 63854
rect 20808 63718 21020 63784
rect 20808 63654 20814 63718
rect 20878 63654 21020 63718
rect 20808 63648 21020 63654
rect 21216 63648 21564 63790
rect 21624 63854 21836 63860
rect 21624 63790 21766 63854
rect 21830 63790 21836 63854
rect 21624 63718 21836 63790
rect 21624 63654 21766 63718
rect 21830 63654 21836 63718
rect 21624 63648 21836 63654
rect 22032 63854 22244 63860
rect 22032 63790 22038 63854
rect 22102 63790 22244 63854
rect 22032 63718 22244 63790
rect 22032 63654 22038 63718
rect 22102 63654 22244 63718
rect 22032 63648 22244 63654
rect 26928 63648 27276 63860
rect 68952 63920 69164 64132
rect 73848 64262 74060 64268
rect 73848 64198 73854 64262
rect 73918 64198 74060 64262
rect 73848 64126 74060 64198
rect 73848 64062 73990 64126
rect 74054 64062 74060 64126
rect 73848 64056 74060 64062
rect 74256 64262 74468 64268
rect 74256 64198 74398 64262
rect 74462 64198 74468 64262
rect 74256 64126 74468 64198
rect 74256 64062 74398 64126
rect 74462 64062 74468 64126
rect 74256 64056 74468 64062
rect 74664 64262 74876 64268
rect 74664 64198 74806 64262
rect 74870 64198 74876 64262
rect 74664 64056 74876 64198
rect 75072 64056 75284 64268
rect 75480 64262 75692 64268
rect 75480 64198 75622 64262
rect 75686 64198 75692 64262
rect 75480 64126 75692 64198
rect 75480 64062 75622 64126
rect 75686 64062 75692 64126
rect 75480 64056 75692 64062
rect 94112 64240 94324 64268
rect 94112 64184 94176 64240
rect 94232 64184 94324 64240
rect 94112 64132 94324 64184
rect 94112 64126 94732 64132
rect 94112 64062 94662 64126
rect 94726 64062 94732 64126
rect 94112 64056 94732 64062
rect 75072 63996 75148 64056
rect 74800 63920 75148 63996
rect 68952 63860 69028 63920
rect 74800 63860 74876 63920
rect 68952 63648 69164 63860
rect 73848 63854 74060 63860
rect 73848 63790 73990 63854
rect 74054 63790 74060 63854
rect 73848 63718 74060 63790
rect 73848 63654 73990 63718
rect 74054 63654 74060 63718
rect 73848 63648 74060 63654
rect 74256 63854 74468 63860
rect 74256 63790 74398 63854
rect 74462 63790 74468 63854
rect 74256 63718 74468 63790
rect 74256 63654 74262 63718
rect 74326 63654 74468 63718
rect 74256 63648 74468 63654
rect 74664 63784 75284 63860
rect 74664 63648 74876 63784
rect 75072 63724 75284 63784
rect 74974 63718 75284 63724
rect 74936 63654 74942 63718
rect 75006 63654 75284 63718
rect 74974 63648 75284 63654
rect 75480 63854 75692 63860
rect 75480 63790 75622 63854
rect 75686 63790 75692 63854
rect 75480 63718 75692 63790
rect 75480 63654 75622 63718
rect 75686 63654 75692 63718
rect 75480 63648 75692 63654
rect 27064 63588 27140 63648
rect 68952 63588 69028 63648
rect 20400 63446 20612 63452
rect 20400 63382 20542 63446
rect 20606 63382 20612 63446
rect 20400 63240 20612 63382
rect 20808 63446 21020 63452
rect 20808 63382 20814 63446
rect 20878 63382 21020 63446
rect 20808 63310 21020 63382
rect 20808 63246 20814 63310
rect 20878 63246 21020 63310
rect 20808 63240 21020 63246
rect 21216 63310 21564 63452
rect 21216 63246 21494 63310
rect 21558 63246 21564 63310
rect 21216 63240 21564 63246
rect 21624 63446 21836 63452
rect 21624 63382 21766 63446
rect 21830 63382 21836 63446
rect 21624 63310 21836 63382
rect 21624 63246 21630 63310
rect 21694 63246 21836 63310
rect 21624 63240 21836 63246
rect 22032 63446 22244 63452
rect 22032 63382 22038 63446
rect 22102 63382 22244 63446
rect 22032 63310 22244 63382
rect 26928 63376 27276 63588
rect 68952 63376 69164 63588
rect 27200 63316 27276 63376
rect 69088 63316 69164 63376
rect 22032 63246 22174 63310
rect 22238 63246 22244 63310
rect 22032 63240 22244 63246
rect 20400 63180 20476 63240
rect 20400 62832 20612 63180
rect 26928 63174 27276 63316
rect 26928 63110 27206 63174
rect 27270 63110 27276 63174
rect 26928 63104 27276 63110
rect 68952 63104 69164 63316
rect 73848 63446 74060 63452
rect 73848 63382 73990 63446
rect 74054 63382 74060 63446
rect 73848 63310 74060 63382
rect 73848 63246 73854 63310
rect 73918 63246 74060 63310
rect 73848 63240 74060 63246
rect 74256 63446 74468 63452
rect 74256 63382 74262 63446
rect 74326 63382 74468 63446
rect 74256 63310 74468 63382
rect 74256 63246 74398 63310
rect 74462 63246 74468 63310
rect 74256 63240 74468 63246
rect 74664 63446 75012 63452
rect 74664 63382 74942 63446
rect 75006 63382 75012 63446
rect 74664 63376 75012 63382
rect 74664 63316 74876 63376
rect 75072 63316 75284 63452
rect 74664 63310 75284 63316
rect 74664 63246 74806 63310
rect 74870 63246 75214 63310
rect 75278 63246 75284 63310
rect 74664 63240 75284 63246
rect 75480 63446 75692 63452
rect 75480 63382 75622 63446
rect 75686 63382 75692 63446
rect 75480 63240 75692 63382
rect 75616 63180 75692 63240
rect 27200 63044 27276 63104
rect 69088 63044 69164 63104
rect 20808 63038 21020 63044
rect 20808 62974 20814 63038
rect 20878 62974 21020 63038
rect 20808 62832 21020 62974
rect 21216 63038 21564 63044
rect 21216 62974 21494 63038
rect 21558 62974 21564 63038
rect 21216 62908 21564 62974
rect 20400 62772 20476 62832
rect 20944 62772 21020 62832
rect 21080 62832 21564 62908
rect 21624 63038 21836 63044
rect 21624 62974 21630 63038
rect 21694 62974 21836 63038
rect 21624 62902 21836 62974
rect 21624 62838 21766 62902
rect 21830 62838 21836 62902
rect 21624 62832 21836 62838
rect 22032 63038 22244 63044
rect 22032 62974 22174 63038
rect 22238 62974 22244 63038
rect 22032 62902 22244 62974
rect 22032 62838 22174 62902
rect 22238 62838 22244 62902
rect 22032 62832 22244 62838
rect 26928 62902 27276 63044
rect 26928 62838 27070 62902
rect 27134 62838 27206 62902
rect 27270 62838 27276 62902
rect 21080 62772 21156 62832
rect 1768 62560 1980 62636
rect 1768 62504 1818 62560
rect 1874 62504 1980 62560
rect 1768 62500 1980 62504
rect 1224 62494 1980 62500
rect 1224 62430 1230 62494
rect 1294 62430 1980 62494
rect 1224 62424 1980 62430
rect 20400 62424 20612 62772
rect 20808 62696 21156 62772
rect 20808 62636 21020 62696
rect 21216 62636 21564 62772
rect 20808 62560 21564 62636
rect 20808 62494 21020 62560
rect 20808 62430 20814 62494
rect 20878 62430 21020 62494
rect 20808 62424 21020 62430
rect 21216 62424 21564 62560
rect 21624 62630 21836 62636
rect 21624 62566 21766 62630
rect 21830 62566 21836 62630
rect 21624 62424 21836 62566
rect 22032 62630 22244 62636
rect 22032 62566 22174 62630
rect 22238 62566 22244 62630
rect 22032 62424 22244 62566
rect 26928 62560 27276 62838
rect 27200 62500 27276 62560
rect 20400 62364 20476 62424
rect 21760 62364 21836 62424
rect 22168 62364 22244 62424
rect 20400 62222 20612 62364
rect 20400 62158 20542 62222
rect 20606 62158 20612 62222
rect 20400 62152 20612 62158
rect 20808 62222 21020 62228
rect 20808 62158 20814 62222
rect 20878 62158 21020 62222
rect 20808 62016 21020 62158
rect 21216 62092 21564 62228
rect 21080 62016 21564 62092
rect 21624 62016 21836 62364
rect 22032 62016 22244 62364
rect 26928 62358 27276 62500
rect 26928 62294 26934 62358
rect 26998 62294 27070 62358
rect 27134 62294 27276 62358
rect 26928 62086 27276 62294
rect 26928 62022 26934 62086
rect 26998 62022 27276 62086
rect 20808 61956 20884 62016
rect 21080 61956 21156 62016
rect 21352 61956 21428 62016
rect 21624 61956 21700 62016
rect 22032 61956 22108 62016
rect 20400 61950 20612 61956
rect 20400 61886 20542 61950
rect 20606 61886 20612 61950
rect 20400 61814 20612 61886
rect 20400 61750 20406 61814
rect 20470 61750 20612 61814
rect 20400 61744 20612 61750
rect 20808 61880 21156 61956
rect 20808 61820 21020 61880
rect 20808 61814 21156 61820
rect 20808 61750 20950 61814
rect 21014 61750 21086 61814
rect 21150 61750 21156 61814
rect 20808 61744 21156 61750
rect 21216 61744 21564 61956
rect 21624 61608 21836 61956
rect 22032 61608 22244 61956
rect 26928 61950 27276 62022
rect 26928 61886 26934 61950
rect 26998 61886 27276 61950
rect 26928 61880 27276 61886
rect 68952 62560 69164 63044
rect 73848 63038 74060 63044
rect 73848 62974 73854 63038
rect 73918 62974 74060 63038
rect 73848 62902 74060 62974
rect 73848 62838 73990 62902
rect 74054 62838 74060 62902
rect 73848 62832 74060 62838
rect 74256 63038 74468 63044
rect 74256 62974 74398 63038
rect 74462 62974 74468 63038
rect 74256 62902 74468 62974
rect 74256 62838 74398 62902
rect 74462 62838 74468 62902
rect 74256 62832 74468 62838
rect 74664 63038 74876 63044
rect 74664 62974 74806 63038
rect 74870 62974 74876 63038
rect 74664 62908 74876 62974
rect 75072 63038 75284 63044
rect 75072 62974 75214 63038
rect 75278 62974 75284 63038
rect 74664 62832 75012 62908
rect 75072 62832 75284 62974
rect 75480 62832 75692 63180
rect 91936 62908 92148 63044
rect 92616 62908 92828 63044
rect 91936 62902 94188 62908
rect 91936 62838 94118 62902
rect 94182 62838 94188 62902
rect 91936 62832 94188 62838
rect 74664 62772 74740 62832
rect 74936 62772 75012 62832
rect 75480 62772 75556 62832
rect 73848 62630 74060 62636
rect 73848 62566 73990 62630
rect 74054 62566 74060 62630
rect 68952 62500 69028 62560
rect 68952 61950 69164 62500
rect 73848 62424 74060 62566
rect 74256 62630 74468 62636
rect 74256 62566 74398 62630
rect 74462 62566 74468 62630
rect 74256 62424 74468 62566
rect 74664 62424 74876 62772
rect 74936 62696 75284 62772
rect 75072 62500 75284 62696
rect 74974 62494 75284 62500
rect 74936 62430 74942 62494
rect 75006 62430 75284 62494
rect 74974 62424 75284 62430
rect 75480 62424 75692 62772
rect 94112 62630 94324 62636
rect 94112 62566 94118 62630
rect 94182 62566 94324 62630
rect 94112 62560 94324 62566
rect 94112 62504 94176 62560
rect 94232 62504 94324 62560
rect 94112 62500 94324 62504
rect 94112 62494 94732 62500
rect 94112 62430 94662 62494
rect 94726 62430 94732 62494
rect 94112 62424 94732 62430
rect 73984 62364 74060 62424
rect 74392 62364 74468 62424
rect 75616 62364 75692 62424
rect 68952 61886 68958 61950
rect 69022 61886 69164 61950
rect 68952 61880 69164 61886
rect 73848 62016 74060 62364
rect 74256 62016 74468 62364
rect 74664 62222 75012 62228
rect 74664 62158 74942 62222
rect 75006 62158 75012 62222
rect 74664 62152 75012 62158
rect 74664 62016 74876 62152
rect 75072 62016 75284 62228
rect 75480 62222 75692 62364
rect 75480 62158 75622 62222
rect 75686 62158 75692 62222
rect 75480 62152 75692 62158
rect 73848 61956 73924 62016
rect 74256 61956 74332 62016
rect 74800 61956 74876 62016
rect 75208 61956 75284 62016
rect 21760 61548 21836 61608
rect 22168 61548 22244 61608
rect 20400 61542 20612 61548
rect 20400 61478 20406 61542
rect 20470 61478 20612 61542
rect 20400 61406 20612 61478
rect 20400 61342 20542 61406
rect 20606 61342 20612 61406
rect 20400 61336 20612 61342
rect 20808 61542 21020 61548
rect 21118 61542 21564 61548
rect 20808 61478 20950 61542
rect 21014 61478 21020 61542
rect 21080 61478 21086 61542
rect 21150 61478 21564 61542
rect 20808 61200 21020 61478
rect 21118 61472 21564 61478
rect 21216 61200 21564 61472
rect 21624 61406 21836 61548
rect 21624 61342 21630 61406
rect 21694 61342 21836 61406
rect 21624 61336 21836 61342
rect 22032 61406 22244 61548
rect 22032 61342 22038 61406
rect 22102 61342 22244 61406
rect 22032 61336 22244 61342
rect 26928 61678 27276 61684
rect 26928 61614 26934 61678
rect 26998 61614 27276 61678
rect 26928 61542 27276 61614
rect 26928 61478 27206 61542
rect 27270 61478 27276 61542
rect 26928 61336 27276 61478
rect 27200 61276 27276 61336
rect 20808 61140 20884 61200
rect 21488 61140 21564 61200
rect 26928 61270 27276 61276
rect 26928 61206 27206 61270
rect 27270 61206 27276 61270
rect 20400 61134 20612 61140
rect 20400 61070 20542 61134
rect 20606 61070 20612 61134
rect 1768 60880 1980 61004
rect 20400 60998 20612 61070
rect 20400 60934 20406 60998
rect 20470 60934 20612 60998
rect 20400 60928 20612 60934
rect 20808 60928 21020 61140
rect 21216 61004 21564 61140
rect 21118 60998 21564 61004
rect 21080 60934 21086 60998
rect 21150 60934 21358 60998
rect 21422 60934 21564 60998
rect 21118 60928 21564 60934
rect 21624 61134 21836 61140
rect 21624 61070 21630 61134
rect 21694 61070 21836 61134
rect 21624 60998 21836 61070
rect 21624 60934 21630 60998
rect 21694 60934 21836 60998
rect 21624 60928 21836 60934
rect 22032 61134 22244 61140
rect 22032 61070 22038 61134
rect 22102 61070 22244 61134
rect 22032 60998 22244 61070
rect 26928 61064 27276 61206
rect 68952 61678 69164 61684
rect 68952 61614 68958 61678
rect 69022 61614 69164 61678
rect 68952 61336 69164 61614
rect 73848 61608 74060 61956
rect 74256 61608 74468 61956
rect 74664 61814 74876 61956
rect 74664 61750 74670 61814
rect 74734 61750 74876 61814
rect 74664 61744 74876 61750
rect 75072 61814 75284 61956
rect 75072 61750 75078 61814
rect 75142 61750 75284 61814
rect 75072 61744 75284 61750
rect 75480 61950 75692 61956
rect 75480 61886 75622 61950
rect 75686 61886 75692 61950
rect 75480 61814 75692 61886
rect 75480 61750 75486 61814
rect 75550 61750 75692 61814
rect 75480 61744 75692 61750
rect 73984 61548 74060 61608
rect 74392 61548 74468 61608
rect 91936 61678 95412 61684
rect 91936 61614 95342 61678
rect 95406 61614 95412 61678
rect 91936 61608 95412 61614
rect 73848 61406 74060 61548
rect 73848 61342 73990 61406
rect 74054 61342 74060 61406
rect 73848 61336 74060 61342
rect 74256 61406 74468 61548
rect 74256 61342 74262 61406
rect 74326 61342 74468 61406
rect 74256 61336 74468 61342
rect 74664 61542 75284 61548
rect 74664 61478 74670 61542
rect 74734 61478 75078 61542
rect 75142 61478 75284 61542
rect 74664 61472 75284 61478
rect 68952 61276 69028 61336
rect 74664 61276 74876 61472
rect 68952 61064 69164 61276
rect 74664 61200 75012 61276
rect 75072 61200 75284 61472
rect 75480 61542 75692 61548
rect 75480 61478 75486 61542
rect 75550 61478 75692 61542
rect 75480 61406 75692 61478
rect 91936 61542 92148 61608
rect 91936 61478 91942 61542
rect 92006 61478 92148 61542
rect 91936 61472 92148 61478
rect 92616 61472 92828 61608
rect 75480 61342 75622 61406
rect 75686 61342 75692 61406
rect 75480 61336 75692 61342
rect 74664 61140 74740 61200
rect 74936 61140 75012 61200
rect 27064 61004 27140 61064
rect 69088 61004 69164 61064
rect 22032 60934 22038 60998
rect 22102 60934 22244 60998
rect 22032 60928 22244 60934
rect 1768 60868 1818 60880
rect 1224 60862 1818 60868
rect 1224 60798 1230 60862
rect 1294 60824 1818 60862
rect 1874 60824 1980 60880
rect 1294 60798 1980 60824
rect 1224 60792 1980 60798
rect 20400 60726 20612 60732
rect 20400 60662 20406 60726
rect 20470 60662 20612 60726
rect 20400 60590 20612 60662
rect 20400 60526 20542 60590
rect 20606 60526 20612 60590
rect 20400 60520 20612 60526
rect 20808 60726 21156 60732
rect 20808 60662 21086 60726
rect 21150 60662 21156 60726
rect 20808 60656 21156 60662
rect 21216 60726 21564 60732
rect 21216 60662 21358 60726
rect 21422 60662 21564 60726
rect 20808 60596 21020 60656
rect 20808 60590 21156 60596
rect 20808 60526 20950 60590
rect 21014 60526 21086 60590
rect 21150 60526 21156 60590
rect 20808 60520 21156 60526
rect 21216 60520 21564 60662
rect 21624 60726 21836 60732
rect 21624 60662 21630 60726
rect 21694 60662 21836 60726
rect 21624 60590 21836 60662
rect 21624 60526 21766 60590
rect 21830 60526 21836 60590
rect 21624 60520 21836 60526
rect 22032 60726 22244 60732
rect 22032 60662 22038 60726
rect 22102 60662 22244 60726
rect 22032 60590 22244 60662
rect 22032 60526 22038 60590
rect 22102 60526 22244 60590
rect 22032 60520 22244 60526
rect 26928 60520 27276 61004
rect 68952 60520 69164 61004
rect 73848 61134 74060 61140
rect 73848 61070 73990 61134
rect 74054 61070 74060 61134
rect 73848 60998 74060 61070
rect 73848 60934 73990 60998
rect 74054 60934 74060 60998
rect 73848 60928 74060 60934
rect 74256 61134 74468 61140
rect 74256 61070 74262 61134
rect 74326 61070 74468 61134
rect 74256 60998 74468 61070
rect 74256 60934 74262 60998
rect 74326 60934 74468 60998
rect 74256 60928 74468 60934
rect 74664 60928 74876 61140
rect 74936 61064 75284 61140
rect 75072 60998 75284 61064
rect 75072 60934 75078 60998
rect 75142 60934 75284 60998
rect 75072 60928 75284 60934
rect 75480 61134 75692 61140
rect 75480 61070 75622 61134
rect 75686 61070 75692 61134
rect 75480 60998 75692 61070
rect 75480 60934 75622 60998
rect 75686 60934 75692 60998
rect 75480 60928 75692 60934
rect 94112 60880 94324 61004
rect 94112 60862 94176 60880
rect 94232 60868 94324 60880
rect 94232 60862 94732 60868
rect 94112 60798 94118 60862
rect 94232 60824 94662 60862
rect 94182 60798 94662 60824
rect 94726 60798 94732 60862
rect 94112 60792 94732 60798
rect 73848 60726 74060 60732
rect 73848 60662 73990 60726
rect 74054 60662 74060 60726
rect 73848 60590 74060 60662
rect 73848 60526 73990 60590
rect 74054 60526 74060 60590
rect 73848 60520 74060 60526
rect 74256 60726 74468 60732
rect 74256 60662 74262 60726
rect 74326 60662 74468 60726
rect 74256 60590 74468 60662
rect 74256 60526 74398 60590
rect 74462 60526 74468 60590
rect 74256 60520 74468 60526
rect 74664 60590 74876 60732
rect 75072 60726 75284 60732
rect 75072 60662 75078 60726
rect 75142 60662 75284 60726
rect 75072 60596 75284 60662
rect 74974 60590 75284 60596
rect 74664 60526 74670 60590
rect 74734 60526 74876 60590
rect 74936 60526 74942 60590
rect 75006 60526 75284 60590
rect 74664 60520 74876 60526
rect 74974 60520 75284 60526
rect 75480 60726 75692 60732
rect 75480 60662 75622 60726
rect 75686 60662 75692 60726
rect 75480 60590 75692 60662
rect 75480 60526 75486 60590
rect 75550 60526 75692 60590
rect 75480 60520 75692 60526
rect 27064 60460 27140 60520
rect 68952 60460 69028 60520
rect 20400 60318 20612 60324
rect 20400 60254 20542 60318
rect 20606 60254 20612 60318
rect 20400 60182 20612 60254
rect 20400 60118 20542 60182
rect 20606 60118 20612 60182
rect 20400 60112 20612 60118
rect 20808 60318 21020 60324
rect 21118 60318 21564 60324
rect 20808 60254 20950 60318
rect 21014 60254 21020 60318
rect 21080 60254 21086 60318
rect 21150 60254 21564 60318
rect 20808 60112 21020 60254
rect 21118 60248 21564 60254
rect 21216 60182 21564 60248
rect 21216 60118 21358 60182
rect 21422 60118 21564 60182
rect 21216 60112 21564 60118
rect 21624 60318 21836 60324
rect 21624 60254 21766 60318
rect 21830 60254 21836 60318
rect 21624 60182 21836 60254
rect 21624 60118 21630 60182
rect 21694 60118 21836 60182
rect 21624 60112 21836 60118
rect 22032 60318 22244 60324
rect 22032 60254 22038 60318
rect 22102 60254 22244 60318
rect 22032 60182 22244 60254
rect 22032 60118 22174 60182
rect 22238 60118 22244 60182
rect 22032 60112 22244 60118
rect 26928 60248 27276 60460
rect 68952 60248 69164 60460
rect 26928 60188 27004 60248
rect 69088 60188 69164 60248
rect 26928 59976 27276 60188
rect 68952 59976 69164 60188
rect 73848 60318 74060 60324
rect 73848 60254 73990 60318
rect 74054 60254 74060 60318
rect 73848 60182 74060 60254
rect 73848 60118 73854 60182
rect 73918 60118 74060 60182
rect 73848 60112 74060 60118
rect 74256 60318 74468 60324
rect 74256 60254 74398 60318
rect 74462 60254 74468 60318
rect 74256 60182 74468 60254
rect 74256 60118 74262 60182
rect 74326 60118 74468 60182
rect 74256 60112 74468 60118
rect 74664 60318 75012 60324
rect 74664 60254 74670 60318
rect 74734 60254 74942 60318
rect 75006 60254 75012 60318
rect 74664 60248 75012 60254
rect 74664 60188 74876 60248
rect 75072 60188 75284 60324
rect 74664 60182 75284 60188
rect 74664 60118 74806 60182
rect 74870 60118 75284 60182
rect 74664 60112 75284 60118
rect 75480 60318 75692 60324
rect 75480 60254 75486 60318
rect 75550 60254 75692 60318
rect 75480 60182 75692 60254
rect 75480 60118 75622 60182
rect 75686 60118 75692 60182
rect 75480 60112 75692 60118
rect 91936 60318 94188 60324
rect 91936 60254 94118 60318
rect 94182 60254 94188 60318
rect 91936 60248 94188 60254
rect 74800 60052 74876 60112
rect 74800 59976 75148 60052
rect 91936 59976 92148 60248
rect 92616 59976 92828 60248
rect 26928 59916 27004 59976
rect 69088 59916 69164 59976
rect 75072 59916 75148 59976
rect 20400 59910 20612 59916
rect 20400 59846 20542 59910
rect 20606 59846 20612 59910
rect 20400 59774 20612 59846
rect 20400 59710 20542 59774
rect 20606 59710 20612 59774
rect 20400 59704 20612 59710
rect 20808 59774 21020 59916
rect 21216 59910 21564 59916
rect 21216 59846 21358 59910
rect 21422 59846 21564 59910
rect 21216 59780 21564 59846
rect 21118 59774 21564 59780
rect 20808 59710 20814 59774
rect 20878 59710 21020 59774
rect 21080 59710 21086 59774
rect 21150 59710 21494 59774
rect 21558 59710 21564 59774
rect 20808 59704 21020 59710
rect 21118 59704 21564 59710
rect 21624 59910 21836 59916
rect 21624 59846 21630 59910
rect 21694 59846 21836 59910
rect 21624 59774 21836 59846
rect 21624 59710 21630 59774
rect 21694 59710 21836 59774
rect 21624 59704 21836 59710
rect 22032 59910 22244 59916
rect 22032 59846 22174 59910
rect 22238 59846 22244 59910
rect 22032 59774 22244 59846
rect 22032 59710 22038 59774
rect 22102 59710 22244 59774
rect 22032 59704 22244 59710
rect 26928 59704 27276 59916
rect 68952 59704 69164 59916
rect 73848 59910 74060 59916
rect 73848 59846 73854 59910
rect 73918 59846 74060 59910
rect 73848 59774 74060 59846
rect 73848 59710 73854 59774
rect 73918 59710 74060 59774
rect 73848 59704 74060 59710
rect 74256 59910 74468 59916
rect 74256 59846 74262 59910
rect 74326 59846 74468 59910
rect 74256 59774 74468 59846
rect 74256 59710 74398 59774
rect 74462 59710 74468 59774
rect 74256 59704 74468 59710
rect 74664 59910 74876 59916
rect 74664 59846 74806 59910
rect 74870 59846 74876 59910
rect 74664 59774 74876 59846
rect 74664 59710 74670 59774
rect 74734 59710 74876 59774
rect 74664 59704 74876 59710
rect 75072 59704 75284 59916
rect 75480 59910 75692 59916
rect 75480 59846 75622 59910
rect 75686 59846 75692 59910
rect 75480 59774 75692 59846
rect 75480 59710 75622 59774
rect 75686 59710 75692 59774
rect 75480 59704 75692 59710
rect 26928 59644 27004 59704
rect 68952 59644 69028 59704
rect 20400 59502 20612 59508
rect 20400 59438 20542 59502
rect 20606 59438 20612 59502
rect 20400 59296 20612 59438
rect 20808 59502 21156 59508
rect 20808 59438 20814 59502
rect 20878 59438 21086 59502
rect 21150 59438 21156 59502
rect 20808 59432 21156 59438
rect 21216 59502 21564 59508
rect 21216 59438 21494 59502
rect 21558 59438 21564 59502
rect 20808 59372 21020 59432
rect 20808 59366 21156 59372
rect 20808 59302 20950 59366
rect 21014 59302 21086 59366
rect 21150 59302 21156 59366
rect 20808 59296 21156 59302
rect 21216 59296 21564 59438
rect 21624 59502 21836 59508
rect 21624 59438 21630 59502
rect 21694 59438 21836 59502
rect 21624 59366 21836 59438
rect 21624 59302 21630 59366
rect 21694 59302 21836 59366
rect 21624 59296 21836 59302
rect 22032 59502 22244 59508
rect 22032 59438 22038 59502
rect 22102 59438 22244 59502
rect 22032 59366 22244 59438
rect 26928 59432 27276 59644
rect 27200 59372 27276 59432
rect 22032 59302 22038 59366
rect 22102 59302 22244 59366
rect 22032 59296 22244 59302
rect 20536 59236 20612 59296
rect 1224 59230 1980 59236
rect 1224 59166 1230 59230
rect 1294 59200 1980 59230
rect 1294 59166 1818 59200
rect 1224 59160 1818 59166
rect 1768 59144 1818 59160
rect 1874 59144 1980 59200
rect 1768 59024 1980 59144
rect 20400 58888 20612 59236
rect 26928 59160 27276 59372
rect 68952 59432 69164 59644
rect 73848 59502 74060 59508
rect 73848 59438 73854 59502
rect 73918 59438 74060 59502
rect 68952 59372 69028 59432
rect 68952 59160 69164 59372
rect 73848 59366 74060 59438
rect 73848 59302 73854 59366
rect 73918 59302 74060 59366
rect 73848 59296 74060 59302
rect 74256 59502 74468 59508
rect 74256 59438 74398 59502
rect 74462 59438 74468 59502
rect 74256 59366 74468 59438
rect 74256 59302 74398 59366
rect 74462 59302 74468 59366
rect 74256 59296 74468 59302
rect 74664 59502 75284 59508
rect 74664 59438 74670 59502
rect 74734 59438 75284 59502
rect 74664 59432 75284 59438
rect 74664 59296 74876 59432
rect 75072 59366 75284 59432
rect 75072 59302 75078 59366
rect 75142 59302 75284 59366
rect 75072 59296 75284 59302
rect 75480 59502 75692 59508
rect 75480 59438 75622 59502
rect 75686 59438 75692 59502
rect 75480 59296 75692 59438
rect 93424 59427 93490 59428
rect 93382 59363 93425 59427
rect 93489 59363 93532 59427
rect 93424 59362 93490 59363
rect 27064 59100 27140 59160
rect 69088 59100 69164 59160
rect 75480 59236 75556 59296
rect 20808 59094 21020 59100
rect 21118 59094 21564 59100
rect 20808 59030 20950 59094
rect 21014 59030 21020 59094
rect 21080 59030 21086 59094
rect 21150 59030 21564 59094
rect 20808 58888 21020 59030
rect 21118 59024 21564 59030
rect 21216 58888 21564 59024
rect 21624 59094 21836 59100
rect 21624 59030 21630 59094
rect 21694 59030 21836 59094
rect 21624 58958 21836 59030
rect 21624 58894 21630 58958
rect 21694 58894 21836 58958
rect 21624 58888 21836 58894
rect 22032 59094 22244 59100
rect 22032 59030 22038 59094
rect 22102 59030 22244 59094
rect 22032 58958 22244 59030
rect 22032 58894 22174 58958
rect 22238 58894 22244 58958
rect 22032 58888 22244 58894
rect 20400 58828 20476 58888
rect 21488 58828 21564 58888
rect 20400 58480 20612 58828
rect 20808 58692 21020 58828
rect 21216 58692 21564 58828
rect 20808 58616 21564 58692
rect 20808 58556 21020 58616
rect 20808 58550 21156 58556
rect 20808 58486 20814 58550
rect 20878 58486 21086 58550
rect 21150 58486 21156 58550
rect 20808 58480 21156 58486
rect 21216 58480 21564 58616
rect 21624 58686 21836 58692
rect 21624 58622 21630 58686
rect 21694 58622 21836 58686
rect 21624 58550 21836 58622
rect 21624 58486 21766 58550
rect 21830 58486 21836 58550
rect 21624 58480 21836 58486
rect 22032 58686 22244 58692
rect 22032 58622 22174 58686
rect 22238 58622 22244 58686
rect 22032 58550 22244 58622
rect 26928 58616 27276 59100
rect 68952 58616 69164 59100
rect 73848 59094 74060 59100
rect 73848 59030 73854 59094
rect 73918 59030 74060 59094
rect 73848 58958 74060 59030
rect 73848 58894 73854 58958
rect 73918 58894 74060 58958
rect 73848 58888 74060 58894
rect 74256 59094 74468 59100
rect 74256 59030 74398 59094
rect 74462 59030 74468 59094
rect 74256 58958 74468 59030
rect 74256 58894 74262 58958
rect 74326 58894 74468 58958
rect 74256 58888 74468 58894
rect 74664 58888 74876 59100
rect 74800 58828 74876 58888
rect 74664 58692 74876 58828
rect 75072 59094 75284 59100
rect 75072 59030 75078 59094
rect 75142 59030 75284 59094
rect 75072 58888 75284 59030
rect 75480 58888 75692 59236
rect 94112 59200 94324 59236
rect 94112 59144 94176 59200
rect 94232 59144 94324 59200
rect 94112 59100 94324 59144
rect 94112 59094 94732 59100
rect 94112 59030 94662 59094
rect 94726 59030 94732 59094
rect 94112 59024 94732 59030
rect 75072 58828 75148 58888
rect 75616 58828 75692 58888
rect 75072 58692 75284 58828
rect 73848 58686 74060 58692
rect 73848 58622 73854 58686
rect 73918 58622 74060 58686
rect 27064 58556 27140 58616
rect 68952 58556 69028 58616
rect 22032 58486 22174 58550
rect 22238 58486 22244 58550
rect 22032 58480 22244 58486
rect 20400 58420 20476 58480
rect 20400 58278 20612 58420
rect 26928 58414 27276 58556
rect 26928 58350 26934 58414
rect 26998 58350 27276 58414
rect 26928 58344 27276 58350
rect 27200 58284 27276 58344
rect 20400 58214 20406 58278
rect 20470 58214 20612 58278
rect 20400 58208 20612 58214
rect 20808 58278 21020 58284
rect 21118 58278 21564 58284
rect 20808 58214 20814 58278
rect 20878 58214 21020 58278
rect 21080 58214 21086 58278
rect 21150 58214 21564 58278
rect 20808 58148 21020 58214
rect 21118 58208 21564 58214
rect 20808 58072 21156 58148
rect 21216 58072 21564 58208
rect 21624 58278 21836 58284
rect 21624 58214 21766 58278
rect 21830 58214 21836 58278
rect 21624 58072 21836 58214
rect 22032 58278 22244 58284
rect 22032 58214 22174 58278
rect 22238 58214 22244 58278
rect 22032 58072 22244 58214
rect 20944 58012 21020 58072
rect 20400 58006 20612 58012
rect 20400 57942 20406 58006
rect 20470 57942 20612 58006
rect 20400 57870 20612 57942
rect 20400 57806 20542 57870
rect 20606 57806 20612 57870
rect 20400 57800 20612 57806
rect 20808 57870 21020 58012
rect 21080 58012 21156 58072
rect 21760 58012 21836 58072
rect 22168 58012 22244 58072
rect 21080 57936 21564 58012
rect 20808 57806 20814 57870
rect 20878 57806 21020 57870
rect 20808 57800 21020 57806
rect 21216 57800 21564 57936
rect 21624 57664 21836 58012
rect 22032 57664 22244 58012
rect 26928 58142 27276 58284
rect 26928 58078 26934 58142
rect 26998 58078 27206 58142
rect 27270 58078 27276 58142
rect 26928 57936 27276 58078
rect 68952 58414 69164 58556
rect 73848 58550 74060 58622
rect 73848 58486 73990 58550
rect 74054 58486 74060 58550
rect 73848 58480 74060 58486
rect 74256 58686 74468 58692
rect 74256 58622 74262 58686
rect 74326 58622 74468 58686
rect 74256 58550 74468 58622
rect 74256 58486 74398 58550
rect 74462 58486 74468 58550
rect 74256 58480 74468 58486
rect 74664 58616 75284 58692
rect 74664 58550 74876 58616
rect 74664 58486 74670 58550
rect 74734 58486 74876 58550
rect 74664 58480 74876 58486
rect 75072 58480 75284 58616
rect 75480 58480 75692 58828
rect 91936 58822 92148 58828
rect 91936 58758 91942 58822
rect 92006 58758 92148 58822
rect 91936 58692 92148 58758
rect 92616 58692 92828 58828
rect 91936 58616 92828 58692
rect 68952 58350 68958 58414
rect 69022 58350 69164 58414
rect 68952 58344 69164 58350
rect 75480 58420 75556 58480
rect 68952 58284 69028 58344
rect 68952 58142 69164 58284
rect 68952 58078 68958 58142
rect 69022 58078 69164 58142
rect 68952 58006 69164 58078
rect 73848 58278 74060 58284
rect 73848 58214 73990 58278
rect 74054 58214 74060 58278
rect 73848 58072 74060 58214
rect 74256 58278 74468 58284
rect 74256 58214 74398 58278
rect 74462 58214 74468 58278
rect 74256 58072 74468 58214
rect 74664 58278 74876 58284
rect 74664 58214 74670 58278
rect 74734 58214 74876 58278
rect 74664 58072 74876 58214
rect 75072 58148 75284 58284
rect 75480 58278 75692 58420
rect 75480 58214 75622 58278
rect 75686 58214 75692 58278
rect 75480 58208 75692 58214
rect 74974 58142 75284 58148
rect 74936 58078 74942 58142
rect 75006 58078 75284 58142
rect 74974 58072 75284 58078
rect 73984 58012 74060 58072
rect 74392 58012 74468 58072
rect 74800 58012 74876 58072
rect 68952 57942 69094 58006
rect 69158 57942 69164 58006
rect 68952 57936 69164 57942
rect 26928 57734 27276 57740
rect 26928 57670 27206 57734
rect 27270 57670 27276 57734
rect 21624 57604 21700 57664
rect 22032 57604 22108 57664
rect 1768 57520 1980 57604
rect 1768 57468 1818 57520
rect 1224 57464 1818 57468
rect 1874 57464 1980 57520
rect 1224 57462 1980 57464
rect 1224 57398 1230 57462
rect 1294 57398 1980 57462
rect 1224 57392 1980 57398
rect 20400 57598 20612 57604
rect 20400 57534 20542 57598
rect 20606 57534 20612 57598
rect 20400 57462 20612 57534
rect 20400 57398 20542 57462
rect 20606 57398 20612 57462
rect 20400 57392 20612 57398
rect 20808 57598 21020 57604
rect 20808 57534 20814 57598
rect 20878 57534 21020 57598
rect 20808 57332 21020 57534
rect 20808 57256 21156 57332
rect 21216 57256 21564 57604
rect 21624 57256 21836 57604
rect 22032 57256 22244 57604
rect 20944 57196 21020 57256
rect 20400 57190 20612 57196
rect 20400 57126 20542 57190
rect 20606 57126 20612 57190
rect 20400 57054 20612 57126
rect 20400 56990 20542 57054
rect 20606 56990 20612 57054
rect 20400 56984 20612 56990
rect 20808 56984 21020 57196
rect 21080 57196 21156 57256
rect 21352 57196 21428 57256
rect 21760 57196 21836 57256
rect 22168 57196 22244 57256
rect 21080 57120 21564 57196
rect 21216 57054 21564 57120
rect 21216 56990 21494 57054
rect 21558 56990 21564 57054
rect 21216 56984 21564 56990
rect 21624 57054 21836 57196
rect 21624 56990 21630 57054
rect 21694 56990 21836 57054
rect 21624 56984 21836 56990
rect 22032 57054 22244 57196
rect 22032 56990 22174 57054
rect 22238 56990 22244 57054
rect 22032 56984 22244 56990
rect 26928 57120 27276 57670
rect 68952 57734 69164 57740
rect 68952 57670 69094 57734
rect 69158 57670 69164 57734
rect 68952 57120 69164 57670
rect 73848 57664 74060 58012
rect 73984 57604 74060 57664
rect 73848 57256 74060 57604
rect 74256 57664 74468 58012
rect 74664 57936 75284 58012
rect 74664 57876 74876 57936
rect 74664 57870 75012 57876
rect 74664 57806 74942 57870
rect 75006 57806 75012 57870
rect 74664 57800 75012 57806
rect 75072 57870 75284 57936
rect 75072 57806 75214 57870
rect 75278 57806 75284 57870
rect 75072 57800 75284 57806
rect 75480 58006 75692 58012
rect 75480 57942 75622 58006
rect 75686 57942 75692 58006
rect 75480 57870 75692 57942
rect 75480 57806 75622 57870
rect 75686 57806 75692 57870
rect 75480 57800 75692 57806
rect 74256 57604 74332 57664
rect 74256 57256 74468 57604
rect 73984 57196 74060 57256
rect 74392 57196 74468 57256
rect 26928 57060 27004 57120
rect 68952 57060 69028 57120
rect 20400 56782 20612 56788
rect 20400 56718 20542 56782
rect 20606 56718 20612 56782
rect 20400 56646 20612 56718
rect 20400 56582 20406 56646
rect 20470 56582 20612 56646
rect 20400 56576 20612 56582
rect 20808 56646 21020 56788
rect 20808 56582 20950 56646
rect 21014 56582 21020 56646
rect 20808 56576 21020 56582
rect 21216 56782 21564 56788
rect 21216 56718 21494 56782
rect 21558 56718 21564 56782
rect 21216 56576 21564 56718
rect 21624 56782 21836 56788
rect 21624 56718 21630 56782
rect 21694 56718 21836 56782
rect 21624 56646 21836 56718
rect 21624 56582 21630 56646
rect 21694 56582 21836 56646
rect 21624 56576 21836 56582
rect 22032 56782 22244 56788
rect 22032 56718 22174 56782
rect 22238 56718 22244 56782
rect 22032 56646 22244 56718
rect 22032 56582 22038 56646
rect 22102 56582 22244 56646
rect 22032 56576 22244 56582
rect 26928 56782 27276 57060
rect 26928 56718 27206 56782
rect 27270 56718 27276 56782
rect 26928 56576 27276 56718
rect 68952 56576 69164 57060
rect 73848 57054 74060 57196
rect 73848 56990 73854 57054
rect 73918 56990 74060 57054
rect 73848 56984 74060 56990
rect 74256 57054 74468 57196
rect 74256 56990 74262 57054
rect 74326 56990 74468 57054
rect 74256 56984 74468 56990
rect 74664 57256 74876 57604
rect 75072 57598 75284 57604
rect 75072 57534 75214 57598
rect 75278 57534 75284 57598
rect 75072 57256 75284 57534
rect 75480 57598 75692 57604
rect 75480 57534 75622 57598
rect 75686 57534 75692 57598
rect 75480 57462 75692 57534
rect 75480 57398 75486 57462
rect 75550 57398 75692 57462
rect 75480 57392 75692 57398
rect 94112 57520 94324 57604
rect 94112 57464 94176 57520
rect 94232 57468 94324 57520
rect 94232 57464 94732 57468
rect 94112 57462 94732 57464
rect 94112 57398 94662 57462
rect 94726 57398 94732 57462
rect 94112 57392 94732 57398
rect 74664 57196 74740 57256
rect 75072 57196 75148 57256
rect 74664 57054 74876 57196
rect 75072 57060 75284 57196
rect 74974 57054 75284 57060
rect 74664 56990 74806 57054
rect 74870 56990 74876 57054
rect 74936 56990 74942 57054
rect 75006 56990 75284 57054
rect 74664 56984 74876 56990
rect 74974 56984 75284 56990
rect 75480 57190 75692 57196
rect 75480 57126 75486 57190
rect 75550 57126 75692 57190
rect 75480 57054 75692 57126
rect 75480 56990 75486 57054
rect 75550 56990 75692 57054
rect 75480 56984 75692 56990
rect 73848 56782 74060 56788
rect 73848 56718 73854 56782
rect 73918 56718 74060 56782
rect 73848 56646 74060 56718
rect 73848 56582 73854 56646
rect 73918 56582 74060 56646
rect 73848 56576 74060 56582
rect 74256 56782 74468 56788
rect 74256 56718 74262 56782
rect 74326 56718 74468 56782
rect 74256 56646 74468 56718
rect 74256 56582 74398 56646
rect 74462 56582 74468 56646
rect 74256 56576 74468 56582
rect 74664 56782 75012 56788
rect 74664 56718 74806 56782
rect 74870 56718 74942 56782
rect 75006 56718 75012 56782
rect 74664 56712 75012 56718
rect 74664 56652 74876 56712
rect 75072 56652 75284 56788
rect 74664 56646 75284 56652
rect 74664 56582 75214 56646
rect 75278 56582 75284 56646
rect 74664 56576 75284 56582
rect 75480 56782 75692 56788
rect 75480 56718 75486 56782
rect 75550 56718 75692 56782
rect 75480 56646 75692 56718
rect 75480 56582 75622 56646
rect 75686 56582 75692 56646
rect 75480 56576 75692 56582
rect 21216 56516 21292 56576
rect 20944 56440 21292 56516
rect 26928 56516 27004 56576
rect 69088 56516 69164 56576
rect 26928 56510 27276 56516
rect 26928 56446 27206 56510
rect 27270 56446 27276 56510
rect 20944 56380 21020 56440
rect 20400 56374 20612 56380
rect 20400 56310 20406 56374
rect 20470 56310 20612 56374
rect 20400 56238 20612 56310
rect 20400 56174 20406 56238
rect 20470 56174 20612 56238
rect 20400 56168 20612 56174
rect 20808 56374 21564 56380
rect 20808 56310 20950 56374
rect 21014 56310 21564 56374
rect 20808 56304 21564 56310
rect 20808 56244 21020 56304
rect 20808 56238 21156 56244
rect 20808 56174 20950 56238
rect 21014 56174 21086 56238
rect 21150 56174 21156 56238
rect 20808 56168 21156 56174
rect 21216 56168 21564 56304
rect 21624 56374 21836 56380
rect 21624 56310 21630 56374
rect 21694 56310 21836 56374
rect 21624 56238 21836 56310
rect 21624 56174 21766 56238
rect 21830 56174 21836 56238
rect 21624 56168 21836 56174
rect 22032 56374 22244 56380
rect 22032 56310 22038 56374
rect 22102 56310 22244 56374
rect 22032 56238 22244 56310
rect 26928 56304 27276 56446
rect 68952 56304 69164 56516
rect 73848 56374 74060 56380
rect 73848 56310 73854 56374
rect 73918 56310 74060 56374
rect 27064 56244 27140 56304
rect 68952 56244 69028 56304
rect 22032 56174 22038 56238
rect 22102 56174 22244 56238
rect 22032 56168 22244 56174
rect 26928 56032 27276 56244
rect 68952 56032 69164 56244
rect 73848 56238 74060 56310
rect 73848 56174 73990 56238
rect 74054 56174 74060 56238
rect 73848 56168 74060 56174
rect 74256 56374 74468 56380
rect 74256 56310 74398 56374
rect 74462 56310 74468 56374
rect 74256 56238 74468 56310
rect 74256 56174 74398 56238
rect 74462 56174 74468 56238
rect 74256 56168 74468 56174
rect 74664 56238 74876 56380
rect 74664 56174 74670 56238
rect 74734 56174 74876 56238
rect 74664 56168 74876 56174
rect 75072 56374 75284 56380
rect 75072 56310 75214 56374
rect 75278 56310 75284 56374
rect 75072 56238 75284 56310
rect 75072 56174 75078 56238
rect 75142 56174 75284 56238
rect 75072 56168 75284 56174
rect 75480 56374 75692 56380
rect 75480 56310 75622 56374
rect 75686 56310 75692 56374
rect 75480 56238 75692 56310
rect 75480 56174 75486 56238
rect 75550 56174 75692 56238
rect 75480 56168 75692 56174
rect 27064 55972 27140 56032
rect 68952 55972 69028 56032
rect 1224 55966 1980 55972
rect 1224 55902 1230 55966
rect 1294 55902 1980 55966
rect 1224 55896 1980 55902
rect 1768 55840 1980 55896
rect 1768 55784 1818 55840
rect 1874 55784 1980 55840
rect 1768 55760 1980 55784
rect 20400 55966 20612 55972
rect 20400 55902 20406 55966
rect 20470 55902 20612 55966
rect 20400 55830 20612 55902
rect 20400 55766 20406 55830
rect 20470 55766 20612 55830
rect 20400 55760 20612 55766
rect 20808 55966 21020 55972
rect 21118 55966 21564 55972
rect 20808 55902 20950 55966
rect 21014 55902 21020 55966
rect 21080 55902 21086 55966
rect 21150 55902 21564 55966
rect 20808 55830 21020 55902
rect 21118 55896 21564 55902
rect 20808 55766 20814 55830
rect 20878 55766 21020 55830
rect 20808 55760 21020 55766
rect 21216 55760 21564 55896
rect 21624 55966 21836 55972
rect 21624 55902 21766 55966
rect 21830 55902 21836 55966
rect 21624 55830 21836 55902
rect 21624 55766 21630 55830
rect 21694 55766 21836 55830
rect 21624 55760 21836 55766
rect 22032 55966 22244 55972
rect 22032 55902 22038 55966
rect 22102 55902 22244 55966
rect 22032 55830 22244 55902
rect 22032 55766 22038 55830
rect 22102 55766 22244 55830
rect 22032 55760 22244 55766
rect 26928 55760 27276 55972
rect 68952 55760 69164 55972
rect 73848 55966 74060 55972
rect 73848 55902 73990 55966
rect 74054 55902 74060 55966
rect 73848 55830 74060 55902
rect 73848 55766 73854 55830
rect 73918 55766 74060 55830
rect 73848 55760 74060 55766
rect 74256 55966 74468 55972
rect 74256 55902 74398 55966
rect 74462 55902 74468 55966
rect 74256 55830 74468 55902
rect 74256 55766 74262 55830
rect 74326 55766 74468 55830
rect 74256 55760 74468 55766
rect 74664 55966 74876 55972
rect 74664 55902 74670 55966
rect 74734 55902 74876 55966
rect 74664 55836 74876 55902
rect 75072 55966 75284 55972
rect 75072 55902 75078 55966
rect 75142 55902 75284 55966
rect 75072 55836 75284 55902
rect 74664 55760 75284 55836
rect 75480 55966 75692 55972
rect 75480 55902 75486 55966
rect 75550 55902 75692 55966
rect 75480 55830 75692 55902
rect 75480 55766 75622 55830
rect 75686 55766 75692 55830
rect 75480 55760 75692 55766
rect 94112 55966 94732 55972
rect 94112 55902 94662 55966
rect 94726 55902 94732 55966
rect 94112 55896 94732 55902
rect 94112 55840 94324 55896
rect 94112 55784 94176 55840
rect 94232 55784 94324 55840
rect 94112 55760 94324 55784
rect 26928 55700 27004 55760
rect 69088 55700 69164 55760
rect 75072 55700 75148 55760
rect 20400 55558 20612 55564
rect 20400 55494 20406 55558
rect 20470 55494 20612 55558
rect 20400 55352 20612 55494
rect 20808 55558 21020 55564
rect 20808 55494 20814 55558
rect 20878 55494 21020 55558
rect 20808 55422 21020 55494
rect 21216 55428 21564 55564
rect 21118 55422 21564 55428
rect 20808 55358 20814 55422
rect 20878 55358 21020 55422
rect 21080 55358 21086 55422
rect 21150 55358 21494 55422
rect 21558 55358 21564 55422
rect 20808 55352 21020 55358
rect 21118 55352 21564 55358
rect 21624 55558 21836 55564
rect 21624 55494 21630 55558
rect 21694 55494 21836 55558
rect 21624 55422 21836 55494
rect 21624 55358 21630 55422
rect 21694 55358 21836 55422
rect 21624 55352 21836 55358
rect 22032 55558 22244 55564
rect 22032 55494 22038 55558
rect 22102 55494 22244 55558
rect 22032 55422 22244 55494
rect 26928 55488 27276 55700
rect 68952 55488 69164 55700
rect 74800 55624 75148 55700
rect 74800 55564 74876 55624
rect 27064 55428 27140 55488
rect 69088 55428 69164 55488
rect 22032 55358 22174 55422
rect 22238 55358 22244 55422
rect 22032 55352 22244 55358
rect 20536 55292 20612 55352
rect 20400 55014 20612 55292
rect 26928 55216 27276 55428
rect 27200 55156 27276 55216
rect 20400 54950 20406 55014
rect 20470 54950 20612 55014
rect 20400 54944 20612 54950
rect 20808 55150 21156 55156
rect 20808 55086 20814 55150
rect 20878 55086 21086 55150
rect 21150 55086 21156 55150
rect 20808 55080 21156 55086
rect 21216 55150 21564 55156
rect 21216 55086 21494 55150
rect 21558 55086 21564 55150
rect 20808 55020 21020 55080
rect 20808 55014 21156 55020
rect 20808 54950 20950 55014
rect 21014 54950 21086 55014
rect 21150 54950 21156 55014
rect 20808 54944 21156 54950
rect 21216 54944 21564 55086
rect 21624 55150 21836 55156
rect 21624 55086 21630 55150
rect 21694 55086 21836 55150
rect 21624 55014 21836 55086
rect 21624 54950 21630 55014
rect 21694 54950 21836 55014
rect 21624 54944 21836 54950
rect 22032 55150 22244 55156
rect 22032 55086 22174 55150
rect 22238 55086 22244 55150
rect 22032 55014 22244 55086
rect 22032 54950 22038 55014
rect 22102 54950 22244 55014
rect 22032 54944 22244 54950
rect 26928 54944 27276 55156
rect 27200 54884 27276 54944
rect 20400 54742 20612 54748
rect 20400 54678 20406 54742
rect 20470 54678 20612 54742
rect 20400 54536 20612 54678
rect 20808 54742 21020 54748
rect 21118 54742 21564 54748
rect 20808 54678 20950 54742
rect 21014 54678 21020 54742
rect 21080 54678 21086 54742
rect 21150 54678 21564 54742
rect 20808 54536 21020 54678
rect 21118 54672 21564 54678
rect 21216 54606 21564 54672
rect 21216 54542 21494 54606
rect 21558 54542 21564 54606
rect 21216 54536 21564 54542
rect 21624 54742 21836 54748
rect 21624 54678 21630 54742
rect 21694 54678 21836 54742
rect 21624 54606 21836 54678
rect 21624 54542 21630 54606
rect 21694 54542 21836 54606
rect 21624 54536 21836 54542
rect 22032 54742 22244 54748
rect 22032 54678 22038 54742
rect 22102 54678 22244 54742
rect 22032 54606 22244 54678
rect 26928 54672 27276 54884
rect 68952 55216 69164 55428
rect 73848 55558 74060 55564
rect 73848 55494 73854 55558
rect 73918 55494 74060 55558
rect 73848 55422 74060 55494
rect 73848 55358 73990 55422
rect 74054 55358 74060 55422
rect 73848 55352 74060 55358
rect 74256 55558 74468 55564
rect 74256 55494 74262 55558
rect 74326 55494 74468 55558
rect 74256 55422 74468 55494
rect 74256 55358 74398 55422
rect 74462 55358 74468 55422
rect 74256 55352 74468 55358
rect 74664 55488 75284 55564
rect 74664 55352 74876 55488
rect 75072 55422 75284 55488
rect 75072 55358 75214 55422
rect 75278 55358 75284 55422
rect 75072 55352 75284 55358
rect 75480 55558 75692 55564
rect 75480 55494 75622 55558
rect 75686 55494 75692 55558
rect 75480 55352 75692 55494
rect 75616 55292 75692 55352
rect 68952 55156 69028 55216
rect 68952 54944 69164 55156
rect 73848 55150 74060 55156
rect 73848 55086 73990 55150
rect 74054 55086 74060 55150
rect 73848 55014 74060 55086
rect 73848 54950 73854 55014
rect 73918 54950 74060 55014
rect 73848 54944 74060 54950
rect 74256 55150 74468 55156
rect 74256 55086 74398 55150
rect 74462 55086 74468 55150
rect 74256 55014 74468 55086
rect 74256 54950 74262 55014
rect 74326 54950 74468 55014
rect 74256 54944 74468 54950
rect 74664 55014 74876 55156
rect 74664 54950 74670 55014
rect 74734 54950 74876 55014
rect 74664 54944 74876 54950
rect 75072 55150 75284 55156
rect 75072 55086 75214 55150
rect 75278 55086 75284 55150
rect 75072 54944 75284 55086
rect 75480 55014 75692 55292
rect 75480 54950 75622 55014
rect 75686 54950 75692 55014
rect 75480 54944 75692 54950
rect 68952 54884 69028 54944
rect 75072 54884 75148 54944
rect 68952 54672 69164 54884
rect 74800 54808 75148 54884
rect 74800 54748 74876 54808
rect 27200 54612 27276 54672
rect 69088 54612 69164 54672
rect 22032 54542 22038 54606
rect 22102 54542 22244 54606
rect 22032 54536 22244 54542
rect 20536 54476 20612 54536
rect 20400 54334 20612 54476
rect 26928 54400 27276 54612
rect 68952 54400 69164 54612
rect 73848 54742 74060 54748
rect 73848 54678 73854 54742
rect 73918 54678 74060 54742
rect 73848 54606 74060 54678
rect 73848 54542 73854 54606
rect 73918 54542 74060 54606
rect 73848 54536 74060 54542
rect 74256 54742 74468 54748
rect 74256 54678 74262 54742
rect 74326 54678 74468 54742
rect 74256 54606 74468 54678
rect 74256 54542 74262 54606
rect 74326 54542 74468 54606
rect 74256 54536 74468 54542
rect 74664 54742 75284 54748
rect 74664 54678 74670 54742
rect 74734 54678 75284 54742
rect 74664 54672 75284 54678
rect 74664 54536 74876 54672
rect 75072 54606 75284 54672
rect 75072 54542 75214 54606
rect 75278 54542 75284 54606
rect 75072 54536 75284 54542
rect 75480 54742 75692 54748
rect 75480 54678 75622 54742
rect 75686 54678 75692 54742
rect 75480 54536 75692 54678
rect 75616 54476 75692 54536
rect 27200 54340 27276 54400
rect 69088 54340 69164 54400
rect 20400 54270 20406 54334
rect 20470 54270 20612 54334
rect 20400 54264 20612 54270
rect 1768 54160 1980 54204
rect 1768 54104 1818 54160
rect 1874 54104 1980 54160
rect 20808 54128 21020 54340
rect 21216 54334 21564 54340
rect 21216 54270 21494 54334
rect 21558 54270 21564 54334
rect 21216 54128 21564 54270
rect 21624 54334 21836 54340
rect 21624 54270 21630 54334
rect 21694 54270 21836 54334
rect 21624 54128 21836 54270
rect 22032 54334 22244 54340
rect 22032 54270 22038 54334
rect 22102 54270 22244 54334
rect 22032 54128 22244 54270
rect 1768 54068 1980 54104
rect 20944 54068 21020 54128
rect 21352 54068 21428 54128
rect 21760 54068 21836 54128
rect 22168 54068 22244 54128
rect 1224 54062 1980 54068
rect 1224 53998 1230 54062
rect 1294 53998 1980 54062
rect 1224 53992 1980 53998
rect 20400 54062 20612 54068
rect 20400 53998 20406 54062
rect 20470 53998 20612 54062
rect 20400 53926 20612 53998
rect 20400 53862 20542 53926
rect 20606 53862 20612 53926
rect 20400 53856 20612 53862
rect 20808 53992 21564 54068
rect 20808 53856 21020 53992
rect 21216 53926 21564 53992
rect 21216 53862 21494 53926
rect 21558 53862 21564 53926
rect 21216 53856 21564 53862
rect 21624 53720 21836 54068
rect 21760 53660 21836 53720
rect 20400 53654 20612 53660
rect 20400 53590 20542 53654
rect 20606 53590 20612 53654
rect 20400 53518 20612 53590
rect 20400 53454 20542 53518
rect 20606 53454 20612 53518
rect 20400 53448 20612 53454
rect 20808 53312 21020 53660
rect 21216 53654 21564 53660
rect 21216 53590 21494 53654
rect 21558 53590 21564 53654
rect 21216 53388 21564 53590
rect 21080 53312 21564 53388
rect 21624 53312 21836 53660
rect 22032 53720 22244 54068
rect 26928 54062 27276 54340
rect 26928 53998 27070 54062
rect 27134 53998 27206 54062
rect 27270 53998 27276 54062
rect 26928 53992 27276 53998
rect 68952 54062 69164 54340
rect 73848 54334 74060 54340
rect 73848 54270 73854 54334
rect 73918 54270 74060 54334
rect 73848 54128 74060 54270
rect 74256 54334 74468 54340
rect 74256 54270 74262 54334
rect 74326 54270 74468 54334
rect 74256 54128 74468 54270
rect 73984 54068 74060 54128
rect 74392 54068 74468 54128
rect 68952 53998 68958 54062
rect 69022 53998 69164 54062
rect 68952 53992 69164 53998
rect 26928 53790 27276 53796
rect 26928 53726 27206 53790
rect 27270 53726 27276 53790
rect 22032 53660 22108 53720
rect 22032 53312 22244 53660
rect 20808 53252 20884 53312
rect 21080 53252 21156 53312
rect 21760 53252 21836 53312
rect 22168 53252 22244 53312
rect 20400 53246 20612 53252
rect 20400 53182 20542 53246
rect 20606 53182 20612 53246
rect 20400 53110 20612 53182
rect 20400 53046 20406 53110
rect 20470 53046 20612 53110
rect 20400 53040 20612 53046
rect 20808 53176 21156 53252
rect 20808 53110 21020 53176
rect 21216 53116 21564 53252
rect 21118 53110 21564 53116
rect 20808 53046 20950 53110
rect 21014 53046 21020 53110
rect 21080 53046 21086 53110
rect 21150 53046 21564 53110
rect 20808 53040 21020 53046
rect 21118 53040 21564 53046
rect 21624 53110 21836 53252
rect 21624 53046 21766 53110
rect 21830 53046 21836 53110
rect 21624 53040 21836 53046
rect 22032 53110 22244 53252
rect 22032 53046 22038 53110
rect 22102 53046 22244 53110
rect 22032 53040 22244 53046
rect 26928 53654 27276 53726
rect 26928 53590 26934 53654
rect 26998 53590 27070 53654
rect 27134 53590 27276 53654
rect 26928 53382 27276 53590
rect 26928 53318 26934 53382
rect 26998 53318 27276 53382
rect 26928 53176 27276 53318
rect 68952 53790 69164 53796
rect 68952 53726 68958 53790
rect 69022 53726 69164 53790
rect 68952 53654 69164 53726
rect 73848 53720 74060 54068
rect 74256 53720 74468 54068
rect 74664 54128 74876 54340
rect 75072 54334 75284 54340
rect 75072 54270 75214 54334
rect 75278 54270 75284 54334
rect 75072 54128 75284 54270
rect 75480 54334 75692 54476
rect 75480 54270 75486 54334
rect 75550 54270 75692 54334
rect 75480 54264 75692 54270
rect 94112 54160 94324 54204
rect 74664 54068 74740 54128
rect 75072 54068 75148 54128
rect 94112 54104 94176 54160
rect 94232 54104 94324 54160
rect 94112 54068 94324 54104
rect 74664 53926 74876 54068
rect 74664 53862 74670 53926
rect 74734 53862 74876 53926
rect 74664 53856 74876 53862
rect 75072 53926 75284 54068
rect 75072 53862 75078 53926
rect 75142 53862 75284 53926
rect 75072 53856 75284 53862
rect 75480 54062 75692 54068
rect 75480 53998 75486 54062
rect 75550 53998 75692 54062
rect 75480 53926 75692 53998
rect 94112 54062 94732 54068
rect 94112 53998 94662 54062
rect 94726 53998 94732 54062
rect 94112 53992 94732 53998
rect 75480 53862 75486 53926
rect 75550 53862 75692 53926
rect 75480 53856 75692 53862
rect 73984 53660 74060 53720
rect 74392 53660 74468 53720
rect 68952 53590 69094 53654
rect 69158 53590 69164 53654
rect 68952 53382 69164 53590
rect 68952 53318 69094 53382
rect 69158 53318 69164 53382
rect 68952 53176 69164 53318
rect 73848 53312 74060 53660
rect 73984 53252 74060 53312
rect 26928 53116 27004 53176
rect 69088 53116 69164 53176
rect 20400 52838 20612 52844
rect 20400 52774 20406 52838
rect 20470 52774 20612 52838
rect 20400 52702 20612 52774
rect 20400 52638 20542 52702
rect 20606 52638 20612 52702
rect 20400 52632 20612 52638
rect 20808 52838 21156 52844
rect 20808 52774 20950 52838
rect 21014 52774 21086 52838
rect 21150 52774 21156 52838
rect 20808 52768 21156 52774
rect 20808 52708 21020 52768
rect 21216 52708 21564 52844
rect 20808 52632 21564 52708
rect 21624 52838 21836 52844
rect 21624 52774 21766 52838
rect 21830 52774 21836 52838
rect 21624 52702 21836 52774
rect 21624 52638 21630 52702
rect 21694 52638 21836 52702
rect 21624 52632 21836 52638
rect 22032 52838 22244 52844
rect 22032 52774 22038 52838
rect 22102 52774 22244 52838
rect 22032 52702 22244 52774
rect 22032 52638 22038 52702
rect 22102 52638 22244 52702
rect 22032 52632 22244 52638
rect 26928 52838 27276 53116
rect 26928 52774 27206 52838
rect 27270 52774 27276 52838
rect 26928 52632 27276 52774
rect 68952 52838 69164 53116
rect 73848 53110 74060 53252
rect 73848 53046 73990 53110
rect 74054 53046 74060 53110
rect 73848 53040 74060 53046
rect 74256 53312 74468 53660
rect 74664 53654 74876 53660
rect 74664 53590 74670 53654
rect 74734 53590 74876 53654
rect 74664 53524 74876 53590
rect 75072 53654 75284 53660
rect 75072 53590 75078 53654
rect 75142 53590 75284 53654
rect 74664 53518 75012 53524
rect 74664 53454 74942 53518
rect 75006 53454 75012 53518
rect 74664 53448 75012 53454
rect 74664 53388 74876 53448
rect 75072 53388 75284 53590
rect 75480 53654 75692 53660
rect 75480 53590 75486 53654
rect 75550 53590 75692 53654
rect 75480 53518 75692 53590
rect 75480 53454 75622 53518
rect 75686 53454 75692 53518
rect 75480 53448 75692 53454
rect 74664 53312 75284 53388
rect 74256 53252 74332 53312
rect 74800 53252 74876 53312
rect 74256 53110 74468 53252
rect 74256 53046 74262 53110
rect 74326 53046 74468 53110
rect 74256 53040 74468 53046
rect 74664 53110 74876 53252
rect 74974 53246 75284 53252
rect 74936 53182 74942 53246
rect 75006 53182 75284 53246
rect 74974 53176 75284 53182
rect 74664 53046 74670 53110
rect 74734 53046 74876 53110
rect 74664 53040 74876 53046
rect 75072 53040 75284 53176
rect 75480 53246 75692 53252
rect 75480 53182 75622 53246
rect 75686 53182 75692 53246
rect 75480 53110 75692 53182
rect 75480 53046 75486 53110
rect 75550 53046 75692 53110
rect 75480 53040 75692 53046
rect 68952 52774 69094 52838
rect 69158 52774 69164 52838
rect 68952 52632 69164 52774
rect 73848 52838 74060 52844
rect 73848 52774 73990 52838
rect 74054 52774 74060 52838
rect 73848 52702 74060 52774
rect 73848 52638 73854 52702
rect 73918 52638 74060 52702
rect 73848 52632 74060 52638
rect 74256 52838 74468 52844
rect 74256 52774 74262 52838
rect 74326 52774 74468 52838
rect 74256 52702 74468 52774
rect 74256 52638 74398 52702
rect 74462 52638 74468 52702
rect 74256 52632 74468 52638
rect 74664 52838 74876 52844
rect 74664 52774 74670 52838
rect 74734 52774 74876 52838
rect 74664 52702 74876 52774
rect 74664 52638 74806 52702
rect 74870 52638 74876 52702
rect 74664 52632 74876 52638
rect 75072 52632 75284 52844
rect 75480 52838 75692 52844
rect 75480 52774 75486 52838
rect 75550 52774 75692 52838
rect 75480 52702 75692 52774
rect 75480 52638 75486 52702
rect 75550 52638 75692 52702
rect 75480 52632 75692 52638
rect 21216 52572 21292 52632
rect 27200 52572 27276 52632
rect 69088 52572 69164 52632
rect 75072 52572 75148 52632
rect 1768 52480 1980 52572
rect 1768 52436 1818 52480
rect 1224 52430 1818 52436
rect 1224 52366 1230 52430
rect 1294 52424 1818 52430
rect 1874 52424 1980 52480
rect 21080 52496 21292 52572
rect 26928 52566 27276 52572
rect 26928 52502 27206 52566
rect 27270 52502 27276 52566
rect 21080 52436 21156 52496
rect 1294 52366 1980 52424
rect 1224 52360 1980 52366
rect 20400 52430 20612 52436
rect 20400 52366 20542 52430
rect 20606 52366 20612 52430
rect 20400 52294 20612 52366
rect 20400 52230 20542 52294
rect 20606 52230 20612 52294
rect 20400 52224 20612 52230
rect 20808 52360 21156 52436
rect 20808 52294 21020 52360
rect 21216 52300 21564 52436
rect 21118 52294 21564 52300
rect 20808 52230 20950 52294
rect 21014 52230 21020 52294
rect 21080 52230 21086 52294
rect 21150 52230 21222 52294
rect 21286 52230 21564 52294
rect 20808 52224 21020 52230
rect 21118 52224 21564 52230
rect 21624 52430 21836 52436
rect 21624 52366 21630 52430
rect 21694 52366 21836 52430
rect 21624 52294 21836 52366
rect 21624 52230 21630 52294
rect 21694 52230 21836 52294
rect 21624 52224 21836 52230
rect 22032 52430 22244 52436
rect 22032 52366 22038 52430
rect 22102 52366 22244 52430
rect 22032 52294 22244 52366
rect 22032 52230 22038 52294
rect 22102 52230 22244 52294
rect 22032 52224 22244 52230
rect 26928 52360 27276 52502
rect 68952 52566 69164 52572
rect 68952 52502 69094 52566
rect 69158 52502 69164 52566
rect 68952 52360 69164 52502
rect 74800 52496 75148 52572
rect 74800 52436 74876 52496
rect 94112 52480 94324 52572
rect 26928 52300 27004 52360
rect 69088 52300 69164 52360
rect 26928 52088 27276 52300
rect 27200 52028 27276 52088
rect 20400 52022 20612 52028
rect 20400 51958 20542 52022
rect 20606 51958 20612 52022
rect 20400 51886 20612 51958
rect 20400 51822 20542 51886
rect 20606 51822 20612 51886
rect 20400 51816 20612 51822
rect 20808 52022 21156 52028
rect 20808 51958 20950 52022
rect 21014 51958 21086 52022
rect 21150 51958 21156 52022
rect 20808 51952 21156 51958
rect 21216 52022 21564 52028
rect 21216 51958 21222 52022
rect 21286 51958 21564 52022
rect 20808 51816 21020 51952
rect 21216 51886 21564 51958
rect 21216 51822 21494 51886
rect 21558 51822 21564 51886
rect 21216 51816 21564 51822
rect 21624 52022 21836 52028
rect 21624 51958 21630 52022
rect 21694 51958 21836 52022
rect 21624 51886 21836 51958
rect 21624 51822 21766 51886
rect 21830 51822 21836 51886
rect 21624 51816 21836 51822
rect 22032 52022 22244 52028
rect 22032 51958 22038 52022
rect 22102 51958 22244 52022
rect 22032 51886 22244 51958
rect 22032 51822 22174 51886
rect 22238 51822 22244 51886
rect 22032 51816 22244 51822
rect 26928 51816 27276 52028
rect 27200 51756 27276 51816
rect 20400 51614 20612 51620
rect 20400 51550 20542 51614
rect 20606 51550 20612 51614
rect 20400 51408 20612 51550
rect 20808 51478 21020 51620
rect 20808 51414 20814 51478
rect 20878 51414 21020 51478
rect 20808 51408 21020 51414
rect 21216 51614 21564 51620
rect 21216 51550 21494 51614
rect 21558 51550 21564 51614
rect 21216 51478 21564 51550
rect 21216 51414 21358 51478
rect 21422 51414 21564 51478
rect 21216 51408 21564 51414
rect 21624 51614 21836 51620
rect 21624 51550 21766 51614
rect 21830 51550 21836 51614
rect 21624 51478 21836 51550
rect 21624 51414 21630 51478
rect 21694 51414 21836 51478
rect 21624 51408 21836 51414
rect 22032 51614 22244 51620
rect 22032 51550 22174 51614
rect 22238 51550 22244 51614
rect 22032 51478 22244 51550
rect 26928 51544 27276 51756
rect 68952 52088 69164 52300
rect 73848 52430 74060 52436
rect 73848 52366 73854 52430
rect 73918 52366 74060 52430
rect 73848 52294 74060 52366
rect 73848 52230 73990 52294
rect 74054 52230 74060 52294
rect 73848 52224 74060 52230
rect 74256 52430 74468 52436
rect 74256 52366 74398 52430
rect 74462 52366 74468 52430
rect 74256 52294 74468 52366
rect 74256 52230 74262 52294
rect 74326 52230 74468 52294
rect 74256 52224 74468 52230
rect 74664 52430 75284 52436
rect 74664 52366 74806 52430
rect 74870 52366 75284 52430
rect 74664 52360 75284 52366
rect 74664 52294 74876 52360
rect 74664 52230 74670 52294
rect 74734 52230 74876 52294
rect 74664 52224 74876 52230
rect 75072 52224 75284 52360
rect 75480 52430 75692 52436
rect 75480 52366 75486 52430
rect 75550 52366 75692 52430
rect 75480 52294 75692 52366
rect 94112 52424 94176 52480
rect 94232 52436 94324 52480
rect 94232 52430 94732 52436
rect 94232 52424 94662 52430
rect 94112 52366 94662 52424
rect 94726 52366 94732 52430
rect 94112 52360 94732 52366
rect 75480 52230 75486 52294
rect 75550 52230 75692 52294
rect 75480 52224 75692 52230
rect 68952 52028 69028 52088
rect 68952 51816 69164 52028
rect 73848 52022 74060 52028
rect 73848 51958 73990 52022
rect 74054 51958 74060 52022
rect 73848 51886 74060 51958
rect 73848 51822 73990 51886
rect 74054 51822 74060 51886
rect 73848 51816 74060 51822
rect 74256 52022 74468 52028
rect 74256 51958 74262 52022
rect 74326 51958 74468 52022
rect 74256 51886 74468 51958
rect 74256 51822 74398 51886
rect 74462 51822 74468 51886
rect 74256 51816 74468 51822
rect 74664 52022 75284 52028
rect 74664 51958 74670 52022
rect 74734 51958 75284 52022
rect 74664 51952 75284 51958
rect 74664 51892 74876 51952
rect 74664 51886 75012 51892
rect 74664 51822 74942 51886
rect 75006 51822 75012 51886
rect 74664 51816 75012 51822
rect 75072 51816 75284 51952
rect 75480 52022 75692 52028
rect 75480 51958 75486 52022
rect 75550 51958 75692 52022
rect 75480 51886 75692 51958
rect 75480 51822 75486 51886
rect 75550 51822 75692 51886
rect 75480 51816 75692 51822
rect 68952 51756 69028 51816
rect 68952 51544 69164 51756
rect 27064 51484 27140 51544
rect 69088 51484 69164 51544
rect 22032 51414 22038 51478
rect 22102 51414 22244 51478
rect 22032 51408 22244 51414
rect 20400 51348 20476 51408
rect 20400 51070 20612 51348
rect 26928 51272 27276 51484
rect 68952 51272 69164 51484
rect 73848 51614 74060 51620
rect 73848 51550 73990 51614
rect 74054 51550 74060 51614
rect 73848 51478 74060 51550
rect 73848 51414 73854 51478
rect 73918 51414 74060 51478
rect 73848 51408 74060 51414
rect 74256 51614 74468 51620
rect 74256 51550 74398 51614
rect 74462 51550 74468 51614
rect 74256 51478 74468 51550
rect 74256 51414 74398 51478
rect 74462 51414 74468 51478
rect 74256 51408 74468 51414
rect 74664 51478 74876 51620
rect 74974 51614 75284 51620
rect 74936 51550 74942 51614
rect 75006 51550 75284 51614
rect 74974 51544 75284 51550
rect 74664 51414 74806 51478
rect 74870 51414 74876 51478
rect 74664 51408 74876 51414
rect 75072 51408 75284 51544
rect 75480 51614 75692 51620
rect 75480 51550 75486 51614
rect 75550 51550 75692 51614
rect 75480 51408 75692 51550
rect 75072 51348 75148 51408
rect 75616 51348 75692 51408
rect 27064 51212 27140 51272
rect 69088 51212 69164 51272
rect 74800 51272 75148 51348
rect 74800 51212 74876 51272
rect 20400 51006 20406 51070
rect 20470 51006 20612 51070
rect 20400 51000 20612 51006
rect 20808 51206 21020 51212
rect 20808 51142 20814 51206
rect 20878 51142 21020 51206
rect 20808 51070 21020 51142
rect 21216 51206 21564 51212
rect 21216 51142 21358 51206
rect 21422 51142 21564 51206
rect 21216 51076 21564 51142
rect 21118 51070 21564 51076
rect 20808 51006 20814 51070
rect 20878 51006 21020 51070
rect 21080 51006 21086 51070
rect 21150 51006 21564 51070
rect 20808 51000 21020 51006
rect 21118 51000 21564 51006
rect 21624 51206 21836 51212
rect 21624 51142 21630 51206
rect 21694 51142 21836 51206
rect 21624 51070 21836 51142
rect 21624 51006 21630 51070
rect 21694 51006 21836 51070
rect 21624 51000 21836 51006
rect 22032 51206 22244 51212
rect 22032 51142 22038 51206
rect 22102 51142 22244 51206
rect 22032 51070 22244 51142
rect 22032 51006 22038 51070
rect 22102 51006 22244 51070
rect 22032 51000 22244 51006
rect 26928 51000 27276 51212
rect 68952 51000 69164 51212
rect 73848 51206 74060 51212
rect 73848 51142 73854 51206
rect 73918 51142 74060 51206
rect 73848 51070 74060 51142
rect 73848 51006 73854 51070
rect 73918 51006 74060 51070
rect 73848 51000 74060 51006
rect 74256 51206 74468 51212
rect 74256 51142 74398 51206
rect 74462 51142 74468 51206
rect 74256 51070 74468 51142
rect 74256 51006 74398 51070
rect 74462 51006 74468 51070
rect 74256 51000 74468 51006
rect 74664 51206 75284 51212
rect 74664 51142 74806 51206
rect 74870 51142 75284 51206
rect 74664 51136 75284 51142
rect 74664 51000 74876 51136
rect 75072 51070 75284 51136
rect 75072 51006 75214 51070
rect 75278 51006 75284 51070
rect 75072 51000 75284 51006
rect 75480 51070 75692 51348
rect 75480 51006 75622 51070
rect 75686 51006 75692 51070
rect 75480 51000 75692 51006
rect 27064 50940 27140 51000
rect 68952 50940 69028 51000
rect 1768 50804 1980 50940
rect 1224 50800 1980 50804
rect 1224 50798 1818 50800
rect 1224 50734 1230 50798
rect 1294 50744 1818 50798
rect 1874 50744 1980 50800
rect 1294 50734 1980 50744
rect 1224 50728 1980 50734
rect 1768 50592 1980 50728
rect 20400 50798 20612 50804
rect 20400 50734 20406 50798
rect 20470 50734 20612 50798
rect 20400 50592 20612 50734
rect 20808 50798 21156 50804
rect 20808 50734 20814 50798
rect 20878 50734 21086 50798
rect 21150 50734 21156 50798
rect 20808 50728 21156 50734
rect 20808 50668 21020 50728
rect 21216 50668 21564 50804
rect 20808 50662 21564 50668
rect 20808 50598 21222 50662
rect 21286 50598 21564 50662
rect 20808 50592 21564 50598
rect 21624 50798 21836 50804
rect 21624 50734 21630 50798
rect 21694 50734 21836 50798
rect 21624 50662 21836 50734
rect 21624 50598 21766 50662
rect 21830 50598 21836 50662
rect 21624 50592 21836 50598
rect 22032 50798 22244 50804
rect 22032 50734 22038 50798
rect 22102 50734 22244 50798
rect 22032 50662 22244 50734
rect 26928 50728 27276 50940
rect 27200 50668 27276 50728
rect 22032 50598 22174 50662
rect 22238 50598 22244 50662
rect 22032 50592 22244 50598
rect 20536 50532 20612 50592
rect 20400 50390 20612 50532
rect 26928 50456 27276 50668
rect 68952 50728 69164 50940
rect 73848 50798 74060 50804
rect 73848 50734 73854 50798
rect 73918 50734 74060 50798
rect 68952 50668 69028 50728
rect 68952 50456 69164 50668
rect 73848 50662 74060 50734
rect 73848 50598 73854 50662
rect 73918 50598 74060 50662
rect 73848 50592 74060 50598
rect 74256 50798 74468 50804
rect 74256 50734 74398 50798
rect 74462 50734 74468 50798
rect 74256 50662 74468 50734
rect 74256 50598 74262 50662
rect 74326 50598 74468 50662
rect 74256 50592 74468 50598
rect 74664 50662 74876 50804
rect 74664 50598 74806 50662
rect 74870 50598 74876 50662
rect 74664 50592 74876 50598
rect 75072 50798 75284 50804
rect 75072 50734 75214 50798
rect 75278 50734 75284 50798
rect 75072 50662 75284 50734
rect 75072 50598 75078 50662
rect 75142 50598 75284 50662
rect 75072 50592 75284 50598
rect 75480 50798 75692 50804
rect 75480 50734 75622 50798
rect 75686 50734 75692 50798
rect 75480 50592 75692 50734
rect 94112 50800 94324 50940
rect 94112 50744 94176 50800
rect 94232 50744 94324 50800
rect 94112 50668 94324 50744
rect 94112 50662 94732 50668
rect 94112 50598 94662 50662
rect 94726 50598 94732 50662
rect 94112 50592 94732 50598
rect 75480 50532 75556 50592
rect 26928 50396 27004 50456
rect 68952 50396 69028 50456
rect 20400 50326 20406 50390
rect 20470 50326 20612 50390
rect 20400 50320 20612 50326
rect 20808 50184 21020 50396
rect 21216 50390 21564 50396
rect 21216 50326 21222 50390
rect 21286 50326 21564 50390
rect 21216 50184 21564 50326
rect 21624 50390 21836 50396
rect 21624 50326 21766 50390
rect 21830 50326 21836 50390
rect 21624 50254 21836 50326
rect 21624 50190 21630 50254
rect 21694 50190 21836 50254
rect 21624 50184 21836 50190
rect 22032 50390 22244 50396
rect 22032 50326 22174 50390
rect 22238 50326 22244 50390
rect 22032 50254 22244 50326
rect 22032 50190 22174 50254
rect 22238 50190 22244 50254
rect 22032 50184 22244 50190
rect 20808 50124 20884 50184
rect 21488 50124 21564 50184
rect 20400 50118 20612 50124
rect 20400 50054 20406 50118
rect 20470 50054 20612 50118
rect 20400 49776 20612 50054
rect 20808 49852 21020 50124
rect 20808 49776 21156 49852
rect 21216 49846 21564 50124
rect 21216 49782 21358 49846
rect 21422 49782 21564 49846
rect 21216 49776 21564 49782
rect 21624 49982 21836 49988
rect 21624 49918 21630 49982
rect 21694 49918 21836 49982
rect 21624 49776 21836 49918
rect 22032 49982 22244 49988
rect 22032 49918 22174 49982
rect 22238 49918 22244 49982
rect 22032 49776 22244 49918
rect 26928 49912 27276 50396
rect 68952 49982 69164 50396
rect 73848 50390 74060 50396
rect 73848 50326 73854 50390
rect 73918 50326 74060 50390
rect 73848 50254 74060 50326
rect 73848 50190 73854 50254
rect 73918 50190 74060 50254
rect 73848 50184 74060 50190
rect 74256 50390 74468 50396
rect 74256 50326 74262 50390
rect 74326 50326 74468 50390
rect 74256 50254 74468 50326
rect 74256 50190 74262 50254
rect 74326 50190 74468 50254
rect 74256 50184 74468 50190
rect 74664 50390 75284 50396
rect 74664 50326 74806 50390
rect 74870 50326 75078 50390
rect 75142 50326 75284 50390
rect 74664 50320 75284 50326
rect 75480 50390 75692 50532
rect 75480 50326 75622 50390
rect 75686 50326 75692 50390
rect 75480 50320 75692 50326
rect 74664 50260 74876 50320
rect 74664 50184 75012 50260
rect 75072 50184 75284 50320
rect 74800 50124 74876 50184
rect 68952 49918 69094 49982
rect 69158 49918 69164 49982
rect 68952 49912 69164 49918
rect 73848 49982 74060 49988
rect 73848 49918 73854 49982
rect 73918 49918 74060 49982
rect 27064 49852 27140 49912
rect 68952 49852 69028 49912
rect 20400 49716 20476 49776
rect 21080 49716 21156 49776
rect 21624 49716 21700 49776
rect 22032 49716 22108 49776
rect 20400 49574 20612 49716
rect 21080 49640 21292 49716
rect 21216 49580 21292 49640
rect 20400 49510 20406 49574
rect 20470 49510 20612 49574
rect 20400 49504 20612 49510
rect 20808 49574 21564 49580
rect 20808 49510 21358 49574
rect 21422 49510 21564 49574
rect 20808 49504 21564 49510
rect 20808 49368 21020 49504
rect 20944 49308 21020 49368
rect 20400 49302 20612 49308
rect 20400 49238 20406 49302
rect 20470 49238 20612 49302
rect 1224 49166 1980 49172
rect 1224 49102 1230 49166
rect 1294 49120 1980 49166
rect 1294 49102 1818 49120
rect 1224 49096 1818 49102
rect 1768 49064 1818 49096
rect 1874 49064 1980 49120
rect 20400 49166 20612 49238
rect 20400 49102 20542 49166
rect 20606 49102 20612 49166
rect 20400 49096 20612 49102
rect 20808 49096 21020 49308
rect 21216 49368 21564 49504
rect 21624 49368 21836 49716
rect 22032 49368 22244 49716
rect 26928 49710 27276 49852
rect 26928 49646 27206 49710
rect 27270 49646 27276 49710
rect 26928 49438 27276 49646
rect 26928 49374 27206 49438
rect 27270 49374 27276 49438
rect 21216 49308 21292 49368
rect 21624 49308 21700 49368
rect 22032 49308 22108 49368
rect 21216 49166 21564 49308
rect 21216 49102 21222 49166
rect 21286 49102 21564 49166
rect 21216 49096 21564 49102
rect 1768 48960 1980 49064
rect 21624 48960 21836 49308
rect 22032 48960 22244 49308
rect 26928 49232 27276 49374
rect 68952 49710 69164 49852
rect 73848 49776 74060 49918
rect 74256 49982 74468 49988
rect 74256 49918 74262 49982
rect 74326 49918 74468 49982
rect 74256 49776 74468 49918
rect 74664 49776 74876 50124
rect 74936 50124 75012 50184
rect 74936 50048 75284 50124
rect 75072 49846 75284 50048
rect 75072 49782 75078 49846
rect 75142 49782 75284 49846
rect 75072 49776 75284 49782
rect 75480 50118 75692 50124
rect 75480 50054 75622 50118
rect 75686 50054 75692 50118
rect 75480 49776 75692 50054
rect 73984 49716 74060 49776
rect 74392 49716 74468 49776
rect 68952 49646 68958 49710
rect 69022 49646 69094 49710
rect 69158 49646 69164 49710
rect 68952 49438 69164 49646
rect 68952 49374 68958 49438
rect 69022 49374 69164 49438
rect 68952 49232 69164 49374
rect 27064 49172 27140 49232
rect 69088 49172 69164 49232
rect 26928 49096 27276 49172
rect 21624 48900 21700 48960
rect 22168 48900 22244 48960
rect 27054 48900 27152 49096
rect 20400 48894 20612 48900
rect 20400 48830 20542 48894
rect 20606 48830 20612 48894
rect 20400 48758 20612 48830
rect 20400 48694 20542 48758
rect 20606 48694 20612 48758
rect 20400 48688 20612 48694
rect 20808 48552 21020 48900
rect 21216 48894 21564 48900
rect 21216 48830 21222 48894
rect 21286 48830 21564 48894
rect 21216 48628 21564 48830
rect 21624 48758 21836 48900
rect 21624 48694 21766 48758
rect 21830 48694 21836 48758
rect 21624 48688 21836 48694
rect 22032 48758 22244 48900
rect 22032 48694 22038 48758
rect 22102 48694 22244 48758
rect 22032 48688 22244 48694
rect 26928 48688 27276 48900
rect 68952 48894 69164 49172
rect 68952 48830 69094 48894
rect 69158 48830 69164 48894
rect 68952 48688 69164 48830
rect 73848 49368 74060 49716
rect 74256 49368 74468 49716
rect 75480 49716 75556 49776
rect 74664 49368 74876 49580
rect 75072 49574 75284 49580
rect 75072 49510 75078 49574
rect 75142 49510 75284 49574
rect 75072 49444 75284 49510
rect 75480 49574 75692 49716
rect 75480 49510 75622 49574
rect 75686 49510 75692 49574
rect 75480 49504 75692 49510
rect 74936 49368 75284 49444
rect 73848 49308 73924 49368
rect 74256 49308 74332 49368
rect 74664 49308 74740 49368
rect 74936 49308 75012 49368
rect 73848 48960 74060 49308
rect 74256 48960 74468 49308
rect 74664 49232 75012 49308
rect 75072 49308 75148 49368
rect 74664 49096 74876 49232
rect 75072 49166 75284 49308
rect 75072 49102 75214 49166
rect 75278 49102 75284 49166
rect 75072 49096 75284 49102
rect 75480 49302 75692 49308
rect 75480 49238 75622 49302
rect 75686 49238 75692 49302
rect 75480 49166 75692 49238
rect 75480 49102 75622 49166
rect 75686 49102 75692 49166
rect 75480 49096 75692 49102
rect 94112 49166 94732 49172
rect 94112 49120 94662 49166
rect 94112 49064 94176 49120
rect 94232 49102 94662 49120
rect 94726 49102 94732 49166
rect 94232 49096 94732 49102
rect 94232 49064 94324 49096
rect 94112 48960 94324 49064
rect 73848 48900 73924 48960
rect 74392 48900 74468 48960
rect 73848 48758 74060 48900
rect 73848 48694 73990 48758
rect 74054 48694 74060 48758
rect 73848 48688 74060 48694
rect 74256 48758 74468 48900
rect 74256 48694 74398 48758
rect 74462 48694 74468 48758
rect 74256 48688 74468 48694
rect 27064 48628 27140 48688
rect 68952 48628 69028 48688
rect 20944 48492 21020 48552
rect 21080 48552 21564 48628
rect 21080 48492 21156 48552
rect 21352 48492 21428 48552
rect 20400 48486 20612 48492
rect 20400 48422 20542 48486
rect 20606 48422 20612 48486
rect 20400 48350 20612 48422
rect 20400 48286 20542 48350
rect 20606 48286 20612 48350
rect 20400 48280 20612 48286
rect 20808 48416 21156 48492
rect 20808 48350 21020 48416
rect 20808 48286 20814 48350
rect 20878 48286 21020 48350
rect 20808 48280 21020 48286
rect 21216 48350 21564 48492
rect 21216 48286 21494 48350
rect 21558 48286 21564 48350
rect 21216 48280 21564 48286
rect 21624 48486 21836 48492
rect 21624 48422 21766 48486
rect 21830 48422 21836 48486
rect 21624 48350 21836 48422
rect 21624 48286 21766 48350
rect 21830 48286 21836 48350
rect 21624 48280 21836 48286
rect 22032 48486 22244 48492
rect 22032 48422 22038 48486
rect 22102 48422 22244 48486
rect 22032 48350 22244 48422
rect 26928 48416 27276 48628
rect 27200 48356 27276 48416
rect 22032 48286 22038 48350
rect 22102 48286 22244 48350
rect 22032 48280 22244 48286
rect 26928 48144 27276 48356
rect 68952 48622 69164 48628
rect 68952 48558 69094 48622
rect 69158 48558 69164 48622
rect 68952 48416 69164 48558
rect 74664 48552 74876 48900
rect 75072 48894 75284 48900
rect 75072 48830 75214 48894
rect 75278 48830 75284 48894
rect 75072 48552 75284 48830
rect 75480 48894 75692 48900
rect 75480 48830 75622 48894
rect 75686 48830 75692 48894
rect 75480 48758 75692 48830
rect 75480 48694 75486 48758
rect 75550 48694 75692 48758
rect 75480 48688 75692 48694
rect 74664 48492 74740 48552
rect 75072 48492 75148 48552
rect 73848 48486 74060 48492
rect 73848 48422 73990 48486
rect 74054 48422 74060 48486
rect 68952 48356 69028 48416
rect 68952 48144 69164 48356
rect 73848 48350 74060 48422
rect 73848 48286 73854 48350
rect 73918 48286 74060 48350
rect 73848 48280 74060 48286
rect 74256 48486 74468 48492
rect 74256 48422 74398 48486
rect 74462 48422 74468 48486
rect 74256 48350 74468 48422
rect 74256 48286 74398 48350
rect 74462 48286 74468 48350
rect 74256 48280 74468 48286
rect 74664 48350 74876 48492
rect 74664 48286 74806 48350
rect 74870 48286 74876 48350
rect 74664 48280 74876 48286
rect 75072 48280 75284 48492
rect 75480 48486 75692 48492
rect 75480 48422 75486 48486
rect 75550 48422 75692 48486
rect 75480 48350 75692 48422
rect 75480 48286 75622 48350
rect 75686 48286 75692 48350
rect 75480 48280 75692 48286
rect 75072 48220 75148 48280
rect 27200 48084 27276 48144
rect 69088 48084 69164 48144
rect 74800 48144 75148 48220
rect 74800 48084 74876 48144
rect 20400 48078 20612 48084
rect 20400 48014 20542 48078
rect 20606 48014 20612 48078
rect 20400 47942 20612 48014
rect 20400 47878 20406 47942
rect 20470 47878 20612 47942
rect 20400 47872 20612 47878
rect 20808 48078 21020 48084
rect 20808 48014 20814 48078
rect 20878 48014 21020 48078
rect 20808 47872 21020 48014
rect 21216 48078 21564 48084
rect 21216 48014 21494 48078
rect 21558 48014 21564 48078
rect 21216 47948 21564 48014
rect 21118 47942 21564 47948
rect 21080 47878 21086 47942
rect 21150 47878 21358 47942
rect 21422 47878 21564 47942
rect 21118 47872 21564 47878
rect 21624 48078 21836 48084
rect 21624 48014 21766 48078
rect 21830 48014 21836 48078
rect 21624 47942 21836 48014
rect 21624 47878 21766 47942
rect 21830 47878 21836 47942
rect 21624 47872 21836 47878
rect 22032 48078 22244 48084
rect 22032 48014 22038 48078
rect 22102 48014 22244 48078
rect 22032 47942 22244 48014
rect 22032 47878 22038 47942
rect 22102 47878 22244 47942
rect 22032 47872 22244 47878
rect 26928 47872 27276 48084
rect 68952 47872 69164 48084
rect 73848 48078 74060 48084
rect 73848 48014 73854 48078
rect 73918 48014 74060 48078
rect 73848 47942 74060 48014
rect 73848 47878 73990 47942
rect 74054 47878 74060 47942
rect 73848 47872 74060 47878
rect 74256 48078 74468 48084
rect 74256 48014 74398 48078
rect 74462 48014 74468 48078
rect 74256 47942 74468 48014
rect 74256 47878 74398 47942
rect 74462 47878 74468 47942
rect 74256 47872 74468 47878
rect 74664 48078 75284 48084
rect 74664 48014 74806 48078
rect 74870 48014 75284 48078
rect 74664 48008 75284 48014
rect 74664 47872 74876 48008
rect 75072 47942 75284 48008
rect 75072 47878 75078 47942
rect 75142 47878 75284 47942
rect 75072 47872 75284 47878
rect 75480 48078 75692 48084
rect 75480 48014 75622 48078
rect 75686 48014 75692 48078
rect 75480 47942 75692 48014
rect 75480 47878 75622 47942
rect 75686 47878 75692 47942
rect 75480 47872 75692 47878
rect 26928 47812 27004 47872
rect 69088 47812 69164 47872
rect 20400 47670 20612 47676
rect 20400 47606 20406 47670
rect 20470 47606 20612 47670
rect 1224 47534 1980 47540
rect 1224 47470 1230 47534
rect 1294 47470 1980 47534
rect 1224 47464 1980 47470
rect 20400 47534 20612 47606
rect 20400 47470 20542 47534
rect 20606 47470 20612 47534
rect 20400 47464 20612 47470
rect 20808 47670 21156 47676
rect 20808 47606 21086 47670
rect 21150 47606 21156 47670
rect 20808 47600 21156 47606
rect 21216 47670 21564 47676
rect 21216 47606 21358 47670
rect 21422 47606 21564 47670
rect 20808 47540 21020 47600
rect 20808 47534 21156 47540
rect 20808 47470 21086 47534
rect 21150 47470 21156 47534
rect 20808 47464 21156 47470
rect 21216 47464 21564 47606
rect 21624 47670 21836 47676
rect 21624 47606 21766 47670
rect 21830 47606 21836 47670
rect 21624 47534 21836 47606
rect 21624 47470 21766 47534
rect 21830 47470 21836 47534
rect 21624 47464 21836 47470
rect 22032 47670 22244 47676
rect 22032 47606 22038 47670
rect 22102 47606 22244 47670
rect 22032 47534 22244 47606
rect 26928 47600 27276 47812
rect 27200 47540 27276 47600
rect 22032 47470 22174 47534
rect 22238 47470 22244 47534
rect 22032 47464 22244 47470
rect 1768 47440 1980 47464
rect 1768 47384 1818 47440
rect 1874 47384 1980 47440
rect 1768 47328 1980 47384
rect 26928 47328 27276 47540
rect 68952 47600 69164 47812
rect 73848 47670 74060 47676
rect 73848 47606 73990 47670
rect 74054 47606 74060 47670
rect 68952 47540 69028 47600
rect 68952 47328 69164 47540
rect 73848 47534 74060 47606
rect 73848 47470 73990 47534
rect 74054 47470 74060 47534
rect 73848 47464 74060 47470
rect 74256 47670 74468 47676
rect 74256 47606 74398 47670
rect 74462 47606 74468 47670
rect 74256 47534 74468 47606
rect 74256 47470 74398 47534
rect 74462 47470 74468 47534
rect 74256 47464 74468 47470
rect 74664 47670 75284 47676
rect 74664 47606 75078 47670
rect 75142 47606 75284 47670
rect 74664 47600 75284 47606
rect 74664 47534 74876 47600
rect 74664 47470 74670 47534
rect 74734 47470 74876 47534
rect 74664 47464 74876 47470
rect 75072 47464 75284 47600
rect 75480 47670 75692 47676
rect 75480 47606 75622 47670
rect 75686 47606 75692 47670
rect 75480 47534 75692 47606
rect 75480 47470 75486 47534
rect 75550 47470 75692 47534
rect 75480 47464 75692 47470
rect 94112 47534 94732 47540
rect 94112 47470 94662 47534
rect 94726 47470 94732 47534
rect 94112 47464 94732 47470
rect 94112 47440 94324 47464
rect 94112 47384 94176 47440
rect 94232 47384 94324 47440
rect 94112 47328 94324 47384
rect 27064 47268 27140 47328
rect 68952 47268 69028 47328
rect 20400 47262 20612 47268
rect 20400 47198 20542 47262
rect 20606 47198 20612 47262
rect 20400 47126 20612 47198
rect 20400 47062 20406 47126
rect 20470 47062 20612 47126
rect 20400 47056 20612 47062
rect 20808 47126 21020 47268
rect 21118 47262 21564 47268
rect 21080 47198 21086 47262
rect 21150 47198 21564 47262
rect 21118 47192 21564 47198
rect 20808 47062 20814 47126
rect 20878 47062 21020 47126
rect 20808 47056 21020 47062
rect 21216 47126 21564 47192
rect 21216 47062 21494 47126
rect 21558 47062 21564 47126
rect 21216 47056 21564 47062
rect 21624 47262 21836 47268
rect 21624 47198 21766 47262
rect 21830 47198 21836 47262
rect 21624 47126 21836 47198
rect 21624 47062 21630 47126
rect 21694 47062 21836 47126
rect 21624 47056 21836 47062
rect 22032 47262 22244 47268
rect 22032 47198 22174 47262
rect 22238 47198 22244 47262
rect 22032 47126 22244 47198
rect 22032 47062 22038 47126
rect 22102 47062 22244 47126
rect 22032 47056 22244 47062
rect 26928 47056 27276 47268
rect 68952 47056 69164 47268
rect 73848 47262 74060 47268
rect 73848 47198 73990 47262
rect 74054 47198 74060 47262
rect 73848 47126 74060 47198
rect 73848 47062 73854 47126
rect 73918 47062 74060 47126
rect 73848 47056 74060 47062
rect 74256 47262 74468 47268
rect 74256 47198 74398 47262
rect 74462 47198 74468 47262
rect 74256 47126 74468 47198
rect 74256 47062 74262 47126
rect 74326 47062 74468 47126
rect 74256 47056 74468 47062
rect 74664 47262 74876 47268
rect 74664 47198 74670 47262
rect 74734 47198 74876 47262
rect 74664 47126 74876 47198
rect 75072 47132 75284 47268
rect 74974 47126 75284 47132
rect 74664 47062 74806 47126
rect 74870 47062 74876 47126
rect 74936 47062 74942 47126
rect 75006 47062 75284 47126
rect 74664 47056 74876 47062
rect 74974 47056 75284 47062
rect 75480 47262 75692 47268
rect 75480 47198 75486 47262
rect 75550 47198 75692 47262
rect 75480 47126 75692 47198
rect 75480 47062 75622 47126
rect 75686 47062 75692 47126
rect 75480 47056 75692 47062
rect 21488 46996 21564 47056
rect 26928 46996 27004 47056
rect 69088 46996 69164 47056
rect 21488 46920 22108 46996
rect 22032 46860 22108 46920
rect 20400 46854 20612 46860
rect 20400 46790 20406 46854
rect 20470 46790 20612 46854
rect 20400 46648 20612 46790
rect 20808 46854 21020 46860
rect 20808 46790 20814 46854
rect 20878 46790 21020 46854
rect 20808 46718 21020 46790
rect 20808 46654 20814 46718
rect 20878 46654 21020 46718
rect 20808 46648 21020 46654
rect 21216 46854 21564 46860
rect 21216 46790 21494 46854
rect 21558 46790 21564 46854
rect 21216 46648 21564 46790
rect 21624 46854 21836 46860
rect 21624 46790 21630 46854
rect 21694 46790 21836 46854
rect 21624 46718 21836 46790
rect 21624 46654 21766 46718
rect 21830 46654 21836 46718
rect 21624 46648 21836 46654
rect 22032 46854 22244 46860
rect 22032 46790 22038 46854
rect 22102 46790 22244 46854
rect 22032 46718 22244 46790
rect 26928 46784 27276 46996
rect 68952 46784 69164 46996
rect 27064 46724 27140 46784
rect 69088 46724 69164 46784
rect 22032 46654 22174 46718
rect 22238 46654 22244 46718
rect 22032 46648 22244 46654
rect 20400 46588 20476 46648
rect 21216 46588 21292 46648
rect 20400 46240 20612 46588
rect 20944 46512 21292 46588
rect 26928 46512 27276 46724
rect 20944 46452 21020 46512
rect 27200 46452 27276 46512
rect 20808 46446 21564 46452
rect 20808 46382 20814 46446
rect 20878 46382 21564 46446
rect 20808 46376 21564 46382
rect 20808 46240 21020 46376
rect 20536 46180 20612 46240
rect 20944 46180 21020 46240
rect 1224 45902 1980 45908
rect 1224 45838 1230 45902
rect 1294 45838 1980 45902
rect 1224 45832 1980 45838
rect 20400 45832 20612 46180
rect 20808 45832 21020 46180
rect 21216 46240 21564 46376
rect 21624 46446 21836 46452
rect 21624 46382 21766 46446
rect 21830 46382 21836 46446
rect 21624 46310 21836 46382
rect 21624 46246 21766 46310
rect 21830 46246 21836 46310
rect 21624 46240 21836 46246
rect 22032 46446 22244 46452
rect 22032 46382 22174 46446
rect 22238 46382 22244 46446
rect 22032 46310 22244 46382
rect 22032 46246 22038 46310
rect 22102 46246 22244 46310
rect 22032 46240 22244 46246
rect 21216 46180 21292 46240
rect 21216 45902 21564 46180
rect 21216 45838 21494 45902
rect 21558 45838 21564 45902
rect 21216 45832 21564 45838
rect 21624 46038 21836 46044
rect 21624 45974 21766 46038
rect 21830 45974 21836 46038
rect 21624 45832 21836 45974
rect 22032 46038 22244 46044
rect 22032 45974 22038 46038
rect 22102 45974 22244 46038
rect 22032 45832 22244 45974
rect 26928 45968 27276 46452
rect 68952 46582 69164 46724
rect 73848 46854 74060 46860
rect 73848 46790 73854 46854
rect 73918 46790 74060 46854
rect 73848 46718 74060 46790
rect 73848 46654 73990 46718
rect 74054 46654 74060 46718
rect 73848 46648 74060 46654
rect 74256 46854 74468 46860
rect 74256 46790 74262 46854
rect 74326 46790 74468 46854
rect 74256 46718 74468 46790
rect 74256 46654 74262 46718
rect 74326 46654 74468 46718
rect 74256 46648 74468 46654
rect 74664 46854 75012 46860
rect 74664 46790 74806 46854
rect 74870 46790 74942 46854
rect 75006 46790 75012 46854
rect 74664 46784 75012 46790
rect 74664 46724 74876 46784
rect 75072 46724 75284 46860
rect 74664 46718 75284 46724
rect 74664 46654 74670 46718
rect 74734 46654 75284 46718
rect 74664 46648 75284 46654
rect 75480 46854 75692 46860
rect 75480 46790 75622 46854
rect 75686 46790 75692 46854
rect 75480 46648 75692 46790
rect 68952 46518 68958 46582
rect 69022 46518 69164 46582
rect 68952 46512 69164 46518
rect 75480 46588 75556 46648
rect 68952 46452 69028 46512
rect 68952 46310 69164 46452
rect 68952 46246 68958 46310
rect 69022 46246 69164 46310
rect 68952 46038 69164 46246
rect 73848 46446 74060 46452
rect 73848 46382 73990 46446
rect 74054 46382 74060 46446
rect 73848 46310 74060 46382
rect 73848 46246 73990 46310
rect 74054 46246 74060 46310
rect 73848 46240 74060 46246
rect 74256 46446 74468 46452
rect 74256 46382 74262 46446
rect 74326 46382 74468 46446
rect 74256 46310 74468 46382
rect 74256 46246 74262 46310
rect 74326 46246 74468 46310
rect 74256 46240 74468 46246
rect 74664 46446 74876 46452
rect 74664 46382 74670 46446
rect 74734 46382 74876 46446
rect 74664 46240 74876 46382
rect 75072 46316 75284 46452
rect 74800 46180 74876 46240
rect 74936 46240 75284 46316
rect 75480 46240 75692 46588
rect 74936 46180 75012 46240
rect 75480 46180 75556 46240
rect 74664 46104 75012 46180
rect 74664 46044 74876 46104
rect 75072 46044 75284 46180
rect 68952 45974 68958 46038
rect 69022 45974 69164 46038
rect 68952 45968 69164 45974
rect 73848 46038 74060 46044
rect 73848 45974 73990 46038
rect 74054 45974 74060 46038
rect 26928 45908 27004 45968
rect 1768 45760 1980 45832
rect 20536 45772 20612 45832
rect 1768 45704 1818 45760
rect 1874 45704 1980 45760
rect 1768 45560 1980 45704
rect 20400 45630 20612 45772
rect 21624 45772 21700 45832
rect 22032 45772 22108 45832
rect 20400 45566 20542 45630
rect 20606 45566 20612 45630
rect 20400 45560 20612 45566
rect 20808 45424 21020 45636
rect 21216 45630 21564 45636
rect 21216 45566 21494 45630
rect 21558 45566 21564 45630
rect 21216 45500 21564 45566
rect 21118 45494 21564 45500
rect 21080 45430 21086 45494
rect 21150 45430 21564 45494
rect 21118 45424 21564 45430
rect 21624 45424 21836 45772
rect 22032 45424 22244 45772
rect 20944 45364 21020 45424
rect 21624 45364 21700 45424
rect 22168 45364 22244 45424
rect 20400 45358 20612 45364
rect 20400 45294 20542 45358
rect 20606 45294 20612 45358
rect 20400 45222 20612 45294
rect 20400 45158 20542 45222
rect 20606 45158 20612 45222
rect 20400 45152 20612 45158
rect 20808 45288 21564 45364
rect 20808 45228 21020 45288
rect 20808 45222 21156 45228
rect 20808 45158 21086 45222
rect 21150 45158 21156 45222
rect 20808 45152 21156 45158
rect 21216 45222 21564 45288
rect 21216 45158 21358 45222
rect 21422 45158 21564 45222
rect 21216 45152 21564 45158
rect 21624 45016 21836 45364
rect 22032 45016 22244 45364
rect 26928 45358 27276 45908
rect 26928 45294 27206 45358
rect 27270 45294 27276 45358
rect 26928 45288 27276 45294
rect 68952 45766 69164 45908
rect 68952 45702 68958 45766
rect 69022 45702 69094 45766
rect 69158 45702 69164 45766
rect 68952 45494 69164 45702
rect 68952 45430 69094 45494
rect 69158 45430 69164 45494
rect 68952 45358 69164 45430
rect 73848 45832 74060 45974
rect 74256 46038 74468 46044
rect 74256 45974 74262 46038
rect 74326 45974 74468 46038
rect 74256 45832 74468 45974
rect 74664 45968 75284 46044
rect 74664 45908 74876 45968
rect 74664 45902 75012 45908
rect 74664 45838 74806 45902
rect 74870 45838 74942 45902
rect 75006 45838 75012 45902
rect 74664 45832 75012 45838
rect 75072 45832 75284 45968
rect 75480 45832 75692 46180
rect 73848 45772 73924 45832
rect 74256 45772 74332 45832
rect 75616 45772 75692 45832
rect 73848 45424 74060 45772
rect 74256 45500 74468 45772
rect 74664 45630 74876 45636
rect 74974 45630 75284 45636
rect 74664 45566 74806 45630
rect 74870 45566 74876 45630
rect 74936 45566 74942 45630
rect 75006 45566 75284 45630
rect 74256 45494 74604 45500
rect 74256 45430 74534 45494
rect 74598 45430 74604 45494
rect 74256 45424 74604 45430
rect 74664 45424 74876 45566
rect 74974 45560 75284 45566
rect 75480 45630 75692 45772
rect 75480 45566 75486 45630
rect 75550 45566 75692 45630
rect 75480 45560 75692 45566
rect 94112 45902 94732 45908
rect 94112 45838 94662 45902
rect 94726 45838 94732 45902
rect 94112 45832 94732 45838
rect 94112 45760 94324 45832
rect 94112 45704 94176 45760
rect 94232 45704 94324 45760
rect 94112 45560 94324 45704
rect 75072 45424 75284 45560
rect 73984 45364 74060 45424
rect 74392 45364 74468 45424
rect 68952 45294 68958 45358
rect 69022 45294 69164 45358
rect 68952 45288 69164 45294
rect 26928 45086 27276 45092
rect 26928 45022 27206 45086
rect 27270 45022 27276 45086
rect 21624 44956 21700 45016
rect 22032 44956 22108 45016
rect 20400 44950 20612 44956
rect 20400 44886 20542 44950
rect 20606 44886 20612 44950
rect 20400 44814 20612 44886
rect 20400 44750 20406 44814
rect 20470 44750 20612 44814
rect 20400 44744 20612 44750
rect 20808 44608 21020 44956
rect 21216 44950 21564 44956
rect 21216 44886 21358 44950
rect 21422 44886 21564 44950
rect 21216 44684 21564 44886
rect 21624 44814 21836 44956
rect 21624 44750 21630 44814
rect 21694 44750 21836 44814
rect 21624 44744 21836 44750
rect 22032 44814 22244 44956
rect 22032 44750 22174 44814
rect 22238 44750 22244 44814
rect 22032 44744 22244 44750
rect 26928 44744 27276 45022
rect 68952 45086 69164 45092
rect 68952 45022 68958 45086
rect 69022 45022 69164 45086
rect 68952 44950 69164 45022
rect 68952 44886 69094 44950
rect 69158 44886 69164 44950
rect 68952 44744 69164 44886
rect 73848 45016 74060 45364
rect 74256 45016 74468 45364
rect 74664 45364 74740 45424
rect 75072 45364 75148 45424
rect 74664 45152 74876 45364
rect 75072 45222 75284 45364
rect 75072 45158 75078 45222
rect 75142 45158 75284 45222
rect 75072 45152 75284 45158
rect 75480 45358 75692 45364
rect 75480 45294 75486 45358
rect 75550 45294 75692 45358
rect 75480 45222 75692 45294
rect 75480 45158 75486 45222
rect 75550 45158 75692 45222
rect 75480 45152 75692 45158
rect 74566 45086 75556 45092
rect 74528 45022 74534 45086
rect 74598 45022 75556 45086
rect 74566 45016 75556 45022
rect 73848 44956 73924 45016
rect 74256 44956 74332 45016
rect 75480 44956 75556 45016
rect 73848 44814 74060 44956
rect 73848 44750 73854 44814
rect 73918 44750 74060 44814
rect 73848 44744 74060 44750
rect 74256 44814 74468 44956
rect 74256 44750 74262 44814
rect 74326 44750 74468 44814
rect 74256 44744 74468 44750
rect 74664 44820 74876 44956
rect 75072 44950 75284 44956
rect 75072 44886 75078 44950
rect 75142 44886 75284 44950
rect 74664 44814 75012 44820
rect 74664 44750 74942 44814
rect 75006 44750 75012 44814
rect 74664 44744 75012 44750
rect 27064 44684 27140 44744
rect 69088 44684 69164 44744
rect 21080 44608 21564 44684
rect 20808 44548 20884 44608
rect 21080 44548 21156 44608
rect 20400 44542 20612 44548
rect 20400 44478 20406 44542
rect 20470 44478 20612 44542
rect 20400 44406 20612 44478
rect 20400 44342 20542 44406
rect 20606 44342 20612 44406
rect 20400 44336 20612 44342
rect 20808 44472 21156 44548
rect 20808 44412 21020 44472
rect 21216 44412 21564 44548
rect 20808 44336 21564 44412
rect 21624 44542 21836 44548
rect 21624 44478 21630 44542
rect 21694 44478 21836 44542
rect 21624 44406 21836 44478
rect 21624 44342 21766 44406
rect 21830 44342 21836 44406
rect 21624 44336 21836 44342
rect 22032 44542 22244 44548
rect 22032 44478 22174 44542
rect 22238 44478 22244 44542
rect 22032 44406 22244 44478
rect 26928 44472 27276 44684
rect 27200 44412 27276 44472
rect 22032 44342 22038 44406
rect 22102 44342 22244 44406
rect 22032 44336 22244 44342
rect 21216 44276 21292 44336
rect 20944 44200 21292 44276
rect 20944 44140 21020 44200
rect 1768 44080 1980 44140
rect 1768 44024 1818 44080
rect 1874 44024 1980 44080
rect 1768 44004 1980 44024
rect 1224 43998 1980 44004
rect 1224 43934 1230 43998
rect 1294 43934 1980 43998
rect 1224 43928 1980 43934
rect 20400 44134 20612 44140
rect 20400 44070 20542 44134
rect 20606 44070 20612 44134
rect 20400 43998 20612 44070
rect 20400 43934 20406 43998
rect 20470 43934 20612 43998
rect 20400 43928 20612 43934
rect 20808 44064 21564 44140
rect 20808 44004 21020 44064
rect 20808 43998 21156 44004
rect 20808 43934 21086 43998
rect 21150 43934 21156 43998
rect 20808 43928 21156 43934
rect 21216 43928 21564 44064
rect 21624 44134 21836 44140
rect 21624 44070 21766 44134
rect 21830 44070 21836 44134
rect 21624 43998 21836 44070
rect 21624 43934 21766 43998
rect 21830 43934 21836 43998
rect 21624 43928 21836 43934
rect 22032 44134 22244 44140
rect 22032 44070 22038 44134
rect 22102 44070 22244 44134
rect 22032 43998 22244 44070
rect 22032 43934 22038 43998
rect 22102 43934 22244 43998
rect 22032 43928 22244 43934
rect 26928 43928 27276 44412
rect 68952 44678 69164 44684
rect 68952 44614 69094 44678
rect 69158 44614 69164 44678
rect 68952 44472 69164 44614
rect 74664 44684 74876 44744
rect 75072 44684 75284 44886
rect 75480 44950 75692 44956
rect 75480 44886 75486 44950
rect 75550 44886 75692 44950
rect 75480 44814 75692 44886
rect 75480 44750 75622 44814
rect 75686 44750 75692 44814
rect 75480 44744 75692 44750
rect 74664 44608 75284 44684
rect 74800 44548 74876 44608
rect 73848 44542 74060 44548
rect 73848 44478 73854 44542
rect 73918 44478 74060 44542
rect 68952 44412 69028 44472
rect 68952 44134 69164 44412
rect 73848 44406 74060 44478
rect 73848 44342 73990 44406
rect 74054 44342 74060 44406
rect 73848 44336 74060 44342
rect 74256 44542 74468 44548
rect 74256 44478 74262 44542
rect 74326 44478 74468 44542
rect 74256 44406 74468 44478
rect 74256 44342 74398 44406
rect 74462 44342 74468 44406
rect 74256 44336 74468 44342
rect 74664 44406 74876 44548
rect 74974 44542 75284 44548
rect 74936 44478 74942 44542
rect 75006 44478 75284 44542
rect 74974 44472 75284 44478
rect 74664 44342 74670 44406
rect 74734 44342 74876 44406
rect 74664 44336 74876 44342
rect 75072 44336 75284 44472
rect 75480 44542 75692 44548
rect 75480 44478 75622 44542
rect 75686 44478 75692 44542
rect 75480 44406 75692 44478
rect 75480 44342 75486 44406
rect 75550 44342 75692 44406
rect 75480 44336 75692 44342
rect 68952 44070 69094 44134
rect 69158 44070 69164 44134
rect 68952 43928 69164 44070
rect 73848 44134 74060 44140
rect 73848 44070 73990 44134
rect 74054 44070 74060 44134
rect 73848 43998 74060 44070
rect 73848 43934 73990 43998
rect 74054 43934 74060 43998
rect 73848 43928 74060 43934
rect 74256 44134 74468 44140
rect 74256 44070 74398 44134
rect 74462 44070 74468 44134
rect 74256 43998 74468 44070
rect 74256 43934 74398 43998
rect 74462 43934 74468 43998
rect 74256 43928 74468 43934
rect 74664 44134 74876 44140
rect 74664 44070 74670 44134
rect 74734 44070 74876 44134
rect 74664 43998 74876 44070
rect 74664 43934 74806 43998
rect 74870 43934 74876 43998
rect 74664 43928 74876 43934
rect 75072 43928 75284 44140
rect 75480 44134 75692 44140
rect 75480 44070 75486 44134
rect 75550 44070 75692 44134
rect 75480 43998 75692 44070
rect 75480 43934 75622 43998
rect 75686 43934 75692 43998
rect 75480 43928 75692 43934
rect 94112 44080 94324 44140
rect 94112 44024 94176 44080
rect 94232 44024 94324 44080
rect 94112 44004 94324 44024
rect 94112 43998 94732 44004
rect 94112 43934 94662 43998
rect 94726 43934 94732 43998
rect 94112 43928 94732 43934
rect 27200 43868 27276 43928
rect 69088 43868 69164 43928
rect 75072 43868 75148 43928
rect 20400 43726 20612 43732
rect 20400 43662 20406 43726
rect 20470 43662 20612 43726
rect 20400 43590 20612 43662
rect 20400 43526 20406 43590
rect 20470 43526 20612 43590
rect 20400 43520 20612 43526
rect 20808 43590 21020 43732
rect 21118 43726 21564 43732
rect 21080 43662 21086 43726
rect 21150 43662 21564 43726
rect 21118 43656 21564 43662
rect 21216 43596 21564 43656
rect 21118 43590 21564 43596
rect 20808 43526 20950 43590
rect 21014 43526 21020 43590
rect 21080 43526 21086 43590
rect 21150 43526 21564 43590
rect 20808 43520 21020 43526
rect 21118 43520 21564 43526
rect 21624 43726 21836 43732
rect 21624 43662 21766 43726
rect 21830 43662 21836 43726
rect 21624 43590 21836 43662
rect 21624 43526 21766 43590
rect 21830 43526 21836 43590
rect 21624 43520 21836 43526
rect 22032 43726 22244 43732
rect 22032 43662 22038 43726
rect 22102 43662 22244 43726
rect 22032 43590 22244 43662
rect 26928 43656 27276 43868
rect 68952 43862 69164 43868
rect 68952 43798 69094 43862
rect 69158 43798 69164 43862
rect 68952 43656 69164 43798
rect 74800 43792 75148 43868
rect 74800 43732 74876 43792
rect 27064 43596 27140 43656
rect 69088 43596 69164 43656
rect 22032 43526 22038 43590
rect 22102 43526 22244 43590
rect 22032 43520 22244 43526
rect 26928 43384 27276 43596
rect 27200 43324 27276 43384
rect 20400 43318 20612 43324
rect 20400 43254 20406 43318
rect 20470 43254 20612 43318
rect 20400 43182 20612 43254
rect 20400 43118 20542 43182
rect 20606 43118 20612 43182
rect 20400 43112 20612 43118
rect 20808 43318 21156 43324
rect 20808 43254 20950 43318
rect 21014 43254 21086 43318
rect 21150 43254 21156 43318
rect 20808 43248 21156 43254
rect 20808 43188 21020 43248
rect 21216 43188 21564 43324
rect 20808 43182 21564 43188
rect 20808 43118 21222 43182
rect 21286 43118 21564 43182
rect 20808 43112 21564 43118
rect 21624 43318 21836 43324
rect 21624 43254 21766 43318
rect 21830 43254 21836 43318
rect 21624 43182 21836 43254
rect 21624 43118 21766 43182
rect 21830 43118 21836 43182
rect 21624 43112 21836 43118
rect 22032 43318 22244 43324
rect 22032 43254 22038 43318
rect 22102 43254 22244 43318
rect 22032 43182 22244 43254
rect 22032 43118 22174 43182
rect 22238 43118 22244 43182
rect 22032 43112 22244 43118
rect 26928 43112 27276 43324
rect 68952 43384 69164 43596
rect 73848 43726 74060 43732
rect 73848 43662 73990 43726
rect 74054 43662 74060 43726
rect 73848 43590 74060 43662
rect 73848 43526 73990 43590
rect 74054 43526 74060 43590
rect 73848 43520 74060 43526
rect 74256 43726 74468 43732
rect 74256 43662 74398 43726
rect 74462 43662 74468 43726
rect 74256 43590 74468 43662
rect 74256 43526 74262 43590
rect 74326 43526 74468 43590
rect 74256 43520 74468 43526
rect 74664 43726 75284 43732
rect 74664 43662 74806 43726
rect 74870 43662 75284 43726
rect 74664 43656 75284 43662
rect 74664 43590 74876 43656
rect 74664 43526 74670 43590
rect 74734 43526 74876 43590
rect 74664 43520 74876 43526
rect 75072 43520 75284 43656
rect 75480 43726 75692 43732
rect 75480 43662 75622 43726
rect 75686 43662 75692 43726
rect 75480 43590 75692 43662
rect 75480 43526 75622 43590
rect 75686 43526 75692 43590
rect 75480 43520 75692 43526
rect 68952 43324 69028 43384
rect 68952 43112 69164 43324
rect 73848 43318 74060 43324
rect 73848 43254 73990 43318
rect 74054 43254 74060 43318
rect 73848 43182 74060 43254
rect 73848 43118 73990 43182
rect 74054 43118 74060 43182
rect 73848 43112 74060 43118
rect 74256 43318 74468 43324
rect 74256 43254 74262 43318
rect 74326 43254 74468 43318
rect 74256 43182 74468 43254
rect 74256 43118 74262 43182
rect 74326 43118 74468 43182
rect 74256 43112 74468 43118
rect 74664 43318 74876 43324
rect 74664 43254 74670 43318
rect 74734 43254 74876 43318
rect 74664 43182 74876 43254
rect 74664 43118 74670 43182
rect 74734 43118 74876 43182
rect 74664 43112 74876 43118
rect 75072 43182 75284 43324
rect 75072 43118 75078 43182
rect 75142 43118 75284 43182
rect 75072 43112 75284 43118
rect 75480 43318 75692 43324
rect 75480 43254 75622 43318
rect 75686 43254 75692 43318
rect 75480 43182 75692 43254
rect 75480 43118 75486 43182
rect 75550 43118 75692 43182
rect 75480 43112 75692 43118
rect 27064 43052 27140 43112
rect 68952 43052 69028 43112
rect 26928 42916 27276 43052
rect 20400 42910 20612 42916
rect 20400 42846 20542 42910
rect 20606 42846 20612 42910
rect 20400 42704 20612 42846
rect 20808 42774 21020 42916
rect 20808 42710 20814 42774
rect 20878 42710 21020 42774
rect 20808 42704 21020 42710
rect 21216 42910 21564 42916
rect 21216 42846 21222 42910
rect 21286 42846 21564 42910
rect 21216 42774 21564 42846
rect 21216 42710 21358 42774
rect 21422 42710 21564 42774
rect 21216 42704 21564 42710
rect 21624 42910 21836 42916
rect 21624 42846 21766 42910
rect 21830 42846 21836 42910
rect 21624 42780 21836 42846
rect 22032 42910 22244 42916
rect 25470 42910 27276 42916
rect 22032 42846 22174 42910
rect 22238 42846 22244 42910
rect 25432 42846 25438 42910
rect 25502 42846 27276 42910
rect 21624 42774 21972 42780
rect 21624 42710 21630 42774
rect 21694 42710 21972 42774
rect 21624 42704 21972 42710
rect 22032 42774 22244 42846
rect 25470 42840 27276 42846
rect 68952 42840 69164 43052
rect 73848 42910 74060 42916
rect 73848 42846 73990 42910
rect 74054 42846 74060 42910
rect 27064 42780 27140 42840
rect 68952 42780 69028 42840
rect 73848 42780 74060 42846
rect 22032 42710 22038 42774
rect 22102 42710 22244 42774
rect 22032 42704 22244 42710
rect 20536 42644 20612 42704
rect 1768 42400 1980 42508
rect 1768 42372 1818 42400
rect 1224 42366 1818 42372
rect 1224 42302 1230 42366
rect 1294 42344 1818 42366
rect 1874 42344 1980 42400
rect 1294 42302 1980 42344
rect 1224 42296 1980 42302
rect 20400 42296 20612 42644
rect 21896 42644 21972 42704
rect 21896 42568 22516 42644
rect 22440 42508 22516 42568
rect 22712 42568 24012 42644
rect 22712 42508 22788 42568
rect 23936 42508 24012 42568
rect 26928 42568 27276 42780
rect 68952 42638 69164 42780
rect 73342 42774 74060 42780
rect 73304 42710 73310 42774
rect 73374 42710 73854 42774
rect 73918 42710 74060 42774
rect 73342 42704 74060 42710
rect 74256 42910 74468 42916
rect 74256 42846 74262 42910
rect 74326 42846 74468 42910
rect 74256 42774 74468 42846
rect 74256 42710 74262 42774
rect 74326 42710 74468 42774
rect 74256 42704 74468 42710
rect 74664 42910 74876 42916
rect 74664 42846 74670 42910
rect 74734 42846 74876 42910
rect 74664 42780 74876 42846
rect 75072 42910 75284 42916
rect 75072 42846 75078 42910
rect 75142 42846 75284 42910
rect 74664 42774 75012 42780
rect 74664 42710 74942 42774
rect 75006 42710 75012 42774
rect 74664 42704 75012 42710
rect 75072 42704 75284 42846
rect 75480 42910 75692 42916
rect 75480 42846 75486 42910
rect 75550 42846 75692 42910
rect 75480 42704 75692 42846
rect 75072 42644 75148 42704
rect 75616 42644 75692 42704
rect 68952 42574 69094 42638
rect 69158 42574 69164 42638
rect 68952 42568 69164 42574
rect 26928 42508 27004 42568
rect 69088 42508 69164 42568
rect 71808 42568 73108 42644
rect 71808 42508 71884 42568
rect 73032 42508 73108 42568
rect 74800 42568 75148 42644
rect 74800 42508 74876 42568
rect 20808 42502 21020 42508
rect 20808 42438 20814 42502
rect 20878 42438 21020 42502
rect 20808 42296 21020 42438
rect 21216 42502 21564 42508
rect 21216 42438 21358 42502
rect 21422 42438 21564 42502
rect 21216 42372 21564 42438
rect 21080 42296 21564 42372
rect 21624 42502 21836 42508
rect 21624 42438 21630 42502
rect 21694 42438 21836 42502
rect 21624 42366 21836 42438
rect 21624 42302 21766 42366
rect 21830 42302 21836 42366
rect 21624 42296 21836 42302
rect 22032 42502 22244 42508
rect 22032 42438 22038 42502
rect 22102 42438 22244 42502
rect 22032 42372 22244 42438
rect 22440 42432 22788 42508
rect 22032 42366 22380 42372
rect 22032 42302 22174 42366
rect 22238 42302 22380 42366
rect 22032 42296 22380 42302
rect 22440 42296 22652 42432
rect 22848 42372 23196 42508
rect 23936 42502 25508 42508
rect 23936 42438 25438 42502
rect 25502 42438 25508 42502
rect 23936 42432 25508 42438
rect 22848 42296 23876 42372
rect 23936 42296 24148 42432
rect 25568 42296 25780 42508
rect 20400 42236 20476 42296
rect 20808 42236 20884 42296
rect 21080 42236 21156 42296
rect 22304 42236 22380 42296
rect 22848 42236 22924 42296
rect 20400 41888 20612 42236
rect 20808 42160 21156 42236
rect 20808 42100 21020 42160
rect 21216 42100 21564 42236
rect 22304 42160 22924 42236
rect 23800 42236 23876 42296
rect 25568 42236 25644 42296
rect 23800 42160 25644 42236
rect 20808 42024 21564 42100
rect 20808 41964 21020 42024
rect 20808 41958 21156 41964
rect 20808 41894 21086 41958
rect 21150 41894 21156 41958
rect 20808 41888 21156 41894
rect 21216 41888 21564 42024
rect 21624 42094 21836 42100
rect 21624 42030 21766 42094
rect 21830 42030 21836 42094
rect 21624 41958 21836 42030
rect 21624 41894 21766 41958
rect 21830 41894 21836 41958
rect 21624 41888 21836 41894
rect 22032 42094 22244 42100
rect 22032 42030 22174 42094
rect 22238 42030 22244 42094
rect 22032 41958 22244 42030
rect 26928 42024 27276 42508
rect 27200 41964 27276 42024
rect 22032 41894 22038 41958
rect 22102 41894 22244 41958
rect 22032 41888 22244 41894
rect 20536 41828 20612 41888
rect 20400 41686 20612 41828
rect 26928 41752 27276 41964
rect 68952 42372 69164 42508
rect 70312 42432 71884 42508
rect 68952 42366 70252 42372
rect 68952 42302 69094 42366
rect 69158 42302 70252 42366
rect 68952 42296 70252 42302
rect 70312 42296 70524 42432
rect 71944 42372 72156 42508
rect 73032 42502 73380 42508
rect 73032 42438 73310 42502
rect 73374 42438 73380 42502
rect 73032 42432 73380 42438
rect 71944 42296 72972 42372
rect 73032 42296 73244 42432
rect 73440 42372 73652 42508
rect 73848 42502 74060 42508
rect 73848 42438 73854 42502
rect 73918 42438 74060 42502
rect 73440 42296 73788 42372
rect 73848 42366 74060 42438
rect 73848 42302 73854 42366
rect 73918 42302 74060 42366
rect 73848 42296 74060 42302
rect 74256 42502 74468 42508
rect 74256 42438 74262 42502
rect 74326 42438 74468 42502
rect 74256 42366 74468 42438
rect 74256 42302 74262 42366
rect 74326 42302 74468 42366
rect 74256 42296 74468 42302
rect 74664 42372 74876 42508
rect 74974 42502 75284 42508
rect 74936 42438 74942 42502
rect 75006 42438 75284 42502
rect 74974 42432 75284 42438
rect 74664 42366 75012 42372
rect 74664 42302 74806 42366
rect 74870 42302 75012 42366
rect 74664 42296 75012 42302
rect 75072 42366 75284 42432
rect 75072 42302 75078 42366
rect 75142 42302 75284 42366
rect 75072 42296 75284 42302
rect 75480 42296 75692 42644
rect 94112 42400 94324 42508
rect 94112 42344 94176 42400
rect 94232 42372 94324 42400
rect 94232 42366 94732 42372
rect 94232 42344 94662 42366
rect 94112 42302 94662 42344
rect 94726 42302 94732 42366
rect 94112 42296 94732 42302
rect 68952 42024 69164 42296
rect 70176 42236 70252 42296
rect 71944 42236 72020 42296
rect 70176 42160 72020 42236
rect 72896 42236 72972 42296
rect 73440 42236 73516 42296
rect 72896 42160 73516 42236
rect 73712 42236 73788 42296
rect 74664 42236 74740 42296
rect 74936 42236 75012 42296
rect 75616 42236 75692 42296
rect 73712 42160 74332 42236
rect 74256 42100 74332 42160
rect 73848 42094 74060 42100
rect 73848 42030 73854 42094
rect 73918 42030 74060 42094
rect 68952 41964 69028 42024
rect 68952 41752 69164 41964
rect 73848 41958 74060 42030
rect 73848 41894 73854 41958
rect 73918 41894 74060 41958
rect 73848 41888 74060 41894
rect 74256 42094 74468 42100
rect 74256 42030 74262 42094
rect 74326 42030 74468 42094
rect 74256 41958 74468 42030
rect 74256 41894 74262 41958
rect 74326 41894 74468 41958
rect 74256 41888 74468 41894
rect 74664 41888 74876 42236
rect 74936 42160 75284 42236
rect 75072 41964 75284 42160
rect 74974 41958 75284 41964
rect 74936 41894 74942 41958
rect 75006 41894 75284 41958
rect 74974 41888 75284 41894
rect 75480 41888 75692 42236
rect 75480 41828 75556 41888
rect 26928 41692 27004 41752
rect 69088 41692 69164 41752
rect 74800 41752 75148 41828
rect 74800 41692 74876 41752
rect 75072 41692 75148 41752
rect 20400 41622 20542 41686
rect 20606 41622 20612 41686
rect 20400 41616 20612 41622
rect 20808 41480 21020 41692
rect 21118 41686 21564 41692
rect 21080 41622 21086 41686
rect 21150 41622 21564 41686
rect 21118 41616 21564 41622
rect 21216 41480 21564 41616
rect 20808 41420 20884 41480
rect 21488 41420 21564 41480
rect 20400 41414 20612 41420
rect 20400 41350 20542 41414
rect 20606 41350 20612 41414
rect 20400 41278 20612 41350
rect 20400 41214 20542 41278
rect 20606 41214 20612 41278
rect 20400 41208 20612 41214
rect 20808 41344 21564 41420
rect 20808 41208 21020 41344
rect 21216 41278 21564 41344
rect 21216 41214 21494 41278
rect 21558 41214 21564 41278
rect 21216 41208 21564 41214
rect 21624 41686 21836 41692
rect 21624 41622 21766 41686
rect 21830 41622 21836 41686
rect 21624 41480 21836 41622
rect 22032 41686 22244 41692
rect 22032 41622 22038 41686
rect 22102 41622 22244 41686
rect 22032 41480 22244 41622
rect 21624 41420 21700 41480
rect 22032 41420 22108 41480
rect 21624 41072 21836 41420
rect 21760 41012 21836 41072
rect 20400 41006 20612 41012
rect 20400 40942 20542 41006
rect 20606 40942 20612 41006
rect 1768 40720 1980 40876
rect 20400 40870 20612 40942
rect 20400 40806 20406 40870
rect 20470 40806 20612 40870
rect 20400 40800 20612 40806
rect 20808 40876 21020 41012
rect 21216 41006 21564 41012
rect 21216 40942 21494 41006
rect 21558 40942 21564 41006
rect 21216 40876 21564 40942
rect 20808 40800 21564 40876
rect 21624 40870 21836 41012
rect 21624 40806 21766 40870
rect 21830 40806 21836 40870
rect 21624 40800 21836 40806
rect 22032 41072 22244 41420
rect 26928 41414 27276 41692
rect 26928 41350 27070 41414
rect 27134 41350 27276 41414
rect 26928 41344 27276 41350
rect 68952 41414 69164 41692
rect 68952 41350 69094 41414
rect 69158 41350 69164 41414
rect 68952 41344 69164 41350
rect 73848 41686 74060 41692
rect 73848 41622 73854 41686
rect 73918 41622 74060 41686
rect 73848 41480 74060 41622
rect 74256 41686 74468 41692
rect 74256 41622 74262 41686
rect 74326 41622 74468 41686
rect 74256 41480 74468 41622
rect 74664 41686 75012 41692
rect 74664 41622 74942 41686
rect 75006 41622 75012 41686
rect 74664 41616 75012 41622
rect 74664 41556 74876 41616
rect 74664 41480 75012 41556
rect 75072 41480 75284 41692
rect 75480 41686 75692 41828
rect 75480 41622 75622 41686
rect 75686 41622 75692 41686
rect 75480 41616 75692 41622
rect 73848 41420 73924 41480
rect 74256 41420 74332 41480
rect 74800 41420 74876 41480
rect 26928 41142 27276 41148
rect 26928 41078 27070 41142
rect 27134 41078 27276 41142
rect 22032 41012 22108 41072
rect 22032 40870 22244 41012
rect 22032 40806 22174 40870
rect 22238 40806 22244 40870
rect 22032 40800 22244 40806
rect 26928 41006 27276 41078
rect 26928 40942 27206 41006
rect 27270 40942 27276 41006
rect 26928 40800 27276 40942
rect 1768 40664 1818 40720
rect 1874 40664 1980 40720
rect 1768 40604 1980 40664
rect 20808 40740 21020 40800
rect 20808 40664 21156 40740
rect 21216 40664 21564 40800
rect 27200 40740 27276 40800
rect 26928 40734 27276 40740
rect 26928 40670 27206 40734
rect 27270 40670 27276 40734
rect 20808 40604 20884 40664
rect 21080 40604 21156 40664
rect 1224 40598 1980 40604
rect 1224 40534 1230 40598
rect 1294 40534 1980 40598
rect 1224 40528 1980 40534
rect 20400 40598 20612 40604
rect 20400 40534 20406 40598
rect 20470 40534 20612 40598
rect 20400 40462 20612 40534
rect 20400 40398 20542 40462
rect 20606 40398 20612 40462
rect 20400 40392 20612 40398
rect 20808 40392 21020 40604
rect 21080 40528 21564 40604
rect 21216 40462 21564 40528
rect 21216 40398 21222 40462
rect 21286 40398 21564 40462
rect 21216 40392 21564 40398
rect 21624 40598 21836 40604
rect 21624 40534 21766 40598
rect 21830 40534 21836 40598
rect 21624 40462 21836 40534
rect 21624 40398 21630 40462
rect 21694 40398 21836 40462
rect 21624 40392 21836 40398
rect 22032 40598 22244 40604
rect 22032 40534 22174 40598
rect 22238 40534 22244 40598
rect 22032 40462 22244 40534
rect 26928 40528 27276 40670
rect 68952 41142 69164 41148
rect 68952 41078 69094 41142
rect 69158 41078 69164 41142
rect 68952 41006 69164 41078
rect 73848 41072 74060 41420
rect 73984 41012 74060 41072
rect 68952 40942 68958 41006
rect 69022 40942 69164 41006
rect 68952 40800 69164 40942
rect 73848 40870 74060 41012
rect 73848 40806 73854 40870
rect 73918 40806 74060 40870
rect 73848 40800 74060 40806
rect 74256 41072 74468 41420
rect 74664 41208 74876 41420
rect 74936 41420 75012 41480
rect 74936 41344 75284 41420
rect 75072 41278 75284 41344
rect 75072 41214 75214 41278
rect 75278 41214 75284 41278
rect 75072 41208 75284 41214
rect 75480 41414 75692 41420
rect 75480 41350 75622 41414
rect 75686 41350 75692 41414
rect 75480 41278 75692 41350
rect 75480 41214 75622 41278
rect 75686 41214 75692 41278
rect 75480 41208 75692 41214
rect 74256 41012 74332 41072
rect 74256 40870 74468 41012
rect 74256 40806 74262 40870
rect 74326 40806 74468 40870
rect 74256 40800 74468 40806
rect 68952 40740 69028 40800
rect 68952 40734 69164 40740
rect 68952 40670 68958 40734
rect 69022 40670 69164 40734
rect 68952 40528 69164 40670
rect 74664 40664 74876 41012
rect 74800 40604 74876 40664
rect 75072 41006 75284 41012
rect 75072 40942 75214 41006
rect 75278 40942 75284 41006
rect 75072 40664 75284 40942
rect 75480 41006 75692 41012
rect 75480 40942 75622 41006
rect 75686 40942 75692 41006
rect 75480 40870 75692 40942
rect 75480 40806 75622 40870
rect 75686 40806 75692 40870
rect 75480 40800 75692 40806
rect 94112 40740 94324 40876
rect 94112 40734 94732 40740
rect 94112 40720 94662 40734
rect 94112 40664 94176 40720
rect 94232 40670 94662 40720
rect 94726 40670 94732 40734
rect 94232 40664 94732 40670
rect 75072 40604 75148 40664
rect 27064 40468 27140 40528
rect 69088 40468 69164 40528
rect 22032 40398 22174 40462
rect 22238 40398 22244 40462
rect 22032 40392 22244 40398
rect 20400 40190 20612 40196
rect 20400 40126 20542 40190
rect 20606 40126 20612 40190
rect 20400 40054 20612 40126
rect 20400 39990 20542 40054
rect 20606 39990 20612 40054
rect 20400 39984 20612 39990
rect 20808 40060 21020 40196
rect 21216 40190 21564 40196
rect 21216 40126 21222 40190
rect 21286 40126 21564 40190
rect 21216 40060 21564 40126
rect 20808 40054 21564 40060
rect 20808 39990 20950 40054
rect 21014 39990 21564 40054
rect 20808 39984 21564 39990
rect 21624 40190 21836 40196
rect 21624 40126 21630 40190
rect 21694 40126 21836 40190
rect 21624 40054 21836 40126
rect 21624 39990 21766 40054
rect 21830 39990 21836 40054
rect 21624 39984 21836 39990
rect 22032 40190 22244 40196
rect 22032 40126 22174 40190
rect 22238 40126 22244 40190
rect 22032 40054 22244 40126
rect 22032 39990 22038 40054
rect 22102 39990 22244 40054
rect 22032 39984 22244 39990
rect 26928 39984 27276 40468
rect 27200 39924 27276 39984
rect 20400 39782 20612 39788
rect 20400 39718 20542 39782
rect 20606 39718 20612 39782
rect 20400 39646 20612 39718
rect 20400 39582 20542 39646
rect 20606 39582 20612 39646
rect 20400 39576 20612 39582
rect 20808 39782 21564 39788
rect 20808 39718 20950 39782
rect 21014 39718 21564 39782
rect 20808 39712 21564 39718
rect 20808 39646 21020 39712
rect 20808 39582 20814 39646
rect 20878 39582 21020 39646
rect 20808 39576 21020 39582
rect 21216 39576 21564 39712
rect 21624 39782 21836 39788
rect 21624 39718 21766 39782
rect 21830 39718 21836 39782
rect 21624 39646 21836 39718
rect 21624 39582 21766 39646
rect 21830 39582 21836 39646
rect 21624 39576 21836 39582
rect 22032 39782 22244 39788
rect 22032 39718 22038 39782
rect 22102 39718 22244 39782
rect 22032 39646 22244 39718
rect 22032 39582 22174 39646
rect 22238 39582 22244 39646
rect 22032 39576 22244 39582
rect 26928 39712 27276 39924
rect 68952 40190 69164 40468
rect 73848 40598 74060 40604
rect 73848 40534 73854 40598
rect 73918 40534 74060 40598
rect 73848 40462 74060 40534
rect 73848 40398 73854 40462
rect 73918 40398 74060 40462
rect 73848 40392 74060 40398
rect 74256 40598 74468 40604
rect 74256 40534 74262 40598
rect 74326 40534 74468 40598
rect 74256 40462 74468 40534
rect 74256 40398 74262 40462
rect 74326 40398 74468 40462
rect 74256 40392 74468 40398
rect 74664 40528 75284 40604
rect 74664 40392 74876 40528
rect 75072 40462 75284 40528
rect 75072 40398 75214 40462
rect 75278 40398 75284 40462
rect 75072 40392 75284 40398
rect 75480 40598 75692 40604
rect 75480 40534 75622 40598
rect 75686 40534 75692 40598
rect 75480 40462 75692 40534
rect 94112 40528 94324 40664
rect 75480 40398 75622 40462
rect 75686 40398 75692 40462
rect 75480 40392 75692 40398
rect 68952 40126 69094 40190
rect 69158 40126 69164 40190
rect 68952 39984 69164 40126
rect 73848 40190 74060 40196
rect 73848 40126 73854 40190
rect 73918 40126 74060 40190
rect 73848 40054 74060 40126
rect 73848 39990 73990 40054
rect 74054 39990 74060 40054
rect 73848 39984 74060 39990
rect 74256 40190 74468 40196
rect 74256 40126 74262 40190
rect 74326 40126 74468 40190
rect 74256 40054 74468 40126
rect 74256 39990 74262 40054
rect 74326 39990 74468 40054
rect 74256 39984 74468 39990
rect 74664 40054 74876 40196
rect 74664 39990 74670 40054
rect 74734 39990 74876 40054
rect 74664 39984 74876 39990
rect 75072 40190 75284 40196
rect 75072 40126 75214 40190
rect 75278 40126 75284 40190
rect 75072 40054 75284 40126
rect 75072 39990 75214 40054
rect 75278 39990 75284 40054
rect 75072 39984 75284 39990
rect 75480 40190 75692 40196
rect 75480 40126 75622 40190
rect 75686 40126 75692 40190
rect 75480 40054 75692 40126
rect 75480 39990 75486 40054
rect 75550 39990 75692 40054
rect 75480 39984 75692 39990
rect 68952 39924 69028 39984
rect 68952 39918 69164 39924
rect 68952 39854 69094 39918
rect 69158 39854 69164 39918
rect 68952 39712 69164 39854
rect 73848 39782 74060 39788
rect 73848 39718 73990 39782
rect 74054 39718 74060 39782
rect 26928 39652 27004 39712
rect 68952 39652 69028 39712
rect 26928 39440 27276 39652
rect 68952 39440 69164 39652
rect 73848 39646 74060 39718
rect 73848 39582 73990 39646
rect 74054 39582 74060 39646
rect 73848 39576 74060 39582
rect 74256 39782 74468 39788
rect 74256 39718 74262 39782
rect 74326 39718 74468 39782
rect 74256 39646 74468 39718
rect 74256 39582 74262 39646
rect 74326 39582 74468 39646
rect 74256 39576 74468 39582
rect 74664 39782 74876 39788
rect 74664 39718 74670 39782
rect 74734 39718 74876 39782
rect 74664 39646 74876 39718
rect 75072 39782 75284 39788
rect 75072 39718 75214 39782
rect 75278 39718 75284 39782
rect 75072 39652 75284 39718
rect 74974 39646 75284 39652
rect 74664 39582 74670 39646
rect 74734 39582 74876 39646
rect 74936 39582 74942 39646
rect 75006 39582 75214 39646
rect 75278 39582 75284 39646
rect 74664 39576 74876 39582
rect 74974 39576 75284 39582
rect 75480 39782 75692 39788
rect 75480 39718 75486 39782
rect 75550 39718 75692 39782
rect 75480 39646 75692 39718
rect 75480 39582 75622 39646
rect 75686 39582 75692 39646
rect 75480 39576 75692 39582
rect 27064 39380 27140 39440
rect 69088 39380 69164 39440
rect 20400 39374 20612 39380
rect 20400 39310 20542 39374
rect 20606 39310 20612 39374
rect 20400 39238 20612 39310
rect 20400 39174 20406 39238
rect 20470 39174 20612 39238
rect 20400 39168 20612 39174
rect 20808 39374 21020 39380
rect 20808 39310 20814 39374
rect 20878 39310 21020 39374
rect 20808 39238 21020 39310
rect 21216 39244 21564 39380
rect 21118 39238 21564 39244
rect 20808 39174 20814 39238
rect 20878 39174 21020 39238
rect 21080 39174 21086 39238
rect 21150 39174 21564 39238
rect 20808 39168 21020 39174
rect 21118 39168 21564 39174
rect 21624 39374 21836 39380
rect 21624 39310 21766 39374
rect 21830 39310 21836 39374
rect 21624 39238 21836 39310
rect 21624 39174 21630 39238
rect 21694 39174 21836 39238
rect 21624 39168 21836 39174
rect 22032 39374 22244 39380
rect 22032 39310 22174 39374
rect 22238 39310 22244 39374
rect 22032 39238 22244 39310
rect 22032 39174 22038 39238
rect 22102 39174 22244 39238
rect 22032 39168 22244 39174
rect 26928 39168 27276 39380
rect 68952 39168 69164 39380
rect 73848 39374 74060 39380
rect 73848 39310 73990 39374
rect 74054 39310 74060 39374
rect 73848 39238 74060 39310
rect 73848 39174 73990 39238
rect 74054 39174 74060 39238
rect 73848 39168 74060 39174
rect 74256 39374 74468 39380
rect 74256 39310 74262 39374
rect 74326 39310 74468 39374
rect 74256 39238 74468 39310
rect 74256 39174 74262 39238
rect 74326 39174 74468 39238
rect 74256 39168 74468 39174
rect 74664 39374 75012 39380
rect 74664 39310 74670 39374
rect 74734 39310 74942 39374
rect 75006 39310 75012 39374
rect 74664 39304 75012 39310
rect 75072 39374 75284 39380
rect 75072 39310 75214 39374
rect 75278 39310 75284 39374
rect 74664 39168 74876 39304
rect 75072 39238 75284 39310
rect 75072 39174 75078 39238
rect 75142 39174 75284 39238
rect 75072 39168 75284 39174
rect 75480 39374 75692 39380
rect 75480 39310 75622 39374
rect 75686 39310 75692 39374
rect 75480 39238 75692 39310
rect 75480 39174 75622 39238
rect 75686 39174 75692 39238
rect 75480 39168 75692 39174
rect 26928 39108 27004 39168
rect 69088 39108 69164 39168
rect 1768 39040 1980 39108
rect 1768 38984 1818 39040
rect 1874 38984 1980 39040
rect 1768 38972 1980 38984
rect 1224 38966 1980 38972
rect 1224 38902 1230 38966
rect 1294 38902 1980 38966
rect 1224 38896 1980 38902
rect 20400 38966 20612 38972
rect 20400 38902 20406 38966
rect 20470 38902 20612 38966
rect 20400 38760 20612 38902
rect 20808 38966 21156 38972
rect 20808 38902 20814 38966
rect 20878 38902 21086 38966
rect 21150 38902 21156 38966
rect 20808 38896 21156 38902
rect 20808 38836 21020 38896
rect 21216 38836 21564 38972
rect 20808 38830 21564 38836
rect 20808 38766 21494 38830
rect 21558 38766 21564 38830
rect 20808 38760 21564 38766
rect 21624 38966 21836 38972
rect 21624 38902 21630 38966
rect 21694 38902 21836 38966
rect 21624 38830 21836 38902
rect 21624 38766 21766 38830
rect 21830 38766 21836 38830
rect 21624 38760 21836 38766
rect 22032 38966 22244 38972
rect 22032 38902 22038 38966
rect 22102 38902 22244 38966
rect 22032 38830 22244 38902
rect 26928 38896 27276 39108
rect 27200 38836 27276 38896
rect 22032 38766 22174 38830
rect 22238 38766 22244 38830
rect 22032 38760 22244 38766
rect 20400 38700 20476 38760
rect 20400 38352 20612 38700
rect 26928 38624 27276 38836
rect 68952 38896 69164 39108
rect 94112 39040 94324 39108
rect 94112 38984 94176 39040
rect 94232 38984 94324 39040
rect 94112 38972 94324 38984
rect 73848 38966 74060 38972
rect 73848 38902 73990 38966
rect 74054 38902 74060 38966
rect 68952 38836 69028 38896
rect 68952 38624 69164 38836
rect 73848 38830 74060 38902
rect 73848 38766 73990 38830
rect 74054 38766 74060 38830
rect 73848 38760 74060 38766
rect 74256 38966 74468 38972
rect 74256 38902 74262 38966
rect 74326 38902 74468 38966
rect 74256 38830 74468 38902
rect 74256 38766 74398 38830
rect 74462 38766 74468 38830
rect 74256 38760 74468 38766
rect 74664 38830 74876 38972
rect 74664 38766 74670 38830
rect 74734 38766 74876 38830
rect 74664 38760 74876 38766
rect 75072 38966 75284 38972
rect 75072 38902 75078 38966
rect 75142 38902 75284 38966
rect 75072 38830 75284 38902
rect 75072 38766 75078 38830
rect 75142 38766 75284 38830
rect 75072 38760 75284 38766
rect 75480 38966 75692 38972
rect 75480 38902 75622 38966
rect 75686 38902 75692 38966
rect 75480 38760 75692 38902
rect 94112 38966 94732 38972
rect 94112 38902 94662 38966
rect 94726 38902 94732 38966
rect 94112 38896 94732 38902
rect 75480 38700 75556 38760
rect 27064 38564 27140 38624
rect 68952 38564 69028 38624
rect 20536 38292 20612 38352
rect 20400 37944 20612 38292
rect 20808 38352 21020 38564
rect 21216 38558 21564 38564
rect 21216 38494 21494 38558
rect 21558 38494 21564 38558
rect 21216 38352 21564 38494
rect 21624 38558 21836 38564
rect 21624 38494 21766 38558
rect 21830 38494 21836 38558
rect 21624 38422 21836 38494
rect 21624 38358 21630 38422
rect 21694 38358 21836 38422
rect 21624 38352 21836 38358
rect 22032 38558 22244 38564
rect 22032 38494 22174 38558
rect 22238 38494 22244 38558
rect 22032 38422 22244 38494
rect 22032 38358 22174 38422
rect 22238 38358 22244 38422
rect 22032 38352 22244 38358
rect 26928 38352 27276 38564
rect 20808 38292 20884 38352
rect 21216 38292 21292 38352
rect 20808 38156 21020 38292
rect 21216 38156 21564 38292
rect 27054 38156 27152 38352
rect 20808 38080 21564 38156
rect 20808 37944 21020 38080
rect 21216 38020 21564 38080
rect 21118 38014 21564 38020
rect 21080 37950 21086 38014
rect 21150 37950 21564 38014
rect 21118 37944 21564 37950
rect 21624 38150 21836 38156
rect 21624 38086 21630 38150
rect 21694 38086 21836 38150
rect 21624 38014 21836 38086
rect 21624 37950 21630 38014
rect 21694 37950 21836 38014
rect 21624 37944 21836 37950
rect 22032 38150 22244 38156
rect 22032 38086 22174 38150
rect 22238 38086 22244 38150
rect 22032 38014 22244 38086
rect 26928 38080 27276 38156
rect 68952 38080 69164 38564
rect 73848 38558 74060 38564
rect 73848 38494 73990 38558
rect 74054 38494 74060 38558
rect 73848 38422 74060 38494
rect 73848 38358 73854 38422
rect 73918 38358 74060 38422
rect 73848 38352 74060 38358
rect 74256 38558 74468 38564
rect 74256 38494 74398 38558
rect 74462 38494 74468 38558
rect 74256 38422 74468 38494
rect 74256 38358 74262 38422
rect 74326 38358 74468 38422
rect 74256 38352 74468 38358
rect 74664 38558 74876 38564
rect 74664 38494 74670 38558
rect 74734 38494 74876 38558
rect 74664 38352 74876 38494
rect 75072 38558 75284 38564
rect 75072 38494 75078 38558
rect 75142 38494 75284 38558
rect 75072 38428 75284 38494
rect 74800 38292 74876 38352
rect 74936 38352 75284 38428
rect 75480 38352 75692 38700
rect 74936 38292 75012 38352
rect 75480 38292 75556 38352
rect 74664 38216 75012 38292
rect 27064 38020 27140 38080
rect 69088 38020 69164 38080
rect 22032 37950 22174 38014
rect 22238 37950 22244 38014
rect 22032 37944 22244 37950
rect 20400 37884 20476 37944
rect 20400 37742 20612 37884
rect 26928 37878 27276 38020
rect 26928 37814 26934 37878
rect 26998 37814 27276 37878
rect 26928 37808 27276 37814
rect 27200 37748 27276 37808
rect 20400 37678 20542 37742
rect 20606 37678 20612 37742
rect 20400 37672 20612 37678
rect 20808 37742 21156 37748
rect 20808 37678 21086 37742
rect 21150 37678 21156 37742
rect 20808 37672 21156 37678
rect 20808 37612 21020 37672
rect 20808 37536 21156 37612
rect 21216 37536 21564 37748
rect 21624 37742 21836 37748
rect 21624 37678 21630 37742
rect 21694 37678 21836 37742
rect 21624 37536 21836 37678
rect 22032 37742 22244 37748
rect 22032 37678 22174 37742
rect 22238 37678 22244 37742
rect 22032 37536 22244 37678
rect 20944 37476 21020 37536
rect 1224 37470 1980 37476
rect 1224 37406 1230 37470
rect 1294 37406 1980 37470
rect 1224 37400 1980 37406
rect 1768 37360 1980 37400
rect 1768 37304 1818 37360
rect 1874 37304 1980 37360
rect 1768 37264 1980 37304
rect 20400 37470 20612 37476
rect 20400 37406 20542 37470
rect 20606 37406 20612 37470
rect 20400 37334 20612 37406
rect 20400 37270 20406 37334
rect 20470 37270 20612 37334
rect 20400 37264 20612 37270
rect 20808 37334 21020 37476
rect 21080 37476 21156 37536
rect 21352 37476 21428 37536
rect 21760 37476 21836 37536
rect 22168 37476 22244 37536
rect 21080 37400 21564 37476
rect 20808 37270 20814 37334
rect 20878 37270 21020 37334
rect 20808 37264 21020 37270
rect 21216 37264 21564 37400
rect 21624 37128 21836 37476
rect 22032 37128 22244 37476
rect 26928 37606 27276 37748
rect 26928 37542 26934 37606
rect 26998 37542 27276 37606
rect 26928 37470 27276 37542
rect 26928 37406 27070 37470
rect 27134 37406 27276 37470
rect 26928 37400 27276 37406
rect 68952 37808 69164 38020
rect 73848 38150 74060 38156
rect 73848 38086 73854 38150
rect 73918 38086 74060 38150
rect 73848 38014 74060 38086
rect 73848 37950 73990 38014
rect 74054 37950 74060 38014
rect 73848 37944 74060 37950
rect 74256 38150 74468 38156
rect 74256 38086 74262 38150
rect 74326 38086 74468 38150
rect 74256 38014 74468 38086
rect 74256 37950 74398 38014
rect 74462 37950 74468 38014
rect 74256 37944 74468 37950
rect 74664 38020 74876 38216
rect 75072 38020 75284 38292
rect 74664 38014 75284 38020
rect 74664 37950 74670 38014
rect 74734 37950 75284 38014
rect 74664 37944 75284 37950
rect 75480 37944 75692 38292
rect 75616 37884 75692 37944
rect 68952 37748 69028 37808
rect 68952 37470 69164 37748
rect 73848 37742 74060 37748
rect 73848 37678 73990 37742
rect 74054 37678 74060 37742
rect 73848 37536 74060 37678
rect 74256 37742 74468 37748
rect 74256 37678 74398 37742
rect 74462 37678 74468 37742
rect 74256 37536 74468 37678
rect 73984 37476 74060 37536
rect 74392 37476 74468 37536
rect 68952 37406 68958 37470
rect 69022 37406 69164 37470
rect 68952 37400 69164 37406
rect 21760 37068 21836 37128
rect 22168 37068 22244 37128
rect 20400 37062 20612 37068
rect 20400 36998 20406 37062
rect 20470 36998 20612 37062
rect 20400 36926 20612 36998
rect 20400 36862 20542 36926
rect 20606 36862 20612 36926
rect 20400 36856 20612 36862
rect 20808 37062 21020 37068
rect 20808 36998 20814 37062
rect 20878 36998 21020 37062
rect 20808 36720 21020 36998
rect 21216 36720 21564 37068
rect 21624 36720 21836 37068
rect 22032 36720 22244 37068
rect 20808 36660 20884 36720
rect 21488 36660 21564 36720
rect 21760 36660 21836 36720
rect 22168 36660 22244 36720
rect 20400 36654 20612 36660
rect 20400 36590 20542 36654
rect 20606 36590 20612 36654
rect 20400 36518 20612 36590
rect 20400 36454 20406 36518
rect 20470 36454 20612 36518
rect 20400 36448 20612 36454
rect 20808 36584 21564 36660
rect 20808 36448 21020 36584
rect 21216 36518 21564 36584
rect 21216 36454 21358 36518
rect 21422 36454 21564 36518
rect 21216 36448 21564 36454
rect 21624 36518 21836 36660
rect 21624 36454 21630 36518
rect 21694 36454 21836 36518
rect 21624 36448 21836 36454
rect 22032 36518 22244 36660
rect 26928 37198 27276 37204
rect 26928 37134 27070 37198
rect 27134 37134 27276 37198
rect 26928 36584 27276 37134
rect 27200 36524 27276 36584
rect 22032 36454 22038 36518
rect 22102 36454 22244 36518
rect 22032 36448 22244 36454
rect 20400 36246 20612 36252
rect 20400 36182 20406 36246
rect 20470 36182 20612 36246
rect 20400 36110 20612 36182
rect 20400 36046 20406 36110
rect 20470 36046 20612 36110
rect 20400 36040 20612 36046
rect 20808 36110 21020 36252
rect 20808 36046 20814 36110
rect 20878 36046 21020 36110
rect 20808 36040 21020 36046
rect 21216 36246 21564 36252
rect 21216 36182 21358 36246
rect 21422 36182 21564 36246
rect 21216 36110 21564 36182
rect 21216 36046 21222 36110
rect 21286 36046 21564 36110
rect 21216 36040 21564 36046
rect 21624 36246 21836 36252
rect 21624 36182 21630 36246
rect 21694 36182 21836 36246
rect 21624 36110 21836 36182
rect 21624 36046 21630 36110
rect 21694 36046 21836 36110
rect 21624 36040 21836 36046
rect 22032 36246 22244 36252
rect 22032 36182 22038 36246
rect 22102 36182 22244 36246
rect 22032 36110 22244 36182
rect 22032 36046 22174 36110
rect 22238 36046 22244 36110
rect 22032 36040 22244 36046
rect 26928 36040 27276 36524
rect 68952 37198 69164 37204
rect 68952 37134 68958 37198
rect 69022 37134 69164 37198
rect 68952 37062 69164 37134
rect 68952 36998 68958 37062
rect 69022 36998 69164 37062
rect 68952 36790 69164 36998
rect 68952 36726 68958 36790
rect 69022 36726 69164 36790
rect 68952 36584 69164 36726
rect 73848 37128 74060 37476
rect 74256 37128 74468 37476
rect 74664 37742 74876 37748
rect 74664 37678 74670 37742
rect 74734 37678 74876 37742
rect 74664 37536 74876 37678
rect 75072 37536 75284 37748
rect 75480 37742 75692 37884
rect 75480 37678 75486 37742
rect 75550 37678 75692 37742
rect 75480 37672 75692 37678
rect 74664 37476 74740 37536
rect 75072 37476 75148 37536
rect 74664 37334 74876 37476
rect 75072 37340 75284 37476
rect 74974 37334 75284 37340
rect 74664 37270 74670 37334
rect 74734 37270 74876 37334
rect 74936 37270 74942 37334
rect 75006 37270 75284 37334
rect 74664 37264 74876 37270
rect 74974 37264 75284 37270
rect 75480 37470 75692 37476
rect 75480 37406 75486 37470
rect 75550 37406 75692 37470
rect 75480 37334 75692 37406
rect 75480 37270 75622 37334
rect 75686 37270 75692 37334
rect 75480 37264 75692 37270
rect 94112 37470 94732 37476
rect 94112 37406 94662 37470
rect 94726 37406 94732 37470
rect 94112 37400 94732 37406
rect 94112 37360 94324 37400
rect 94112 37304 94176 37360
rect 94232 37304 94324 37360
rect 94112 37264 94324 37304
rect 73848 37068 73924 37128
rect 74392 37068 74468 37128
rect 73848 36720 74060 37068
rect 73984 36660 74060 36720
rect 68952 36524 69028 36584
rect 68952 36246 69164 36524
rect 73848 36518 74060 36660
rect 73848 36454 73854 36518
rect 73918 36454 74060 36518
rect 73848 36448 74060 36454
rect 74256 36720 74468 37068
rect 74664 37062 75012 37068
rect 74664 36998 74670 37062
rect 74734 36998 74942 37062
rect 75006 36998 75012 37062
rect 74664 36992 75012 36998
rect 74664 36932 74876 36992
rect 75072 36932 75284 37068
rect 74664 36856 75284 36932
rect 75480 37062 75692 37068
rect 75480 36998 75622 37062
rect 75686 36998 75692 37062
rect 75480 36926 75692 36998
rect 75480 36862 75622 36926
rect 75686 36862 75692 36926
rect 75480 36856 75692 36862
rect 74664 36720 74876 36856
rect 75072 36720 75284 36856
rect 74256 36660 74332 36720
rect 74664 36660 74740 36720
rect 75072 36660 75148 36720
rect 74256 36518 74468 36660
rect 74256 36454 74262 36518
rect 74326 36454 74468 36518
rect 74256 36448 74468 36454
rect 74664 36448 74876 36660
rect 75072 36524 75284 36660
rect 74974 36518 75284 36524
rect 74936 36454 74942 36518
rect 75006 36454 75078 36518
rect 75142 36454 75284 36518
rect 74974 36448 75284 36454
rect 75480 36654 75692 36660
rect 75480 36590 75622 36654
rect 75686 36590 75692 36654
rect 75480 36518 75692 36590
rect 75480 36454 75622 36518
rect 75686 36454 75692 36518
rect 75480 36448 75692 36454
rect 68952 36182 69094 36246
rect 69158 36182 69164 36246
rect 68952 36040 69164 36182
rect 73848 36246 74060 36252
rect 73848 36182 73854 36246
rect 73918 36182 74060 36246
rect 73848 36110 74060 36182
rect 73848 36046 73854 36110
rect 73918 36046 74060 36110
rect 73848 36040 74060 36046
rect 74256 36246 74468 36252
rect 74256 36182 74262 36246
rect 74326 36182 74468 36246
rect 74256 36110 74468 36182
rect 74256 36046 74398 36110
rect 74462 36046 74468 36110
rect 74256 36040 74468 36046
rect 74664 36246 75012 36252
rect 74664 36182 74942 36246
rect 75006 36182 75012 36246
rect 74664 36176 75012 36182
rect 75072 36246 75284 36252
rect 75072 36182 75078 36246
rect 75142 36182 75284 36246
rect 74664 36040 74876 36176
rect 75072 36110 75284 36182
rect 75072 36046 75078 36110
rect 75142 36046 75284 36110
rect 75072 36040 75284 36046
rect 75480 36246 75692 36252
rect 75480 36182 75622 36246
rect 75686 36182 75692 36246
rect 75480 36110 75692 36182
rect 75480 36046 75622 36110
rect 75686 36046 75692 36110
rect 75480 36040 75692 36046
rect 27064 35980 27140 36040
rect 69088 35980 69164 36040
rect 20400 35838 20612 35844
rect 20400 35774 20406 35838
rect 20470 35774 20612 35838
rect 1768 35680 1980 35708
rect 1768 35624 1818 35680
rect 1874 35624 1980 35680
rect 20400 35702 20612 35774
rect 20400 35638 20542 35702
rect 20606 35638 20612 35702
rect 20400 35632 20612 35638
rect 20808 35838 21020 35844
rect 20808 35774 20814 35838
rect 20878 35774 21020 35838
rect 20808 35708 21020 35774
rect 21216 35838 21564 35844
rect 21216 35774 21222 35838
rect 21286 35774 21564 35838
rect 21216 35708 21564 35774
rect 20808 35702 21564 35708
rect 20808 35638 20950 35702
rect 21014 35638 21564 35702
rect 20808 35632 21564 35638
rect 21624 35838 21836 35844
rect 21624 35774 21630 35838
rect 21694 35774 21836 35838
rect 21624 35702 21836 35774
rect 21624 35638 21766 35702
rect 21830 35638 21836 35702
rect 21624 35632 21836 35638
rect 22032 35838 22244 35844
rect 22032 35774 22174 35838
rect 22238 35774 22244 35838
rect 22032 35702 22244 35774
rect 26928 35768 27276 35980
rect 68952 35974 69164 35980
rect 68952 35910 69094 35974
rect 69158 35910 69164 35974
rect 68952 35768 69164 35910
rect 27200 35708 27276 35768
rect 69088 35708 69164 35768
rect 22032 35638 22038 35702
rect 22102 35638 22244 35702
rect 22032 35632 22244 35638
rect 1768 35572 1980 35624
rect 1224 35566 1980 35572
rect 1224 35502 1230 35566
rect 1294 35502 1980 35566
rect 1224 35496 1980 35502
rect 20944 35572 21020 35632
rect 20944 35496 21292 35572
rect 26928 35496 27276 35708
rect 68952 35496 69164 35708
rect 73848 35838 74060 35844
rect 73848 35774 73854 35838
rect 73918 35774 74060 35838
rect 73848 35702 74060 35774
rect 73848 35638 73990 35702
rect 74054 35638 74060 35702
rect 73848 35632 74060 35638
rect 74256 35838 74468 35844
rect 74256 35774 74398 35838
rect 74462 35774 74468 35838
rect 74256 35702 74468 35774
rect 74256 35638 74262 35702
rect 74326 35638 74468 35702
rect 74256 35632 74468 35638
rect 74664 35702 74876 35844
rect 74664 35638 74670 35702
rect 74734 35638 74876 35702
rect 74664 35632 74876 35638
rect 75072 35838 75284 35844
rect 75072 35774 75078 35838
rect 75142 35774 75284 35838
rect 75072 35702 75284 35774
rect 75072 35638 75078 35702
rect 75142 35638 75284 35702
rect 75072 35632 75284 35638
rect 75480 35838 75692 35844
rect 75480 35774 75622 35838
rect 75686 35774 75692 35838
rect 75480 35702 75692 35774
rect 75480 35638 75486 35702
rect 75550 35638 75692 35702
rect 75480 35632 75692 35638
rect 94112 35680 94324 35708
rect 94112 35624 94176 35680
rect 94232 35624 94324 35680
rect 94112 35572 94324 35624
rect 94112 35566 94732 35572
rect 94112 35502 94662 35566
rect 94726 35502 94732 35566
rect 94112 35496 94732 35502
rect 21216 35436 21292 35496
rect 27064 35436 27140 35496
rect 68952 35436 69028 35496
rect 20400 35430 20612 35436
rect 20400 35366 20542 35430
rect 20606 35366 20612 35430
rect 20400 35294 20612 35366
rect 20400 35230 20406 35294
rect 20470 35230 20612 35294
rect 20400 35224 20612 35230
rect 20808 35430 21020 35436
rect 20808 35366 20950 35430
rect 21014 35366 21020 35430
rect 20808 35294 21020 35366
rect 20808 35230 20814 35294
rect 20878 35230 21020 35294
rect 20808 35224 21020 35230
rect 21216 35224 21564 35436
rect 21624 35430 21836 35436
rect 21624 35366 21766 35430
rect 21830 35366 21836 35430
rect 21624 35294 21836 35366
rect 21624 35230 21766 35294
rect 21830 35230 21836 35294
rect 21624 35224 21836 35230
rect 22032 35430 22244 35436
rect 22032 35366 22038 35430
rect 22102 35366 22244 35430
rect 22032 35294 22244 35366
rect 22032 35230 22038 35294
rect 22102 35230 22244 35294
rect 22032 35224 22244 35230
rect 26928 35224 27276 35436
rect 27200 35164 27276 35224
rect 13600 34886 13812 35028
rect 13600 34822 13742 34886
rect 13806 34822 13812 34886
rect 13600 34816 13812 34822
rect 20400 35022 20612 35028
rect 20400 34958 20406 35022
rect 20470 34958 20612 35022
rect 20400 34816 20612 34958
rect 20808 35022 21020 35028
rect 20808 34958 20814 35022
rect 20878 34958 21020 35022
rect 20808 34886 21020 34958
rect 21216 34892 21564 35028
rect 21118 34886 21564 34892
rect 20808 34822 20950 34886
rect 21014 34822 21020 34886
rect 21080 34822 21086 34886
rect 21150 34822 21564 34886
rect 20808 34816 21020 34822
rect 21118 34816 21564 34822
rect 21624 35022 21836 35028
rect 21624 34958 21766 35022
rect 21830 34958 21836 35022
rect 21624 34886 21836 34958
rect 21624 34822 21766 34886
rect 21830 34822 21836 34886
rect 21624 34816 21836 34822
rect 22032 35022 22244 35028
rect 22032 34958 22038 35022
rect 22102 34958 22244 35022
rect 22032 34886 22244 34958
rect 26928 34952 27276 35164
rect 68952 35224 69164 35436
rect 73848 35430 74060 35436
rect 73848 35366 73990 35430
rect 74054 35366 74060 35430
rect 73848 35294 74060 35366
rect 73848 35230 73990 35294
rect 74054 35230 74060 35294
rect 73848 35224 74060 35230
rect 74256 35430 74468 35436
rect 74256 35366 74262 35430
rect 74326 35366 74468 35430
rect 74256 35294 74468 35366
rect 74256 35230 74262 35294
rect 74326 35230 74468 35294
rect 74256 35224 74468 35230
rect 74664 35430 74876 35436
rect 74664 35366 74670 35430
rect 74734 35366 74876 35430
rect 74664 35294 74876 35366
rect 75072 35430 75284 35436
rect 75072 35366 75078 35430
rect 75142 35366 75284 35430
rect 75072 35300 75284 35366
rect 74974 35294 75284 35300
rect 74664 35230 74806 35294
rect 74870 35230 74876 35294
rect 74936 35230 74942 35294
rect 75006 35230 75284 35294
rect 74664 35224 74876 35230
rect 74974 35224 75284 35230
rect 75480 35430 75692 35436
rect 75480 35366 75486 35430
rect 75550 35366 75692 35430
rect 75480 35294 75692 35366
rect 75480 35230 75622 35294
rect 75686 35230 75692 35294
rect 75480 35224 75692 35230
rect 68952 35164 69028 35224
rect 68952 34952 69164 35164
rect 27064 34892 27140 34952
rect 69088 34892 69164 34952
rect 22032 34822 22038 34886
rect 22102 34822 22244 34886
rect 22032 34816 22244 34822
rect 20536 34756 20612 34816
rect 20400 34478 20612 34756
rect 26928 34680 27276 34892
rect 27200 34620 27276 34680
rect 20400 34414 20542 34478
rect 20606 34414 20612 34478
rect 20400 34408 20612 34414
rect 20808 34614 21156 34620
rect 20808 34550 20950 34614
rect 21014 34550 21086 34614
rect 21150 34550 21156 34614
rect 20808 34544 21156 34550
rect 20808 34484 21020 34544
rect 21216 34484 21564 34620
rect 20808 34478 21564 34484
rect 20808 34414 21494 34478
rect 21558 34414 21564 34478
rect 20808 34408 21564 34414
rect 21624 34614 21836 34620
rect 21624 34550 21766 34614
rect 21830 34550 21836 34614
rect 21624 34478 21836 34550
rect 21624 34414 21766 34478
rect 21830 34414 21836 34478
rect 21624 34408 21836 34414
rect 22032 34614 22244 34620
rect 22032 34550 22038 34614
rect 22102 34550 22244 34614
rect 22032 34478 22244 34550
rect 22032 34414 22038 34478
rect 22102 34414 22244 34478
rect 22032 34408 22244 34414
rect 26928 34408 27276 34620
rect 68952 34680 69164 34892
rect 73848 35022 74060 35028
rect 73848 34958 73990 35022
rect 74054 34958 74060 35022
rect 73848 34886 74060 34958
rect 73848 34822 73990 34886
rect 74054 34822 74060 34886
rect 73848 34816 74060 34822
rect 74256 35022 74468 35028
rect 74256 34958 74262 35022
rect 74326 34958 74468 35022
rect 74256 34886 74468 34958
rect 74256 34822 74262 34886
rect 74326 34822 74468 34886
rect 74256 34816 74468 34822
rect 74664 35022 75012 35028
rect 74664 34958 74806 35022
rect 74870 34958 74942 35022
rect 75006 34958 75012 35022
rect 74664 34952 75012 34958
rect 74664 34892 74876 34952
rect 75072 34892 75284 35028
rect 74664 34886 75284 34892
rect 74664 34822 75078 34886
rect 75142 34822 75284 34886
rect 74664 34816 75284 34822
rect 75480 35022 75692 35028
rect 75480 34958 75622 35022
rect 75686 34958 75692 35022
rect 75480 34816 75692 34958
rect 75616 34756 75692 34816
rect 68952 34620 69028 34680
rect 68952 34408 69164 34620
rect 73848 34614 74060 34620
rect 73848 34550 73990 34614
rect 74054 34550 74060 34614
rect 73848 34478 74060 34550
rect 73848 34414 73990 34478
rect 74054 34414 74060 34478
rect 73848 34408 74060 34414
rect 74256 34614 74468 34620
rect 74256 34550 74262 34614
rect 74326 34550 74468 34614
rect 74256 34478 74468 34550
rect 74256 34414 74398 34478
rect 74462 34414 74468 34478
rect 74256 34408 74468 34414
rect 74664 34478 74876 34620
rect 74664 34414 74670 34478
rect 74734 34414 74876 34478
rect 74664 34408 74876 34414
rect 75072 34614 75284 34620
rect 75072 34550 75078 34614
rect 75142 34550 75284 34614
rect 75072 34478 75284 34550
rect 75072 34414 75214 34478
rect 75278 34414 75284 34478
rect 75072 34408 75284 34414
rect 75480 34478 75692 34756
rect 75480 34414 75486 34478
rect 75550 34414 75692 34478
rect 75480 34408 75692 34414
rect 27064 34348 27140 34408
rect 68952 34348 69028 34408
rect 0 34136 13404 34212
rect 20400 34206 20612 34212
rect 14200 34199 14266 34202
rect 14934 34199 15000 34202
rect 14200 34197 15000 34199
rect 14200 34141 14205 34197
rect 14261 34141 14939 34197
rect 14995 34141 15000 34197
rect 14200 34139 15000 34141
rect 14200 34136 14266 34139
rect 14934 34136 15000 34139
rect 20400 34142 20542 34206
rect 20606 34142 20612 34206
rect 13192 34126 13404 34136
rect 1768 34000 1980 34076
rect 13192 34070 13260 34126
rect 13316 34070 13404 34126
rect 13192 34000 13404 34070
rect 20400 34000 20612 34142
rect 20808 34206 21564 34212
rect 20808 34142 21494 34206
rect 21558 34142 21564 34206
rect 20808 34136 21564 34142
rect 20808 34000 21020 34136
rect 21216 34070 21564 34136
rect 21216 34006 21358 34070
rect 21422 34006 21564 34070
rect 21216 34000 21564 34006
rect 21624 34206 21836 34212
rect 21624 34142 21766 34206
rect 21830 34142 21836 34206
rect 21624 34070 21836 34142
rect 21624 34006 21630 34070
rect 21694 34006 21836 34070
rect 21624 34000 21836 34006
rect 22032 34206 22244 34212
rect 22032 34142 22038 34206
rect 22102 34142 22244 34206
rect 22032 34070 22244 34142
rect 26928 34136 27276 34348
rect 68952 34136 69164 34348
rect 73848 34206 74060 34212
rect 73848 34142 73990 34206
rect 74054 34142 74060 34206
rect 27064 34076 27140 34136
rect 68952 34076 69028 34136
rect 22032 34006 22174 34070
rect 22238 34006 22244 34070
rect 22032 34000 22244 34006
rect 1768 33944 1818 34000
rect 1874 33944 1980 34000
rect 1768 33940 1980 33944
rect 1224 33934 1980 33940
rect 1224 33870 1230 33934
rect 1294 33870 1980 33934
rect 1224 33864 1980 33870
rect 20400 33940 20476 34000
rect 20400 33798 20612 33940
rect 26928 33864 27276 34076
rect 68952 33864 69164 34076
rect 73848 34070 74060 34142
rect 73848 34006 73854 34070
rect 73918 34006 74060 34070
rect 73848 34000 74060 34006
rect 74256 34206 74468 34212
rect 74256 34142 74398 34206
rect 74462 34142 74468 34206
rect 74256 34070 74468 34142
rect 74256 34006 74262 34070
rect 74326 34006 74468 34070
rect 74256 34000 74468 34006
rect 74664 34206 74876 34212
rect 74664 34142 74670 34206
rect 74734 34142 74876 34206
rect 74664 34070 74876 34142
rect 75072 34206 75284 34212
rect 75072 34142 75214 34206
rect 75278 34142 75284 34206
rect 75072 34076 75284 34142
rect 74974 34070 75284 34076
rect 74664 34006 74806 34070
rect 74870 34006 74876 34070
rect 74936 34006 74942 34070
rect 75006 34006 75284 34070
rect 74664 34000 74876 34006
rect 74974 34000 75284 34006
rect 75480 34206 75692 34212
rect 75480 34142 75486 34206
rect 75550 34142 75692 34206
rect 75480 34000 75692 34142
rect 75616 33940 75692 34000
rect 27064 33804 27140 33864
rect 69088 33804 69164 33864
rect 20400 33734 20406 33798
rect 20470 33734 20612 33798
rect 20400 33728 20612 33734
rect 13600 33526 13812 33668
rect 20808 33592 21020 33804
rect 21216 33798 21564 33804
rect 21216 33734 21358 33798
rect 21422 33734 21564 33798
rect 21216 33592 21564 33734
rect 21624 33798 21836 33804
rect 21624 33734 21630 33798
rect 21694 33734 21836 33798
rect 21624 33662 21836 33734
rect 21624 33598 21766 33662
rect 21830 33598 21836 33662
rect 21624 33592 21836 33598
rect 22032 33798 22244 33804
rect 22032 33734 22174 33798
rect 22238 33734 22244 33798
rect 22032 33662 22244 33734
rect 22032 33598 22174 33662
rect 22238 33598 22244 33662
rect 22032 33592 22244 33598
rect 20808 33532 20884 33592
rect 21216 33532 21292 33592
rect 13600 33462 13606 33526
rect 13670 33462 13812 33526
rect 13600 33456 13812 33462
rect 20400 33526 20612 33532
rect 20400 33462 20406 33526
rect 20470 33462 20612 33526
rect 20400 33184 20612 33462
rect 20808 33260 21020 33532
rect 21216 33260 21564 33532
rect 20808 33184 21564 33260
rect 21624 33390 21836 33396
rect 21624 33326 21766 33390
rect 21830 33326 21836 33390
rect 21624 33184 21836 33326
rect 22032 33390 22244 33396
rect 22032 33326 22174 33390
rect 22238 33326 22244 33390
rect 22032 33184 22244 33326
rect 26928 33320 27276 33804
rect 27200 33260 27276 33320
rect 20536 33124 20612 33184
rect 13192 32998 13404 33124
rect 13192 32988 13260 32998
rect 0 32942 13260 32988
rect 13316 32942 13404 32998
rect 0 32912 13404 32942
rect 20400 32982 20612 33124
rect 20944 33124 21020 33184
rect 21760 33124 21836 33184
rect 22168 33124 22244 33184
rect 20944 33048 21292 33124
rect 21216 32988 21292 33048
rect 14200 32929 14266 32932
rect 14854 32929 14920 32932
rect 14200 32927 14920 32929
rect 14200 32871 14205 32927
rect 14261 32871 14859 32927
rect 14915 32871 14920 32927
rect 20400 32918 20542 32982
rect 20606 32918 20612 32982
rect 20400 32912 20612 32918
rect 14200 32869 14920 32871
rect 14200 32866 14266 32869
rect 14854 32866 14920 32869
rect 20808 32776 21020 32988
rect 21216 32776 21564 32988
rect 20808 32716 20884 32776
rect 21488 32716 21564 32776
rect 20400 32710 20612 32716
rect 20400 32646 20542 32710
rect 20606 32646 20612 32710
rect 20400 32574 20612 32646
rect 20400 32510 20542 32574
rect 20606 32510 20612 32574
rect 20400 32504 20612 32510
rect 20808 32574 21020 32716
rect 20808 32510 20814 32574
rect 20878 32510 21020 32574
rect 20808 32504 21020 32510
rect 21216 32504 21564 32716
rect 21624 32776 21836 33124
rect 22032 32776 22244 33124
rect 21624 32716 21700 32776
rect 22168 32716 22244 32776
rect 21624 32574 21836 32716
rect 21624 32510 21630 32574
rect 21694 32510 21836 32574
rect 21624 32504 21836 32510
rect 22032 32574 22244 32716
rect 26928 33118 27276 33260
rect 26928 33054 27206 33118
rect 27270 33054 27276 33118
rect 26928 32846 27276 33054
rect 26928 32782 27206 32846
rect 27270 32782 27276 32846
rect 26928 32640 27276 32782
rect 68952 33320 69164 33804
rect 73848 33798 74060 33804
rect 73848 33734 73854 33798
rect 73918 33734 74060 33798
rect 73848 33662 74060 33734
rect 73848 33598 73854 33662
rect 73918 33598 74060 33662
rect 73848 33592 74060 33598
rect 74256 33798 74468 33804
rect 74256 33734 74262 33798
rect 74326 33734 74468 33798
rect 74256 33662 74468 33734
rect 74256 33598 74262 33662
rect 74326 33598 74468 33662
rect 74256 33592 74468 33598
rect 74664 33798 75012 33804
rect 74664 33734 74806 33798
rect 74870 33734 74942 33798
rect 75006 33734 75012 33798
rect 74664 33728 75012 33734
rect 74664 33668 74876 33728
rect 75072 33668 75284 33804
rect 75480 33798 75692 33940
rect 94112 34000 94324 34076
rect 94112 33944 94176 34000
rect 94232 33944 94324 34000
rect 94112 33940 94324 33944
rect 94112 33934 94732 33940
rect 94112 33870 94662 33934
rect 94726 33870 94732 33934
rect 94112 33864 94732 33870
rect 75480 33734 75486 33798
rect 75550 33734 75692 33798
rect 75480 33728 75692 33734
rect 74664 33592 75284 33668
rect 74800 33532 74876 33592
rect 73848 33390 74060 33396
rect 73848 33326 73854 33390
rect 73918 33326 74060 33390
rect 68952 33260 69028 33320
rect 68952 33118 69164 33260
rect 73848 33184 74060 33326
rect 74256 33390 74468 33396
rect 74256 33326 74262 33390
rect 74326 33326 74468 33390
rect 74256 33184 74468 33326
rect 74664 33254 74876 33532
rect 75072 33260 75284 33532
rect 74974 33254 75284 33260
rect 74664 33190 74806 33254
rect 74870 33190 74876 33254
rect 74936 33190 74942 33254
rect 75006 33190 75284 33254
rect 74664 33184 74876 33190
rect 74974 33184 75284 33190
rect 75480 33526 75692 33532
rect 75480 33462 75486 33526
rect 75550 33462 75692 33526
rect 75480 33184 75692 33462
rect 73984 33124 74060 33184
rect 74392 33124 74468 33184
rect 75480 33124 75556 33184
rect 68952 33054 68958 33118
rect 69022 33054 69164 33118
rect 68952 32846 69164 33054
rect 68952 32782 68958 32846
rect 69022 32782 69164 32846
rect 68952 32640 69164 32782
rect 27200 32580 27276 32640
rect 69088 32580 69164 32640
rect 22032 32510 22174 32574
rect 22238 32510 22244 32574
rect 22032 32504 22244 32510
rect 21216 32444 21292 32504
rect 1768 32320 1980 32444
rect 1768 32308 1818 32320
rect 1224 32302 1818 32308
rect 1224 32238 1230 32302
rect 1294 32264 1818 32302
rect 1874 32264 1980 32320
rect 20944 32368 21292 32444
rect 20944 32308 21020 32368
rect 1294 32238 1980 32264
rect 1224 32232 1980 32238
rect 20400 32302 20612 32308
rect 20400 32238 20542 32302
rect 20606 32238 20612 32302
rect 13600 32166 13812 32172
rect 13600 32102 13742 32166
rect 13806 32102 13812 32166
rect 13600 32030 13812 32102
rect 20400 32166 20612 32238
rect 20400 32102 20406 32166
rect 20470 32102 20612 32166
rect 20400 32096 20612 32102
rect 20808 32302 21564 32308
rect 20808 32238 20814 32302
rect 20878 32238 21564 32302
rect 20808 32232 21564 32238
rect 20808 32166 21020 32232
rect 20808 32102 20950 32166
rect 21014 32102 21020 32166
rect 20808 32096 21020 32102
rect 21216 32166 21564 32232
rect 21216 32102 21494 32166
rect 21558 32102 21564 32166
rect 21216 32096 21564 32102
rect 21624 32302 21836 32308
rect 21624 32238 21630 32302
rect 21694 32238 21836 32302
rect 21624 32166 21836 32238
rect 21624 32102 21630 32166
rect 21694 32102 21836 32166
rect 21624 32096 21836 32102
rect 22032 32302 22244 32308
rect 22032 32238 22174 32302
rect 22238 32238 22244 32302
rect 22032 32166 22244 32238
rect 22032 32102 22038 32166
rect 22102 32102 22244 32166
rect 22032 32096 22244 32102
rect 26928 32302 27276 32580
rect 26928 32238 27206 32302
rect 27270 32238 27276 32302
rect 26928 32096 27276 32238
rect 27200 32036 27276 32096
rect 13600 31966 13742 32030
rect 13806 31966 13812 32030
rect 13600 31960 13812 31966
rect 26928 32030 27276 32036
rect 26928 31966 27206 32030
rect 27270 31966 27276 32030
rect 20400 31894 20612 31900
rect 20400 31830 20406 31894
rect 20470 31830 20612 31894
rect 20400 31758 20612 31830
rect 20400 31694 20542 31758
rect 20606 31694 20612 31758
rect 20400 31688 20612 31694
rect 20808 31894 21020 31900
rect 20808 31830 20950 31894
rect 21014 31830 21020 31894
rect 20808 31688 21020 31830
rect 21216 31894 21564 31900
rect 21216 31830 21494 31894
rect 21558 31830 21564 31894
rect 21216 31758 21564 31830
rect 21216 31694 21222 31758
rect 21286 31694 21564 31758
rect 21216 31688 21564 31694
rect 21624 31894 21836 31900
rect 21624 31830 21630 31894
rect 21694 31830 21836 31894
rect 21624 31758 21836 31830
rect 21624 31694 21630 31758
rect 21694 31694 21836 31758
rect 21624 31688 21836 31694
rect 22032 31894 22244 31900
rect 22032 31830 22038 31894
rect 22102 31830 22244 31894
rect 22032 31758 22244 31830
rect 26928 31824 27276 31966
rect 68952 32096 69164 32580
rect 73848 32776 74060 33124
rect 74256 32776 74468 33124
rect 74800 33048 75148 33124
rect 74800 32988 74876 33048
rect 75072 32988 75148 33048
rect 74664 32982 75012 32988
rect 74664 32918 74806 32982
rect 74870 32918 74942 32982
rect 75006 32918 75012 32982
rect 74664 32912 75012 32918
rect 74664 32852 74876 32912
rect 74664 32776 75012 32852
rect 75072 32776 75284 32988
rect 75480 32982 75692 33124
rect 75480 32918 75622 32982
rect 75686 32918 75692 32982
rect 75480 32912 75692 32918
rect 73848 32716 73924 32776
rect 74392 32716 74468 32776
rect 74800 32716 74876 32776
rect 73848 32574 74060 32716
rect 73848 32510 73990 32574
rect 74054 32510 74060 32574
rect 73848 32504 74060 32510
rect 74256 32574 74468 32716
rect 74256 32510 74398 32574
rect 74462 32510 74468 32574
rect 74256 32504 74468 32510
rect 74664 32574 74876 32716
rect 74936 32716 75012 32776
rect 74936 32640 75284 32716
rect 74664 32510 74670 32574
rect 74734 32510 74876 32574
rect 74664 32504 74876 32510
rect 75072 32504 75284 32640
rect 75480 32710 75692 32716
rect 75480 32646 75622 32710
rect 75686 32646 75692 32710
rect 75480 32574 75692 32646
rect 75480 32510 75486 32574
rect 75550 32510 75692 32574
rect 75480 32504 75692 32510
rect 94112 32320 94324 32444
rect 73848 32302 74060 32308
rect 73848 32238 73990 32302
rect 74054 32238 74060 32302
rect 73848 32166 74060 32238
rect 73848 32102 73990 32166
rect 74054 32102 74060 32166
rect 73848 32096 74060 32102
rect 74256 32302 74468 32308
rect 74256 32238 74398 32302
rect 74462 32238 74468 32302
rect 74256 32166 74468 32238
rect 74256 32102 74262 32166
rect 74326 32102 74468 32166
rect 74256 32096 74468 32102
rect 74664 32302 74876 32308
rect 74664 32238 74670 32302
rect 74734 32238 74876 32302
rect 74664 32166 74876 32238
rect 74664 32102 74806 32166
rect 74870 32102 74876 32166
rect 74664 32096 74876 32102
rect 75072 32096 75284 32308
rect 75480 32302 75692 32308
rect 75480 32238 75486 32302
rect 75550 32238 75692 32302
rect 75480 32166 75692 32238
rect 94112 32264 94176 32320
rect 94232 32308 94324 32320
rect 94232 32302 94732 32308
rect 94232 32264 94662 32302
rect 94112 32238 94662 32264
rect 94726 32238 94732 32302
rect 94112 32232 94732 32238
rect 75480 32102 75486 32166
rect 75550 32102 75692 32166
rect 75480 32096 75692 32102
rect 68952 32036 69028 32096
rect 75072 32036 75148 32096
rect 68952 31824 69164 32036
rect 74800 31960 75148 32036
rect 74800 31900 74876 31960
rect 27064 31764 27140 31824
rect 69088 31764 69164 31824
rect 22032 31694 22174 31758
rect 22238 31694 22244 31758
rect 22032 31688 22244 31694
rect 26928 31552 27276 31764
rect 68952 31552 69164 31764
rect 73848 31894 74060 31900
rect 73848 31830 73990 31894
rect 74054 31830 74060 31894
rect 73848 31758 74060 31830
rect 73848 31694 73854 31758
rect 73918 31694 74060 31758
rect 73848 31688 74060 31694
rect 74256 31894 74468 31900
rect 74256 31830 74262 31894
rect 74326 31830 74468 31894
rect 74256 31758 74468 31830
rect 74256 31694 74398 31758
rect 74462 31694 74468 31758
rect 74256 31688 74468 31694
rect 74664 31894 75284 31900
rect 74664 31830 74806 31894
rect 74870 31830 75284 31894
rect 74664 31824 75284 31830
rect 74664 31758 74876 31824
rect 74664 31694 74806 31758
rect 74870 31694 74876 31758
rect 74664 31688 74876 31694
rect 75072 31758 75284 31824
rect 75072 31694 75214 31758
rect 75278 31694 75284 31758
rect 75072 31688 75284 31694
rect 75480 31894 75692 31900
rect 75480 31830 75486 31894
rect 75550 31830 75692 31894
rect 75480 31758 75692 31830
rect 75480 31694 75622 31758
rect 75686 31694 75692 31758
rect 75480 31688 75692 31694
rect 26928 31492 27004 31552
rect 69088 31492 69164 31552
rect 20400 31486 20612 31492
rect 20400 31422 20542 31486
rect 20606 31422 20612 31486
rect 14200 31371 14266 31374
rect 14774 31371 14840 31374
rect 14200 31369 14840 31371
rect 13192 31298 13404 31356
rect 14200 31313 14205 31369
rect 14261 31313 14779 31369
rect 14835 31313 14840 31369
rect 14200 31311 14840 31313
rect 14200 31308 14266 31311
rect 14774 31308 14840 31311
rect 20400 31350 20612 31422
rect 13192 31242 13260 31298
rect 13316 31242 13404 31298
rect 20400 31286 20406 31350
rect 20470 31286 20612 31350
rect 20400 31280 20612 31286
rect 20808 31486 21564 31492
rect 20808 31422 21222 31486
rect 21286 31422 21564 31486
rect 20808 31416 21564 31422
rect 20808 31356 21020 31416
rect 20808 31350 21156 31356
rect 20808 31286 20950 31350
rect 21014 31286 21086 31350
rect 21150 31286 21156 31350
rect 20808 31280 21156 31286
rect 21216 31280 21564 31416
rect 21624 31486 21836 31492
rect 21624 31422 21630 31486
rect 21694 31422 21836 31486
rect 21624 31350 21836 31422
rect 21624 31286 21766 31350
rect 21830 31286 21836 31350
rect 21624 31280 21836 31286
rect 22032 31486 22244 31492
rect 22032 31422 22174 31486
rect 22238 31422 22244 31486
rect 22032 31350 22244 31422
rect 22032 31286 22038 31350
rect 22102 31286 22244 31350
rect 22032 31280 22244 31286
rect 26928 31280 27276 31492
rect 13192 31220 13404 31242
rect 27200 31220 27276 31280
rect 0 31144 13404 31220
rect 20400 31078 20612 31084
rect 20400 31014 20406 31078
rect 20470 31014 20612 31078
rect 20400 30942 20612 31014
rect 20400 30878 20406 30942
rect 20470 30878 20612 30942
rect 20400 30872 20612 30878
rect 20808 31078 21020 31084
rect 21118 31078 21564 31084
rect 20808 31014 20950 31078
rect 21014 31014 21020 31078
rect 21080 31014 21086 31078
rect 21150 31014 21564 31078
rect 20808 30942 21020 31014
rect 21118 31008 21564 31014
rect 20808 30878 20814 30942
rect 20878 30878 21020 30942
rect 20808 30872 21020 30878
rect 21216 30942 21564 31008
rect 21216 30878 21494 30942
rect 21558 30878 21564 30942
rect 21216 30872 21564 30878
rect 21624 31078 21836 31084
rect 21624 31014 21766 31078
rect 21830 31014 21836 31078
rect 21624 30942 21836 31014
rect 21624 30878 21766 30942
rect 21830 30878 21836 30942
rect 21624 30872 21836 30878
rect 22032 31078 22244 31084
rect 22032 31014 22038 31078
rect 22102 31014 22244 31078
rect 22032 30942 22244 31014
rect 22032 30878 22174 30942
rect 22238 30878 22244 30942
rect 22032 30872 22244 30878
rect 26928 31008 27276 31220
rect 68952 31280 69164 31492
rect 73848 31486 74060 31492
rect 73848 31422 73854 31486
rect 73918 31422 74060 31486
rect 73848 31350 74060 31422
rect 73848 31286 73990 31350
rect 74054 31286 74060 31350
rect 73848 31280 74060 31286
rect 74256 31486 74468 31492
rect 74256 31422 74398 31486
rect 74462 31422 74468 31486
rect 74256 31350 74468 31422
rect 74256 31286 74398 31350
rect 74462 31286 74468 31350
rect 74256 31280 74468 31286
rect 74664 31486 74876 31492
rect 74664 31422 74806 31486
rect 74870 31422 74876 31486
rect 74664 31280 74876 31422
rect 75072 31486 75284 31492
rect 75072 31422 75214 31486
rect 75278 31422 75284 31486
rect 75072 31350 75284 31422
rect 75072 31286 75078 31350
rect 75142 31286 75284 31350
rect 75072 31280 75284 31286
rect 75480 31486 75692 31492
rect 75480 31422 75622 31486
rect 75686 31422 75692 31486
rect 75480 31350 75692 31422
rect 75480 31286 75486 31350
rect 75550 31286 75692 31350
rect 75480 31280 75692 31286
rect 68952 31220 69028 31280
rect 68952 31008 69164 31220
rect 73848 31078 74060 31084
rect 73848 31014 73990 31078
rect 74054 31014 74060 31078
rect 26928 30948 27004 31008
rect 68952 30948 69028 31008
rect 13600 30806 13812 30812
rect 13600 30742 13606 30806
rect 13670 30742 13812 30806
rect 13600 30676 13812 30742
rect 26928 30736 27276 30948
rect 68952 30736 69164 30948
rect 73848 30942 74060 31014
rect 73848 30878 73854 30942
rect 73918 30878 74060 30942
rect 73848 30872 74060 30878
rect 74256 31078 74468 31084
rect 74256 31014 74398 31078
rect 74462 31014 74468 31078
rect 74256 30942 74468 31014
rect 74256 30878 74398 30942
rect 74462 30878 74468 30942
rect 74256 30872 74468 30878
rect 74664 30942 74876 31084
rect 74664 30878 74670 30942
rect 74734 30878 74876 30942
rect 74664 30872 74876 30878
rect 75072 31078 75284 31084
rect 75072 31014 75078 31078
rect 75142 31014 75284 31078
rect 75072 30872 75284 31014
rect 75480 31078 75692 31084
rect 75480 31014 75486 31078
rect 75550 31014 75692 31078
rect 75480 30942 75692 31014
rect 75480 30878 75622 30942
rect 75686 30878 75692 30942
rect 75480 30872 75692 30878
rect 75072 30812 75148 30872
rect 27064 30676 27140 30736
rect 69088 30676 69164 30736
rect 74800 30736 75148 30812
rect 74800 30676 74876 30736
rect 1224 30670 1980 30676
rect 1224 30606 1230 30670
rect 1294 30640 1980 30670
rect 1294 30606 1818 30640
rect 1224 30600 1818 30606
rect 1768 30584 1818 30600
rect 1874 30584 1980 30640
rect 13464 30670 13812 30676
rect 13464 30606 13470 30670
rect 13534 30606 13812 30670
rect 13464 30600 13812 30606
rect 20400 30670 20612 30676
rect 20400 30606 20406 30670
rect 20470 30606 20612 30670
rect 1768 30464 1980 30584
rect 20400 30534 20612 30606
rect 20400 30470 20406 30534
rect 20470 30470 20612 30534
rect 20400 30464 20612 30470
rect 20808 30670 21020 30676
rect 20808 30606 20814 30670
rect 20878 30606 21020 30670
rect 20808 30464 21020 30606
rect 21216 30670 21564 30676
rect 21216 30606 21494 30670
rect 21558 30606 21564 30670
rect 21216 30464 21564 30606
rect 21624 30670 21836 30676
rect 21624 30606 21766 30670
rect 21830 30606 21836 30670
rect 21624 30534 21836 30606
rect 21624 30470 21766 30534
rect 21830 30470 21836 30534
rect 21624 30464 21836 30470
rect 22032 30670 22244 30676
rect 22032 30606 22174 30670
rect 22238 30606 22244 30670
rect 22032 30534 22244 30606
rect 22032 30470 22038 30534
rect 22102 30470 22244 30534
rect 22032 30464 22244 30470
rect 26928 30464 27276 30676
rect 68952 30464 69164 30676
rect 73848 30670 74060 30676
rect 73848 30606 73854 30670
rect 73918 30606 74060 30670
rect 73848 30534 74060 30606
rect 73848 30470 73854 30534
rect 73918 30470 74060 30534
rect 73848 30464 74060 30470
rect 74256 30670 74468 30676
rect 74256 30606 74398 30670
rect 74462 30606 74468 30670
rect 74256 30534 74468 30606
rect 74256 30470 74262 30534
rect 74326 30470 74468 30534
rect 74256 30464 74468 30470
rect 74664 30670 75284 30676
rect 74664 30606 74670 30670
rect 74734 30606 75284 30670
rect 74664 30600 75284 30606
rect 74664 30534 74876 30600
rect 74664 30470 74806 30534
rect 74870 30470 74876 30534
rect 74664 30464 74876 30470
rect 75072 30464 75284 30600
rect 75480 30670 75692 30676
rect 75480 30606 75622 30670
rect 75686 30606 75692 30670
rect 75480 30534 75692 30606
rect 75480 30470 75486 30534
rect 75550 30470 75692 30534
rect 75480 30464 75692 30470
rect 94112 30670 94732 30676
rect 94112 30640 94662 30670
rect 94112 30584 94176 30640
rect 94232 30606 94662 30640
rect 94726 30606 94732 30670
rect 94232 30600 94732 30606
rect 94232 30584 94324 30600
rect 94112 30464 94324 30584
rect 21216 30404 21292 30464
rect 20944 30328 21292 30404
rect 26928 30404 27004 30464
rect 69088 30404 69164 30464
rect 20944 30268 21020 30328
rect 13192 30170 13404 30268
rect 13192 30132 13260 30170
rect 0 30114 13260 30132
rect 13316 30114 13404 30170
rect 0 30056 13404 30114
rect 20400 30262 20612 30268
rect 20400 30198 20406 30262
rect 20470 30198 20612 30262
rect 14200 30101 14266 30104
rect 14694 30101 14760 30104
rect 14200 30099 14760 30101
rect 14200 30043 14205 30099
rect 14261 30043 14699 30099
rect 14755 30043 14760 30099
rect 14200 30041 14760 30043
rect 14200 30038 14266 30041
rect 14694 30038 14760 30041
rect 20400 30056 20612 30198
rect 20808 30192 21564 30268
rect 20808 30056 21020 30192
rect 21216 30126 21564 30192
rect 21216 30062 21222 30126
rect 21286 30062 21564 30126
rect 21216 30056 21564 30062
rect 21624 30262 21836 30268
rect 21624 30198 21766 30262
rect 21830 30198 21836 30262
rect 21624 30126 21836 30198
rect 21624 30062 21766 30126
rect 21830 30062 21836 30126
rect 21624 30056 21836 30062
rect 22032 30262 22244 30268
rect 22032 30198 22038 30262
rect 22102 30198 22244 30262
rect 22032 30126 22244 30198
rect 26928 30192 27276 30404
rect 27200 30132 27276 30192
rect 22032 30062 22038 30126
rect 22102 30062 22244 30126
rect 22032 30056 22244 30062
rect 20400 29996 20476 30056
rect 20400 29854 20612 29996
rect 26928 29920 27276 30132
rect 68952 30192 69164 30404
rect 73848 30262 74060 30268
rect 73848 30198 73854 30262
rect 73918 30198 74060 30262
rect 68952 30132 69028 30192
rect 68952 29920 69164 30132
rect 73848 30126 74060 30198
rect 73848 30062 73990 30126
rect 74054 30062 74060 30126
rect 73848 30056 74060 30062
rect 74256 30262 74468 30268
rect 74256 30198 74262 30262
rect 74326 30198 74468 30262
rect 74256 30126 74468 30198
rect 74256 30062 74262 30126
rect 74326 30062 74468 30126
rect 74256 30056 74468 30062
rect 74664 30262 74876 30268
rect 74664 30198 74806 30262
rect 74870 30198 74876 30262
rect 74664 30126 74876 30198
rect 75072 30132 75284 30268
rect 74974 30126 75284 30132
rect 74664 30062 74670 30126
rect 74734 30062 74876 30126
rect 74936 30062 74942 30126
rect 75006 30062 75284 30126
rect 74664 30056 74876 30062
rect 74974 30056 75284 30062
rect 75480 30262 75692 30268
rect 75480 30198 75486 30262
rect 75550 30198 75692 30262
rect 75480 30056 75692 30198
rect 75480 29996 75556 30056
rect 27064 29860 27140 29920
rect 68952 29860 69028 29920
rect 20400 29790 20542 29854
rect 20606 29790 20612 29854
rect 20400 29784 20612 29790
rect 20808 29648 21020 29860
rect 20944 29588 21020 29648
rect 20400 29582 20612 29588
rect 20400 29518 20542 29582
rect 20606 29518 20612 29582
rect 13600 29446 13812 29452
rect 13600 29382 13742 29446
rect 13806 29382 13812 29446
rect 13600 29310 13812 29382
rect 13600 29246 13606 29310
rect 13670 29246 13812 29310
rect 13600 29240 13812 29246
rect 20400 29240 20612 29518
rect 20808 29452 21020 29588
rect 21216 29854 21564 29860
rect 21216 29790 21222 29854
rect 21286 29790 21564 29854
rect 21216 29648 21564 29790
rect 21624 29854 21836 29860
rect 21624 29790 21766 29854
rect 21830 29790 21836 29854
rect 21624 29718 21836 29790
rect 21624 29654 21630 29718
rect 21694 29654 21836 29718
rect 21624 29648 21836 29654
rect 22032 29854 22244 29860
rect 22032 29790 22038 29854
rect 22102 29790 22244 29854
rect 22032 29718 22244 29790
rect 22032 29654 22174 29718
rect 22238 29654 22244 29718
rect 22032 29648 22244 29654
rect 21216 29588 21292 29648
rect 21216 29452 21564 29588
rect 20808 29376 21564 29452
rect 20808 29240 21020 29376
rect 21216 29316 21564 29376
rect 21118 29310 21564 29316
rect 21080 29246 21086 29310
rect 21150 29246 21564 29310
rect 21118 29240 21564 29246
rect 21624 29446 21836 29452
rect 21624 29382 21630 29446
rect 21694 29382 21836 29446
rect 21624 29240 21836 29382
rect 22032 29446 22244 29452
rect 22032 29382 22174 29446
rect 22238 29382 22244 29446
rect 22032 29240 22244 29382
rect 26928 29376 27276 29860
rect 68952 29376 69164 29860
rect 73848 29854 74060 29860
rect 73848 29790 73990 29854
rect 74054 29790 74060 29854
rect 73848 29718 74060 29790
rect 73848 29654 73854 29718
rect 73918 29654 74060 29718
rect 73848 29648 74060 29654
rect 74256 29854 74468 29860
rect 74256 29790 74262 29854
rect 74326 29790 74468 29854
rect 74256 29718 74468 29790
rect 74256 29654 74398 29718
rect 74462 29654 74468 29718
rect 74256 29648 74468 29654
rect 74664 29854 75012 29860
rect 74664 29790 74670 29854
rect 74734 29790 74942 29854
rect 75006 29790 75012 29854
rect 74664 29784 75012 29790
rect 74664 29648 74876 29784
rect 75072 29724 75284 29860
rect 75480 29854 75692 29996
rect 75480 29790 75622 29854
rect 75686 29790 75692 29854
rect 75480 29784 75692 29790
rect 74800 29588 74876 29648
rect 74936 29648 75284 29724
rect 74936 29588 75012 29648
rect 75208 29588 75284 29648
rect 74664 29512 75012 29588
rect 27064 29316 27140 29376
rect 69088 29316 69164 29376
rect 20400 29180 20476 29240
rect 21624 29180 21700 29240
rect 22032 29180 22108 29240
rect 1224 29038 1980 29044
rect 1224 28974 1230 29038
rect 1294 28974 1980 29038
rect 1224 28968 1980 28974
rect 20400 29038 20612 29180
rect 20400 28974 20406 29038
rect 20470 28974 20612 29038
rect 20400 28968 20612 28974
rect 20808 29038 21156 29044
rect 20808 28974 21086 29038
rect 21150 28974 21156 29038
rect 20808 28968 21156 28974
rect 1768 28960 1980 28968
rect 1768 28904 1818 28960
rect 1874 28904 1980 28960
rect 1768 28832 1980 28904
rect 20808 28908 21020 28968
rect 21216 28908 21564 29044
rect 20808 28902 21564 28908
rect 20808 28838 20950 28902
rect 21014 28838 21564 28902
rect 20808 28832 21564 28838
rect 21624 28832 21836 29180
rect 22032 28832 22244 29180
rect 20944 28772 21020 28832
rect 21760 28772 21836 28832
rect 22168 28772 22244 28832
rect 20400 28766 20612 28772
rect 20400 28702 20406 28766
rect 20470 28702 20612 28766
rect 20400 28630 20612 28702
rect 20400 28566 20542 28630
rect 20606 28566 20612 28630
rect 20400 28560 20612 28566
rect 20808 28630 21020 28772
rect 21118 28766 21564 28772
rect 21080 28702 21086 28766
rect 21150 28702 21564 28766
rect 21118 28696 21564 28702
rect 20808 28566 20814 28630
rect 20878 28566 21020 28630
rect 20808 28560 21020 28566
rect 21216 28560 21564 28696
rect 14200 28543 14266 28546
rect 14614 28543 14680 28546
rect 14200 28541 14680 28543
rect 0 28470 13404 28500
rect 14200 28485 14205 28541
rect 14261 28485 14619 28541
rect 14675 28485 14680 28541
rect 14200 28483 14680 28485
rect 14200 28480 14266 28483
rect 14614 28480 14680 28483
rect 0 28424 13260 28470
rect 13192 28414 13260 28424
rect 13316 28414 13404 28470
rect 21624 28424 21836 28772
rect 22032 28424 22244 28772
rect 26928 29174 27276 29316
rect 26928 29110 27206 29174
rect 27270 29110 27276 29174
rect 26928 28902 27276 29110
rect 26928 28838 27206 28902
rect 27270 28838 27276 28902
rect 26928 28766 27276 28838
rect 26928 28702 27070 28766
rect 27134 28702 27276 28766
rect 26928 28696 27276 28702
rect 68952 29174 69164 29316
rect 68952 29110 68958 29174
rect 69022 29110 69164 29174
rect 68952 28902 69164 29110
rect 68952 28838 68958 28902
rect 69022 28838 69164 28902
rect 68952 28766 69164 28838
rect 73848 29446 74060 29452
rect 73848 29382 73854 29446
rect 73918 29382 74060 29446
rect 73848 29240 74060 29382
rect 74256 29446 74468 29452
rect 74256 29382 74398 29446
rect 74462 29382 74468 29446
rect 74256 29240 74468 29382
rect 74664 29310 74876 29512
rect 74664 29246 74670 29310
rect 74734 29246 74876 29310
rect 74664 29240 74876 29246
rect 75072 29240 75284 29588
rect 75480 29582 75692 29588
rect 75480 29518 75622 29582
rect 75686 29518 75692 29582
rect 75480 29240 75692 29518
rect 73848 29180 73924 29240
rect 74392 29180 74468 29240
rect 75616 29180 75692 29240
rect 73848 28832 74060 29180
rect 74256 28832 74468 29180
rect 73984 28772 74060 28832
rect 74392 28772 74468 28832
rect 68952 28702 68958 28766
rect 69022 28702 69094 28766
rect 69158 28702 69164 28766
rect 68952 28696 69164 28702
rect 13192 28288 13404 28414
rect 21760 28364 21836 28424
rect 22168 28364 22244 28424
rect 20400 28358 20612 28364
rect 20400 28294 20542 28358
rect 20606 28294 20612 28358
rect 20400 28222 20612 28294
rect 20400 28158 20542 28222
rect 20606 28158 20612 28222
rect 20400 28152 20612 28158
rect 20808 28358 21020 28364
rect 20808 28294 20814 28358
rect 20878 28294 21020 28358
rect 20808 28092 21020 28294
rect 20808 28016 21156 28092
rect 21216 28016 21564 28364
rect 21624 28222 21836 28364
rect 21624 28158 21766 28222
rect 21830 28158 21836 28222
rect 21624 28152 21836 28158
rect 22032 28222 22244 28364
rect 22032 28158 22038 28222
rect 22102 28158 22244 28222
rect 22032 28152 22244 28158
rect 26928 28494 27276 28500
rect 26928 28430 27070 28494
rect 27134 28430 27276 28494
rect 26928 28152 27276 28430
rect 68952 28494 69164 28500
rect 68952 28430 68958 28494
rect 69022 28430 69164 28494
rect 68952 28358 69164 28430
rect 73848 28424 74060 28772
rect 74256 28424 74468 28772
rect 74664 29038 74876 29044
rect 74664 28974 74670 29038
rect 74734 28974 74876 29038
rect 74664 28832 74876 28974
rect 75072 28908 75284 29044
rect 75480 29038 75692 29180
rect 75480 28974 75486 29038
rect 75550 28974 75692 29038
rect 75480 28968 75692 28974
rect 94112 29038 94732 29044
rect 94112 28974 94662 29038
rect 94726 28974 94732 29038
rect 94112 28968 94732 28974
rect 74936 28832 75284 28908
rect 94112 28960 94324 28968
rect 94112 28904 94176 28960
rect 94232 28904 94324 28960
rect 94112 28832 94324 28904
rect 74664 28772 74740 28832
rect 74936 28772 75012 28832
rect 74664 28696 75012 28772
rect 75072 28772 75148 28832
rect 74664 28636 74876 28696
rect 74664 28630 75012 28636
rect 74664 28566 74942 28630
rect 75006 28566 75012 28630
rect 74664 28560 75012 28566
rect 75072 28560 75284 28772
rect 75480 28766 75692 28772
rect 75480 28702 75486 28766
rect 75550 28702 75692 28766
rect 75480 28630 75692 28702
rect 75480 28566 75622 28630
rect 75686 28566 75692 28630
rect 75480 28560 75692 28566
rect 73984 28364 74060 28424
rect 74392 28364 74468 28424
rect 68952 28294 69094 28358
rect 69158 28294 69164 28358
rect 68952 28152 69164 28294
rect 73848 28222 74060 28364
rect 73848 28158 73990 28222
rect 74054 28158 74060 28222
rect 73848 28152 74060 28158
rect 74256 28222 74468 28364
rect 74256 28158 74262 28222
rect 74326 28158 74468 28222
rect 74256 28152 74468 28158
rect 74664 28228 74876 28364
rect 74974 28358 75284 28364
rect 74936 28294 74942 28358
rect 75006 28294 75284 28358
rect 74974 28288 75284 28294
rect 75072 28228 75284 28288
rect 74664 28152 75284 28228
rect 75480 28358 75692 28364
rect 75480 28294 75622 28358
rect 75686 28294 75692 28358
rect 75480 28222 75692 28294
rect 75480 28158 75622 28222
rect 75686 28158 75692 28222
rect 75480 28152 75692 28158
rect 27064 28092 27140 28152
rect 68952 28092 69028 28152
rect 20944 27956 21020 28016
rect 13502 27950 13812 27956
rect 13464 27886 13470 27950
rect 13534 27886 13812 27950
rect 13502 27880 13812 27886
rect 13600 27814 13812 27880
rect 13600 27750 13742 27814
rect 13806 27750 13812 27814
rect 13600 27744 13812 27750
rect 20400 27950 20612 27956
rect 20400 27886 20542 27950
rect 20606 27886 20612 27950
rect 20400 27814 20612 27886
rect 20400 27750 20406 27814
rect 20470 27750 20612 27814
rect 20400 27744 20612 27750
rect 20808 27744 21020 27956
rect 21080 27956 21156 28016
rect 21352 27956 21428 28016
rect 21080 27880 21564 27956
rect 21216 27814 21564 27880
rect 21216 27750 21494 27814
rect 21558 27750 21564 27814
rect 21216 27744 21564 27750
rect 21624 27950 21836 27956
rect 21624 27886 21766 27950
rect 21830 27886 21836 27950
rect 21624 27814 21836 27886
rect 21624 27750 21630 27814
rect 21694 27750 21836 27814
rect 21624 27744 21836 27750
rect 22032 27950 22244 27956
rect 22032 27886 22038 27950
rect 22102 27886 22244 27950
rect 22032 27814 22244 27886
rect 26928 27880 27276 28092
rect 27200 27820 27276 27880
rect 22032 27750 22038 27814
rect 22102 27750 22244 27814
rect 22032 27744 22244 27750
rect 26928 27744 27276 27820
rect 68952 27880 69164 28092
rect 74664 28016 74876 28152
rect 75072 28016 75284 28152
rect 75072 27956 75148 28016
rect 73848 27950 74060 27956
rect 73848 27886 73990 27950
rect 74054 27886 74060 27950
rect 68952 27820 69028 27880
rect 27054 27548 27152 27744
rect 0 27472 2116 27548
rect 2040 27412 2116 27472
rect 20400 27542 20612 27548
rect 20400 27478 20406 27542
rect 20470 27478 20612 27542
rect 1224 27406 1844 27412
rect 1224 27342 1230 27406
rect 1294 27342 1844 27406
rect 1224 27336 1844 27342
rect 2040 27342 13404 27412
rect 2040 27336 13260 27342
rect 1768 27301 1844 27336
rect 1768 27280 1895 27301
rect 1768 27224 1818 27280
rect 1874 27276 1895 27280
rect 13192 27286 13260 27336
rect 13316 27286 13404 27342
rect 20400 27406 20612 27478
rect 20400 27342 20542 27406
rect 20606 27342 20612 27406
rect 20400 27336 20612 27342
rect 20808 27406 21020 27548
rect 21216 27542 21564 27548
rect 21216 27478 21494 27542
rect 21558 27478 21564 27542
rect 21216 27412 21564 27478
rect 21118 27406 21564 27412
rect 20808 27342 20814 27406
rect 20878 27342 21020 27406
rect 21080 27342 21086 27406
rect 21150 27342 21564 27406
rect 20808 27336 21020 27342
rect 21118 27336 21564 27342
rect 21624 27542 21836 27548
rect 21624 27478 21630 27542
rect 21694 27478 21836 27542
rect 21624 27406 21836 27478
rect 21624 27342 21630 27406
rect 21694 27342 21836 27406
rect 21624 27336 21836 27342
rect 22032 27542 22244 27548
rect 22032 27478 22038 27542
rect 22102 27478 22244 27542
rect 22032 27406 22244 27478
rect 22032 27342 22038 27406
rect 22102 27342 22244 27406
rect 22032 27336 22244 27342
rect 26928 27542 27276 27548
rect 26928 27478 27070 27542
rect 27134 27478 27276 27542
rect 26928 27336 27276 27478
rect 68952 27542 69164 27820
rect 73848 27814 74060 27886
rect 73848 27750 73990 27814
rect 74054 27750 74060 27814
rect 73848 27744 74060 27750
rect 74256 27950 74468 27956
rect 74256 27886 74262 27950
rect 74326 27886 74468 27950
rect 74256 27814 74468 27886
rect 74256 27750 74262 27814
rect 74326 27750 74468 27814
rect 74256 27744 74468 27750
rect 74664 27814 74876 27956
rect 74664 27750 74670 27814
rect 74734 27750 74876 27814
rect 74664 27744 74876 27750
rect 75072 27744 75284 27956
rect 75480 27950 75692 27956
rect 75480 27886 75622 27950
rect 75686 27886 75692 27950
rect 75480 27814 75692 27886
rect 75480 27750 75486 27814
rect 75550 27750 75692 27814
rect 75480 27744 75692 27750
rect 75072 27684 75148 27744
rect 74800 27608 75148 27684
rect 74800 27548 74876 27608
rect 68952 27478 69094 27542
rect 69158 27478 69164 27542
rect 68952 27336 69164 27478
rect 73848 27542 74060 27548
rect 73848 27478 73990 27542
rect 74054 27478 74060 27542
rect 73848 27406 74060 27478
rect 73848 27342 73854 27406
rect 73918 27342 74060 27406
rect 73848 27336 74060 27342
rect 74256 27542 74468 27548
rect 74256 27478 74262 27542
rect 74326 27478 74468 27542
rect 74256 27406 74468 27478
rect 74256 27342 74262 27406
rect 74326 27342 74468 27406
rect 74256 27336 74468 27342
rect 74664 27542 75284 27548
rect 74664 27478 74670 27542
rect 74734 27478 75284 27542
rect 74664 27472 75284 27478
rect 74664 27336 74876 27472
rect 75072 27406 75284 27472
rect 75072 27342 75214 27406
rect 75278 27342 75284 27406
rect 75072 27336 75284 27342
rect 75480 27542 75692 27548
rect 75480 27478 75486 27542
rect 75550 27478 75692 27542
rect 75480 27406 75692 27478
rect 75480 27342 75622 27406
rect 75686 27342 75692 27406
rect 75480 27336 75692 27342
rect 94112 27406 94732 27412
rect 94112 27342 94662 27406
rect 94726 27342 94732 27406
rect 94112 27336 94732 27342
rect 1874 27224 1980 27276
rect 1768 27200 1980 27224
rect 13192 27200 13404 27286
rect 21624 27276 21700 27336
rect 27064 27276 27140 27336
rect 69088 27276 69164 27336
rect 14200 27273 14266 27276
rect 14534 27273 14600 27276
rect 14200 27271 14600 27273
rect 14200 27215 14205 27271
rect 14261 27215 14539 27271
rect 14595 27215 14600 27271
rect 14200 27213 14600 27215
rect 14200 27210 14266 27213
rect 14534 27210 14600 27213
rect 20672 27200 21700 27276
rect 26928 27270 27276 27276
rect 26928 27206 27070 27270
rect 27134 27206 27276 27270
rect 20672 27140 20748 27200
rect 20400 27134 20748 27140
rect 20400 27070 20542 27134
rect 20606 27070 20748 27134
rect 20400 27064 20748 27070
rect 20808 27134 21156 27140
rect 20808 27070 20814 27134
rect 20878 27070 21086 27134
rect 21150 27070 21156 27134
rect 20808 27064 21156 27070
rect 20400 26998 20612 27064
rect 20400 26934 20406 26998
rect 20470 26934 20612 26998
rect 20400 26928 20612 26934
rect 20808 27004 21020 27064
rect 20808 26998 21156 27004
rect 20808 26934 20950 26998
rect 21014 26934 21086 26998
rect 21150 26934 21156 26998
rect 20808 26928 21156 26934
rect 21216 26928 21564 27140
rect 21624 27134 21836 27140
rect 21624 27070 21630 27134
rect 21694 27070 21836 27134
rect 21624 26998 21836 27070
rect 21624 26934 21766 26998
rect 21830 26934 21836 26998
rect 21624 26928 21836 26934
rect 22032 27134 22244 27140
rect 22032 27070 22038 27134
rect 22102 27070 22244 27134
rect 22032 26998 22244 27070
rect 22032 26934 22038 26998
rect 22102 26934 22244 26998
rect 22032 26928 22244 26934
rect 26928 27064 27276 27206
rect 68952 27270 69164 27276
rect 68952 27206 69094 27270
rect 69158 27206 69164 27270
rect 68952 27064 69164 27206
rect 94112 27280 94324 27336
rect 94112 27224 94176 27280
rect 94232 27224 94324 27280
rect 94112 27200 94324 27224
rect 73848 27134 74060 27140
rect 73848 27070 73854 27134
rect 73918 27070 74060 27134
rect 26928 27004 27004 27064
rect 68952 27004 69028 27064
rect 20944 26868 21020 26928
rect 21216 26868 21292 26928
rect 20944 26792 21292 26868
rect 26928 26792 27276 27004
rect 68952 26792 69164 27004
rect 73848 26998 74060 27070
rect 73848 26934 73990 26998
rect 74054 26934 74060 26998
rect 73848 26928 74060 26934
rect 74256 27134 74468 27140
rect 74256 27070 74262 27134
rect 74326 27070 74468 27134
rect 74256 26998 74468 27070
rect 74256 26934 74262 26998
rect 74326 26934 74468 26998
rect 74256 26928 74468 26934
rect 74664 26998 74876 27140
rect 74664 26934 74670 26998
rect 74734 26934 74876 26998
rect 74664 26928 74876 26934
rect 75072 27134 75284 27140
rect 75072 27070 75214 27134
rect 75278 27070 75284 27134
rect 75072 26998 75284 27070
rect 75072 26934 75078 26998
rect 75142 26934 75284 26998
rect 75072 26928 75284 26934
rect 75480 27134 75692 27140
rect 75480 27070 75622 27134
rect 75686 27070 75692 27134
rect 75480 26998 75692 27070
rect 75480 26934 75486 26998
rect 75550 26934 75692 26998
rect 75480 26928 75692 26934
rect 26928 26732 27004 26792
rect 68952 26732 69028 26792
rect 20400 26726 20612 26732
rect 20400 26662 20406 26726
rect 20470 26662 20612 26726
rect 13600 26590 13812 26596
rect 13600 26526 13606 26590
rect 13670 26526 13812 26590
rect 13600 26460 13812 26526
rect 20400 26590 20612 26662
rect 20400 26526 20542 26590
rect 20606 26526 20612 26590
rect 20400 26520 20612 26526
rect 20808 26726 21020 26732
rect 21118 26726 21564 26732
rect 20808 26662 20950 26726
rect 21014 26662 21020 26726
rect 21080 26662 21086 26726
rect 21150 26662 21564 26726
rect 20808 26590 21020 26662
rect 21118 26656 21564 26662
rect 20808 26526 20814 26590
rect 20878 26526 21020 26590
rect 20808 26520 21020 26526
rect 21216 26590 21564 26656
rect 21216 26526 21494 26590
rect 21558 26526 21564 26590
rect 21216 26520 21564 26526
rect 21624 26726 21836 26732
rect 21624 26662 21766 26726
rect 21830 26662 21836 26726
rect 21624 26590 21836 26662
rect 21624 26526 21766 26590
rect 21830 26526 21836 26590
rect 21624 26520 21836 26526
rect 22032 26726 22244 26732
rect 22032 26662 22038 26726
rect 22102 26662 22244 26726
rect 22032 26590 22244 26662
rect 22032 26526 22038 26590
rect 22102 26526 22244 26590
rect 22032 26520 22244 26526
rect 26928 26520 27276 26732
rect 68952 26520 69164 26732
rect 73848 26726 74060 26732
rect 73848 26662 73990 26726
rect 74054 26662 74060 26726
rect 73848 26590 74060 26662
rect 73848 26526 73854 26590
rect 73918 26526 74060 26590
rect 73848 26520 74060 26526
rect 74256 26726 74468 26732
rect 74256 26662 74262 26726
rect 74326 26662 74468 26726
rect 74256 26590 74468 26662
rect 74256 26526 74262 26590
rect 74326 26526 74468 26590
rect 74256 26520 74468 26526
rect 74664 26726 74876 26732
rect 74664 26662 74670 26726
rect 74734 26662 74876 26726
rect 74664 26590 74876 26662
rect 75072 26726 75284 26732
rect 75072 26662 75078 26726
rect 75142 26662 75284 26726
rect 75072 26596 75284 26662
rect 74974 26590 75284 26596
rect 74664 26526 74670 26590
rect 74734 26526 74876 26590
rect 74936 26526 74942 26590
rect 75006 26526 75284 26590
rect 74664 26520 74876 26526
rect 74974 26520 75284 26526
rect 75480 26726 75692 26732
rect 75480 26662 75486 26726
rect 75550 26662 75692 26726
rect 75480 26590 75692 26662
rect 75480 26526 75622 26590
rect 75686 26526 75692 26590
rect 75480 26520 75692 26526
rect 27200 26460 27276 26520
rect 69088 26460 69164 26520
rect 13600 26454 17484 26460
rect 13600 26390 17414 26454
rect 17478 26390 17484 26454
rect 13600 26384 17484 26390
rect 20400 26318 20612 26324
rect 20400 26254 20542 26318
rect 20606 26254 20612 26318
rect 20400 26112 20612 26254
rect 20808 26318 21020 26324
rect 20808 26254 20814 26318
rect 20878 26254 21020 26318
rect 20808 26112 21020 26254
rect 21216 26318 21564 26324
rect 21216 26254 21494 26318
rect 21558 26254 21564 26318
rect 21216 26112 21564 26254
rect 21624 26318 21836 26324
rect 21624 26254 21766 26318
rect 21830 26254 21836 26318
rect 21624 26182 21836 26254
rect 21624 26118 21766 26182
rect 21830 26118 21836 26182
rect 21624 26112 21836 26118
rect 22032 26318 22244 26324
rect 22032 26254 22038 26318
rect 22102 26254 22244 26318
rect 22032 26182 22244 26254
rect 22032 26118 22174 26182
rect 22238 26118 22244 26182
rect 22032 26112 22244 26118
rect 26928 26248 27276 26460
rect 68952 26248 69164 26460
rect 26928 26188 27004 26248
rect 69088 26188 69164 26248
rect 20536 26052 20612 26112
rect 21216 26052 21292 26112
rect 0 25704 13404 25780
rect 1768 25600 1980 25644
rect 1768 25544 1818 25600
rect 1874 25544 1980 25600
rect 13192 25642 13404 25704
rect 14200 25715 14266 25718
rect 14454 25715 14520 25718
rect 14200 25713 14520 25715
rect 14200 25657 14205 25713
rect 14261 25657 14459 25713
rect 14515 25657 14520 25713
rect 20400 25704 20612 26052
rect 20944 25976 21292 26052
rect 26928 26046 27276 26188
rect 26928 25982 27206 26046
rect 27270 25982 27276 26046
rect 26928 25976 27276 25982
rect 20944 25916 21020 25976
rect 27200 25916 27276 25976
rect 20808 25840 21564 25916
rect 20808 25780 21020 25840
rect 20808 25704 21156 25780
rect 21216 25704 21564 25840
rect 21624 25910 21836 25916
rect 21624 25846 21766 25910
rect 21830 25846 21836 25910
rect 21624 25774 21836 25846
rect 21624 25710 21766 25774
rect 21830 25710 21836 25774
rect 21624 25704 21836 25710
rect 22032 25910 22244 25916
rect 22032 25846 22174 25910
rect 22238 25846 22244 25910
rect 22032 25774 22244 25846
rect 22032 25710 22174 25774
rect 22238 25710 22244 25774
rect 22032 25704 22244 25710
rect 26928 25774 27276 25916
rect 26928 25710 27206 25774
rect 27270 25710 27276 25774
rect 14200 25655 14520 25657
rect 14200 25652 14266 25655
rect 14454 25652 14520 25655
rect 20536 25644 20612 25704
rect 20944 25644 21020 25704
rect 13192 25586 13260 25642
rect 13316 25586 13404 25642
rect 13192 25568 13404 25586
rect 13239 25565 13337 25568
rect 1768 25508 1980 25544
rect 1224 25502 1980 25508
rect 1224 25438 1230 25502
rect 1294 25438 1980 25502
rect 1224 25432 1980 25438
rect 14286 25391 14370 25395
rect 14286 25386 14403 25391
rect 14286 25330 14342 25386
rect 14398 25330 14403 25386
rect 14286 25325 14403 25330
rect 14286 25321 14370 25325
rect 20400 25296 20612 25644
rect 20808 25366 21020 25644
rect 21080 25644 21156 25704
rect 21080 25568 21564 25644
rect 20808 25302 20814 25366
rect 20878 25302 21020 25366
rect 20808 25296 21020 25302
rect 21216 25366 21564 25568
rect 21216 25302 21358 25366
rect 21422 25302 21564 25366
rect 21216 25296 21564 25302
rect 21624 25502 21836 25508
rect 21624 25438 21766 25502
rect 21830 25438 21836 25502
rect 21624 25366 21836 25438
rect 21624 25302 21630 25366
rect 21694 25302 21836 25366
rect 21624 25296 21836 25302
rect 22032 25502 22244 25508
rect 22032 25438 22174 25502
rect 22238 25438 22244 25502
rect 22032 25366 22244 25438
rect 22032 25302 22038 25366
rect 22102 25302 22244 25366
rect 22032 25296 22244 25302
rect 26928 25432 27276 25710
rect 68952 25976 69164 26188
rect 73848 26318 74060 26324
rect 73848 26254 73854 26318
rect 73918 26254 74060 26318
rect 73848 26182 74060 26254
rect 73848 26118 73854 26182
rect 73918 26118 74060 26182
rect 73848 26112 74060 26118
rect 74256 26318 74468 26324
rect 74256 26254 74262 26318
rect 74326 26254 74468 26318
rect 74256 26182 74468 26254
rect 74256 26118 74262 26182
rect 74326 26118 74468 26182
rect 74256 26112 74468 26118
rect 74664 26318 75012 26324
rect 74664 26254 74670 26318
rect 74734 26254 74942 26318
rect 75006 26254 75012 26318
rect 74664 26248 75012 26254
rect 74664 26188 74876 26248
rect 75072 26188 75284 26324
rect 74664 26182 75284 26188
rect 74664 26118 75078 26182
rect 75142 26118 75284 26182
rect 74664 26112 75284 26118
rect 75480 26318 75692 26324
rect 75480 26254 75622 26318
rect 75686 26254 75692 26318
rect 75480 26112 75692 26254
rect 75616 26052 75692 26112
rect 68952 25916 69028 25976
rect 68952 25432 69164 25916
rect 73848 25910 74060 25916
rect 73848 25846 73854 25910
rect 73918 25846 74060 25910
rect 73848 25774 74060 25846
rect 73848 25710 73990 25774
rect 74054 25710 74060 25774
rect 73848 25704 74060 25710
rect 74256 25910 74468 25916
rect 74256 25846 74262 25910
rect 74326 25846 74468 25910
rect 74256 25774 74468 25846
rect 74256 25710 74262 25774
rect 74326 25710 74468 25774
rect 74256 25704 74468 25710
rect 74664 25704 74876 25916
rect 75072 25910 75284 25916
rect 75072 25846 75078 25910
rect 75142 25846 75284 25910
rect 75072 25704 75284 25846
rect 75480 25704 75692 26052
rect 74664 25644 74740 25704
rect 75072 25644 75148 25704
rect 75480 25644 75556 25704
rect 73848 25502 74060 25508
rect 73848 25438 73990 25502
rect 74054 25438 74060 25502
rect 26928 25372 27004 25432
rect 68952 25372 69028 25432
rect 20536 25236 20612 25296
rect 13600 25094 13812 25100
rect 13600 25030 13742 25094
rect 13806 25030 13812 25094
rect 13600 24964 13812 25030
rect 20400 25094 20612 25236
rect 26928 25160 27276 25372
rect 68952 25160 69164 25372
rect 73848 25366 74060 25438
rect 73848 25302 73854 25366
rect 73918 25302 74060 25366
rect 73848 25296 74060 25302
rect 74256 25502 74468 25508
rect 74256 25438 74262 25502
rect 74326 25438 74468 25502
rect 74256 25366 74468 25438
rect 74256 25302 74398 25366
rect 74462 25302 74468 25366
rect 74256 25296 74468 25302
rect 74664 25366 74876 25644
rect 75072 25372 75284 25644
rect 74974 25366 75284 25372
rect 74664 25302 74806 25366
rect 74870 25302 74876 25366
rect 74936 25302 74942 25366
rect 75006 25302 75284 25366
rect 74664 25296 74876 25302
rect 74974 25296 75284 25302
rect 75480 25296 75692 25644
rect 94112 25600 94324 25644
rect 94112 25544 94176 25600
rect 94232 25544 94324 25600
rect 94112 25508 94324 25544
rect 94112 25502 94732 25508
rect 94112 25438 94662 25502
rect 94726 25438 94732 25502
rect 94112 25432 94732 25438
rect 27064 25100 27140 25160
rect 69088 25100 69164 25160
rect 75480 25236 75556 25296
rect 20400 25030 20406 25094
rect 20470 25030 20612 25094
rect 20400 25024 20612 25030
rect 13600 24958 15580 24964
rect 13600 24894 15510 24958
rect 15574 24894 15580 24958
rect 13600 24888 15580 24894
rect 20808 24888 21020 25100
rect 21216 25094 21564 25100
rect 21216 25030 21358 25094
rect 21422 25030 21564 25094
rect 21216 24964 21564 25030
rect 21080 24888 21564 24964
rect 21624 25094 21836 25100
rect 21624 25030 21630 25094
rect 21694 25030 21836 25094
rect 21624 24888 21836 25030
rect 22032 25094 22244 25100
rect 22032 25030 22038 25094
rect 22102 25030 22244 25094
rect 22032 24888 22244 25030
rect 20808 24828 20884 24888
rect 21080 24828 21156 24888
rect 17000 24686 17212 24828
rect 17000 24622 17142 24686
rect 17206 24622 17212 24686
rect 17000 24616 17212 24622
rect 17408 24822 17620 24828
rect 17408 24758 17414 24822
rect 17478 24758 17620 24822
rect 17408 24692 17620 24758
rect 17816 24692 18028 24828
rect 17408 24686 18028 24692
rect 17408 24622 17958 24686
rect 18022 24622 18028 24686
rect 17408 24616 18028 24622
rect 18224 24550 18436 24828
rect 18224 24486 18366 24550
rect 18430 24486 18436 24550
rect 18224 24480 18436 24486
rect 18632 24556 18844 24828
rect 20400 24822 20612 24828
rect 20400 24758 20406 24822
rect 20470 24758 20612 24822
rect 20400 24686 20612 24758
rect 20400 24622 20542 24686
rect 20606 24622 20612 24686
rect 20400 24616 20612 24622
rect 20808 24752 21156 24828
rect 21216 24828 21292 24888
rect 21624 24828 21700 24888
rect 22032 24828 22108 24888
rect 20808 24616 21020 24752
rect 21216 24686 21564 24828
rect 21216 24622 21494 24686
rect 21558 24622 21564 24686
rect 21216 24616 21564 24622
rect 18632 24550 20884 24556
rect 18632 24486 18638 24550
rect 18702 24486 20814 24550
rect 20878 24486 20884 24550
rect 18632 24480 20884 24486
rect 21624 24480 21836 24828
rect 21760 24420 21836 24480
rect 20400 24414 20612 24420
rect 20400 24350 20542 24414
rect 20606 24350 20612 24414
rect 17310 24278 18300 24284
rect 17272 24214 17278 24278
rect 17342 24214 18230 24278
rect 18294 24214 18300 24278
rect 17310 24208 18300 24214
rect 20400 24278 20612 24350
rect 20400 24214 20406 24278
rect 20470 24214 20612 24278
rect 20400 24208 20612 24214
rect 18088 24072 18708 24148
rect 18088 24012 18164 24072
rect 18632 24012 18708 24072
rect 20808 24072 21020 24420
rect 21216 24414 21564 24420
rect 21216 24350 21494 24414
rect 21558 24350 21564 24414
rect 21216 24072 21564 24350
rect 21624 24278 21836 24420
rect 21624 24214 21630 24278
rect 21694 24214 21836 24278
rect 21624 24208 21836 24214
rect 22032 24480 22244 24828
rect 26928 24822 27276 25100
rect 26928 24758 26934 24822
rect 26998 24758 27276 24822
rect 26928 24752 27276 24758
rect 68952 24822 69164 25100
rect 68952 24758 68958 24822
rect 69022 24758 69164 24822
rect 68952 24752 69164 24758
rect 73848 25094 74060 25100
rect 73848 25030 73854 25094
rect 73918 25030 74060 25094
rect 73848 24888 74060 25030
rect 74256 25094 74468 25100
rect 74256 25030 74398 25094
rect 74462 25030 74468 25094
rect 74256 24888 74468 25030
rect 74664 25094 75012 25100
rect 74664 25030 74806 25094
rect 74870 25030 74942 25094
rect 75006 25030 75012 25094
rect 74664 25024 75012 25030
rect 74664 24964 74876 25024
rect 74664 24888 75012 24964
rect 73848 24828 73924 24888
rect 74256 24828 74332 24888
rect 74800 24828 74876 24888
rect 26928 24550 27276 24556
rect 26928 24486 26934 24550
rect 26998 24486 27276 24550
rect 22032 24420 22108 24480
rect 22032 24278 22244 24420
rect 22032 24214 22174 24278
rect 22238 24214 22244 24278
rect 22032 24208 22244 24214
rect 26928 24208 27276 24486
rect 68952 24550 69164 24556
rect 68952 24486 68958 24550
rect 69022 24486 69164 24550
rect 68952 24414 69164 24486
rect 73848 24480 74060 24828
rect 73984 24420 74060 24480
rect 68952 24350 68958 24414
rect 69022 24350 69164 24414
rect 68952 24208 69164 24350
rect 73848 24278 74060 24420
rect 73848 24214 73854 24278
rect 73918 24214 74060 24278
rect 73848 24208 74060 24214
rect 74256 24480 74468 24828
rect 74664 24686 74876 24828
rect 74936 24828 75012 24888
rect 75072 24888 75284 25100
rect 75480 25094 75692 25236
rect 75480 25030 75622 25094
rect 75686 25030 75692 25094
rect 75480 25024 75692 25030
rect 75072 24828 75148 24888
rect 74936 24752 75284 24828
rect 74664 24622 74670 24686
rect 74734 24622 74876 24686
rect 74664 24616 74876 24622
rect 75072 24616 75284 24752
rect 75480 24822 75692 24828
rect 75480 24758 75622 24822
rect 75686 24758 75692 24822
rect 75480 24686 75692 24758
rect 75480 24622 75486 24686
rect 75550 24622 75692 24686
rect 75480 24616 75692 24622
rect 77248 24550 77460 24828
rect 77248 24486 77254 24550
rect 77318 24486 77460 24550
rect 77248 24480 77460 24486
rect 77656 24550 77868 24828
rect 78064 24692 78276 24828
rect 78472 24692 78684 24828
rect 78064 24686 78684 24692
rect 78064 24622 78070 24686
rect 78134 24622 78684 24686
rect 78064 24616 78684 24622
rect 78880 24686 79228 24828
rect 78880 24622 79022 24686
rect 79086 24622 79228 24686
rect 78880 24616 79228 24622
rect 77656 24486 77798 24550
rect 77862 24486 77868 24550
rect 77656 24480 77868 24486
rect 74256 24420 74332 24480
rect 74256 24278 74468 24420
rect 74256 24214 74398 24278
rect 74462 24214 74468 24278
rect 74256 24208 74468 24214
rect 74664 24414 74876 24420
rect 74664 24350 74670 24414
rect 74734 24350 74876 24414
rect 20808 24012 20884 24072
rect 21488 24012 21564 24072
rect 26928 24148 27004 24208
rect 69088 24148 69164 24208
rect 1768 23920 1980 24012
rect 1768 23876 1818 23920
rect 1224 23870 1818 23876
rect 1224 23806 1230 23870
rect 1294 23864 1818 23870
rect 1874 23864 1980 23920
rect 1294 23806 1980 23864
rect 1224 23800 1980 23806
rect 17000 24006 17348 24012
rect 17000 23942 17142 24006
rect 17206 23942 17278 24006
rect 17342 23942 17348 24006
rect 17000 23936 17348 23942
rect 17000 23870 17212 23936
rect 17000 23806 17142 23870
rect 17206 23806 17212 23870
rect 17000 23800 17212 23806
rect 17408 23876 17620 24012
rect 17816 24006 18164 24012
rect 17816 23942 17958 24006
rect 18022 23942 18164 24006
rect 17816 23936 18164 23942
rect 18224 24006 18436 24012
rect 18224 23942 18230 24006
rect 18294 23942 18366 24006
rect 18430 23942 18436 24006
rect 17816 23876 18028 23936
rect 17408 23800 18028 23876
rect 18224 23870 18436 23942
rect 18224 23806 18366 23870
rect 18430 23806 18436 23870
rect 18224 23800 18436 23806
rect 18632 24006 18844 24012
rect 18632 23942 18638 24006
rect 18702 23942 18844 24006
rect 18632 23800 18844 23942
rect 20400 24006 20612 24012
rect 20400 23942 20406 24006
rect 20470 23942 20612 24006
rect 20400 23870 20612 23942
rect 20400 23806 20542 23870
rect 20606 23806 20612 23870
rect 20400 23800 20612 23806
rect 20808 23870 21020 24012
rect 20808 23806 20814 23870
rect 20878 23806 21020 23870
rect 20808 23800 21020 23806
rect 21216 23800 21564 24012
rect 21624 24006 21836 24012
rect 21624 23942 21630 24006
rect 21694 23942 21836 24006
rect 21624 23870 21836 23942
rect 21624 23806 21766 23870
rect 21830 23806 21836 23870
rect 21624 23800 21836 23806
rect 22032 24006 22244 24012
rect 22032 23942 22174 24006
rect 22238 23942 22244 24006
rect 22032 23870 22244 23942
rect 26928 24006 27276 24148
rect 26928 23942 27070 24006
rect 27134 23942 27276 24006
rect 26928 23936 27276 23942
rect 68952 24142 69164 24148
rect 68952 24078 68958 24142
rect 69022 24078 69164 24142
rect 68952 23936 69164 24078
rect 74664 24072 74876 24350
rect 75072 24148 75284 24420
rect 75480 24414 75692 24420
rect 75480 24350 75486 24414
rect 75550 24350 75692 24414
rect 75480 24278 75692 24350
rect 75480 24214 75622 24278
rect 75686 24214 75692 24278
rect 75480 24208 75692 24214
rect 74974 24142 75284 24148
rect 74936 24078 74942 24142
rect 75006 24078 75284 24142
rect 74974 24072 75284 24078
rect 77928 24072 78956 24148
rect 74800 24012 74876 24072
rect 77928 24012 78004 24072
rect 78880 24012 78956 24072
rect 27200 23876 27276 23936
rect 69088 23876 69164 23936
rect 22032 23806 22038 23870
rect 22102 23806 22244 23870
rect 22032 23800 22244 23806
rect 17544 23740 17620 23800
rect 21216 23740 21292 23800
rect 17544 23734 17892 23740
rect 17544 23670 17822 23734
rect 17886 23670 17892 23734
rect 17544 23664 17892 23670
rect 20944 23664 21292 23740
rect 20944 23604 21020 23664
rect 20400 23598 20612 23604
rect 20400 23534 20542 23598
rect 20606 23534 20612 23598
rect 544 23462 3476 23468
rect 544 23398 550 23462
rect 614 23398 3476 23462
rect 544 23392 3476 23398
rect 3128 23332 3476 23392
rect 3944 23332 4156 23468
rect 20400 23462 20612 23534
rect 20400 23398 20406 23462
rect 20470 23398 20612 23462
rect 20400 23392 20612 23398
rect 20808 23598 21564 23604
rect 20808 23534 20814 23598
rect 20878 23534 21564 23598
rect 20808 23528 21564 23534
rect 20808 23462 21020 23528
rect 20808 23398 20950 23462
rect 21014 23398 21020 23462
rect 20808 23392 21020 23398
rect 21216 23462 21564 23528
rect 21216 23398 21494 23462
rect 21558 23398 21564 23462
rect 21216 23392 21564 23398
rect 21624 23598 21836 23604
rect 21624 23534 21766 23598
rect 21830 23534 21836 23598
rect 21624 23462 21836 23534
rect 21624 23398 21766 23462
rect 21830 23398 21836 23462
rect 21624 23392 21836 23398
rect 22032 23598 22244 23604
rect 22032 23534 22038 23598
rect 22102 23534 22244 23598
rect 22032 23462 22244 23534
rect 22032 23398 22038 23462
rect 22102 23398 22244 23462
rect 22032 23392 22244 23398
rect 26928 23598 27276 23876
rect 26928 23534 27070 23598
rect 27134 23534 27276 23598
rect 26928 23392 27276 23534
rect 27200 23332 27276 23392
rect 3128 23256 4156 23332
rect 18088 23256 18708 23332
rect 18088 23196 18164 23256
rect 18632 23196 18708 23256
rect 17000 23190 17212 23196
rect 17000 23126 17142 23190
rect 17206 23126 17212 23190
rect 17000 23054 17212 23126
rect 17000 22990 17006 23054
rect 17070 22990 17212 23054
rect 17000 22984 17212 22990
rect 17408 23190 18164 23196
rect 17408 23126 17822 23190
rect 17886 23126 18164 23190
rect 17408 23120 18164 23126
rect 18224 23190 18436 23196
rect 18224 23126 18366 23190
rect 18430 23126 18436 23190
rect 17408 22984 17620 23120
rect 17816 23060 18028 23120
rect 17718 23054 18028 23060
rect 17680 22990 17686 23054
rect 17750 22990 18028 23054
rect 17718 22984 18028 22990
rect 18224 23054 18436 23126
rect 18224 22990 18366 23054
rect 18430 22990 18436 23054
rect 18224 22984 18436 22990
rect 18632 23054 18844 23196
rect 18632 22990 18774 23054
rect 18838 22990 18844 23054
rect 18632 22984 18844 22990
rect 20400 23190 20612 23196
rect 20400 23126 20406 23190
rect 20470 23126 20612 23190
rect 20400 23054 20612 23126
rect 20400 22990 20542 23054
rect 20606 22990 20612 23054
rect 20400 22984 20612 22990
rect 20808 23190 21020 23196
rect 20808 23126 20950 23190
rect 21014 23126 21020 23190
rect 20808 23054 21020 23126
rect 20808 22990 20814 23054
rect 20878 22990 21020 23054
rect 20808 22984 21020 22990
rect 21216 23190 21564 23196
rect 21216 23126 21494 23190
rect 21558 23126 21564 23190
rect 21216 22984 21564 23126
rect 21624 23190 21836 23196
rect 21624 23126 21766 23190
rect 21830 23126 21836 23190
rect 21624 23054 21836 23126
rect 21624 22990 21630 23054
rect 21694 22990 21836 23054
rect 21624 22984 21836 22990
rect 22032 23190 22244 23196
rect 22032 23126 22038 23190
rect 22102 23126 22244 23190
rect 22032 23054 22244 23126
rect 26928 23120 27276 23332
rect 68952 23598 69164 23876
rect 73848 24006 74060 24012
rect 73848 23942 73854 24006
rect 73918 23942 74060 24006
rect 73848 23870 74060 23942
rect 73848 23806 73990 23870
rect 74054 23806 74060 23870
rect 73848 23800 74060 23806
rect 74256 24006 74468 24012
rect 74256 23942 74398 24006
rect 74462 23942 74468 24006
rect 74256 23870 74468 23942
rect 74256 23806 74398 23870
rect 74462 23806 74468 23870
rect 74256 23800 74468 23806
rect 74664 23936 75284 24012
rect 74664 23876 74876 23936
rect 74664 23870 75012 23876
rect 74664 23806 74942 23870
rect 75006 23806 75012 23870
rect 74664 23800 75012 23806
rect 75072 23870 75284 23936
rect 75072 23806 75214 23870
rect 75278 23806 75284 23870
rect 75072 23800 75284 23806
rect 75480 24006 75692 24012
rect 75480 23942 75622 24006
rect 75686 23942 75692 24006
rect 75480 23870 75692 23942
rect 75480 23806 75486 23870
rect 75550 23806 75692 23870
rect 75480 23800 75692 23806
rect 77248 24006 77460 24012
rect 77248 23942 77254 24006
rect 77318 23942 77460 24006
rect 77248 23876 77460 23942
rect 77656 24006 78004 24012
rect 77656 23942 77798 24006
rect 77862 23942 78004 24006
rect 77656 23936 78004 23942
rect 78064 24006 78684 24012
rect 78064 23942 78070 24006
rect 78134 23942 78684 24006
rect 78064 23936 78684 23942
rect 77248 23800 77596 23876
rect 77656 23870 77868 23936
rect 77656 23806 77662 23870
rect 77726 23806 77798 23870
rect 77862 23806 77868 23870
rect 77656 23800 77868 23806
rect 78064 23876 78276 23936
rect 78064 23870 78412 23876
rect 78064 23806 78342 23870
rect 78406 23806 78412 23870
rect 78064 23800 78412 23806
rect 78472 23800 78684 23936
rect 78880 24006 79228 24012
rect 78880 23942 79022 24006
rect 79086 23942 79228 24006
rect 78880 23870 79228 23942
rect 78880 23806 79022 23870
rect 79086 23806 79228 23870
rect 78880 23800 79228 23806
rect 94112 23920 94324 24012
rect 94112 23864 94176 23920
rect 94232 23876 94324 23920
rect 94232 23870 94732 23876
rect 94232 23864 94662 23870
rect 94112 23806 94662 23864
rect 94726 23806 94732 23870
rect 94112 23800 94732 23806
rect 77520 23740 77596 23800
rect 78064 23740 78140 23800
rect 77520 23664 78140 23740
rect 68952 23534 68958 23598
rect 69022 23534 69164 23598
rect 68952 23392 69164 23534
rect 73848 23598 74060 23604
rect 73848 23534 73990 23598
rect 74054 23534 74060 23598
rect 73848 23468 74060 23534
rect 74256 23598 74468 23604
rect 74256 23534 74398 23598
rect 74462 23534 74468 23598
rect 73848 23462 74196 23468
rect 73848 23398 73990 23462
rect 74054 23398 74196 23462
rect 73848 23392 74196 23398
rect 74256 23462 74468 23534
rect 74256 23398 74262 23462
rect 74326 23398 74468 23462
rect 74256 23392 74468 23398
rect 74664 23462 74876 23604
rect 74664 23398 74806 23462
rect 74870 23398 74876 23462
rect 74664 23392 74876 23398
rect 75072 23598 75284 23604
rect 75072 23534 75214 23598
rect 75278 23534 75284 23598
rect 75072 23392 75284 23534
rect 75480 23598 75692 23604
rect 75480 23534 75486 23598
rect 75550 23534 75692 23598
rect 75480 23462 75692 23534
rect 75480 23398 75486 23462
rect 75550 23398 75692 23462
rect 75480 23392 75692 23398
rect 68952 23332 69028 23392
rect 74120 23332 74196 23392
rect 74664 23332 74740 23392
rect 75072 23332 75148 23392
rect 68952 23326 69164 23332
rect 68952 23262 68958 23326
rect 69022 23262 69164 23326
rect 68952 23120 69164 23262
rect 74120 23256 74740 23332
rect 74800 23256 75148 23332
rect 77112 23326 77732 23332
rect 77112 23262 77662 23326
rect 77726 23262 77732 23326
rect 77112 23256 77732 23262
rect 74800 23196 74876 23256
rect 77112 23196 77188 23256
rect 27064 23060 27140 23120
rect 69088 23060 69164 23120
rect 22032 22990 22038 23054
rect 22102 22990 22244 23054
rect 22032 22984 22244 22990
rect 26928 22848 27276 23060
rect 68952 22848 69164 23060
rect 73848 23190 74060 23196
rect 73848 23126 73990 23190
rect 74054 23126 74060 23190
rect 73848 23054 74060 23126
rect 73848 22990 73854 23054
rect 73918 22990 74060 23054
rect 73848 22984 74060 22990
rect 74256 23190 74468 23196
rect 74256 23126 74262 23190
rect 74326 23126 74468 23190
rect 74256 23054 74468 23126
rect 74256 22990 74398 23054
rect 74462 22990 74468 23054
rect 74256 22984 74468 22990
rect 74664 23190 75284 23196
rect 74664 23126 74806 23190
rect 74870 23126 75284 23190
rect 74664 23120 75284 23126
rect 74664 22984 74876 23120
rect 75072 23054 75284 23120
rect 75072 22990 75214 23054
rect 75278 22990 75284 23054
rect 75072 22984 75284 22990
rect 75480 23190 77188 23196
rect 75480 23126 75486 23190
rect 75550 23126 77188 23190
rect 75480 23120 77188 23126
rect 75480 23054 75692 23120
rect 75480 22990 75622 23054
rect 75686 22990 75692 23054
rect 75480 22984 75692 22990
rect 77248 23060 77460 23196
rect 77656 23190 77868 23196
rect 77656 23126 77798 23190
rect 77862 23126 77868 23190
rect 77248 23054 77596 23060
rect 77248 22990 77254 23054
rect 77318 22990 77596 23054
rect 77248 22984 77596 22990
rect 77656 23054 77868 23126
rect 77656 22990 77798 23054
rect 77862 22990 77868 23054
rect 77656 22984 77868 22990
rect 78064 23060 78276 23196
rect 78374 23190 78684 23196
rect 78336 23126 78342 23190
rect 78406 23126 78684 23190
rect 78374 23120 78684 23126
rect 78472 23060 78684 23120
rect 78064 23054 78684 23060
rect 78064 22990 78614 23054
rect 78678 22990 78684 23054
rect 78064 22984 78684 22990
rect 78880 23190 79228 23196
rect 78880 23126 79022 23190
rect 79086 23126 79228 23190
rect 78880 23054 79228 23126
rect 78880 22990 78886 23054
rect 78950 22990 79228 23054
rect 78880 22984 79228 22990
rect 77520 22924 77596 22984
rect 78064 22924 78140 22984
rect 77520 22848 78140 22924
rect 26928 22788 27004 22848
rect 69088 22788 69164 22848
rect 20400 22782 20612 22788
rect 20400 22718 20542 22782
rect 20606 22718 20612 22782
rect 2560 22669 2626 22670
rect 2518 22605 2561 22669
rect 2625 22605 2668 22669
rect 20400 22646 20612 22718
rect 2560 22604 2626 22605
rect 20400 22582 20406 22646
rect 20470 22582 20612 22646
rect 20400 22576 20612 22582
rect 20808 22782 21020 22788
rect 20808 22718 20814 22782
rect 20878 22718 21020 22782
rect 20808 22652 21020 22718
rect 21216 22652 21564 22788
rect 20808 22576 21564 22652
rect 21624 22782 21836 22788
rect 21624 22718 21630 22782
rect 21694 22718 21836 22782
rect 21624 22646 21836 22718
rect 21624 22582 21766 22646
rect 21830 22582 21836 22646
rect 21624 22576 21836 22582
rect 22032 22782 22244 22788
rect 22032 22718 22038 22782
rect 22102 22718 22244 22782
rect 22032 22646 22244 22718
rect 22032 22582 22038 22646
rect 22102 22582 22244 22646
rect 22032 22576 22244 22582
rect 26928 22576 27276 22788
rect 68952 22576 69164 22788
rect 73848 22782 74060 22788
rect 73848 22718 73854 22782
rect 73918 22718 74060 22782
rect 73848 22646 74060 22718
rect 73848 22582 73990 22646
rect 74054 22582 74060 22646
rect 73848 22576 74060 22582
rect 74256 22782 74468 22788
rect 74256 22718 74398 22782
rect 74462 22718 74468 22782
rect 74256 22646 74468 22718
rect 74256 22582 74262 22646
rect 74326 22582 74468 22646
rect 74256 22576 74468 22582
rect 74664 22646 74876 22788
rect 74664 22582 74670 22646
rect 74734 22582 74876 22646
rect 74664 22576 74876 22582
rect 75072 22782 75284 22788
rect 75072 22718 75214 22782
rect 75278 22718 75284 22782
rect 75072 22646 75284 22718
rect 75072 22582 75078 22646
rect 75142 22582 75284 22646
rect 75072 22576 75284 22582
rect 75480 22782 75692 22788
rect 75480 22718 75622 22782
rect 75686 22718 75692 22782
rect 75480 22646 75692 22718
rect 75480 22582 75486 22646
rect 75550 22582 75692 22646
rect 75480 22576 75692 22582
rect 21216 22516 21292 22576
rect 27064 22516 27140 22576
rect 68952 22516 69028 22576
rect 16864 22440 17484 22516
rect 16864 22380 16940 22440
rect 17408 22380 17484 22440
rect 20944 22440 21292 22516
rect 20944 22380 21020 22440
rect 1768 22244 1980 22380
rect 1224 22240 1980 22244
rect 1224 22238 1818 22240
rect 1224 22174 1230 22238
rect 1294 22184 1818 22238
rect 1874 22184 1980 22240
rect 1294 22174 1980 22184
rect 1224 22168 1980 22174
rect 15504 22374 15716 22380
rect 15504 22310 15510 22374
rect 15574 22310 15716 22374
rect 15504 22244 15716 22310
rect 15912 22304 16940 22380
rect 17000 22374 17212 22380
rect 17000 22310 17006 22374
rect 17070 22310 17212 22374
rect 15504 22168 15852 22244
rect 15912 22168 16124 22304
rect 17000 22244 17212 22310
rect 17408 22374 17756 22380
rect 17408 22310 17686 22374
rect 17750 22310 17756 22374
rect 17408 22304 17756 22310
rect 17408 22244 17620 22304
rect 17816 22244 18028 22380
rect 17000 22238 17348 22244
rect 17000 22174 17278 22238
rect 17342 22174 17348 22238
rect 17000 22168 17348 22174
rect 17408 22168 18028 22244
rect 18224 22374 18436 22380
rect 18224 22310 18366 22374
rect 18430 22310 18436 22374
rect 18224 22244 18436 22310
rect 18632 22374 18844 22380
rect 18632 22310 18774 22374
rect 18838 22310 18844 22374
rect 18224 22238 18572 22244
rect 18224 22174 18502 22238
rect 18566 22174 18572 22238
rect 18224 22168 18572 22174
rect 18632 22238 18844 22310
rect 18632 22174 18638 22238
rect 18702 22174 18844 22238
rect 18632 22168 18844 22174
rect 20400 22374 20612 22380
rect 20400 22310 20406 22374
rect 20470 22310 20612 22374
rect 20400 22168 20612 22310
rect 20808 22304 21564 22380
rect 20808 22238 21020 22304
rect 20808 22174 20814 22238
rect 20878 22174 21020 22238
rect 20808 22168 21020 22174
rect 21216 22238 21564 22304
rect 21216 22174 21494 22238
rect 21558 22174 21564 22238
rect 21216 22168 21564 22174
rect 21624 22374 21836 22380
rect 21624 22310 21766 22374
rect 21830 22310 21836 22374
rect 21624 22238 21836 22310
rect 21624 22174 21766 22238
rect 21830 22174 21836 22238
rect 21624 22168 21836 22174
rect 22032 22374 22244 22380
rect 22032 22310 22038 22374
rect 22102 22310 22244 22374
rect 22032 22238 22244 22310
rect 22032 22174 22174 22238
rect 22238 22174 22244 22238
rect 22032 22168 22244 22174
rect 26928 22304 27276 22516
rect 68952 22304 69164 22516
rect 78744 22440 80044 22516
rect 78744 22380 78820 22440
rect 79968 22380 80044 22440
rect 73848 22374 74060 22380
rect 73848 22310 73990 22374
rect 74054 22310 74060 22374
rect 26928 22244 27004 22304
rect 68952 22244 69028 22304
rect 1768 22108 1980 22168
rect 15776 22108 15852 22168
rect 17000 22108 17076 22168
rect 20536 22108 20612 22168
rect 1768 22032 3204 22108
rect 15776 22032 17076 22108
rect 3128 21972 3204 22032
rect 3128 21896 4156 21972
rect 3128 21760 3476 21896
rect 3944 21760 4156 21896
rect 20400 21760 20612 22108
rect 26928 22102 27276 22244
rect 26928 22038 26934 22102
rect 26998 22038 27276 22102
rect 26928 22032 27276 22038
rect 68952 22032 69164 22244
rect 73848 22238 74060 22310
rect 73848 22174 73854 22238
rect 73918 22174 74060 22238
rect 73848 22168 74060 22174
rect 74256 22374 74468 22380
rect 74256 22310 74262 22374
rect 74326 22310 74468 22374
rect 74256 22238 74468 22310
rect 74256 22174 74262 22238
rect 74326 22174 74468 22238
rect 74256 22168 74468 22174
rect 74664 22374 74876 22380
rect 74664 22310 74670 22374
rect 74734 22310 74876 22374
rect 74664 22238 74876 22310
rect 75072 22374 75284 22380
rect 75072 22310 75078 22374
rect 75142 22310 75284 22374
rect 75072 22244 75284 22310
rect 74974 22238 75284 22244
rect 74664 22174 74806 22238
rect 74870 22174 74876 22238
rect 74936 22174 74942 22238
rect 75006 22174 75214 22238
rect 75278 22174 75284 22238
rect 74664 22168 74876 22174
rect 74974 22168 75284 22174
rect 75480 22374 75692 22380
rect 75480 22310 75486 22374
rect 75550 22310 75692 22374
rect 75480 22168 75692 22310
rect 77248 22374 77460 22380
rect 77248 22310 77254 22374
rect 77318 22310 77460 22374
rect 77248 22238 77460 22310
rect 77248 22174 77390 22238
rect 77454 22174 77460 22238
rect 77248 22168 77460 22174
rect 77656 22374 77868 22380
rect 77656 22310 77798 22374
rect 77862 22310 77868 22374
rect 77656 22244 77868 22310
rect 78064 22244 78276 22380
rect 78472 22374 78820 22380
rect 78472 22310 78614 22374
rect 78678 22310 78820 22374
rect 78472 22304 78820 22310
rect 78880 22374 79228 22380
rect 78880 22310 78886 22374
rect 78950 22310 79228 22374
rect 78472 22244 78684 22304
rect 77656 22168 78004 22244
rect 78064 22168 78684 22244
rect 78880 22244 79228 22310
rect 78880 22168 79908 22244
rect 79968 22168 80180 22380
rect 80376 22168 80588 22380
rect 94112 22374 94732 22380
rect 94112 22310 94662 22374
rect 94726 22310 94732 22374
rect 94112 22304 94732 22310
rect 94112 22240 94324 22304
rect 94112 22184 94176 22240
rect 94232 22184 94324 22240
rect 27064 21972 27140 22032
rect 69088 21972 69164 22032
rect 75480 22108 75556 22168
rect 77928 22108 78004 22168
rect 79832 22108 79908 22168
rect 80376 22108 80452 22168
rect 20808 21966 21020 21972
rect 20808 21902 20814 21966
rect 20878 21902 21020 21966
rect 20808 21760 21020 21902
rect 21216 21966 21564 21972
rect 21216 21902 21494 21966
rect 21558 21902 21564 21966
rect 21216 21760 21564 21902
rect 21624 21966 21836 21972
rect 21624 21902 21766 21966
rect 21830 21902 21836 21966
rect 21624 21830 21836 21902
rect 21624 21766 21766 21830
rect 21830 21766 21836 21830
rect 21624 21760 21836 21766
rect 22032 21966 22244 21972
rect 22032 21902 22174 21966
rect 22238 21902 22244 21966
rect 22032 21830 22244 21902
rect 22032 21766 22038 21830
rect 22102 21766 22244 21830
rect 22032 21760 22244 21766
rect 26928 21830 27276 21972
rect 26928 21766 26934 21830
rect 26998 21766 27276 21830
rect 20536 21700 20612 21760
rect 20944 21700 21020 21760
rect 21488 21700 21564 21760
rect 18534 21694 20612 21700
rect 18496 21630 18502 21694
rect 18566 21630 20612 21694
rect 18534 21624 20612 21630
rect 20400 21352 20612 21624
rect 20808 21428 21020 21700
rect 20808 21422 21156 21428
rect 20808 21358 21086 21422
rect 21150 21358 21156 21422
rect 20808 21352 21156 21358
rect 21216 21352 21564 21700
rect 21624 21558 21836 21564
rect 21624 21494 21766 21558
rect 21830 21494 21836 21558
rect 21624 21422 21836 21494
rect 21624 21358 21766 21422
rect 21830 21358 21836 21422
rect 21624 21352 21836 21358
rect 22032 21558 22244 21564
rect 22032 21494 22038 21558
rect 22102 21494 22244 21558
rect 22032 21422 22244 21494
rect 26928 21488 27276 21766
rect 68952 21830 69164 21972
rect 68952 21766 69094 21830
rect 69158 21766 69164 21830
rect 68952 21558 69164 21766
rect 73848 21966 74060 21972
rect 73848 21902 73854 21966
rect 73918 21902 74060 21966
rect 73848 21830 74060 21902
rect 73848 21766 73854 21830
rect 73918 21766 74060 21830
rect 73848 21760 74060 21766
rect 74256 21966 74468 21972
rect 74256 21902 74262 21966
rect 74326 21902 74468 21966
rect 74256 21830 74468 21902
rect 74256 21766 74398 21830
rect 74462 21766 74468 21830
rect 74256 21760 74468 21766
rect 74664 21966 75012 21972
rect 74664 21902 74806 21966
rect 74870 21902 74942 21966
rect 75006 21902 75012 21966
rect 74664 21896 75012 21902
rect 75072 21966 75284 21972
rect 75072 21902 75214 21966
rect 75278 21902 75284 21966
rect 74664 21760 74876 21896
rect 75072 21760 75284 21902
rect 75208 21700 75284 21760
rect 68952 21494 68958 21558
rect 69022 21494 69164 21558
rect 68952 21488 69164 21494
rect 73848 21558 74060 21564
rect 73848 21494 73854 21558
rect 73918 21494 74060 21558
rect 27200 21428 27276 21488
rect 22032 21358 22038 21422
rect 22102 21358 22244 21422
rect 22032 21352 22244 21358
rect 20536 21292 20612 21352
rect 20400 21150 20612 21292
rect 26928 21216 27276 21428
rect 68952 21422 69164 21428
rect 68952 21358 69094 21422
rect 69158 21358 69164 21422
rect 68952 21216 69164 21358
rect 73848 21422 74060 21494
rect 73848 21358 73990 21422
rect 74054 21358 74060 21422
rect 73848 21352 74060 21358
rect 74256 21558 74468 21564
rect 74256 21494 74398 21558
rect 74462 21494 74468 21558
rect 74256 21422 74468 21494
rect 74256 21358 74398 21422
rect 74462 21358 74468 21422
rect 74256 21352 74468 21358
rect 74664 21428 74876 21700
rect 75072 21428 75284 21700
rect 74664 21422 75284 21428
rect 74664 21358 75078 21422
rect 75142 21358 75284 21422
rect 74664 21352 75284 21358
rect 75480 21760 75692 22108
rect 77928 22102 78548 22108
rect 77928 22038 78478 22102
rect 78542 22038 78548 22102
rect 77928 22032 78548 22038
rect 79832 22032 80452 22108
rect 94112 22032 94324 22184
rect 75480 21700 75556 21760
rect 75480 21352 75692 21700
rect 75480 21292 75556 21352
rect 27064 21156 27140 21216
rect 68952 21156 69028 21216
rect 20400 21086 20542 21150
rect 20606 21086 20612 21150
rect 20400 21080 20612 21086
rect 17680 20944 18300 21020
rect 17680 20884 17756 20944
rect 18224 20884 18300 20944
rect 20808 20944 21020 21156
rect 21118 21150 21564 21156
rect 21080 21086 21086 21150
rect 21150 21086 21564 21150
rect 21118 21080 21564 21086
rect 21216 20944 21564 21080
rect 21624 21150 21836 21156
rect 21624 21086 21766 21150
rect 21830 21086 21836 21150
rect 21624 20944 21836 21086
rect 22032 21150 22244 21156
rect 22032 21086 22038 21150
rect 22102 21086 22244 21150
rect 22032 20944 22244 21086
rect 20808 20884 20884 20944
rect 21352 20884 21428 20944
rect 21624 20884 21700 20944
rect 22032 20884 22108 20944
rect 17310 20878 17756 20884
rect 17272 20814 17278 20878
rect 17342 20814 17756 20878
rect 17310 20808 17756 20814
rect 17408 20612 17620 20808
rect 1768 20560 1980 20612
rect 1768 20504 1818 20560
rect 1874 20504 1980 20560
rect 1768 20476 1980 20504
rect 1224 20470 1980 20476
rect 1224 20406 1230 20470
rect 1294 20406 1980 20470
rect 1224 20400 1980 20406
rect 3128 20536 4156 20612
rect 16494 20606 17620 20612
rect 16456 20542 16462 20606
rect 16526 20542 17414 20606
rect 17478 20542 17620 20606
rect 16494 20536 17620 20542
rect 17816 20612 18028 20884
rect 17816 20606 18164 20612
rect 17816 20542 17822 20606
rect 17886 20542 18164 20606
rect 17816 20536 18164 20542
rect 18224 20606 18436 20884
rect 18224 20542 18366 20606
rect 18430 20542 18436 20606
rect 18224 20536 18436 20542
rect 18632 20878 18844 20884
rect 18632 20814 18638 20878
rect 18702 20814 18844 20878
rect 18632 20606 18844 20814
rect 20400 20878 20612 20884
rect 20400 20814 20542 20878
rect 20606 20814 20612 20878
rect 20400 20742 20612 20814
rect 20400 20678 20406 20742
rect 20470 20678 20612 20742
rect 20400 20672 20612 20678
rect 20808 20808 21564 20884
rect 20808 20672 21020 20808
rect 21216 20742 21564 20808
rect 21216 20678 21494 20742
rect 21558 20678 21564 20742
rect 21216 20672 21564 20678
rect 18632 20542 18774 20606
rect 18838 20542 18844 20606
rect 18632 20536 18844 20542
rect 21624 20536 21836 20884
rect 22032 20536 22244 20884
rect 26928 20878 27276 21156
rect 26928 20814 27206 20878
rect 27270 20814 27276 20878
rect 26928 20808 27276 20814
rect 68952 21150 69164 21156
rect 68952 21086 68958 21150
rect 69022 21086 69164 21150
rect 68952 20878 69164 21086
rect 68952 20814 69094 20878
rect 69158 20814 69164 20878
rect 68952 20808 69164 20814
rect 73848 21150 74060 21156
rect 73848 21086 73990 21150
rect 74054 21086 74060 21150
rect 73848 20944 74060 21086
rect 74256 21150 74468 21156
rect 74256 21086 74398 21150
rect 74462 21086 74468 21150
rect 74256 20944 74468 21086
rect 74664 21020 74876 21156
rect 75072 21150 75284 21156
rect 75072 21086 75078 21150
rect 75142 21086 75284 21150
rect 74664 20944 75012 21020
rect 75072 20944 75284 21086
rect 75480 21150 75692 21292
rect 75480 21086 75486 21150
rect 75550 21086 75692 21150
rect 75480 21080 75692 21086
rect 73848 20884 73924 20944
rect 74256 20884 74332 20944
rect 74800 20884 74876 20944
rect 3128 20400 3476 20536
rect 3944 20476 4156 20536
rect 3846 20470 4156 20476
rect 3808 20406 3814 20470
rect 3878 20406 4156 20470
rect 3846 20400 4156 20406
rect 18088 20476 18164 20536
rect 18632 20476 18708 20536
rect 21624 20476 21700 20536
rect 22032 20476 22108 20536
rect 18088 20400 18708 20476
rect 20400 20470 20612 20476
rect 20400 20406 20406 20470
rect 20470 20406 20612 20470
rect 20400 20334 20612 20406
rect 20400 20270 20406 20334
rect 20470 20270 20612 20334
rect 20400 20264 20612 20270
rect 17272 20128 17892 20204
rect 20808 20128 21020 20476
rect 21216 20470 21564 20476
rect 21216 20406 21494 20470
rect 21558 20406 21564 20470
rect 21216 20128 21564 20406
rect 21624 20128 21836 20476
rect 22032 20128 22244 20476
rect 17272 20068 17348 20128
rect 17816 20068 17892 20128
rect 20944 20068 21020 20128
rect 21352 20068 21428 20128
rect 21624 20068 21700 20128
rect 22168 20068 22244 20128
rect 16184 20062 16532 20068
rect 16184 19998 16462 20062
rect 16526 19998 16532 20062
rect 16184 19992 16532 19998
rect 16592 19992 17348 20068
rect 17408 20062 17620 20068
rect 17408 19998 17414 20062
rect 17478 19998 17620 20062
rect 16184 19856 16396 19992
rect 16592 19856 16804 19992
rect 17408 19856 17620 19998
rect 17816 20062 18028 20068
rect 17816 19998 17822 20062
rect 17886 19998 18028 20062
rect 17816 19856 18028 19998
rect 18224 20062 18436 20068
rect 18224 19998 18366 20062
rect 18430 19998 18436 20062
rect 18224 19926 18436 19998
rect 18224 19862 18230 19926
rect 18294 19862 18436 19926
rect 18224 19856 18436 19862
rect 18632 20062 18844 20068
rect 18632 19998 18774 20062
rect 18838 19998 18844 20062
rect 18632 19926 18844 19998
rect 18632 19862 18638 19926
rect 18702 19862 18844 19926
rect 18632 19856 18844 19862
rect 20400 20062 20612 20068
rect 20400 19998 20406 20062
rect 20470 19998 20612 20062
rect 20400 19926 20612 19998
rect 20400 19862 20406 19926
rect 20470 19862 20612 19926
rect 20400 19856 20612 19862
rect 20808 19926 21020 20068
rect 20808 19862 20814 19926
rect 20878 19862 21020 19926
rect 20808 19856 21020 19862
rect 21216 19926 21564 20068
rect 21216 19862 21494 19926
rect 21558 19862 21564 19926
rect 21216 19856 21564 19862
rect 21624 19926 21836 20068
rect 21624 19862 21630 19926
rect 21694 19862 21836 19926
rect 21624 19856 21836 19862
rect 22032 19926 22244 20068
rect 22032 19862 22038 19926
rect 22102 19862 22244 19926
rect 22032 19856 22244 19862
rect 26928 20470 27276 20612
rect 26928 20406 26934 20470
rect 26998 20406 27206 20470
rect 27270 20406 27276 20470
rect 26928 20198 27276 20406
rect 26928 20134 26934 20198
rect 26998 20134 27070 20198
rect 27134 20134 27276 20198
rect 26928 19992 27276 20134
rect 68952 20606 69164 20612
rect 68952 20542 69094 20606
rect 69158 20542 69164 20606
rect 68952 20062 69164 20542
rect 68952 19998 69094 20062
rect 69158 19998 69164 20062
rect 68952 19992 69164 19998
rect 73848 20536 74060 20884
rect 74256 20536 74468 20884
rect 74664 20742 74876 20884
rect 74936 20884 75012 20944
rect 75208 20884 75284 20944
rect 77928 20944 78548 21020
rect 77928 20884 78004 20944
rect 78472 20884 78548 20944
rect 74936 20808 75284 20884
rect 74664 20678 74670 20742
rect 74734 20678 74876 20742
rect 74664 20672 74876 20678
rect 75072 20672 75284 20808
rect 75480 20878 75692 20884
rect 75480 20814 75486 20878
rect 75550 20814 75692 20878
rect 75480 20742 75692 20814
rect 75480 20678 75486 20742
rect 75550 20678 75692 20742
rect 75480 20672 75692 20678
rect 77248 20878 77460 20884
rect 77248 20814 77390 20878
rect 77454 20814 77460 20878
rect 77248 20612 77460 20814
rect 77656 20808 78004 20884
rect 77248 20536 77596 20612
rect 77656 20606 77868 20808
rect 77656 20542 77662 20606
rect 77726 20542 77868 20606
rect 77656 20536 77868 20542
rect 78064 20612 78276 20884
rect 78472 20878 78684 20884
rect 78472 20814 78478 20878
rect 78542 20814 78684 20878
rect 78064 20606 78412 20612
rect 78064 20542 78206 20606
rect 78270 20542 78412 20606
rect 78064 20536 78412 20542
rect 78472 20606 78684 20814
rect 78472 20542 78614 20606
rect 78678 20542 78684 20606
rect 78472 20536 78684 20542
rect 94112 20560 94324 20612
rect 73848 20476 73924 20536
rect 74256 20476 74332 20536
rect 77520 20476 77596 20536
rect 78064 20476 78140 20536
rect 73848 20128 74060 20476
rect 74256 20128 74468 20476
rect 74664 20470 75284 20476
rect 74664 20406 74670 20470
rect 74734 20406 75284 20470
rect 74664 20400 75284 20406
rect 74664 20128 74876 20400
rect 75072 20204 75284 20400
rect 75480 20470 75692 20476
rect 75480 20406 75486 20470
rect 75550 20406 75692 20470
rect 75480 20334 75692 20406
rect 77520 20400 78140 20476
rect 78336 20476 78412 20536
rect 94112 20504 94176 20560
rect 94232 20504 94324 20560
rect 94112 20476 94324 20504
rect 78336 20470 79500 20476
rect 78336 20406 79430 20470
rect 79494 20406 79500 20470
rect 78336 20400 79500 20406
rect 94112 20470 94732 20476
rect 94112 20406 94662 20470
rect 94726 20406 94732 20470
rect 94112 20400 94732 20406
rect 75480 20270 75486 20334
rect 75550 20270 75692 20334
rect 75480 20264 75692 20270
rect 74936 20128 75284 20204
rect 79288 20128 79908 20204
rect 73848 20068 73924 20128
rect 74256 20068 74332 20128
rect 74936 20068 75012 20128
rect 79288 20068 79364 20128
rect 79832 20068 79908 20128
rect 26928 19932 27004 19992
rect 68952 19932 69028 19992
rect 26928 19926 27276 19932
rect 26928 19862 27070 19926
rect 27134 19862 27276 19926
rect 20400 19654 20612 19660
rect 20400 19590 20406 19654
rect 20470 19590 20612 19654
rect 20400 19518 20612 19590
rect 20400 19454 20406 19518
rect 20470 19454 20612 19518
rect 20400 19448 20612 19454
rect 20808 19654 21020 19660
rect 20808 19590 20814 19654
rect 20878 19590 21020 19654
rect 20808 19518 21020 19590
rect 20808 19454 20950 19518
rect 21014 19454 21020 19518
rect 20808 19448 21020 19454
rect 21216 19654 21564 19660
rect 21216 19590 21494 19654
rect 21558 19590 21564 19654
rect 21216 19448 21564 19590
rect 21624 19654 21836 19660
rect 21624 19590 21630 19654
rect 21694 19590 21836 19654
rect 21624 19518 21836 19590
rect 21624 19454 21630 19518
rect 21694 19454 21836 19518
rect 21624 19448 21836 19454
rect 22032 19654 22244 19660
rect 22032 19590 22038 19654
rect 22102 19590 22244 19654
rect 22032 19518 22244 19590
rect 22032 19454 22174 19518
rect 22238 19454 22244 19518
rect 22032 19448 22244 19454
rect 26928 19448 27276 19862
rect 68952 19654 69164 19932
rect 73848 19926 74060 20068
rect 73848 19862 73854 19926
rect 73918 19862 74060 19926
rect 73848 19856 74060 19862
rect 74256 19926 74468 20068
rect 74256 19862 74262 19926
rect 74326 19862 74468 19926
rect 74256 19856 74468 19862
rect 74664 19992 75012 20068
rect 74664 19932 74876 19992
rect 75072 19932 75284 20068
rect 74664 19856 75284 19932
rect 75480 20062 75692 20068
rect 75480 19998 75486 20062
rect 75550 19998 75692 20062
rect 75480 19926 75692 19998
rect 75480 19862 75622 19926
rect 75686 19862 75692 19926
rect 75480 19856 75692 19862
rect 77248 19932 77460 20068
rect 77656 20062 77868 20068
rect 77656 19998 77662 20062
rect 77726 19998 77868 20062
rect 77248 19856 77596 19932
rect 77656 19856 77868 19998
rect 78064 20062 78276 20068
rect 78064 19998 78206 20062
rect 78270 19998 78276 20062
rect 78064 19926 78276 19998
rect 78064 19862 78206 19926
rect 78270 19862 78276 19926
rect 78064 19856 78276 19862
rect 78472 20062 79364 20068
rect 78472 19998 78614 20062
rect 78678 19998 79364 20062
rect 78472 19992 79364 19998
rect 79424 20062 79636 20068
rect 79424 19998 79430 20062
rect 79494 19998 79636 20062
rect 78472 19926 78684 19992
rect 78472 19862 78614 19926
rect 78678 19862 78684 19926
rect 78472 19856 78684 19862
rect 79424 19856 79636 19998
rect 79832 19856 80044 20068
rect 74800 19796 74876 19856
rect 77248 19796 77324 19856
rect 74800 19720 75148 19796
rect 75072 19660 75148 19720
rect 75344 19720 77324 19796
rect 77520 19796 77596 19856
rect 78064 19796 78140 19856
rect 77520 19720 78140 19796
rect 75344 19660 75420 19720
rect 68952 19590 69094 19654
rect 69158 19590 69164 19654
rect 68952 19448 69164 19590
rect 73848 19654 74060 19660
rect 73848 19590 73854 19654
rect 73918 19590 74060 19654
rect 73848 19518 74060 19590
rect 73848 19454 73854 19518
rect 73918 19454 74060 19518
rect 73848 19448 74060 19454
rect 74256 19654 74468 19660
rect 74256 19590 74262 19654
rect 74326 19590 74468 19654
rect 74256 19518 74468 19590
rect 74256 19454 74262 19518
rect 74326 19454 74468 19518
rect 74256 19448 74468 19454
rect 74664 19584 75420 19660
rect 75480 19654 75692 19660
rect 75480 19590 75622 19654
rect 75686 19590 75692 19654
rect 74664 19448 74876 19584
rect 75072 19518 75284 19584
rect 75072 19454 75214 19518
rect 75278 19454 75284 19518
rect 75072 19448 75284 19454
rect 75480 19518 75692 19590
rect 75480 19454 75486 19518
rect 75550 19454 75692 19518
rect 75480 19448 75692 19454
rect 21216 19388 21292 19448
rect 27064 19388 27140 19448
rect 69088 19388 69164 19448
rect 20944 19312 21292 19388
rect 20944 19252 21020 19312
rect 20400 19246 20612 19252
rect 20400 19182 20406 19246
rect 20470 19182 20612 19246
rect 3128 18980 3476 19116
rect 3944 18980 4156 19116
rect 20400 19110 20612 19182
rect 20400 19046 20406 19110
rect 20470 19046 20612 19110
rect 20400 19040 20612 19046
rect 20808 19246 21564 19252
rect 20808 19182 20950 19246
rect 21014 19182 21564 19246
rect 20808 19176 21564 19182
rect 20808 19040 21020 19176
rect 21216 19110 21564 19176
rect 21216 19046 21358 19110
rect 21422 19046 21564 19110
rect 21216 19040 21564 19046
rect 21624 19246 21836 19252
rect 21624 19182 21630 19246
rect 21694 19182 21836 19246
rect 21624 19110 21836 19182
rect 21624 19046 21630 19110
rect 21694 19046 21836 19110
rect 21624 19040 21836 19046
rect 22032 19246 22244 19252
rect 22032 19182 22174 19246
rect 22238 19182 22244 19246
rect 22032 19110 22244 19182
rect 26928 19176 27276 19388
rect 27200 19116 27276 19176
rect 22032 19046 22038 19110
rect 22102 19046 22244 19110
rect 22032 19040 22244 19046
rect 1224 18974 4156 18980
rect 1224 18910 1230 18974
rect 1294 18910 4156 18974
rect 1224 18904 4156 18910
rect 26928 18904 27276 19116
rect 1768 18880 1980 18904
rect 1768 18824 1818 18880
rect 1874 18824 1980 18880
rect 27200 18844 27276 18904
rect 1768 18768 1980 18824
rect 20400 18838 20612 18844
rect 20400 18774 20406 18838
rect 20470 18774 20612 18838
rect 20400 18702 20612 18774
rect 20400 18638 20406 18702
rect 20470 18638 20612 18702
rect 20400 18632 20612 18638
rect 20808 18702 21020 18844
rect 20808 18638 20814 18702
rect 20878 18638 21020 18702
rect 20808 18632 21020 18638
rect 21216 18838 21564 18844
rect 21216 18774 21358 18838
rect 21422 18774 21564 18838
rect 21216 18702 21564 18774
rect 21216 18638 21222 18702
rect 21286 18638 21564 18702
rect 21216 18632 21564 18638
rect 21624 18838 21836 18844
rect 21624 18774 21630 18838
rect 21694 18774 21836 18838
rect 21624 18702 21836 18774
rect 21624 18638 21630 18702
rect 21694 18638 21836 18702
rect 21624 18632 21836 18638
rect 22032 18838 22244 18844
rect 22032 18774 22038 18838
rect 22102 18774 22244 18838
rect 22032 18702 22244 18774
rect 22032 18638 22038 18702
rect 22102 18638 22244 18702
rect 22032 18632 22244 18638
rect 26928 18632 27276 18844
rect 68952 19176 69164 19388
rect 73848 19246 74060 19252
rect 73848 19182 73854 19246
rect 73918 19182 74060 19246
rect 68952 19116 69028 19176
rect 68952 18904 69164 19116
rect 73848 19110 74060 19182
rect 73848 19046 73854 19110
rect 73918 19046 74060 19110
rect 73848 19040 74060 19046
rect 74256 19246 74468 19252
rect 74256 19182 74262 19246
rect 74326 19182 74468 19246
rect 74256 19110 74468 19182
rect 74256 19046 74262 19110
rect 74326 19046 74468 19110
rect 74256 19040 74468 19046
rect 74664 19110 74876 19252
rect 74664 19046 74806 19110
rect 74870 19046 74876 19110
rect 74664 19040 74876 19046
rect 75072 19246 75284 19252
rect 75072 19182 75214 19246
rect 75278 19182 75284 19246
rect 75072 19040 75284 19182
rect 75480 19246 75692 19252
rect 75480 19182 75486 19246
rect 75550 19182 75692 19246
rect 75480 19110 75692 19182
rect 75480 19046 75486 19110
rect 75550 19046 75692 19110
rect 75480 19040 75692 19046
rect 75072 18980 75148 19040
rect 74800 18904 75148 18980
rect 68952 18844 69028 18904
rect 74800 18844 74876 18904
rect 94112 18880 94324 18980
rect 68952 18632 69164 18844
rect 73848 18838 74060 18844
rect 73848 18774 73854 18838
rect 73918 18774 74060 18838
rect 73848 18702 74060 18774
rect 73848 18638 73854 18702
rect 73918 18638 74060 18702
rect 73848 18632 74060 18638
rect 74256 18838 74468 18844
rect 74256 18774 74262 18838
rect 74326 18774 74468 18838
rect 74256 18702 74468 18774
rect 74256 18638 74262 18702
rect 74326 18638 74468 18702
rect 74256 18632 74468 18638
rect 74664 18838 75284 18844
rect 74664 18774 74806 18838
rect 74870 18774 75284 18838
rect 74664 18768 75284 18774
rect 74664 18632 74876 18768
rect 75072 18702 75284 18768
rect 75072 18638 75078 18702
rect 75142 18638 75284 18702
rect 75072 18632 75284 18638
rect 75480 18838 75692 18844
rect 75480 18774 75486 18838
rect 75550 18774 75692 18838
rect 75480 18702 75692 18774
rect 94112 18824 94176 18880
rect 94232 18844 94324 18880
rect 94232 18838 94732 18844
rect 94232 18824 94662 18838
rect 94112 18774 94662 18824
rect 94726 18774 94732 18838
rect 94112 18768 94732 18774
rect 77966 18702 78548 18708
rect 75480 18638 75622 18702
rect 75686 18638 75692 18702
rect 77928 18638 77934 18702
rect 77998 18638 78478 18702
rect 78542 18638 78548 18702
rect 75480 18632 75692 18638
rect 77966 18632 78548 18638
rect 27064 18572 27140 18632
rect 69088 18572 69164 18632
rect 18088 18496 18708 18572
rect 18088 18436 18164 18496
rect 18632 18436 18708 18496
rect 17408 18294 17620 18436
rect 17408 18230 17550 18294
rect 17614 18230 17620 18294
rect 17408 18224 17620 18230
rect 17816 18360 18164 18436
rect 18224 18430 18436 18436
rect 18224 18366 18230 18430
rect 18294 18366 18436 18430
rect 17816 18224 18028 18360
rect 18224 18294 18436 18366
rect 18224 18230 18230 18294
rect 18294 18230 18436 18294
rect 18224 18224 18436 18230
rect 18632 18430 18844 18436
rect 18632 18366 18638 18430
rect 18702 18366 18844 18430
rect 18632 18294 18844 18366
rect 18632 18230 18774 18294
rect 18838 18230 18844 18294
rect 18632 18224 18844 18230
rect 20400 18430 20612 18436
rect 20400 18366 20406 18430
rect 20470 18366 20612 18430
rect 20400 18224 20612 18366
rect 20808 18430 21020 18436
rect 20808 18366 20814 18430
rect 20878 18366 21020 18430
rect 20808 18300 21020 18366
rect 21216 18430 21564 18436
rect 21216 18366 21222 18430
rect 21286 18366 21564 18430
rect 21216 18300 21564 18366
rect 20808 18294 21564 18300
rect 20808 18230 20950 18294
rect 21014 18230 21564 18294
rect 20808 18224 21564 18230
rect 21624 18430 21836 18436
rect 21624 18366 21630 18430
rect 21694 18366 21836 18430
rect 21624 18294 21836 18366
rect 21624 18230 21766 18294
rect 21830 18230 21836 18294
rect 21624 18224 21836 18230
rect 22032 18430 22244 18436
rect 22032 18366 22038 18430
rect 22102 18366 22244 18430
rect 22032 18294 22244 18366
rect 26928 18360 27276 18572
rect 68952 18360 69164 18572
rect 77520 18496 78140 18572
rect 77520 18436 77596 18496
rect 78064 18436 78140 18496
rect 27200 18300 27276 18360
rect 69088 18300 69164 18360
rect 22032 18230 22174 18294
rect 22238 18230 22244 18294
rect 22032 18224 22244 18230
rect 20400 18164 20476 18224
rect 20944 18164 21020 18224
rect 20400 17886 20612 18164
rect 20944 18088 21292 18164
rect 26928 18088 27276 18300
rect 68952 18088 69164 18300
rect 73848 18430 74060 18436
rect 73848 18366 73854 18430
rect 73918 18366 74060 18430
rect 73848 18294 74060 18366
rect 73848 18230 73990 18294
rect 74054 18230 74060 18294
rect 73848 18224 74060 18230
rect 74256 18430 74468 18436
rect 74256 18366 74262 18430
rect 74326 18366 74468 18430
rect 74256 18294 74468 18366
rect 74256 18230 74398 18294
rect 74462 18230 74468 18294
rect 74256 18224 74468 18230
rect 74664 18294 74876 18436
rect 74664 18230 74670 18294
rect 74734 18230 74876 18294
rect 74664 18224 74876 18230
rect 75072 18430 75284 18436
rect 75072 18366 75078 18430
rect 75142 18366 75284 18430
rect 75072 18294 75284 18366
rect 75072 18230 75078 18294
rect 75142 18230 75284 18294
rect 75072 18224 75284 18230
rect 75480 18430 75692 18436
rect 75480 18366 75622 18430
rect 75686 18366 75692 18430
rect 75480 18224 75692 18366
rect 77248 18360 77596 18436
rect 77656 18430 78004 18436
rect 77656 18366 77934 18430
rect 77998 18366 78004 18430
rect 77656 18360 78004 18366
rect 78064 18430 78276 18436
rect 78064 18366 78206 18430
rect 78270 18366 78276 18430
rect 77248 18294 77460 18360
rect 77248 18230 77390 18294
rect 77454 18230 77460 18294
rect 77248 18224 77460 18230
rect 77656 18224 77868 18360
rect 78064 18300 78276 18366
rect 78472 18430 78684 18436
rect 78472 18366 78478 18430
rect 78542 18366 78614 18430
rect 78678 18366 78684 18430
rect 78064 18224 78412 18300
rect 78472 18294 78684 18366
rect 78472 18230 78614 18294
rect 78678 18230 78684 18294
rect 78472 18224 78684 18230
rect 75480 18164 75556 18224
rect 78336 18164 78412 18224
rect 21216 18028 21292 18088
rect 27064 18028 27140 18088
rect 68952 18028 69028 18088
rect 20400 17822 20542 17886
rect 20606 17822 20612 17886
rect 20400 17816 20612 17822
rect 20808 18022 21020 18028
rect 20808 17958 20950 18022
rect 21014 17958 21020 18022
rect 20808 17816 21020 17958
rect 21216 17816 21564 18028
rect 21624 18022 21836 18028
rect 21624 17958 21766 18022
rect 21830 17958 21836 18022
rect 21624 17886 21836 17958
rect 21624 17822 21630 17886
rect 21694 17822 21836 17886
rect 21624 17816 21836 17822
rect 22032 18022 22244 18028
rect 22032 17958 22174 18022
rect 22238 17958 22244 18022
rect 22032 17886 22244 17958
rect 22032 17822 22174 17886
rect 22238 17822 22244 17886
rect 22032 17816 22244 17822
rect 26928 17816 27276 18028
rect 21216 17756 21292 17816
rect 27200 17756 27276 17816
rect 3128 17750 3884 17756
rect 3128 17686 3814 17750
rect 3878 17686 3884 17750
rect 3128 17680 3884 17686
rect 3128 17620 3476 17680
rect 3944 17620 4156 17756
rect 16456 17680 17484 17756
rect 16456 17620 16532 17680
rect 17408 17620 17484 17680
rect 17680 17680 18300 17756
rect 17680 17620 17756 17680
rect 18224 17620 18300 17680
rect 20944 17680 21292 17756
rect 20944 17620 21020 17680
rect 3128 17544 3748 17620
rect 3846 17614 4156 17620
rect 3808 17550 3814 17614
rect 3878 17550 4156 17614
rect 3846 17544 4156 17550
rect 16184 17544 16532 17620
rect 3672 17484 3748 17544
rect 3944 17484 4020 17544
rect 3672 17408 4020 17484
rect 16184 17478 16396 17544
rect 16184 17414 16190 17478
rect 16254 17414 16396 17478
rect 16184 17408 16396 17414
rect 16592 17484 16804 17620
rect 17408 17614 17756 17620
rect 17408 17550 17550 17614
rect 17614 17550 17756 17614
rect 17408 17544 17756 17550
rect 16592 17478 17348 17484
rect 16592 17414 16598 17478
rect 16662 17414 17348 17478
rect 16592 17408 17348 17414
rect 17408 17408 17620 17544
rect 17816 17484 18028 17620
rect 18224 17614 18436 17620
rect 18224 17550 18230 17614
rect 18294 17550 18436 17614
rect 17816 17408 18164 17484
rect 18224 17408 18436 17550
rect 18632 17614 18844 17620
rect 18632 17550 18774 17614
rect 18838 17550 18844 17614
rect 18632 17408 18844 17550
rect 20400 17614 20612 17620
rect 20400 17550 20542 17614
rect 20606 17550 20612 17614
rect 20400 17484 20612 17550
rect 20808 17544 21564 17620
rect 20400 17478 20748 17484
rect 20400 17414 20678 17478
rect 20742 17414 20748 17478
rect 20400 17408 20748 17414
rect 20808 17408 21020 17544
rect 21216 17408 21564 17544
rect 21624 17614 21836 17620
rect 21624 17550 21630 17614
rect 21694 17550 21836 17614
rect 21624 17408 21836 17550
rect 22032 17614 22244 17620
rect 22032 17550 22174 17614
rect 22238 17550 22244 17614
rect 22032 17484 22244 17550
rect 26928 17544 27276 17756
rect 68952 17816 69164 18028
rect 73848 18022 74060 18028
rect 73848 17958 73990 18022
rect 74054 17958 74060 18022
rect 73848 17886 74060 17958
rect 73848 17822 73854 17886
rect 73918 17822 74060 17886
rect 73848 17816 74060 17822
rect 74256 18022 74468 18028
rect 74256 17958 74398 18022
rect 74462 17958 74468 18022
rect 74256 17886 74468 17958
rect 74256 17822 74262 17886
rect 74326 17822 74468 17886
rect 74256 17816 74468 17822
rect 74664 18022 74876 18028
rect 74664 17958 74670 18022
rect 74734 17958 74876 18022
rect 74664 17886 74876 17958
rect 75072 18022 75284 18028
rect 75072 17958 75078 18022
rect 75142 17958 75284 18022
rect 75072 17892 75284 17958
rect 74974 17886 75284 17892
rect 74664 17822 74806 17886
rect 74870 17822 74876 17886
rect 74936 17822 74942 17886
rect 75006 17822 75284 17886
rect 74664 17816 74876 17822
rect 74974 17816 75284 17822
rect 75480 17886 75692 18164
rect 78336 18158 79500 18164
rect 78336 18094 79430 18158
rect 79494 18094 79500 18158
rect 78336 18088 79500 18094
rect 75480 17822 75622 17886
rect 75686 17822 75692 17886
rect 75480 17816 75692 17822
rect 68952 17756 69028 17816
rect 68952 17544 69164 17756
rect 77520 17680 78140 17756
rect 77520 17620 77596 17680
rect 78064 17620 78140 17680
rect 79288 17680 79908 17756
rect 79288 17620 79364 17680
rect 79832 17620 79908 17680
rect 26928 17484 27004 17544
rect 69088 17484 69164 17544
rect 22032 17478 22924 17484
rect 22032 17414 22038 17478
rect 22102 17414 22854 17478
rect 22918 17414 22924 17478
rect 22032 17408 22924 17414
rect 17272 17348 17348 17408
rect 17816 17348 17892 17408
rect 1224 17342 1980 17348
rect 1224 17278 1230 17342
rect 1294 17278 1980 17342
rect 1224 17272 1980 17278
rect 17272 17272 17892 17348
rect 18088 17348 18164 17408
rect 18632 17348 18708 17408
rect 18088 17272 18708 17348
rect 26928 17272 27276 17484
rect 68952 17272 69164 17484
rect 73848 17614 74060 17620
rect 73848 17550 73854 17614
rect 73918 17550 74060 17614
rect 73848 17408 74060 17550
rect 74256 17614 74468 17620
rect 74256 17550 74262 17614
rect 74326 17550 74468 17614
rect 74256 17408 74468 17550
rect 74664 17614 75012 17620
rect 74664 17550 74806 17614
rect 74870 17550 74942 17614
rect 75006 17550 75012 17614
rect 74664 17544 75012 17550
rect 74664 17484 74876 17544
rect 75072 17484 75284 17620
rect 74664 17408 75284 17484
rect 75480 17614 75692 17620
rect 75480 17550 75622 17614
rect 75686 17550 75692 17614
rect 75480 17408 75692 17550
rect 77248 17614 77596 17620
rect 77248 17550 77390 17614
rect 77454 17550 77596 17614
rect 77248 17544 77596 17550
rect 77248 17408 77460 17544
rect 77656 17484 77868 17620
rect 77656 17408 78004 17484
rect 78064 17408 78276 17620
rect 78472 17614 79364 17620
rect 78472 17550 78614 17614
rect 78678 17550 79364 17614
rect 78472 17544 79364 17550
rect 79424 17614 79636 17620
rect 79424 17550 79430 17614
rect 79494 17550 79636 17614
rect 78472 17408 78684 17544
rect 79424 17484 79636 17550
rect 79832 17484 80044 17620
rect 79424 17478 79772 17484
rect 79424 17414 79702 17478
rect 79766 17414 79772 17478
rect 79424 17408 79772 17414
rect 79832 17478 82492 17484
rect 79832 17414 82422 17478
rect 82486 17414 82492 17478
rect 79832 17408 82492 17414
rect 77928 17348 78004 17408
rect 78472 17348 78548 17408
rect 77928 17272 78548 17348
rect 1768 17200 1980 17272
rect 27200 17212 27276 17272
rect 69088 17212 69164 17272
rect 1768 17144 1818 17200
rect 1874 17144 1980 17200
rect 1768 17000 1980 17144
rect 26928 17076 27276 17212
rect 68952 17076 69164 17212
rect 82416 17206 82628 17212
rect 82416 17142 82422 17206
rect 82486 17142 82628 17206
rect 22032 17070 22244 17076
rect 22032 17006 22038 17070
rect 22102 17006 22244 17070
rect 22032 16934 22244 17006
rect 22032 16870 22038 16934
rect 22102 16870 22244 16934
rect 22032 16864 22244 16870
rect 22848 17070 23196 17076
rect 22848 17006 22854 17070
rect 22918 17006 23196 17070
rect 22848 16940 23196 17006
rect 25568 16940 25780 17076
rect 26656 17070 28636 17076
rect 26656 17006 28566 17070
rect 28630 17006 28636 17070
rect 26656 17000 28636 17006
rect 68952 17000 69572 17076
rect 82416 17070 82628 17142
rect 82416 17006 82422 17070
rect 82486 17006 82628 17070
rect 82416 17000 82628 17006
rect 94112 17200 94324 17348
rect 94112 17144 94176 17200
rect 94232 17144 94324 17200
rect 94112 17076 94324 17144
rect 94112 17070 94732 17076
rect 94112 17006 94662 17070
rect 94726 17006 94732 17070
rect 94112 17000 94732 17006
rect 22848 16934 26596 16940
rect 22848 16870 26526 16934
rect 26590 16870 26596 16934
rect 22848 16864 26596 16870
rect 26656 16864 26868 17000
rect 69360 16864 69572 17000
rect 81872 16875 81956 16879
rect 81839 16870 81956 16875
rect 81839 16814 81844 16870
rect 81900 16814 81956 16870
rect 81839 16809 81956 16814
rect 81872 16805 81956 16809
rect 26558 16662 27956 16668
rect 26520 16598 26526 16662
rect 26590 16598 27956 16662
rect 26558 16592 27956 16598
rect 27744 16532 27956 16592
rect 28288 16532 28500 16668
rect 28968 16592 30404 16668
rect 30502 16662 31628 16668
rect 30464 16598 30470 16662
rect 30534 16598 31628 16662
rect 30502 16592 31628 16598
rect 28968 16532 29180 16592
rect 29512 16532 29724 16592
rect 27744 16526 29180 16532
rect 29278 16526 29724 16532
rect 27744 16462 28294 16526
rect 28358 16462 29180 16526
rect 29240 16462 29246 16526
rect 29310 16462 29724 16526
rect 27744 16456 29180 16462
rect 29278 16456 29724 16462
rect 30192 16532 30404 16592
rect 30736 16532 31084 16592
rect 30192 16456 31084 16532
rect 31416 16526 31628 16592
rect 31416 16462 31558 16526
rect 31622 16462 31628 16526
rect 31416 16456 31628 16462
rect 32096 16532 32308 16668
rect 32640 16532 32852 16668
rect 32096 16526 32852 16532
rect 32096 16462 32102 16526
rect 32166 16462 32782 16526
rect 32846 16462 32852 16526
rect 32096 16456 32852 16462
rect 33320 16592 34212 16668
rect 33320 16526 33532 16592
rect 33320 16462 33326 16526
rect 33390 16462 33532 16526
rect 33320 16456 33532 16462
rect 33864 16526 34212 16592
rect 33864 16462 34142 16526
rect 34206 16462 34212 16526
rect 33864 16456 34212 16462
rect 34544 16532 34756 16668
rect 35224 16592 36660 16668
rect 35224 16532 35436 16592
rect 34544 16526 35436 16532
rect 34544 16462 34550 16526
rect 34614 16462 35436 16526
rect 34544 16456 35436 16462
rect 35768 16526 35980 16592
rect 35768 16462 35774 16526
rect 35838 16462 35980 16526
rect 35768 16456 35980 16462
rect 36448 16532 36660 16592
rect 36992 16532 37340 16668
rect 37672 16592 38564 16668
rect 37672 16532 37884 16592
rect 36448 16526 37884 16532
rect 36448 16462 36590 16526
rect 36654 16462 37884 16526
rect 36448 16456 37884 16462
rect 38352 16532 38564 16592
rect 38896 16532 39108 16668
rect 38352 16526 39108 16532
rect 38352 16462 38358 16526
rect 38422 16462 39038 16526
rect 39102 16462 39108 16526
rect 38352 16456 39108 16462
rect 39576 16592 40332 16668
rect 39576 16526 39788 16592
rect 39576 16462 39582 16526
rect 39646 16462 39788 16526
rect 39576 16456 39788 16462
rect 40120 16526 40332 16592
rect 40120 16462 40262 16526
rect 40326 16462 40332 16526
rect 40120 16456 40332 16462
rect 40800 16532 41012 16668
rect 41344 16532 41692 16668
rect 42024 16592 42916 16668
rect 42024 16532 42236 16592
rect 40800 16526 42236 16532
rect 40800 16462 40806 16526
rect 40870 16462 42030 16526
rect 42094 16462 42236 16526
rect 40800 16456 42236 16462
rect 42704 16532 42916 16592
rect 43248 16532 43460 16668
rect 43928 16592 44820 16668
rect 43928 16532 44140 16592
rect 42704 16526 44140 16532
rect 42704 16462 42846 16526
rect 42910 16462 44140 16526
rect 42704 16456 44140 16462
rect 44472 16532 44820 16592
rect 45152 16532 45364 16668
rect 44472 16526 45364 16532
rect 44472 16462 44614 16526
rect 44678 16462 45294 16526
rect 45358 16462 45364 16526
rect 44472 16456 45364 16462
rect 45832 16592 46588 16668
rect 45832 16526 46044 16592
rect 45832 16462 45838 16526
rect 45902 16462 46044 16526
rect 45832 16456 46044 16462
rect 46376 16526 46588 16592
rect 46376 16462 46518 16526
rect 46582 16462 46588 16526
rect 46376 16456 46588 16462
rect 47056 16532 47268 16668
rect 47600 16532 47948 16668
rect 47056 16526 47948 16532
rect 47056 16462 47062 16526
rect 47126 16462 47742 16526
rect 47806 16462 47948 16526
rect 47056 16456 47948 16462
rect 48280 16592 49716 16668
rect 48280 16526 48492 16592
rect 48280 16462 48286 16526
rect 48350 16462 48492 16526
rect 48280 16456 48492 16462
rect 48960 16532 49172 16592
rect 49504 16532 49716 16592
rect 50184 16532 50396 16668
rect 48960 16526 49444 16532
rect 48960 16462 49374 16526
rect 49438 16462 49444 16526
rect 48960 16456 49444 16462
rect 49504 16526 50396 16532
rect 49504 16462 50326 16526
rect 50390 16462 50396 16526
rect 49504 16456 50396 16462
rect 50728 16592 51620 16668
rect 50728 16526 50940 16592
rect 50728 16462 50734 16526
rect 50798 16462 50940 16526
rect 50728 16456 50940 16462
rect 51408 16526 51620 16592
rect 51408 16462 51550 16526
rect 51614 16462 51620 16526
rect 51408 16456 51620 16462
rect 51952 16532 52300 16668
rect 52632 16592 53524 16668
rect 52632 16532 52844 16592
rect 51952 16526 52844 16532
rect 51952 16462 51958 16526
rect 52022 16462 52844 16526
rect 51952 16456 52844 16462
rect 53312 16532 53524 16592
rect 53856 16532 54068 16668
rect 53312 16526 54068 16532
rect 53312 16462 53318 16526
rect 53382 16462 53998 16526
rect 54062 16462 54068 16526
rect 53312 16456 54068 16462
rect 54536 16592 55428 16668
rect 54536 16526 54748 16592
rect 54536 16462 54542 16526
rect 54606 16462 54748 16526
rect 54536 16456 54748 16462
rect 55080 16526 55428 16592
rect 55080 16462 55358 16526
rect 55422 16462 55428 16526
rect 55080 16456 55428 16462
rect 55760 16532 55972 16668
rect 56440 16532 56652 16668
rect 55760 16526 56652 16532
rect 55760 16462 55766 16526
rect 55830 16462 56446 16526
rect 56510 16462 56652 16526
rect 55760 16456 56652 16462
rect 56984 16592 57876 16668
rect 56984 16526 57196 16592
rect 56984 16462 56990 16526
rect 57054 16462 57196 16526
rect 56984 16456 57196 16462
rect 57664 16526 57876 16592
rect 58208 16592 59100 16668
rect 58208 16532 58556 16592
rect 57974 16526 58556 16532
rect 57664 16462 57806 16526
rect 57870 16462 57876 16526
rect 57936 16462 57942 16526
rect 58006 16462 58556 16526
rect 57664 16456 57876 16462
rect 57974 16456 58556 16462
rect 58888 16526 59100 16592
rect 58888 16462 59030 16526
rect 59094 16462 59100 16526
rect 58888 16456 59100 16462
rect 59568 16532 59780 16668
rect 60112 16532 60324 16668
rect 59568 16526 60324 16532
rect 59568 16462 59574 16526
rect 59638 16462 60254 16526
rect 60318 16462 60324 16526
rect 59568 16456 60324 16462
rect 60792 16592 62228 16668
rect 60792 16526 61004 16592
rect 60792 16462 60798 16526
rect 60862 16462 61004 16526
rect 60792 16456 61004 16462
rect 61336 16456 61548 16592
rect 62016 16532 62228 16592
rect 62560 16592 64132 16668
rect 64230 16662 64676 16668
rect 64192 16598 64198 16662
rect 64262 16598 64676 16662
rect 64230 16592 64676 16598
rect 62560 16532 62908 16592
rect 62016 16526 62908 16532
rect 62016 16462 62022 16526
rect 62086 16462 62908 16526
rect 62016 16456 62908 16462
rect 63240 16526 63452 16592
rect 63240 16462 63246 16526
rect 63310 16462 63452 16526
rect 63240 16456 63452 16462
rect 63920 16532 64132 16592
rect 64464 16532 64676 16592
rect 65144 16532 65356 16668
rect 63920 16526 65356 16532
rect 63920 16462 65286 16526
rect 65350 16462 65356 16526
rect 63920 16456 65356 16462
rect 65688 16532 66036 16668
rect 66368 16532 66580 16668
rect 65688 16526 66580 16532
rect 65688 16462 65694 16526
rect 65758 16462 66510 16526
rect 66574 16462 66580 16526
rect 65688 16456 66580 16462
rect 67048 16592 67804 16668
rect 67048 16526 67260 16592
rect 67048 16462 67054 16526
rect 67118 16462 67260 16526
rect 67048 16456 67260 16462
rect 67592 16526 67804 16592
rect 67592 16462 67734 16526
rect 67798 16462 67804 16526
rect 67592 16456 67804 16462
rect 68272 16526 68484 16668
rect 82824 16614 95956 16668
rect 82824 16558 82926 16614
rect 82982 16592 95956 16614
rect 82982 16558 83036 16592
rect 68272 16462 68278 16526
rect 68342 16462 68484 16526
rect 81638 16545 81704 16548
rect 81976 16545 82042 16548
rect 81638 16543 82042 16545
rect 81638 16487 81643 16543
rect 81699 16487 81981 16543
rect 82037 16487 82042 16543
rect 81638 16485 82042 16487
rect 81638 16482 81704 16485
rect 81976 16482 82042 16485
rect 68272 16456 68484 16462
rect 82824 16456 83036 16558
rect 3128 16260 3476 16396
rect 3944 16260 4156 16396
rect 2350 16254 4156 16260
rect 2312 16190 2318 16254
rect 2382 16190 4156 16254
rect 2350 16184 4156 16190
rect 14144 16390 16260 16396
rect 14144 16326 16190 16390
rect 16254 16326 16260 16390
rect 14144 16320 16260 16326
rect 14144 16254 14356 16320
rect 14144 16190 14286 16254
rect 14350 16190 14356 16254
rect 14144 16184 14356 16190
rect 27744 15988 28092 16124
rect 28152 16118 28364 16124
rect 28152 16054 28294 16118
rect 28358 16054 28364 16118
rect 28152 15988 28364 16054
rect 27744 15912 28364 15988
rect 29104 16118 29316 16124
rect 29104 16054 29246 16118
rect 29310 16054 29316 16118
rect 29104 15988 29316 16054
rect 29376 15988 29724 16124
rect 29104 15912 29724 15988
rect 30328 16118 30948 16124
rect 30328 16054 30470 16118
rect 30534 16054 30948 16118
rect 30328 16048 30948 16054
rect 30328 15912 30540 16048
rect 30736 15912 30948 16048
rect 31552 16118 31764 16124
rect 31552 16054 31558 16118
rect 31622 16054 31764 16118
rect 31552 15988 31764 16054
rect 31960 16118 32172 16124
rect 31960 16054 32102 16118
rect 32166 16054 32172 16118
rect 31960 15988 32172 16054
rect 31552 15912 32172 15988
rect 32776 16118 33396 16124
rect 32776 16054 32782 16118
rect 32846 16054 33326 16118
rect 33390 16054 33396 16118
rect 32776 16048 33396 16054
rect 32776 15912 32988 16048
rect 33184 15912 33396 16048
rect 34000 16118 34212 16124
rect 34000 16054 34142 16118
rect 34206 16054 34212 16118
rect 34000 15988 34212 16054
rect 34408 16118 34620 16124
rect 34408 16054 34550 16118
rect 34614 16054 34620 16118
rect 34408 15988 34620 16054
rect 34000 15912 34620 15988
rect 35224 16118 35844 16124
rect 35224 16054 35774 16118
rect 35838 16054 35844 16118
rect 35224 16048 35844 16054
rect 35224 15912 35572 16048
rect 35632 15912 35844 16048
rect 36584 16118 37204 16124
rect 36584 16054 36590 16118
rect 36654 16054 37204 16118
rect 36584 16048 37204 16054
rect 36584 15912 36796 16048
rect 36856 15912 37204 16048
rect 37808 15988 38020 16124
rect 38216 16118 38428 16124
rect 38216 16054 38358 16118
rect 38422 16054 38428 16118
rect 38216 15988 38428 16054
rect 37808 15912 38428 15988
rect 39032 16118 39652 16124
rect 39032 16054 39038 16118
rect 39102 16054 39582 16118
rect 39646 16054 39652 16118
rect 39032 16048 39652 16054
rect 39032 15912 39244 16048
rect 39440 15912 39652 16048
rect 40256 16118 40468 16124
rect 40256 16054 40262 16118
rect 40326 16054 40468 16118
rect 40256 15988 40468 16054
rect 40664 16118 40876 16124
rect 40664 16054 40806 16118
rect 40870 16054 40876 16118
rect 40664 15988 40876 16054
rect 40256 15912 40876 15988
rect 41480 16118 42100 16124
rect 41480 16054 42030 16118
rect 42094 16054 42100 16118
rect 41480 16048 42100 16054
rect 41480 15912 41828 16048
rect 41888 15912 42100 16048
rect 42840 16118 43460 16124
rect 42840 16054 42846 16118
rect 42910 16054 43460 16118
rect 42840 16048 43460 16054
rect 42840 15912 43052 16048
rect 43112 15912 43460 16048
rect 44064 15988 44276 16124
rect 44472 16118 44684 16124
rect 44472 16054 44614 16118
rect 44678 16054 44684 16118
rect 44472 15988 44684 16054
rect 44064 15912 44684 15988
rect 45288 16118 45908 16124
rect 45288 16054 45294 16118
rect 45358 16054 45838 16118
rect 45902 16054 45908 16118
rect 45288 16048 45908 16054
rect 45288 15912 45500 16048
rect 45696 15912 45908 16048
rect 46512 16118 46724 16124
rect 46512 16054 46518 16118
rect 46582 16054 46724 16118
rect 46512 15988 46724 16054
rect 46920 16118 47132 16124
rect 46920 16054 47062 16118
rect 47126 16054 47132 16118
rect 46920 15988 47132 16054
rect 46512 15912 47132 15988
rect 47736 16118 48356 16124
rect 47736 16054 47742 16118
rect 47806 16054 48286 16118
rect 48350 16054 48356 16118
rect 47736 16048 48356 16054
rect 47736 15912 47948 16048
rect 48144 15912 48356 16048
rect 48960 15988 49308 16124
rect 49368 16118 49580 16124
rect 49368 16054 49374 16118
rect 49438 16054 49580 16118
rect 49368 15988 49580 16054
rect 48960 15912 49580 15988
rect 50320 16118 50532 16124
rect 50320 16054 50326 16118
rect 50390 16054 50532 16118
rect 50320 15988 50532 16054
rect 50592 16118 50940 16124
rect 50592 16054 50734 16118
rect 50798 16054 50940 16118
rect 50592 15988 50940 16054
rect 50320 15912 50940 15988
rect 51544 16118 52164 16124
rect 51544 16054 51550 16118
rect 51614 16054 51958 16118
rect 52022 16054 52164 16118
rect 51544 16048 52164 16054
rect 51544 15912 51756 16048
rect 51952 15912 52164 16048
rect 52768 15988 52980 16124
rect 53176 16118 53388 16124
rect 53176 16054 53318 16118
rect 53382 16054 53388 16118
rect 53176 15988 53388 16054
rect 52768 15912 53388 15988
rect 53992 16118 54612 16124
rect 53992 16054 53998 16118
rect 54062 16054 54542 16118
rect 54606 16054 54612 16118
rect 53992 16048 54612 16054
rect 53992 15912 54204 16048
rect 54400 15912 54612 16048
rect 55216 16118 55428 16124
rect 55216 16054 55358 16118
rect 55422 16054 55428 16118
rect 55216 15988 55428 16054
rect 55624 16118 55836 16124
rect 55624 16054 55766 16118
rect 55830 16054 55836 16118
rect 55624 15988 55836 16054
rect 55216 15912 55836 15988
rect 56440 16118 56788 16124
rect 56440 16054 56446 16118
rect 56510 16054 56788 16118
rect 56440 15988 56788 16054
rect 56848 16118 57060 16124
rect 56848 16054 56990 16118
rect 57054 16054 57060 16118
rect 56848 15988 57060 16054
rect 56440 15912 57060 15988
rect 57800 16118 58420 16124
rect 57800 16054 57806 16118
rect 57870 16054 57942 16118
rect 58006 16054 58420 16118
rect 57800 16048 58420 16054
rect 57800 15912 58012 16048
rect 58072 15982 58420 16048
rect 58072 15918 58078 15982
rect 58142 15918 58420 15982
rect 58072 15912 58420 15918
rect 59024 16118 59236 16124
rect 59024 16054 59030 16118
rect 59094 16054 59236 16118
rect 59024 15988 59236 16054
rect 59432 16118 59644 16124
rect 59432 16054 59574 16118
rect 59638 16054 59644 16118
rect 59432 15988 59644 16054
rect 59024 15912 59644 15988
rect 60248 16118 60868 16124
rect 60248 16054 60254 16118
rect 60318 16054 60798 16118
rect 60862 16054 60868 16118
rect 60248 16048 60868 16054
rect 60248 15912 60460 16048
rect 60656 15912 60868 16048
rect 61472 15988 61684 16124
rect 61880 16118 62092 16124
rect 61880 16054 62022 16118
rect 62086 16054 62092 16118
rect 61880 15988 62092 16054
rect 61472 15912 62092 15988
rect 62696 16118 63316 16124
rect 62696 16054 63246 16118
rect 63310 16054 63316 16118
rect 62696 16048 63316 16054
rect 62696 15912 63044 16048
rect 63104 15912 63316 16048
rect 64056 16118 64676 16124
rect 64056 16054 64198 16118
rect 64262 16054 64676 16118
rect 64056 16048 64676 16054
rect 64056 15912 64268 16048
rect 64328 15912 64676 16048
rect 65280 16118 65492 16124
rect 65280 16054 65286 16118
rect 65350 16054 65492 16118
rect 65280 15988 65492 16054
rect 65688 16118 65900 16124
rect 65688 16054 65694 16118
rect 65758 16054 65900 16118
rect 65688 15988 65900 16054
rect 65280 15912 65900 15988
rect 66504 16118 67124 16124
rect 66504 16054 66510 16118
rect 66574 16054 67054 16118
rect 67118 16054 67124 16118
rect 66504 16048 67124 16054
rect 66504 15912 66716 16048
rect 66912 15912 67124 16048
rect 67728 16118 68348 16124
rect 67728 16054 67734 16118
rect 67798 16054 68278 16118
rect 68342 16054 68348 16118
rect 67728 16048 68348 16054
rect 67728 15912 67940 16048
rect 79734 15846 82628 15852
rect 79696 15782 79702 15846
rect 79766 15782 82628 15846
rect 79734 15776 82628 15782
rect 82416 15710 82628 15776
rect 82416 15646 82558 15710
rect 82622 15646 82628 15710
rect 82416 15640 82628 15646
rect 1768 15574 2388 15580
rect 1768 15520 2318 15574
rect 1768 15464 1818 15520
rect 1874 15510 2318 15520
rect 2382 15510 2388 15574
rect 1874 15504 2388 15510
rect 14253 15559 14319 15562
rect 22395 15559 22461 15562
rect 14253 15557 22461 15559
rect 1874 15464 1980 15504
rect 14253 15501 14258 15557
rect 14314 15501 22400 15557
rect 22456 15501 22461 15557
rect 14253 15499 22461 15501
rect 14253 15496 14319 15499
rect 22395 15496 22461 15499
rect 94112 15520 94324 15580
rect 1768 15444 1980 15464
rect 1224 15438 1980 15444
rect 1224 15374 1230 15438
rect 1294 15374 1980 15438
rect 1224 15368 1980 15374
rect 94112 15464 94176 15520
rect 94232 15464 94324 15520
rect 94112 15444 94324 15464
rect 94112 15438 94732 15444
rect 94112 15374 94662 15438
rect 94726 15374 94732 15438
rect 94112 15368 94732 15374
rect 2555 15198 2561 15262
rect 2625 15260 2631 15262
rect 2625 15200 28031 15260
rect 2625 15198 2631 15200
rect 81558 14987 81624 14990
rect 81976 14987 82042 14990
rect 81558 14985 82042 14987
rect 81558 14929 81563 14985
rect 81619 14929 81981 14985
rect 82037 14929 82042 14985
rect 81558 14927 82042 14929
rect 81558 14924 81624 14927
rect 81976 14924 82042 14927
rect 82824 14960 95956 15036
rect 82824 14914 83036 14960
rect 3128 14824 4156 14900
rect 3128 14764 3476 14824
rect 3128 14758 3884 14764
rect 3128 14694 3814 14758
rect 3878 14694 3884 14758
rect 3128 14688 3884 14694
rect 3944 14758 4156 14824
rect 3944 14694 3950 14758
rect 4014 14694 4156 14758
rect 3944 14688 4156 14694
rect 14144 14894 16668 14900
rect 14144 14830 16598 14894
rect 16662 14830 16668 14894
rect 14144 14824 16668 14830
rect 82824 14858 82926 14914
rect 82982 14858 83036 14914
rect 82824 14824 83036 14858
rect 14144 14758 14356 14824
rect 20710 14758 21292 14764
rect 14144 14694 14150 14758
rect 14214 14694 14356 14758
rect 20672 14694 20678 14758
rect 20742 14694 21292 14758
rect 14144 14688 14356 14694
rect 20710 14688 21292 14694
rect 21080 14622 21292 14688
rect 21080 14558 21086 14622
rect 21150 14558 21292 14622
rect 21080 14552 21292 14558
rect 28560 14622 28908 14628
rect 28560 14558 28566 14622
rect 28630 14558 28908 14622
rect 28560 14492 28908 14558
rect 29920 14552 32580 14628
rect 29920 14492 30132 14552
rect 28560 14416 30132 14492
rect 28560 14280 28908 14416
rect 29920 14280 30132 14416
rect 31144 14350 31356 14552
rect 31144 14286 31150 14350
rect 31214 14286 31356 14350
rect 31144 14280 31356 14286
rect 32368 14356 32580 14552
rect 33592 14356 33804 14628
rect 34816 14552 37612 14628
rect 34816 14356 35028 14552
rect 32368 14280 35028 14356
rect 36040 14280 36388 14552
rect 37400 14492 37612 14552
rect 38624 14552 41284 14628
rect 38624 14492 38836 14552
rect 37400 14416 38836 14492
rect 37400 14280 37612 14416
rect 38624 14280 38836 14416
rect 39848 14280 40060 14552
rect 41072 14356 41284 14552
rect 42296 14356 42644 14628
rect 43656 14552 46316 14628
rect 43656 14356 43868 14552
rect 41072 14280 43868 14356
rect 44880 14280 45092 14552
rect 46104 14492 46316 14552
rect 47328 14552 51348 14628
rect 47328 14492 47540 14552
rect 46104 14416 47540 14492
rect 46104 14280 46316 14416
rect 47328 14280 47540 14416
rect 48552 14280 48764 14552
rect 49776 14280 50124 14552
rect 51136 14356 51348 14552
rect 52360 14552 55020 14628
rect 52360 14356 52572 14552
rect 51136 14280 52572 14356
rect 53584 14280 53796 14552
rect 54808 14492 55020 14552
rect 56032 14552 57604 14628
rect 56032 14492 56244 14552
rect 54808 14416 56244 14492
rect 54808 14280 55020 14416
rect 56032 14280 56244 14416
rect 57256 14492 57604 14552
rect 58616 14552 60052 14628
rect 58616 14492 58828 14552
rect 57256 14416 58828 14492
rect 57256 14280 57604 14416
rect 58616 14280 58828 14416
rect 59840 14356 60052 14552
rect 61064 14552 65084 14628
rect 61064 14356 61276 14552
rect 59840 14280 61276 14356
rect 62288 14280 62500 14552
rect 63512 14280 63860 14552
rect 64872 14492 65084 14552
rect 66096 14492 66308 14628
rect 67320 14492 67532 14628
rect 64872 14416 67532 14492
rect 64872 14280 65084 14416
rect 66096 14280 66308 14416
rect 67320 14280 67532 14416
rect 82416 14486 82628 14492
rect 82416 14422 82422 14486
rect 82486 14422 82628 14486
rect 82416 14220 82628 14422
rect 82280 14214 82628 14220
rect 82280 14150 82286 14214
rect 82350 14150 82628 14214
rect 82280 14144 82628 14150
rect 1768 13840 1980 13948
rect 94112 13942 94732 13948
rect 94112 13878 94662 13942
rect 94726 13878 94732 13942
rect 94112 13872 94732 13878
rect 1768 13812 1818 13840
rect 1224 13806 1818 13812
rect 1224 13742 1230 13806
rect 1294 13784 1818 13806
rect 1874 13812 1980 13840
rect 94155 13840 94253 13872
rect 1874 13806 3204 13812
rect 1874 13784 3134 13806
rect 1294 13742 3134 13784
rect 3198 13742 3204 13806
rect 1224 13736 3204 13742
rect 82824 13786 83036 13812
rect 82824 13730 82926 13786
rect 82982 13730 83036 13786
rect 94155 13784 94176 13840
rect 94232 13784 94253 13840
rect 94155 13763 94253 13784
rect 81478 13717 81544 13720
rect 81976 13717 82042 13720
rect 81478 13715 82042 13717
rect 81478 13659 81483 13715
rect 81539 13659 81981 13715
rect 82037 13659 82042 13715
rect 81478 13657 82042 13659
rect 81478 13654 81544 13657
rect 81976 13654 82042 13657
rect 82824 13676 83036 13730
rect 82824 13600 95956 13676
rect 3128 13534 3476 13540
rect 3128 13470 3134 13534
rect 3198 13470 3476 13534
rect 3128 13404 3476 13470
rect 3944 13404 4156 13540
rect 14144 13534 14356 13540
rect 14144 13470 14286 13534
rect 14350 13470 14356 13534
rect 14144 13404 14356 13470
rect 3128 13328 4156 13404
rect 14046 13398 14356 13404
rect 14008 13334 14014 13398
rect 14078 13334 14356 13398
rect 14046 13328 14356 13334
rect 21080 13262 22108 13268
rect 21080 13198 22038 13262
rect 22102 13198 22108 13262
rect 21080 13192 22108 13198
rect 21080 13056 21292 13192
rect 82416 12990 82628 12996
rect 82416 12926 82558 12990
rect 82622 12926 82628 12990
rect 82416 12854 82628 12926
rect 82416 12790 82422 12854
rect 82486 12790 82628 12854
rect 82416 12784 82628 12790
rect 14253 12731 14319 12734
rect 26098 12731 26164 12734
rect 14253 12729 26164 12731
rect 14253 12673 14258 12729
rect 14314 12673 26103 12729
rect 26159 12673 26164 12729
rect 28513 12724 28611 12749
rect 29761 12724 29859 12749
rect 31009 12724 31107 12749
rect 32257 12724 32355 12749
rect 33505 12724 33603 12749
rect 34753 12724 34851 12749
rect 36001 12724 36099 12749
rect 37249 12724 37347 12749
rect 38497 12724 38595 12749
rect 39745 12724 39843 12749
rect 40993 12724 41091 12749
rect 42241 12724 42339 12749
rect 43489 12724 43587 12749
rect 44737 12724 44835 12749
rect 45985 12724 46083 12749
rect 47233 12724 47331 12749
rect 48481 12724 48579 12749
rect 49729 12724 49827 12749
rect 50977 12724 51075 12749
rect 52225 12724 52323 12749
rect 53473 12724 53571 12749
rect 54721 12724 54819 12749
rect 55969 12724 56067 12749
rect 57217 12724 57315 12749
rect 58465 12724 58563 12749
rect 59713 12724 59811 12749
rect 60961 12724 61059 12749
rect 62209 12724 62307 12749
rect 63457 12724 63555 12749
rect 64705 12724 64803 12749
rect 65953 12724 66051 12749
rect 67201 12724 67299 12749
rect 14253 12671 26164 12673
rect 14253 12668 14319 12671
rect 26098 12668 26164 12671
rect 28424 12718 67396 12724
rect 28424 12654 31150 12718
rect 31214 12654 64606 12718
rect 64670 12654 67396 12718
rect 28424 12648 67396 12654
rect 1768 12160 1980 12316
rect 94112 12310 94732 12316
rect 94112 12246 94662 12310
rect 94726 12246 94732 12310
rect 94112 12240 94732 12246
rect 1768 12104 1818 12160
rect 1874 12104 1980 12160
rect 1768 12044 1980 12104
rect 81398 12159 81464 12162
rect 81976 12159 82042 12162
rect 81398 12157 82042 12159
rect 81398 12101 81403 12157
rect 81459 12101 81981 12157
rect 82037 12101 82042 12157
rect 81398 12099 82042 12101
rect 81398 12096 81464 12099
rect 81976 12096 82042 12099
rect 82824 12086 83036 12180
rect 1224 12038 1980 12044
rect 1224 11974 1230 12038
rect 1294 11974 1980 12038
rect 1224 11968 1980 11974
rect 3128 12038 3884 12044
rect 3128 11974 3814 12038
rect 3878 11974 3884 12038
rect 3128 11968 3884 11974
rect 3128 11908 3476 11968
rect 3944 11908 4156 12044
rect 544 11902 4156 11908
rect 544 11838 550 11902
rect 614 11838 4156 11902
rect 544 11832 4156 11838
rect 14144 12038 14356 12044
rect 14144 11974 14150 12038
rect 14214 11974 14356 12038
rect 14144 11902 14356 11974
rect 14144 11838 14286 11902
rect 14350 11838 14356 11902
rect 14144 11832 14356 11838
rect 21080 11902 21292 11908
rect 21080 11838 21086 11902
rect 21150 11838 21292 11902
rect 21080 11696 21292 11838
rect 28424 11902 28636 12044
rect 28424 11838 28430 11902
rect 28494 11838 28636 11902
rect 28424 11832 28636 11838
rect 29648 11908 29860 12044
rect 30872 11908 31084 12044
rect 29648 11902 31084 11908
rect 29648 11838 29790 11902
rect 29854 11838 31014 11902
rect 31078 11838 31084 11902
rect 29648 11832 31084 11838
rect 32096 11902 32308 12044
rect 32096 11838 32102 11902
rect 32166 11838 32308 11902
rect 32096 11832 32308 11838
rect 33320 11968 34892 12044
rect 33320 11902 33532 11968
rect 33320 11838 33462 11902
rect 33526 11838 33532 11902
rect 33320 11832 33532 11838
rect 34544 11902 34892 11968
rect 34544 11838 34686 11902
rect 34750 11838 34892 11902
rect 34544 11832 34892 11838
rect 35904 11908 36116 12044
rect 37128 11908 37340 12044
rect 35904 11902 37340 11908
rect 35904 11838 36046 11902
rect 36110 11838 37134 11902
rect 37198 11838 37340 11902
rect 35904 11832 37340 11838
rect 38352 11908 38564 12044
rect 39576 11908 39788 12044
rect 38352 11902 39788 11908
rect 38352 11838 38494 11902
rect 38558 11838 39718 11902
rect 39782 11838 39788 11902
rect 38352 11832 39788 11838
rect 40800 11902 41012 12044
rect 40800 11838 40806 11902
rect 40870 11838 41012 11902
rect 40800 11832 41012 11838
rect 42024 11968 44820 12044
rect 42024 11902 42372 11968
rect 42024 11838 42166 11902
rect 42230 11838 42372 11902
rect 42024 11832 42372 11838
rect 43384 11902 43596 11968
rect 43384 11838 43390 11902
rect 43454 11838 43596 11902
rect 43384 11832 43596 11838
rect 44608 11908 44820 11968
rect 45832 11968 47268 12044
rect 45832 11908 46044 11968
rect 44608 11902 46044 11908
rect 44608 11838 44750 11902
rect 44814 11838 45838 11902
rect 45902 11838 46044 11902
rect 44608 11832 46044 11838
rect 47056 11908 47268 11968
rect 48280 11968 51076 12044
rect 48280 11908 48628 11968
rect 47056 11902 48628 11908
rect 47056 11838 47198 11902
rect 47262 11838 48422 11902
rect 48486 11838 48628 11902
rect 47056 11832 48628 11838
rect 49640 11902 49852 11968
rect 49640 11838 49782 11902
rect 49846 11838 49852 11902
rect 49640 11832 49852 11838
rect 50864 11908 51076 11968
rect 52088 11908 52300 12044
rect 50864 11902 52300 11908
rect 50864 11838 51006 11902
rect 51070 11838 52094 11902
rect 52158 11838 52300 11902
rect 50864 11832 52300 11838
rect 53312 11902 53524 12044
rect 53312 11838 53454 11902
rect 53518 11838 53524 11902
rect 53312 11832 53524 11838
rect 54536 11968 56108 12044
rect 54536 11902 54748 11968
rect 54536 11838 54542 11902
rect 54606 11838 54748 11902
rect 54536 11832 54748 11838
rect 55760 11902 56108 11968
rect 55760 11838 56038 11902
rect 56102 11838 56108 11902
rect 55760 11832 56108 11838
rect 57120 12038 58148 12044
rect 57120 11974 58078 12038
rect 58142 11974 58148 12038
rect 57120 11968 58148 11974
rect 57120 11908 57332 11968
rect 58344 11908 58556 12044
rect 57120 11902 58556 11908
rect 57120 11838 57126 11902
rect 57190 11838 58486 11902
rect 58550 11838 58556 11902
rect 57120 11832 58556 11838
rect 59568 11908 59780 12044
rect 60792 11908 61004 12044
rect 59568 11902 61004 11908
rect 59568 11838 59710 11902
rect 59774 11838 60798 11902
rect 60862 11838 61004 11902
rect 59568 11832 61004 11838
rect 62016 11908 62228 12044
rect 63240 11908 63588 12044
rect 62016 11902 63588 11908
rect 62016 11838 62158 11902
rect 62222 11838 63382 11902
rect 63446 11838 63588 11902
rect 62016 11832 63588 11838
rect 64600 11902 64812 12044
rect 64600 11838 64742 11902
rect 64806 11838 64812 11902
rect 64600 11832 64812 11838
rect 65824 11902 66036 12044
rect 65824 11838 65830 11902
rect 65894 11838 66036 11902
rect 65824 11832 66036 11838
rect 67048 11902 67260 12044
rect 82824 12030 82926 12086
rect 82982 12044 83036 12086
rect 94112 12160 94324 12240
rect 94112 12104 94176 12160
rect 94232 12104 94324 12160
rect 82982 12038 83172 12044
rect 82982 12030 83102 12038
rect 82824 11974 83102 12030
rect 83166 11974 83172 12038
rect 82824 11968 83172 11974
rect 94112 11968 94324 12104
rect 67048 11838 67190 11902
rect 67254 11838 67260 11902
rect 67048 11832 67260 11838
rect 82318 11630 82628 11636
rect 82280 11566 82286 11630
rect 82350 11566 82628 11630
rect 82318 11560 82628 11566
rect 82416 11494 82628 11560
rect 82416 11430 82558 11494
rect 82622 11430 82628 11494
rect 82416 11424 82628 11430
rect 14253 11317 14319 11320
rect 26346 11317 26412 11320
rect 14253 11315 26412 11317
rect 14253 11259 14258 11315
rect 14314 11259 26351 11315
rect 26407 11259 26412 11315
rect 14253 11257 26412 11259
rect 14253 11254 14319 11257
rect 26346 11254 26412 11257
rect 28424 11222 29860 11228
rect 28424 11158 28430 11222
rect 28494 11158 29790 11222
rect 29854 11158 29860 11222
rect 28424 11152 29860 11158
rect 28443 11039 28636 11152
rect 29691 11039 29860 11152
rect 28560 11016 28636 11039
rect 29784 11016 29860 11039
rect 30872 11222 33668 11228
rect 30872 11158 31014 11222
rect 31078 11158 32102 11222
rect 32166 11158 33462 11222
rect 33526 11158 33668 11222
rect 30872 11152 33668 11158
rect 34680 11222 36116 11228
rect 34680 11158 34686 11222
rect 34750 11158 36046 11222
rect 36110 11158 36116 11222
rect 34680 11152 36116 11158
rect 30872 11016 31084 11152
rect 32187 11039 32308 11152
rect 33435 11039 33668 11152
rect 34683 11039 34892 11152
rect 35931 11039 36116 11152
rect 32232 11016 32308 11039
rect 33592 11016 33668 11039
rect 34816 11016 34892 11039
rect 36040 11016 36116 11039
rect 37128 11222 38564 11228
rect 37128 11158 37134 11222
rect 37198 11158 38494 11222
rect 38558 11158 38564 11222
rect 37128 11152 38564 11158
rect 39576 11222 42372 11228
rect 39576 11158 39718 11222
rect 39782 11158 40806 11222
rect 40870 11158 42166 11222
rect 42230 11158 42372 11222
rect 39576 11152 42372 11158
rect 43384 11222 43596 11228
rect 43384 11158 43390 11222
rect 43454 11158 43596 11222
rect 43384 11152 43596 11158
rect 44608 11222 44820 11228
rect 44608 11158 44750 11222
rect 44814 11158 44820 11222
rect 44608 11152 44820 11158
rect 45832 11222 46044 11228
rect 45832 11158 45838 11222
rect 45902 11158 46044 11222
rect 45832 11152 46044 11158
rect 47056 11222 47268 11228
rect 47056 11158 47198 11222
rect 47262 11158 47268 11222
rect 47056 11152 47268 11158
rect 48280 11222 48628 11228
rect 48280 11158 48422 11222
rect 48486 11158 48628 11222
rect 48280 11152 48628 11158
rect 37128 11016 37340 11152
rect 38427 11086 38564 11152
rect 38427 11039 38494 11086
rect 38488 11022 38494 11039
rect 38558 11022 38564 11086
rect 39675 11039 39773 11152
rect 40923 11039 41148 11152
rect 42171 11039 42372 11152
rect 43419 11039 43596 11152
rect 44667 11039 44820 11152
rect 45915 11039 46044 11152
rect 47163 11039 47268 11152
rect 48411 11039 48628 11152
rect 38488 11016 38564 11022
rect 40936 11016 41148 11039
rect 42296 11016 42372 11039
rect 43520 11016 43596 11039
rect 44744 11016 44820 11039
rect 45968 11016 46044 11039
rect 47192 11016 47268 11039
rect 48552 11016 48628 11039
rect 49640 11222 49852 11228
rect 49640 11158 49782 11222
rect 49846 11158 49852 11222
rect 49640 11016 49852 11158
rect 50864 11222 51076 11228
rect 50864 11158 51006 11222
rect 51070 11158 51076 11222
rect 50864 11152 51076 11158
rect 52088 11222 54884 11228
rect 52088 11158 52094 11222
rect 52158 11158 53454 11222
rect 53518 11158 54542 11222
rect 54606 11158 54884 11222
rect 52088 11152 54884 11158
rect 50907 11039 51076 11152
rect 52155 11039 52300 11152
rect 53403 11039 53524 11152
rect 54651 11039 54884 11152
rect 51000 11016 51076 11039
rect 52224 11016 52300 11039
rect 53448 11016 53524 11039
rect 54808 11016 54884 11039
rect 55896 11222 57332 11228
rect 55896 11158 56038 11222
rect 56102 11158 57126 11222
rect 57190 11158 57332 11222
rect 55896 11152 57332 11158
rect 58344 11222 59780 11228
rect 58344 11158 58486 11222
rect 58550 11158 59710 11222
rect 59774 11158 59780 11222
rect 58344 11152 59780 11158
rect 60792 11222 62364 11228
rect 60792 11158 60798 11222
rect 60862 11158 62158 11222
rect 62222 11158 62364 11222
rect 60792 11152 62364 11158
rect 63376 11222 67260 11228
rect 63376 11158 63382 11222
rect 63446 11158 64742 11222
rect 64806 11158 65830 11222
rect 65894 11158 67190 11222
rect 67254 11158 67260 11222
rect 63376 11152 67260 11158
rect 55896 11016 56108 11152
rect 57147 11039 57332 11152
rect 58395 11039 58556 11152
rect 59643 11039 59780 11152
rect 60891 11039 60989 11152
rect 62139 11039 62364 11152
rect 63387 11039 63588 11152
rect 64635 11039 64812 11152
rect 65883 11039 66036 11152
rect 57256 11016 57332 11039
rect 58480 11016 58556 11039
rect 59704 11016 59780 11039
rect 62288 11016 62364 11039
rect 63512 11016 63588 11039
rect 64736 11016 64812 11039
rect 65960 11016 66036 11039
rect 67048 11016 67260 11152
rect 82824 10958 83036 11092
rect 82824 10956 82926 10958
rect 28152 10813 28364 10956
rect 28560 10815 28636 10820
rect 28152 10757 28210 10813
rect 28266 10757 28364 10813
rect 28152 10684 28364 10757
rect 28443 10717 28636 10815
rect 3128 10608 4156 10684
rect 14008 10678 14356 10684
rect 14008 10614 14014 10678
rect 14078 10614 14356 10678
rect 14008 10608 14356 10614
rect 27880 10678 28364 10684
rect 27880 10614 27886 10678
rect 27950 10614 28364 10678
rect 27880 10608 28364 10614
rect 28560 10678 28636 10717
rect 29376 10813 29588 10956
rect 29784 10815 29860 10820
rect 29376 10757 29458 10813
rect 29514 10757 29588 10813
rect 29376 10684 29588 10757
rect 29691 10717 29860 10815
rect 28560 10614 28566 10678
rect 28630 10614 28636 10678
rect 28560 10608 28636 10614
rect 29240 10678 29588 10684
rect 29240 10614 29246 10678
rect 29310 10614 29588 10678
rect 29240 10608 29588 10614
rect 29784 10678 29860 10717
rect 30600 10813 30812 10956
rect 30600 10757 30706 10813
rect 30762 10757 30812 10813
rect 30600 10684 30812 10757
rect 29784 10614 29790 10678
rect 29854 10614 29860 10678
rect 29784 10608 29860 10614
rect 30328 10678 30812 10684
rect 30328 10614 30334 10678
rect 30398 10614 30812 10678
rect 30328 10608 30812 10614
rect 30872 10678 31084 10820
rect 30872 10614 30878 10678
rect 30942 10614 31084 10678
rect 30872 10608 31084 10614
rect 31824 10813 32036 10956
rect 33048 10880 33396 10956
rect 32232 10815 32308 10820
rect 31824 10757 31954 10813
rect 32010 10757 32036 10813
rect 31824 10678 32036 10757
rect 32187 10717 32308 10815
rect 31824 10614 31966 10678
rect 32030 10614 32036 10678
rect 31824 10608 32036 10614
rect 32232 10678 32308 10717
rect 32232 10614 32238 10678
rect 32302 10614 32308 10678
rect 32232 10608 32308 10614
rect 33048 10813 33279 10880
rect 33592 10815 33668 10820
rect 33048 10757 33202 10813
rect 33258 10757 33279 10813
rect 33048 10736 33279 10757
rect 33048 10678 33260 10736
rect 33435 10717 33668 10815
rect 33048 10614 33190 10678
rect 33254 10614 33260 10678
rect 33048 10608 33260 10614
rect 33456 10678 33668 10717
rect 33456 10614 33462 10678
rect 33526 10614 33668 10678
rect 33456 10608 33668 10614
rect 34408 10813 34620 10956
rect 34816 10815 34892 10820
rect 34408 10757 34450 10813
rect 34506 10757 34620 10813
rect 34408 10678 34620 10757
rect 34683 10717 34892 10815
rect 34408 10614 34414 10678
rect 34478 10614 34620 10678
rect 34408 10608 34620 10614
rect 34816 10678 34892 10717
rect 34816 10614 34822 10678
rect 34886 10614 34892 10678
rect 34816 10608 34892 10614
rect 35632 10813 35844 10956
rect 36040 10815 36116 10820
rect 35632 10757 35698 10813
rect 35754 10757 35844 10813
rect 35632 10678 35844 10757
rect 35931 10717 36116 10815
rect 35632 10614 35638 10678
rect 35702 10614 35844 10678
rect 35632 10608 35844 10614
rect 36040 10678 36116 10717
rect 36040 10614 36046 10678
rect 36110 10614 36116 10678
rect 36040 10608 36116 10614
rect 36856 10813 37068 10956
rect 36856 10757 36946 10813
rect 37002 10757 37068 10813
rect 36856 10678 37068 10757
rect 36856 10614 36862 10678
rect 36926 10614 37068 10678
rect 36856 10608 37068 10614
rect 37128 10678 37340 10820
rect 38080 10813 38292 10956
rect 39304 10880 39652 10956
rect 40664 10880 40876 10956
rect 38488 10815 38564 10820
rect 38080 10757 38194 10813
rect 38250 10757 38292 10813
rect 38080 10684 38292 10757
rect 38427 10717 38564 10815
rect 37128 10614 37134 10678
rect 37198 10614 37340 10678
rect 37128 10608 37340 10614
rect 37808 10678 38292 10684
rect 37808 10614 37814 10678
rect 37878 10614 38292 10678
rect 37808 10608 38292 10614
rect 38488 10684 38564 10717
rect 39304 10813 39519 10880
rect 39304 10757 39442 10813
rect 39498 10757 39519 10813
rect 39304 10736 39519 10757
rect 38488 10678 38662 10684
rect 39304 10678 39516 10736
rect 38488 10614 38630 10678
rect 38694 10614 38700 10678
rect 39304 10614 39310 10678
rect 39374 10614 39516 10678
rect 39675 10684 39773 10815
rect 40664 10813 40767 10880
rect 40936 10815 41148 10820
rect 40664 10757 40690 10813
rect 40746 10757 40767 10813
rect 40664 10736 40767 10757
rect 39675 10678 39788 10684
rect 39675 10646 39718 10678
rect 38488 10608 38662 10614
rect 39304 10608 39516 10614
rect 39712 10614 39718 10646
rect 39782 10614 39788 10678
rect 39712 10608 39788 10614
rect 40664 10678 40740 10736
rect 40923 10717 41148 10815
rect 40664 10614 40670 10678
rect 40734 10614 40740 10678
rect 40664 10608 40740 10614
rect 40936 10684 41148 10717
rect 41888 10813 42100 10956
rect 42296 10815 42372 10820
rect 41888 10757 41938 10813
rect 41994 10757 42100 10813
rect 40936 10678 41828 10684
rect 40936 10614 40942 10678
rect 41006 10614 41758 10678
rect 41822 10614 41828 10678
rect 40936 10608 41828 10614
rect 41888 10678 42100 10757
rect 42171 10717 42372 10815
rect 41888 10614 41894 10678
rect 41958 10614 42100 10678
rect 41888 10608 42100 10614
rect 42296 10678 42372 10717
rect 42296 10614 42302 10678
rect 42366 10614 42372 10678
rect 42296 10608 42372 10614
rect 43112 10813 43324 10956
rect 43520 10815 43596 10820
rect 43112 10757 43186 10813
rect 43242 10757 43324 10813
rect 43112 10678 43324 10757
rect 43419 10717 43596 10815
rect 43112 10614 43118 10678
rect 43182 10614 43324 10678
rect 43112 10608 43324 10614
rect 43520 10678 43596 10717
rect 43520 10614 43526 10678
rect 43590 10614 43596 10678
rect 43520 10608 43596 10614
rect 44336 10813 44548 10956
rect 44744 10815 44820 10820
rect 44336 10757 44434 10813
rect 44490 10757 44548 10813
rect 44336 10678 44548 10757
rect 44667 10717 44820 10815
rect 44336 10614 44342 10678
rect 44406 10614 44548 10678
rect 44336 10608 44548 10614
rect 44744 10684 44820 10717
rect 45560 10813 45772 10956
rect 46784 10880 47132 10956
rect 48144 10880 48356 10956
rect 45968 10815 46044 10820
rect 45560 10757 45682 10813
rect 45738 10757 45772 10813
rect 44744 10678 45364 10684
rect 44744 10614 44750 10678
rect 44814 10614 45294 10678
rect 45358 10614 45364 10678
rect 44744 10608 45364 10614
rect 45560 10678 45772 10757
rect 45915 10717 46044 10815
rect 45560 10614 45566 10678
rect 45630 10614 45772 10678
rect 45560 10608 45772 10614
rect 45968 10678 46044 10717
rect 46784 10813 47007 10880
rect 47192 10815 47268 10820
rect 46784 10757 46930 10813
rect 46986 10757 47007 10813
rect 46784 10736 47007 10757
rect 46784 10684 46996 10736
rect 47163 10717 47268 10815
rect 45968 10614 45974 10678
rect 46038 10614 46044 10678
rect 45968 10608 46044 10614
rect 46648 10678 46996 10684
rect 46648 10614 46654 10678
rect 46718 10614 46996 10678
rect 46648 10608 46996 10614
rect 47192 10684 47268 10717
rect 48144 10813 48255 10880
rect 48552 10815 48628 10820
rect 48144 10757 48178 10813
rect 48234 10757 48255 10813
rect 48144 10736 48255 10757
rect 48144 10684 48220 10736
rect 48411 10717 48628 10815
rect 47192 10678 47812 10684
rect 47192 10614 47198 10678
rect 47262 10614 47742 10678
rect 47806 10614 47812 10678
rect 47192 10608 47812 10614
rect 47872 10678 48220 10684
rect 47872 10614 47878 10678
rect 47942 10614 48220 10678
rect 47872 10608 48220 10614
rect 48416 10684 48628 10717
rect 49368 10813 49580 10956
rect 49368 10757 49426 10813
rect 49482 10757 49580 10813
rect 49368 10684 49580 10757
rect 48416 10678 49036 10684
rect 48416 10614 48422 10678
rect 48486 10614 48966 10678
rect 49030 10614 49036 10678
rect 48416 10608 49036 10614
rect 49096 10678 49580 10684
rect 49096 10614 49102 10678
rect 49166 10614 49580 10678
rect 49096 10608 49580 10614
rect 49640 10678 49852 10820
rect 49640 10614 49646 10678
rect 49710 10614 49782 10678
rect 49846 10614 49852 10678
rect 49640 10608 49852 10614
rect 50592 10813 50804 10956
rect 51000 10815 51076 10820
rect 50592 10757 50674 10813
rect 50730 10757 50804 10813
rect 50592 10678 50804 10757
rect 50907 10717 51076 10815
rect 50592 10614 50598 10678
rect 50662 10614 50804 10678
rect 50592 10608 50804 10614
rect 51000 10678 51076 10717
rect 51816 10813 52028 10956
rect 52224 10815 52300 10820
rect 51816 10757 51922 10813
rect 51978 10757 52028 10813
rect 51816 10684 52028 10757
rect 52155 10717 52300 10815
rect 51000 10614 51006 10678
rect 51070 10614 51076 10678
rect 51000 10608 51076 10614
rect 51408 10678 52028 10684
rect 51408 10614 51414 10678
rect 51478 10614 52028 10678
rect 51408 10608 52028 10614
rect 52224 10678 52300 10717
rect 52224 10614 52230 10678
rect 52294 10614 52300 10678
rect 52224 10608 52300 10614
rect 53040 10813 53252 10956
rect 54264 10880 54612 10956
rect 53448 10815 53524 10820
rect 53040 10757 53170 10813
rect 53226 10757 53252 10813
rect 53040 10678 53252 10757
rect 53403 10717 53524 10815
rect 53040 10614 53182 10678
rect 53246 10614 53252 10678
rect 53040 10608 53252 10614
rect 53448 10678 53524 10717
rect 53448 10614 53454 10678
rect 53518 10614 53524 10678
rect 53448 10608 53524 10614
rect 54264 10813 54495 10880
rect 54808 10815 54884 10820
rect 54264 10757 54418 10813
rect 54474 10757 54495 10813
rect 54264 10736 54495 10757
rect 54264 10678 54476 10736
rect 54651 10717 54884 10815
rect 54264 10614 54406 10678
rect 54470 10614 54476 10678
rect 54264 10608 54476 10614
rect 54672 10678 54884 10717
rect 54672 10614 54678 10678
rect 54742 10614 54884 10678
rect 54672 10608 54884 10614
rect 55624 10813 55836 10956
rect 55624 10757 55666 10813
rect 55722 10757 55836 10813
rect 55624 10678 55836 10757
rect 55624 10614 55630 10678
rect 55694 10614 55836 10678
rect 55624 10608 55836 10614
rect 55896 10678 56108 10820
rect 55896 10614 55902 10678
rect 55966 10614 56108 10678
rect 55896 10608 56108 10614
rect 56848 10813 57060 10956
rect 57256 10815 57332 10820
rect 56848 10757 56914 10813
rect 56970 10757 57060 10813
rect 56848 10678 57060 10757
rect 57147 10717 57332 10815
rect 56848 10614 56854 10678
rect 56918 10614 57060 10678
rect 56848 10608 57060 10614
rect 57256 10678 57332 10717
rect 58072 10813 58284 10956
rect 58480 10815 58556 10820
rect 58072 10757 58162 10813
rect 58218 10757 58284 10813
rect 58072 10684 58284 10757
rect 58395 10717 58556 10815
rect 57256 10614 57262 10678
rect 57326 10614 57332 10678
rect 57256 10608 57332 10614
rect 57800 10678 58284 10684
rect 57800 10614 57806 10678
rect 57870 10614 58284 10678
rect 57800 10608 58284 10614
rect 58480 10684 58556 10717
rect 59296 10813 59508 10956
rect 60520 10880 60868 10956
rect 61880 10880 62092 10956
rect 59704 10815 59780 10820
rect 59296 10757 59410 10813
rect 59466 10757 59508 10813
rect 58480 10678 59236 10684
rect 58480 10614 58486 10678
rect 58550 10614 59166 10678
rect 59230 10614 59236 10678
rect 58480 10608 59236 10614
rect 59296 10678 59508 10757
rect 59643 10717 59780 10815
rect 59296 10614 59302 10678
rect 59366 10614 59508 10678
rect 59296 10608 59508 10614
rect 59704 10678 59780 10717
rect 59704 10614 59710 10678
rect 59774 10614 59780 10678
rect 59704 10608 59780 10614
rect 60520 10813 60735 10880
rect 60520 10757 60658 10813
rect 60714 10757 60735 10813
rect 60520 10736 60735 10757
rect 60520 10678 60732 10736
rect 60520 10614 60526 10678
rect 60590 10614 60732 10678
rect 60891 10684 60989 10815
rect 61880 10813 61983 10880
rect 62288 10815 62364 10820
rect 61880 10757 61906 10813
rect 61962 10757 61983 10813
rect 61880 10736 61983 10757
rect 60891 10678 61820 10684
rect 60891 10646 60934 10678
rect 60520 10608 60732 10614
rect 60928 10614 60934 10646
rect 60998 10614 61750 10678
rect 61814 10614 61820 10678
rect 60928 10608 61820 10614
rect 61880 10678 61956 10736
rect 62139 10684 62364 10815
rect 63104 10813 63316 10956
rect 63512 10815 63588 10820
rect 63104 10757 63154 10813
rect 63210 10757 63316 10813
rect 61880 10614 61886 10678
rect 61950 10614 61956 10678
rect 61880 10608 61956 10614
rect 62152 10678 63044 10684
rect 62152 10614 62158 10678
rect 62222 10614 62974 10678
rect 63038 10614 63044 10678
rect 62152 10608 63044 10614
rect 63104 10678 63316 10757
rect 63387 10717 63588 10815
rect 63104 10614 63110 10678
rect 63174 10614 63316 10678
rect 63104 10608 63316 10614
rect 63512 10678 63588 10717
rect 63512 10614 63518 10678
rect 63582 10614 63588 10678
rect 63512 10608 63588 10614
rect 64328 10813 64540 10956
rect 64736 10815 64812 10820
rect 64328 10757 64402 10813
rect 64458 10757 64540 10813
rect 64328 10678 64540 10757
rect 64635 10814 64812 10815
rect 64635 10750 64742 10814
rect 64806 10750 64812 10814
rect 64635 10717 64812 10750
rect 64328 10614 64334 10678
rect 64398 10614 64540 10678
rect 64328 10608 64540 10614
rect 64736 10684 64812 10717
rect 65552 10813 65764 10956
rect 65960 10815 66036 10820
rect 65552 10757 65650 10813
rect 65706 10757 65764 10813
rect 64736 10678 65492 10684
rect 64736 10614 64742 10678
rect 64806 10614 65422 10678
rect 65486 10614 65492 10678
rect 64736 10608 65492 10614
rect 65552 10678 65764 10757
rect 65883 10717 66036 10815
rect 65552 10614 65558 10678
rect 65622 10614 65764 10678
rect 65552 10608 65764 10614
rect 65960 10678 66036 10717
rect 65960 10614 65966 10678
rect 66030 10614 66036 10678
rect 65960 10608 66036 10614
rect 66776 10813 66988 10956
rect 82688 10950 82926 10956
rect 81318 10889 81384 10892
rect 81976 10889 82042 10892
rect 81318 10887 82042 10889
rect 81318 10831 81323 10887
rect 81379 10831 81981 10887
rect 82037 10831 82042 10887
rect 82688 10886 82694 10950
rect 82758 10902 82926 10950
rect 82982 10902 83036 10958
rect 82758 10886 83036 10902
rect 82688 10880 83036 10886
rect 81318 10829 82042 10831
rect 81318 10826 81384 10829
rect 81976 10826 82042 10829
rect 66776 10757 66898 10813
rect 66954 10757 66988 10813
rect 66776 10678 66988 10757
rect 66776 10614 66782 10678
rect 66846 10614 66988 10678
rect 66776 10608 66988 10614
rect 67048 10678 67260 10820
rect 67048 10614 67054 10678
rect 67118 10614 67260 10678
rect 67048 10608 67260 10614
rect 3128 10548 3476 10608
rect 1224 10542 3476 10548
rect 1224 10478 1230 10542
rect 1294 10480 3476 10542
rect 1294 10478 1818 10480
rect 1224 10472 1818 10478
rect 1768 10424 1818 10472
rect 1874 10472 3476 10480
rect 3944 10472 4156 10608
rect 14144 10548 14356 10608
rect 14008 10542 14356 10548
rect 14008 10478 14014 10542
rect 14078 10478 14356 10542
rect 14008 10472 14356 10478
rect 94112 10542 94732 10548
rect 94112 10480 94662 10542
rect 1874 10424 1980 10472
rect 1768 10336 1980 10424
rect 94112 10424 94176 10480
rect 94232 10478 94662 10480
rect 94726 10478 94732 10542
rect 94232 10472 94732 10478
rect 94232 10424 94324 10472
rect 48998 10406 49716 10412
rect 48960 10342 48966 10406
rect 49030 10342 49646 10406
rect 49710 10342 49716 10406
rect 48998 10336 49716 10342
rect 94112 10336 94324 10424
rect 28288 10134 28636 10140
rect 28288 10070 28566 10134
rect 28630 10070 28636 10134
rect 28288 10064 28636 10070
rect 29512 10134 29860 10140
rect 29512 10070 29790 10134
rect 29854 10070 29860 10134
rect 29512 10064 29860 10070
rect 30736 10134 30948 10140
rect 30736 10070 30878 10134
rect 30942 10070 30948 10134
rect 14253 9903 14319 9906
rect 26222 9903 26288 9906
rect 14253 9901 26288 9903
rect 14253 9845 14258 9901
rect 14314 9845 26227 9901
rect 26283 9845 26288 9901
rect 14253 9843 26288 9845
rect 14253 9840 14319 9843
rect 26222 9840 26288 9843
rect 28288 9862 28500 10064
rect 28288 9798 28430 9862
rect 28494 9798 28500 9862
rect 28288 9792 28500 9798
rect 29512 9868 29724 10064
rect 29512 9862 29860 9868
rect 29512 9798 29790 9862
rect 29854 9798 29860 9862
rect 29512 9792 29860 9798
rect 30736 9862 30948 10070
rect 30736 9798 30878 9862
rect 30942 9798 30948 9862
rect 30736 9792 30948 9798
rect 31960 10134 32308 10140
rect 31960 10070 32238 10134
rect 32302 10070 32308 10134
rect 31960 10064 32308 10070
rect 33320 10134 33532 10140
rect 33320 10070 33462 10134
rect 33526 10070 33532 10134
rect 31960 9868 32172 10064
rect 33320 10004 33532 10070
rect 34544 10134 34892 10140
rect 34544 10070 34822 10134
rect 34886 10070 34892 10134
rect 34544 10064 34892 10070
rect 35768 10134 36116 10140
rect 35768 10070 36046 10134
rect 36110 10070 36116 10134
rect 35768 10064 36116 10070
rect 36992 10134 37204 10140
rect 36992 10070 37134 10134
rect 37198 10070 37204 10134
rect 34544 10004 34756 10064
rect 33320 9928 34756 10004
rect 33320 9868 33532 9928
rect 34544 9868 34756 9928
rect 35768 9868 35980 10064
rect 36992 9868 37204 10070
rect 38216 10134 38700 10140
rect 38216 10070 38630 10134
rect 38694 10070 38700 10134
rect 38216 10064 38700 10070
rect 39440 10134 39788 10140
rect 39440 10070 39718 10134
rect 39782 10070 39788 10134
rect 31960 9862 32444 9868
rect 31960 9798 32374 9862
rect 32438 9798 32444 9862
rect 31960 9792 32444 9798
rect 33320 9862 33668 9868
rect 33320 9798 33598 9862
rect 33662 9798 33668 9862
rect 33320 9792 33668 9798
rect 34544 9862 34892 9868
rect 34544 9798 34822 9862
rect 34886 9798 34892 9862
rect 34544 9792 34892 9798
rect 35768 9862 36116 9868
rect 35768 9798 36046 9862
rect 36110 9798 36116 9862
rect 35768 9792 36116 9798
rect 36992 9862 37340 9868
rect 36992 9798 37270 9862
rect 37334 9798 37340 9862
rect 36992 9792 37340 9798
rect 38216 9862 38428 10064
rect 38216 9798 38222 9862
rect 38286 9798 38428 9862
rect 38216 9792 38428 9798
rect 39440 9862 39788 10070
rect 39440 9798 39718 9862
rect 39782 9798 39788 9862
rect 39440 9792 39788 9798
rect 40800 10134 41012 10140
rect 41790 10134 42372 10140
rect 40800 10070 40942 10134
rect 41006 10070 41012 10134
rect 41752 10070 41758 10134
rect 41822 10070 42302 10134
rect 42366 10070 42372 10134
rect 40800 9868 41012 10070
rect 41790 10064 42372 10070
rect 43248 10134 43596 10140
rect 43248 10070 43526 10134
rect 43590 10070 43596 10134
rect 43248 10064 43596 10070
rect 44472 10134 44820 10140
rect 45326 10134 46044 10140
rect 44472 10070 44750 10134
rect 44814 10070 44820 10134
rect 45288 10070 45294 10134
rect 45358 10070 45974 10134
rect 46038 10070 46044 10134
rect 44472 10064 44820 10070
rect 45326 10064 46044 10070
rect 46920 10134 47268 10140
rect 47774 10134 48492 10140
rect 46920 10070 47198 10134
rect 47262 10070 47268 10134
rect 47736 10070 47742 10134
rect 47806 10070 48422 10134
rect 48486 10070 48492 10134
rect 42024 9868 42236 10064
rect 43248 9868 43460 10064
rect 44472 9868 44684 10064
rect 45696 9868 45908 10064
rect 40800 9862 41148 9868
rect 40800 9798 41078 9862
rect 41142 9798 41148 9862
rect 40800 9792 41148 9798
rect 42024 9862 42372 9868
rect 42024 9798 42302 9862
rect 42366 9798 42372 9862
rect 42024 9792 42372 9798
rect 43248 9862 43558 9868
rect 44472 9862 44820 9868
rect 43248 9798 43526 9862
rect 43590 9798 43596 9862
rect 44472 9798 44750 9862
rect 44814 9798 44820 9862
rect 43248 9792 43558 9798
rect 44472 9792 44820 9798
rect 45696 9862 46044 9868
rect 45696 9798 45974 9862
rect 46038 9798 46044 9862
rect 45696 9792 46044 9798
rect 46920 9862 47268 10070
rect 47774 10064 48492 10070
rect 46920 9798 47198 9862
rect 47262 9798 47268 9862
rect 46920 9792 47268 9798
rect 48280 9862 48492 10064
rect 48280 9798 48422 9862
rect 48486 9798 48492 9862
rect 48280 9792 48492 9798
rect 49504 10134 49852 10140
rect 49504 10070 49782 10134
rect 49846 10070 49852 10134
rect 49504 10064 49852 10070
rect 50728 10134 51076 10140
rect 50728 10070 51006 10134
rect 51070 10070 51076 10134
rect 50728 10064 51076 10070
rect 51952 10134 52300 10140
rect 51952 10070 52230 10134
rect 52294 10070 52300 10134
rect 51952 10064 52300 10070
rect 53176 10134 53524 10140
rect 53176 10070 53454 10134
rect 53518 10070 53524 10134
rect 53176 10064 53524 10070
rect 54536 10134 54748 10140
rect 54536 10070 54678 10134
rect 54742 10070 54748 10134
rect 49504 9868 49716 10064
rect 49504 9862 49852 9868
rect 49504 9798 49782 9862
rect 49846 9798 49852 9862
rect 49504 9792 49852 9798
rect 50728 9862 50940 10064
rect 50728 9798 50870 9862
rect 50934 9798 50940 9862
rect 50728 9792 50940 9798
rect 51952 9862 52164 10064
rect 51952 9798 52094 9862
rect 52158 9798 52164 9862
rect 51952 9792 52164 9798
rect 53176 9868 53388 10064
rect 53176 9862 53660 9868
rect 53176 9798 53590 9862
rect 53654 9798 53660 9862
rect 53176 9792 53660 9798
rect 54536 9862 54748 10070
rect 54536 9798 54678 9862
rect 54742 9798 54748 9862
rect 54536 9792 54748 9798
rect 55760 10134 55972 10140
rect 55760 10070 55902 10134
rect 55966 10070 55972 10134
rect 55760 9868 55972 10070
rect 56984 10134 57332 10140
rect 56984 10070 57262 10134
rect 57326 10070 57332 10134
rect 56984 10064 57332 10070
rect 58208 10134 58556 10140
rect 59198 10134 59780 10140
rect 58208 10070 58486 10134
rect 58550 10070 58556 10134
rect 59160 10070 59166 10134
rect 59230 10070 59710 10134
rect 59774 10070 59780 10134
rect 58208 10064 58556 10070
rect 59198 10064 59780 10070
rect 60656 10134 61004 10140
rect 61782 10134 62228 10140
rect 63006 10134 63588 10140
rect 60656 10070 60934 10134
rect 60998 10070 61004 10134
rect 61744 10070 61750 10134
rect 61814 10070 62158 10134
rect 62222 10070 62228 10134
rect 62968 10070 62974 10134
rect 63038 10070 63518 10134
rect 63582 10070 63588 10134
rect 56984 9868 57196 10064
rect 55760 9862 56108 9868
rect 56750 9862 57196 9868
rect 55760 9798 56038 9862
rect 56102 9798 56108 9862
rect 56712 9798 56718 9862
rect 56782 9798 57126 9862
rect 57190 9798 57196 9862
rect 55760 9792 56108 9798
rect 56750 9792 57196 9798
rect 58208 9868 58420 10064
rect 59432 9868 59644 10064
rect 58208 9862 58556 9868
rect 58208 9798 58486 9862
rect 58550 9798 58556 9862
rect 58208 9792 58556 9798
rect 59432 9862 59780 9868
rect 59432 9798 59710 9862
rect 59774 9798 59780 9862
rect 59432 9792 59780 9798
rect 60656 9862 61004 10070
rect 61782 10064 62228 10070
rect 63006 10064 63588 10070
rect 64464 10134 64812 10140
rect 65454 10134 66036 10140
rect 64464 10070 64742 10134
rect 64806 10070 64812 10134
rect 65416 10070 65422 10134
rect 65486 10070 65966 10134
rect 66030 10070 66036 10134
rect 64464 10064 64812 10070
rect 65454 10064 66036 10070
rect 66912 10134 67124 10140
rect 66912 10070 67054 10134
rect 67118 10070 67124 10134
rect 60656 9798 60934 9862
rect 60998 9798 61004 9862
rect 60656 9792 61004 9798
rect 62016 9868 62228 10064
rect 63240 9868 63452 10064
rect 64464 9868 64676 10064
rect 62016 9862 62364 9868
rect 62016 9798 62294 9862
rect 62358 9798 62364 9862
rect 62016 9792 62364 9798
rect 63240 9862 63588 9868
rect 63240 9798 63518 9862
rect 63582 9798 63588 9862
rect 63240 9792 63588 9798
rect 64464 9862 64774 9868
rect 65688 9862 65900 10064
rect 64464 9798 64742 9862
rect 64806 9798 64812 9862
rect 65688 9798 65830 9862
rect 65894 9798 65900 9862
rect 64464 9792 64774 9798
rect 65688 9792 65900 9798
rect 66912 9868 67124 10070
rect 82416 10134 82628 10140
rect 82416 10070 82422 10134
rect 82486 10070 82628 10134
rect 82416 9998 82628 10070
rect 82416 9934 82422 9998
rect 82486 9934 82628 9998
rect 82416 9928 82628 9934
rect 66912 9862 67260 9868
rect 66912 9798 67190 9862
rect 67254 9798 67260 9862
rect 66912 9792 67260 9798
rect 28288 9454 28500 9596
rect 28288 9390 28294 9454
rect 28358 9390 28500 9454
rect 28288 9384 28500 9390
rect 29512 9520 30948 9596
rect 29512 9454 29724 9520
rect 29512 9390 29654 9454
rect 29718 9390 29724 9454
rect 29512 9384 29724 9390
rect 30736 9454 30948 9520
rect 30736 9390 30742 9454
rect 30806 9390 30948 9454
rect 30736 9384 30948 9390
rect 31960 9460 32172 9596
rect 31960 9454 32308 9460
rect 31960 9390 32238 9454
rect 32302 9390 32308 9454
rect 31960 9384 32308 9390
rect 33184 9454 33532 9596
rect 33184 9390 33462 9454
rect 33526 9390 33532 9454
rect 33184 9384 33532 9390
rect 34544 9454 34756 9596
rect 34544 9390 34686 9454
rect 34750 9390 34756 9454
rect 34544 9384 34756 9390
rect 35768 9520 37204 9596
rect 35768 9454 35980 9520
rect 35768 9390 35910 9454
rect 35974 9390 35980 9454
rect 35768 9384 35980 9390
rect 36992 9454 37204 9520
rect 36992 9390 37134 9454
rect 37198 9390 37204 9454
rect 36992 9384 37204 9390
rect 38216 9590 38564 9596
rect 38216 9526 38494 9590
rect 38558 9526 38564 9590
rect 38216 9520 38564 9526
rect 38216 9460 38428 9520
rect 39440 9460 39652 9596
rect 38216 9454 39652 9460
rect 38216 9390 38358 9454
rect 38422 9390 39582 9454
rect 39646 9390 39652 9454
rect 38216 9384 39652 9390
rect 40664 9520 42236 9596
rect 40664 9454 41012 9520
rect 40664 9390 40942 9454
rect 41006 9390 41012 9454
rect 40664 9384 41012 9390
rect 42024 9454 42236 9520
rect 42024 9390 42166 9454
rect 42230 9390 42236 9454
rect 42024 9384 42236 9390
rect 43248 9454 43460 9596
rect 43248 9390 43390 9454
rect 43454 9390 43460 9454
rect 43248 9384 43460 9390
rect 44472 9520 45908 9596
rect 44472 9454 44684 9520
rect 44472 9390 44614 9454
rect 44678 9390 44684 9454
rect 44472 9384 44684 9390
rect 45696 9460 45908 9520
rect 46920 9460 47268 9596
rect 45696 9454 47268 9460
rect 45696 9390 45838 9454
rect 45902 9390 47062 9454
rect 47126 9390 47268 9454
rect 45696 9384 47268 9390
rect 48280 9454 48492 9596
rect 48280 9390 48286 9454
rect 48350 9390 48492 9454
rect 48280 9384 48492 9390
rect 49504 9460 49716 9596
rect 50728 9460 50940 9596
rect 49504 9454 50940 9460
rect 49504 9390 49646 9454
rect 49710 9390 50734 9454
rect 50798 9390 50940 9454
rect 49504 9384 50940 9390
rect 51952 9454 52164 9596
rect 51952 9390 51958 9454
rect 52022 9390 52164 9454
rect 51952 9384 52164 9390
rect 53176 9520 54748 9596
rect 53176 9460 53388 9520
rect 54400 9460 54748 9520
rect 55760 9460 55972 9596
rect 53176 9454 53524 9460
rect 53176 9390 53454 9454
rect 53518 9390 53524 9454
rect 53176 9384 53524 9390
rect 54400 9454 55972 9460
rect 54400 9390 54542 9454
rect 54606 9390 55902 9454
rect 55966 9390 55972 9454
rect 54400 9384 55972 9390
rect 56984 9454 57196 9596
rect 56984 9390 56990 9454
rect 57054 9390 57196 9454
rect 56984 9384 57196 9390
rect 58208 9460 58420 9596
rect 59432 9460 59644 9596
rect 58208 9454 59644 9460
rect 58208 9390 58350 9454
rect 58414 9390 59574 9454
rect 59638 9390 59644 9454
rect 58208 9384 59644 9390
rect 60656 9460 60868 9596
rect 61880 9460 62228 9596
rect 60656 9454 62228 9460
rect 60656 9390 60798 9454
rect 60862 9390 62158 9454
rect 62222 9390 62228 9454
rect 60656 9384 62228 9390
rect 63240 9520 64676 9596
rect 63240 9454 63452 9520
rect 63240 9390 63382 9454
rect 63446 9390 63452 9454
rect 63240 9384 63452 9390
rect 64464 9454 64676 9520
rect 64464 9390 64606 9454
rect 64670 9390 64676 9454
rect 64464 9384 64676 9390
rect 65688 9454 65900 9596
rect 65688 9390 65694 9454
rect 65758 9390 65900 9454
rect 65688 9384 65900 9390
rect 66912 9454 67124 9596
rect 66912 9390 67054 9454
rect 67118 9390 67124 9454
rect 66912 9384 67124 9390
rect 81238 9331 81304 9334
rect 81976 9331 82042 9334
rect 81238 9329 82042 9331
rect 14144 9318 14356 9324
rect 14144 9254 14286 9318
rect 14350 9254 14356 9318
rect 14144 9182 14356 9254
rect 14144 9118 14150 9182
rect 14214 9118 14356 9182
rect 14144 9112 14356 9118
rect 28424 9318 28636 9324
rect 28424 9254 28430 9318
rect 28494 9254 28636 9318
rect 28424 9188 28636 9254
rect 29648 9318 29860 9324
rect 29648 9254 29790 9318
rect 29854 9254 29860 9318
rect 29648 9188 29860 9254
rect 30872 9318 31084 9324
rect 30872 9254 30878 9318
rect 30942 9254 31084 9318
rect 30872 9188 31084 9254
rect 32096 9318 32406 9324
rect 33320 9318 33630 9324
rect 34544 9318 34892 9324
rect 32096 9254 32374 9318
rect 32438 9254 32444 9318
rect 33320 9254 33598 9318
rect 33662 9254 33668 9318
rect 34544 9254 34822 9318
rect 34886 9254 34892 9318
rect 32096 9248 32406 9254
rect 33320 9248 33630 9254
rect 32096 9188 32308 9248
rect 28424 9112 29588 9188
rect 28424 9052 28500 9112
rect 28288 8916 28500 9052
rect 1224 8910 1980 8916
rect 27782 8910 28500 8916
rect 1224 8846 1230 8910
rect 1294 8846 1980 8910
rect 27744 8846 27750 8910
rect 27814 8846 28500 8910
rect 1224 8840 1980 8846
rect 27782 8840 28500 8846
rect 29512 9052 29588 9112
rect 29648 9112 30812 9188
rect 29648 9052 29724 9112
rect 29512 8840 29724 9052
rect 30736 9052 30812 9112
rect 30872 9112 32036 9188
rect 30872 9052 30948 9112
rect 30736 8840 30948 9052
rect 31960 9052 32036 9112
rect 32096 9112 33260 9188
rect 33320 9112 33532 9248
rect 32096 9052 32172 9112
rect 31960 8840 32172 9052
rect 33184 9052 33260 9112
rect 33456 9052 33532 9112
rect 33184 8840 33532 9052
rect 34544 9188 34892 9254
rect 35904 9318 36116 9324
rect 35904 9254 36046 9318
rect 36110 9254 36116 9318
rect 35904 9188 36116 9254
rect 37128 9318 37340 9324
rect 38254 9318 38564 9324
rect 37128 9254 37270 9318
rect 37334 9254 37340 9318
rect 38216 9254 38222 9318
rect 38286 9254 38564 9318
rect 37128 9188 37340 9254
rect 38254 9248 38564 9254
rect 38352 9188 38564 9248
rect 39576 9318 39788 9324
rect 39576 9254 39718 9318
rect 39782 9254 39788 9318
rect 34544 9112 35844 9188
rect 34544 9052 34620 9112
rect 35768 9052 35844 9112
rect 35904 9112 37068 9188
rect 35904 9052 35980 9112
rect 34544 8840 34756 9052
rect 35768 8840 35980 9052
rect 36992 9052 37068 9112
rect 37128 9112 38292 9188
rect 37128 9052 37204 9112
rect 36992 8840 37204 9052
rect 38216 9052 38292 9112
rect 38352 9112 39516 9188
rect 38352 9052 38428 9112
rect 38216 8840 38428 9052
rect 39440 9052 39516 9112
rect 39576 9112 39788 9254
rect 40800 9318 41148 9324
rect 40800 9254 41078 9318
rect 41142 9254 41148 9318
rect 40800 9188 41148 9254
rect 40664 9112 41148 9188
rect 42160 9318 42372 9324
rect 42160 9254 42302 9318
rect 42366 9254 42372 9318
rect 42160 9188 42372 9254
rect 43384 9188 43596 9324
rect 44608 9318 44820 9324
rect 44608 9254 44750 9318
rect 44814 9254 44820 9318
rect 42160 9112 43324 9188
rect 39576 9052 39652 9112
rect 40664 9052 40740 9112
rect 39440 8976 40740 9052
rect 40800 9052 40876 9112
rect 42160 9052 42236 9112
rect 39440 8840 39788 8976
rect 40800 8840 41012 9052
rect 42024 8840 42236 9052
rect 43248 9052 43324 9112
rect 43384 9112 44548 9188
rect 43384 9052 43460 9112
rect 44472 9052 44548 9112
rect 44608 9112 44820 9254
rect 45832 9318 46044 9324
rect 45832 9254 45974 9318
rect 46038 9254 46044 9318
rect 45832 9188 46044 9254
rect 47056 9318 47268 9324
rect 47056 9254 47198 9318
rect 47262 9254 47268 9318
rect 45832 9112 46996 9188
rect 47056 9112 47268 9254
rect 48280 9318 48628 9324
rect 48280 9254 48422 9318
rect 48486 9254 48628 9318
rect 48280 9112 48628 9254
rect 49640 9318 49852 9324
rect 49640 9254 49782 9318
rect 49846 9254 49852 9318
rect 49640 9188 49852 9254
rect 50864 9318 51076 9324
rect 50864 9254 50870 9318
rect 50934 9254 51076 9318
rect 50864 9188 51076 9254
rect 52088 9188 52300 9324
rect 53312 9318 53622 9324
rect 54536 9318 54748 9324
rect 53312 9254 53590 9318
rect 53654 9254 53660 9318
rect 54536 9254 54678 9318
rect 54742 9254 54748 9318
rect 53312 9248 53622 9254
rect 53312 9188 53524 9248
rect 54536 9188 54748 9254
rect 55760 9318 56788 9324
rect 55760 9254 56038 9318
rect 56102 9254 56718 9318
rect 56782 9254 56788 9318
rect 55760 9248 56788 9254
rect 57120 9318 57332 9324
rect 57120 9254 57126 9318
rect 57190 9254 57332 9318
rect 49640 9112 50804 9188
rect 44608 9052 44684 9112
rect 45832 9052 45908 9112
rect 43248 9046 43596 9052
rect 43248 8982 43526 9046
rect 43590 8982 43596 9046
rect 43248 8976 43596 8982
rect 43248 8840 43460 8976
rect 44472 8840 44684 9052
rect 45696 8840 45908 9052
rect 46920 9052 46996 9112
rect 47192 9052 47268 9112
rect 48416 9052 48492 9112
rect 49640 9052 49716 9112
rect 46920 8840 47268 9052
rect 48280 8840 48492 9052
rect 49504 8840 49716 9052
rect 50728 9052 50804 9112
rect 50864 9112 52028 9188
rect 50864 9052 50940 9112
rect 50728 8840 50940 9052
rect 51952 9052 52028 9112
rect 52088 9112 53252 9188
rect 52088 9052 52164 9112
rect 51952 9046 52164 9052
rect 51952 8982 52094 9046
rect 52158 8982 52164 9046
rect 51952 8840 52164 8982
rect 53176 9052 53252 9112
rect 53312 9112 54476 9188
rect 54536 9112 55700 9188
rect 53312 9052 53388 9112
rect 53176 8840 53388 9052
rect 54400 9052 54476 9112
rect 54672 9052 54748 9112
rect 54400 8840 54748 9052
rect 55624 9052 55700 9112
rect 55760 9112 56108 9248
rect 57120 9188 57332 9254
rect 58344 9318 58556 9324
rect 58344 9254 58486 9318
rect 58550 9254 58556 9318
rect 57120 9112 58284 9188
rect 55760 9052 55836 9112
rect 57120 9052 57196 9112
rect 55624 8976 55972 9052
rect 55760 8840 55972 8976
rect 56984 8840 57196 9052
rect 58208 9052 58284 9112
rect 58344 9112 58556 9254
rect 59568 9318 59780 9324
rect 59568 9254 59710 9318
rect 59774 9254 59780 9318
rect 59568 9188 59780 9254
rect 60792 9318 61004 9324
rect 60792 9254 60934 9318
rect 60998 9254 61004 9318
rect 59568 9112 60732 9188
rect 58344 9052 58420 9112
rect 59568 9052 59644 9112
rect 58208 8840 58420 9052
rect 59432 8840 59644 9052
rect 60656 9052 60732 9112
rect 60792 9112 61004 9254
rect 62016 9318 62364 9324
rect 62016 9254 62294 9318
rect 62358 9254 62364 9318
rect 62016 9112 62364 9254
rect 63376 9318 63588 9324
rect 63376 9254 63518 9318
rect 63582 9254 63588 9318
rect 63376 9188 63588 9254
rect 63376 9112 64540 9188
rect 60792 9052 60868 9112
rect 62152 9052 62228 9112
rect 63376 9052 63452 9112
rect 60656 8840 61004 9052
rect 62016 8840 62228 9052
rect 63240 8840 63452 9052
rect 64464 9052 64540 9112
rect 64600 9112 64812 9324
rect 65824 9318 66036 9324
rect 65824 9254 65830 9318
rect 65894 9254 66036 9318
rect 65824 9188 66036 9254
rect 67048 9318 67260 9324
rect 67048 9254 67190 9318
rect 67254 9254 67260 9318
rect 81238 9273 81243 9329
rect 81299 9273 81981 9329
rect 82037 9273 82042 9329
rect 81238 9271 82042 9273
rect 81238 9268 81304 9271
rect 81976 9268 82042 9271
rect 65824 9112 66988 9188
rect 64600 9052 64676 9112
rect 65824 9052 65900 9112
rect 64464 9046 64812 9052
rect 64464 8982 64742 9046
rect 64806 8982 64812 9046
rect 64464 8976 64812 8982
rect 64464 8840 64676 8976
rect 65688 8840 65900 9052
rect 66912 9052 66988 9112
rect 67048 9112 67260 9254
rect 82824 9258 83036 9324
rect 82824 9202 82926 9258
rect 82982 9202 83036 9258
rect 82824 9182 83036 9202
rect 82824 9118 82830 9182
rect 82894 9118 83036 9182
rect 82824 9112 83036 9118
rect 67048 9052 67124 9112
rect 66912 8916 67124 9052
rect 66912 8910 68076 8916
rect 66912 8846 68006 8910
rect 68070 8846 68076 8910
rect 66912 8840 68076 8846
rect 94112 8910 94732 8916
rect 94112 8846 94662 8910
rect 94726 8846 94732 8910
rect 94112 8840 94732 8846
rect 1768 8800 1980 8840
rect 1768 8744 1818 8800
rect 1874 8744 1980 8800
rect 94112 8800 94324 8840
rect 1768 8704 1980 8744
rect 82416 8774 82628 8780
rect 82416 8710 82558 8774
rect 82622 8710 82628 8774
rect 28190 8638 29724 8644
rect 28152 8574 28158 8638
rect 28222 8574 28294 8638
rect 28358 8574 29654 8638
rect 29718 8574 29724 8638
rect 28190 8568 29724 8574
rect 30736 8638 35980 8644
rect 30736 8574 30742 8638
rect 30806 8574 32238 8638
rect 32302 8574 33462 8638
rect 33526 8574 34686 8638
rect 34750 8574 35910 8638
rect 35974 8574 35980 8638
rect 30736 8568 35980 8574
rect 36992 8638 38428 8644
rect 36992 8574 37134 8638
rect 37198 8574 38358 8638
rect 38422 8574 38428 8638
rect 36992 8568 38428 8574
rect 39440 8638 41012 8644
rect 39440 8574 39582 8638
rect 39646 8574 40942 8638
rect 41006 8574 41012 8638
rect 39440 8568 41012 8574
rect 42024 8638 44684 8644
rect 42024 8574 42166 8638
rect 42230 8574 43390 8638
rect 43454 8574 44614 8638
rect 44678 8574 44684 8638
rect 42024 8568 44684 8574
rect 45696 8638 46044 8644
rect 45696 8574 45838 8638
rect 45902 8574 46044 8638
rect 45696 8568 46044 8574
rect 47056 8638 49716 8644
rect 47056 8574 47062 8638
rect 47126 8574 48286 8638
rect 48350 8574 49646 8638
rect 49710 8574 49716 8638
rect 47056 8568 49716 8574
rect 50728 8638 53524 8644
rect 50728 8574 50734 8638
rect 50798 8574 51958 8638
rect 52022 8574 53454 8638
rect 53518 8574 53524 8638
rect 50728 8568 53524 8574
rect 54536 8638 54748 8644
rect 54536 8574 54542 8638
rect 54606 8574 54748 8638
rect 54536 8568 54748 8574
rect 55760 8638 58420 8644
rect 55760 8574 55902 8638
rect 55966 8574 56990 8638
rect 57054 8574 58350 8638
rect 58414 8574 58420 8638
rect 55760 8568 58420 8574
rect 59432 8638 61004 8644
rect 59432 8574 59574 8638
rect 59638 8574 60798 8638
rect 60862 8574 61004 8638
rect 59432 8568 61004 8574
rect 62016 8638 63452 8644
rect 62016 8574 62158 8638
rect 62222 8574 63382 8638
rect 63446 8574 63452 8638
rect 62016 8568 63452 8574
rect 64464 8638 67940 8644
rect 64464 8574 64606 8638
rect 64670 8574 65694 8638
rect 65758 8574 67054 8638
rect 67118 8574 67870 8638
rect 67934 8574 67940 8638
rect 64464 8568 67940 8574
rect 82416 8568 82628 8710
rect 94112 8744 94176 8800
rect 94232 8744 94324 8800
rect 94112 8704 94324 8744
rect 28338 8537 28436 8568
rect 29586 8537 29684 8568
rect 30834 8537 30932 8568
rect 32082 8537 32180 8568
rect 33330 8537 33428 8568
rect 34578 8537 34676 8568
rect 35826 8537 35924 8568
rect 37074 8537 37172 8568
rect 38322 8537 38420 8568
rect 39570 8537 39668 8568
rect 40818 8537 40916 8568
rect 42066 8537 42164 8568
rect 43314 8537 43412 8568
rect 44562 8537 44660 8568
rect 45810 8537 45908 8568
rect 47058 8537 47156 8568
rect 48306 8537 48404 8568
rect 49554 8537 49652 8568
rect 50802 8537 50900 8568
rect 52050 8537 52148 8568
rect 53298 8537 53396 8568
rect 54546 8537 54644 8568
rect 55794 8537 55892 8568
rect 57042 8537 57140 8568
rect 58290 8537 58388 8568
rect 59538 8537 59636 8568
rect 60786 8537 60884 8568
rect 62034 8537 62132 8568
rect 63282 8537 63380 8568
rect 64530 8537 64628 8568
rect 65778 8537 65876 8568
rect 67026 8537 67124 8568
rect 26656 8230 28228 8236
rect 26656 8166 28158 8230
rect 28222 8166 28228 8230
rect 26656 8160 28228 8166
rect 67864 8230 68212 8236
rect 67864 8166 67870 8230
rect 67934 8166 68212 8230
rect 26656 8024 26868 8160
rect 67864 8024 68212 8166
rect 82824 8130 83036 8236
rect 82824 8074 82926 8130
rect 82982 8094 83036 8130
rect 81158 8061 81224 8064
rect 81976 8061 82042 8064
rect 81158 8059 82042 8061
rect 81158 8003 81163 8059
rect 81219 8003 81981 8059
rect 82037 8003 82042 8059
rect 82824 8030 82966 8074
rect 83030 8030 83036 8094
rect 82824 8024 83036 8030
rect 81158 8001 82042 8003
rect 81158 7998 81224 8001
rect 81976 7998 82042 8001
rect 2584 7692 2796 7828
rect 14046 7822 14356 7828
rect 14008 7758 14014 7822
rect 14078 7758 14356 7822
rect 14046 7752 14356 7758
rect 544 7686 2796 7692
rect 544 7622 550 7686
rect 614 7622 2796 7686
rect 544 7616 2796 7622
rect 14144 7686 14356 7752
rect 14144 7622 14286 7686
rect 14350 7622 14356 7686
rect 14144 7616 14356 7622
rect 82416 7414 82628 7420
rect 82416 7350 82422 7414
rect 82486 7350 82628 7414
rect 0 7216 2932 7284
rect 0 7208 2778 7216
rect 2720 7160 2778 7208
rect 2834 7160 2932 7216
rect 1768 7120 1980 7148
rect 1768 7064 1818 7120
rect 1874 7064 1980 7120
rect 2720 7072 2932 7160
rect 26656 7142 27820 7148
rect 26656 7078 27750 7142
rect 27814 7078 27820 7142
rect 26656 7072 27820 7078
rect 67864 7142 68212 7148
rect 67864 7078 68006 7142
rect 68070 7078 68212 7142
rect 1768 7012 1980 7064
rect 1224 7006 2660 7012
rect 1224 6942 1230 7006
rect 1294 6942 2590 7006
rect 2654 6942 2660 7006
rect 1224 6936 2660 6942
rect 26656 6936 26868 7072
rect 67864 6936 68212 7078
rect 82416 7072 82628 7350
rect 94112 7120 94324 7148
rect 94112 7064 94176 7120
rect 94232 7064 94324 7120
rect 94112 7012 94324 7064
rect 94112 7006 94732 7012
rect 94112 6942 94662 7006
rect 94726 6942 94732 7006
rect 94112 6936 94732 6942
rect 2584 6462 2796 6468
rect 2584 6398 2590 6462
rect 2654 6398 2796 6462
rect 2584 6256 2796 6398
rect 14144 6462 14356 6468
rect 14144 6398 14150 6462
rect 14214 6398 14356 6462
rect 14144 6332 14356 6398
rect 14144 6326 15988 6332
rect 14144 6262 15918 6326
rect 15982 6262 15988 6326
rect 14144 6256 15988 6262
rect 0 5576 2932 5652
rect 2720 5516 2932 5576
rect 1797 5440 1895 5461
rect 1797 5384 1818 5440
rect 1874 5384 1895 5440
rect 1797 5380 1895 5384
rect 2720 5460 2778 5516
rect 2834 5460 2932 5516
rect 1224 5374 1980 5380
rect 1224 5310 1230 5374
rect 1294 5310 1980 5374
rect 1224 5304 1980 5310
rect 2720 5304 2932 5460
rect 5848 5621 6196 5652
rect 5848 5565 5999 5621
rect 6055 5565 6196 5621
rect 5848 5510 6196 5565
rect 5848 5446 5854 5510
rect 5918 5446 6196 5510
rect 5848 5440 6196 5446
rect 94112 5440 94324 5516
rect 94112 5384 94176 5440
rect 94232 5384 94324 5440
rect 94112 5380 94324 5384
rect 94112 5374 94732 5380
rect 94112 5310 94662 5374
rect 94726 5310 94732 5374
rect 94112 5304 94732 5310
rect 544 5102 2796 5108
rect 544 5038 550 5102
rect 614 5038 2796 5102
rect 544 5032 2796 5038
rect 2584 4760 2796 5032
rect 14144 5102 14356 5108
rect 14144 5038 14286 5102
rect 14350 5038 14356 5102
rect 14144 4836 14356 5038
rect 14144 4830 16124 4836
rect 14144 4766 16054 4830
rect 16118 4766 16124 4830
rect 14144 4760 16124 4766
rect 1768 3760 1980 3884
rect 1768 3748 1818 3760
rect 1224 3742 1818 3748
rect 1224 3678 1230 3742
rect 1294 3704 1818 3742
rect 1874 3704 1980 3760
rect 1294 3678 1980 3704
rect 1224 3672 1980 3678
rect 15912 3878 17348 3884
rect 15912 3814 15918 3878
rect 15982 3814 17348 3878
rect 15912 3808 17348 3814
rect 15912 3672 16124 3808
rect 17136 3748 17348 3808
rect 18224 3748 18436 3884
rect 19448 3808 21972 3884
rect 19448 3748 19660 3808
rect 17136 3742 19660 3748
rect 17136 3678 17278 3742
rect 17342 3678 19660 3742
rect 17136 3672 19660 3678
rect 20536 3672 20884 3808
rect 21760 3748 21972 3808
rect 22984 3808 25508 3884
rect 22984 3748 23196 3808
rect 21760 3672 23196 3748
rect 24072 3672 24284 3808
rect 25296 3748 25508 3808
rect 26384 3808 29044 3884
rect 26384 3748 26732 3808
rect 25296 3672 26732 3748
rect 27608 3672 27820 3808
rect 28832 3748 29044 3808
rect 29920 3748 30132 3884
rect 31144 3808 33668 3884
rect 31144 3748 31356 3808
rect 28832 3672 31356 3748
rect 32232 3672 32444 3808
rect 33456 3748 33668 3808
rect 34544 3748 34892 3884
rect 35768 3808 37204 3884
rect 35768 3748 35980 3808
rect 33456 3672 35980 3748
rect 36992 3748 37204 3808
rect 38080 3748 38292 3884
rect 39304 3808 41828 3884
rect 39304 3748 39516 3808
rect 36992 3672 39516 3748
rect 40392 3672 40740 3808
rect 41616 3748 41828 3808
rect 42840 3808 45364 3884
rect 42840 3748 43052 3808
rect 41616 3672 43052 3748
rect 43928 3672 44140 3808
rect 45152 3748 45364 3808
rect 46240 3748 46588 3884
rect 47464 3808 48900 3884
rect 47464 3748 47676 3808
rect 45152 3672 47676 3748
rect 48688 3748 48900 3808
rect 49776 3748 49988 3884
rect 51000 3808 53524 3884
rect 51000 3748 51212 3808
rect 48688 3672 51212 3748
rect 52088 3672 52300 3808
rect 53312 3748 53524 3808
rect 54400 3748 54748 3884
rect 55624 3808 57060 3884
rect 55624 3748 55836 3808
rect 53312 3672 55836 3748
rect 56848 3748 57060 3808
rect 57936 3748 58148 3884
rect 56848 3672 58148 3748
rect 94112 3760 94324 3884
rect 94112 3704 94176 3760
rect 94232 3748 94324 3760
rect 94232 3742 94732 3748
rect 94232 3704 94662 3742
rect 94112 3678 94662 3704
rect 94726 3678 94732 3742
rect 94112 3672 94732 3678
rect 15504 2980 15716 3068
rect 15504 2926 15596 2980
rect 15504 2862 15510 2926
rect 15574 2924 15596 2926
rect 15652 2924 15716 2980
rect 15574 2862 15716 2924
rect 15504 2856 15716 2862
rect 16728 2980 16940 3068
rect 17952 3001 18028 3068
rect 19176 3001 19252 3068
rect 20264 3001 20476 3068
rect 21488 3001 21564 3068
rect 16728 2926 16764 2980
rect 16728 2862 16734 2926
rect 16820 2924 16940 2980
rect 17911 2980 18028 3001
rect 17911 2932 17932 2980
rect 16798 2862 16940 2924
rect 16728 2856 16940 2862
rect 17816 2926 17932 2932
rect 17816 2862 17822 2926
rect 17886 2924 17932 2926
rect 17988 2924 18028 2980
rect 19079 2980 19252 3001
rect 19079 2932 19100 2980
rect 17886 2862 18028 2924
rect 17816 2856 18028 2862
rect 19040 2924 19100 2932
rect 19156 2926 19252 2980
rect 20247 2980 20476 3001
rect 20247 2932 20268 2980
rect 19156 2924 19182 2926
rect 19040 2862 19182 2924
rect 19246 2862 19252 2926
rect 19040 2856 19252 2862
rect 20128 2926 20268 2932
rect 20128 2862 20134 2926
rect 20198 2924 20268 2926
rect 20324 2924 20476 2980
rect 21415 2980 21564 3001
rect 21415 2932 21436 2980
rect 20198 2862 20476 2924
rect 20128 2856 20476 2862
rect 21352 2926 21436 2932
rect 21352 2862 21358 2926
rect 21422 2924 21436 2926
rect 21492 2924 21564 2980
rect 21422 2862 21564 2924
rect 21352 2856 21564 2862
rect 22576 2980 22788 3068
rect 23800 3001 23876 3068
rect 22576 2926 22604 2980
rect 22576 2862 22582 2926
rect 22660 2924 22788 2980
rect 23751 2980 23876 3001
rect 23751 2932 23772 2980
rect 22646 2862 22788 2924
rect 22576 2856 22788 2862
rect 23664 2926 23772 2932
rect 23664 2862 23670 2926
rect 23734 2924 23772 2926
rect 23828 2924 23876 2980
rect 23734 2862 23876 2924
rect 23664 2856 23876 2862
rect 24888 2980 25100 3068
rect 26112 3001 26188 3068
rect 27336 3001 27412 3068
rect 28424 3001 28636 3068
rect 29648 3001 29724 3068
rect 24888 2924 24940 2980
rect 24996 2926 25100 2980
rect 26087 2980 26188 3001
rect 26087 2932 26108 2980
rect 24996 2924 25030 2926
rect 24888 2862 25030 2924
rect 25094 2862 25100 2926
rect 24888 2856 25100 2862
rect 25976 2924 26108 2932
rect 26164 2926 26188 2980
rect 27255 2980 27412 3001
rect 27255 2932 27276 2980
rect 25976 2862 26118 2924
rect 26182 2862 26188 2926
rect 25976 2856 26188 2862
rect 27200 2926 27276 2932
rect 27200 2862 27206 2926
rect 27270 2924 27276 2926
rect 27332 2924 27412 2980
rect 28423 2980 28636 3001
rect 28423 2932 28444 2980
rect 27270 2862 27412 2924
rect 27200 2856 27412 2862
rect 28288 2926 28444 2932
rect 28288 2862 28294 2926
rect 28358 2924 28444 2926
rect 28500 2924 28636 2980
rect 29591 2980 29724 3001
rect 29591 2932 29612 2980
rect 28358 2862 28636 2924
rect 28288 2856 28636 2862
rect 29512 2924 29612 2932
rect 29668 2926 29724 2980
rect 29512 2862 29654 2924
rect 29718 2862 29724 2926
rect 29512 2856 29724 2862
rect 30736 2980 30948 3068
rect 31960 3001 32036 3068
rect 33184 3001 33260 3068
rect 34272 3001 34484 3068
rect 35496 3001 35572 3068
rect 30736 2926 30780 2980
rect 30736 2862 30742 2926
rect 30836 2924 30948 2980
rect 31927 2980 32036 3001
rect 31927 2932 31948 2980
rect 30806 2862 30948 2924
rect 30736 2856 30948 2862
rect 31824 2926 31948 2932
rect 31824 2862 31830 2926
rect 31894 2924 31948 2926
rect 32004 2924 32036 2980
rect 33095 2980 33260 3001
rect 33095 2932 33116 2980
rect 31894 2862 32036 2924
rect 31824 2856 32036 2862
rect 33048 2926 33116 2932
rect 33048 2862 33054 2926
rect 33172 2924 33260 2980
rect 34263 2980 34484 3001
rect 34263 2932 34284 2980
rect 33118 2862 33260 2924
rect 33048 2856 33260 2862
rect 34136 2926 34284 2932
rect 34136 2862 34142 2926
rect 34206 2924 34284 2926
rect 34340 2924 34484 2980
rect 35431 2980 35572 3001
rect 35431 2932 35452 2980
rect 34206 2862 34484 2924
rect 34136 2856 34484 2862
rect 35360 2924 35452 2932
rect 35508 2926 35572 2980
rect 35360 2862 35502 2924
rect 35566 2862 35572 2926
rect 35360 2856 35572 2862
rect 36584 2980 36796 3068
rect 37808 3001 37884 3068
rect 39032 3001 39108 3068
rect 40120 3001 40332 3068
rect 41344 3001 41420 3068
rect 36584 2926 36620 2980
rect 36584 2862 36590 2926
rect 36676 2924 36796 2980
rect 37767 2980 37884 3001
rect 37767 2932 37788 2980
rect 36654 2862 36796 2924
rect 36584 2856 36796 2862
rect 37672 2926 37788 2932
rect 37672 2862 37678 2926
rect 37742 2924 37788 2926
rect 37844 2924 37884 2980
rect 38935 2980 39108 3001
rect 38935 2932 38956 2980
rect 37742 2862 37884 2924
rect 37672 2856 37884 2862
rect 38896 2926 38956 2932
rect 38896 2862 38902 2926
rect 39012 2924 39108 2980
rect 40103 2980 40332 3001
rect 40103 2932 40124 2980
rect 38966 2862 39108 2924
rect 38896 2856 39108 2862
rect 39984 2924 40124 2932
rect 40180 2926 40332 2980
rect 41271 2980 41420 3001
rect 41271 2932 41292 2980
rect 40180 2924 40262 2926
rect 39984 2862 40262 2924
rect 40326 2862 40332 2926
rect 39984 2856 40332 2862
rect 41208 2924 41292 2932
rect 41348 2926 41420 2980
rect 41348 2924 41350 2926
rect 41208 2862 41350 2924
rect 41414 2862 41420 2926
rect 41208 2856 41420 2862
rect 42432 2980 42644 3068
rect 43656 3001 43732 3068
rect 42432 2926 42460 2980
rect 42432 2862 42438 2926
rect 42516 2924 42644 2980
rect 43607 2980 43732 3001
rect 43607 2932 43628 2980
rect 42502 2862 42644 2924
rect 42432 2856 42644 2862
rect 43520 2926 43628 2932
rect 43520 2862 43526 2926
rect 43590 2924 43628 2926
rect 43684 2924 43732 2980
rect 43590 2862 43732 2924
rect 43520 2856 43732 2862
rect 44744 2980 44956 3068
rect 45968 3001 46044 3068
rect 47192 3001 47268 3068
rect 48280 3001 48492 3068
rect 49504 3001 49580 3068
rect 44744 2924 44796 2980
rect 44852 2926 44956 2980
rect 45943 2980 46044 3001
rect 45943 2932 45964 2980
rect 44852 2924 44886 2926
rect 44744 2862 44886 2924
rect 44950 2862 44956 2926
rect 44744 2856 44956 2862
rect 45832 2924 45964 2932
rect 46020 2926 46044 2980
rect 47111 2980 47268 3001
rect 47111 2932 47132 2980
rect 45832 2862 45974 2924
rect 46038 2862 46044 2926
rect 45832 2856 46044 2862
rect 47056 2926 47132 2932
rect 47056 2862 47062 2926
rect 47126 2924 47132 2926
rect 47188 2924 47268 2980
rect 48279 2980 48492 3001
rect 48279 2932 48300 2980
rect 47126 2862 47268 2924
rect 47056 2856 47268 2862
rect 48144 2926 48300 2932
rect 48144 2862 48286 2926
rect 48356 2924 48492 2980
rect 49447 2980 49580 3001
rect 49447 2932 49468 2980
rect 48350 2862 48492 2924
rect 48144 2856 48492 2862
rect 49368 2926 49468 2932
rect 49368 2862 49374 2926
rect 49438 2924 49468 2926
rect 49524 2924 49580 2980
rect 49438 2862 49580 2924
rect 49368 2856 49580 2862
rect 50592 2980 50804 3068
rect 51816 3001 51892 3068
rect 53040 3001 53116 3068
rect 54128 3001 54340 3068
rect 55352 3001 55428 3068
rect 50592 2924 50636 2980
rect 50692 2926 50804 2980
rect 51783 2980 51892 3001
rect 51783 2932 51804 2980
rect 50692 2924 50734 2926
rect 50592 2862 50734 2924
rect 50798 2862 50804 2926
rect 50592 2856 50804 2862
rect 51680 2924 51804 2932
rect 51860 2926 51892 2980
rect 52951 2980 53116 3001
rect 52951 2932 52972 2980
rect 51680 2862 51822 2924
rect 51886 2862 51892 2926
rect 51680 2856 51892 2862
rect 52904 2926 52972 2932
rect 52904 2862 52910 2926
rect 53028 2924 53116 2980
rect 54119 2980 54340 3001
rect 54119 2932 54140 2980
rect 52974 2862 53116 2924
rect 52904 2856 53116 2862
rect 53992 2926 54140 2932
rect 53992 2862 53998 2926
rect 54062 2924 54140 2926
rect 54196 2924 54340 2980
rect 55287 2980 55428 3001
rect 55287 2932 55308 2980
rect 54062 2862 54340 2924
rect 53992 2856 54340 2862
rect 55216 2926 55308 2932
rect 55216 2862 55222 2926
rect 55286 2924 55308 2926
rect 55364 2924 55428 2980
rect 55286 2862 55428 2924
rect 55216 2856 55428 2862
rect 56440 2980 56652 3068
rect 57664 3001 57740 3068
rect 56440 2924 56476 2980
rect 56532 2926 56652 2980
rect 57623 2980 57740 3001
rect 57623 2932 57644 2980
rect 56532 2924 56582 2926
rect 56440 2862 56582 2924
rect 56646 2862 56652 2926
rect 56440 2856 56652 2862
rect 57528 2924 57644 2932
rect 57700 2926 57740 2980
rect 57528 2862 57670 2924
rect 57734 2862 57740 2926
rect 57528 2856 57740 2862
rect 14337 2726 14403 2729
rect 14337 2724 16038 2726
rect 14337 2668 14342 2724
rect 14398 2668 16038 2724
rect 14337 2666 16038 2668
rect 14337 2663 14403 2666
rect 15912 2518 17348 2524
rect 15912 2454 16054 2518
rect 16118 2454 17348 2518
rect 15912 2448 17348 2454
rect 15912 2312 16124 2448
rect 17136 2388 17348 2448
rect 18224 2388 18436 2524
rect 19448 2448 21972 2524
rect 19448 2388 19660 2448
rect 17136 2312 19660 2388
rect 20536 2312 20884 2448
rect 21760 2388 21972 2448
rect 22984 2448 25508 2524
rect 22984 2388 23196 2448
rect 21760 2312 23196 2388
rect 24072 2312 24284 2448
rect 25296 2388 25508 2448
rect 26384 2388 26732 2524
rect 27608 2448 29044 2524
rect 27608 2388 27820 2448
rect 25296 2382 27820 2388
rect 25296 2318 26662 2382
rect 26726 2318 27820 2382
rect 25296 2312 27820 2318
rect 28832 2388 29044 2448
rect 29920 2388 30132 2524
rect 31144 2448 33668 2524
rect 31144 2388 31356 2448
rect 28832 2312 31356 2388
rect 32232 2312 32444 2448
rect 33456 2388 33668 2448
rect 34544 2388 34892 2524
rect 35768 2448 37204 2524
rect 35768 2388 35980 2448
rect 33456 2312 35980 2388
rect 36992 2388 37204 2448
rect 38080 2388 38292 2524
rect 39304 2448 41828 2524
rect 39304 2388 39516 2448
rect 36992 2312 39516 2388
rect 40392 2312 40740 2448
rect 41616 2388 41828 2448
rect 42840 2448 45364 2524
rect 42840 2388 43052 2448
rect 41616 2312 43052 2388
rect 43928 2312 44140 2448
rect 45152 2388 45364 2448
rect 46240 2388 46588 2524
rect 47464 2448 48900 2524
rect 47464 2388 47676 2448
rect 45152 2312 47676 2388
rect 48688 2388 48900 2448
rect 49776 2388 49988 2524
rect 51000 2448 53524 2524
rect 51000 2388 51212 2448
rect 48688 2312 51212 2388
rect 52088 2312 52300 2448
rect 53312 2388 53524 2448
rect 54400 2448 57060 2524
rect 54400 2388 54748 2448
rect 53312 2312 54748 2388
rect 55624 2312 55836 2448
rect 56848 2388 57060 2448
rect 57936 2388 58148 2524
rect 56848 2312 58148 2388
rect 1768 2080 1980 2116
rect 1768 2024 1818 2080
rect 1874 2024 1980 2080
rect 1768 1980 1980 2024
rect 94112 2080 94324 2116
rect 94112 2024 94176 2080
rect 94232 2024 94324 2080
rect 94112 1980 94324 2024
rect 1768 1904 2116 1980
rect 94112 1974 94732 1980
rect 94112 1910 94662 1974
rect 94726 1910 94732 1974
rect 94112 1904 94732 1910
rect 2040 1844 2116 1904
rect 2040 1744 2252 1844
rect 2040 1688 2154 1744
rect 2210 1702 2252 1744
rect 2040 1638 2182 1688
rect 2246 1638 2252 1702
rect 2040 1632 2252 1638
rect 3808 1744 4020 1844
rect 3808 1688 3834 1744
rect 3890 1702 4020 1744
rect 3890 1688 3950 1702
rect 3808 1638 3950 1688
rect 4014 1638 4020 1702
rect 3808 1632 4020 1638
rect 5440 1744 5652 1844
rect 5440 1702 5514 1744
rect 5440 1638 5446 1702
rect 5510 1688 5514 1702
rect 5570 1688 5652 1744
rect 5510 1638 5652 1688
rect 5440 1632 5652 1638
rect 7072 1744 7284 1844
rect 7072 1688 7194 1744
rect 7250 1702 7284 1744
rect 7072 1638 7214 1688
rect 7278 1638 7284 1702
rect 7072 1632 7284 1638
rect 8840 1744 9052 1844
rect 8840 1688 8874 1744
rect 8930 1702 9052 1744
rect 8930 1688 8982 1702
rect 8840 1638 8982 1688
rect 9046 1638 9052 1702
rect 8840 1632 9052 1638
rect 10472 1744 10684 1844
rect 10472 1702 10554 1744
rect 10472 1638 10478 1702
rect 10542 1688 10554 1702
rect 10610 1688 10684 1744
rect 10542 1638 10684 1688
rect 10472 1632 10684 1638
rect 12104 1744 12316 1844
rect 12104 1688 12234 1744
rect 12290 1702 12316 1744
rect 12104 1638 12246 1688
rect 12310 1638 12316 1702
rect 12104 1632 12316 1638
rect 13872 1744 14084 1844
rect 13872 1688 13914 1744
rect 13970 1702 14084 1744
rect 13970 1688 14014 1702
rect 13872 1638 14014 1688
rect 14078 1638 14084 1702
rect 13872 1632 14084 1638
rect 15504 1744 15716 1844
rect 15504 1688 15594 1744
rect 15650 1708 15716 1744
rect 17136 1838 17484 1844
rect 17136 1774 17278 1838
rect 17342 1774 17484 1838
rect 17136 1744 17484 1774
rect 15650 1702 15852 1708
rect 15650 1688 15782 1702
rect 15504 1638 15782 1688
rect 15846 1638 15852 1702
rect 15504 1632 15852 1638
rect 17136 1688 17274 1744
rect 17330 1702 17484 1744
rect 17330 1688 17414 1702
rect 17136 1638 17414 1688
rect 17478 1638 17484 1702
rect 17136 1632 17484 1638
rect 18904 1744 19116 1844
rect 18904 1702 18954 1744
rect 18904 1638 18910 1702
rect 19010 1688 19116 1744
rect 18974 1638 19116 1688
rect 18904 1632 19116 1638
rect 20536 1744 20748 1844
rect 20536 1688 20634 1744
rect 20690 1702 20748 1744
rect 20536 1638 20678 1688
rect 20742 1638 20748 1702
rect 20536 1632 20748 1638
rect 22168 1744 22516 1844
rect 22168 1688 22314 1744
rect 22370 1702 22516 1744
rect 22370 1688 22446 1702
rect 22168 1638 22446 1688
rect 22510 1638 22516 1702
rect 22168 1632 22516 1638
rect 23936 1744 24148 1844
rect 23936 1702 23994 1744
rect 23936 1638 23942 1702
rect 24050 1688 24148 1744
rect 24006 1638 24148 1688
rect 23936 1632 24148 1638
rect 25568 1744 25780 1844
rect 25568 1688 25674 1744
rect 25730 1702 25780 1744
rect 25568 1638 25710 1688
rect 25774 1638 25780 1702
rect 25568 1632 25780 1638
rect 27200 1744 27548 1844
rect 27200 1688 27354 1744
rect 27410 1702 27548 1744
rect 27410 1688 27478 1702
rect 27200 1638 27478 1688
rect 27542 1638 27548 1702
rect 27200 1632 27548 1638
rect 28968 1744 29180 1844
rect 28968 1702 29034 1744
rect 28968 1638 28974 1702
rect 29090 1688 29180 1744
rect 29038 1638 29180 1688
rect 28968 1632 29180 1638
rect 30600 1744 30812 1844
rect 30600 1702 30714 1744
rect 30600 1638 30606 1702
rect 30670 1688 30714 1702
rect 30770 1688 30812 1744
rect 30670 1638 30812 1688
rect 30600 1632 30812 1638
rect 32368 1744 32580 1844
rect 32368 1702 32394 1744
rect 32368 1638 32374 1702
rect 32450 1688 32580 1744
rect 32438 1638 32580 1688
rect 32368 1632 32580 1638
rect 34000 1744 34212 1844
rect 34000 1702 34074 1744
rect 34000 1638 34006 1702
rect 34070 1688 34074 1702
rect 34130 1688 34212 1744
rect 34070 1638 34212 1688
rect 34000 1632 34212 1638
rect 35632 1744 35844 1844
rect 35632 1688 35754 1744
rect 35810 1702 35844 1744
rect 35632 1638 35774 1688
rect 35838 1638 35844 1702
rect 35632 1632 35844 1638
rect 37400 1744 37612 1844
rect 37400 1702 37434 1744
rect 37400 1638 37406 1702
rect 37490 1688 37612 1744
rect 37470 1638 37612 1688
rect 37400 1632 37612 1638
rect 39032 1744 39244 1844
rect 39032 1688 39114 1744
rect 39170 1702 39244 1744
rect 40664 1744 40876 1844
rect 40664 1708 40794 1744
rect 39170 1688 39174 1702
rect 39032 1638 39174 1688
rect 39238 1638 39244 1702
rect 39032 1632 39244 1638
rect 40528 1702 40794 1708
rect 40528 1638 40534 1702
rect 40598 1688 40794 1702
rect 40850 1688 40876 1744
rect 42432 1744 42644 1844
rect 42432 1708 42474 1744
rect 40598 1638 40876 1688
rect 40528 1632 40876 1638
rect 42296 1702 42474 1708
rect 42296 1638 42302 1702
rect 42366 1688 42474 1702
rect 42530 1688 42644 1744
rect 42366 1638 42644 1688
rect 42296 1632 42644 1638
rect 44064 1744 44276 1844
rect 44064 1688 44154 1744
rect 44210 1702 44276 1744
rect 44064 1638 44206 1688
rect 44270 1638 44276 1702
rect 44064 1632 44276 1638
rect 45696 1744 46044 1844
rect 45696 1688 45834 1744
rect 45890 1702 46044 1744
rect 45696 1638 45838 1688
rect 45902 1638 46044 1702
rect 45696 1632 46044 1638
rect 47464 1744 47676 1844
rect 47464 1702 47514 1744
rect 47464 1638 47470 1702
rect 47570 1688 47676 1744
rect 49096 1744 49308 1844
rect 49096 1708 49194 1744
rect 47534 1638 47676 1688
rect 47464 1632 47676 1638
rect 48960 1702 49194 1708
rect 48960 1638 48966 1702
rect 49030 1688 49194 1702
rect 49250 1688 49308 1744
rect 49030 1638 49308 1688
rect 48960 1632 49308 1638
rect 50728 1744 51076 1844
rect 50728 1688 50874 1744
rect 50930 1702 51076 1744
rect 50930 1688 51006 1702
rect 50728 1638 51006 1688
rect 51070 1638 51076 1702
rect 50728 1632 51076 1638
rect 52496 1744 52708 1844
rect 52496 1688 52554 1744
rect 52610 1702 52708 1744
rect 52610 1688 52638 1702
rect 52496 1638 52638 1688
rect 52702 1638 52708 1702
rect 52496 1632 52708 1638
rect 54128 1744 54340 1844
rect 54128 1688 54234 1744
rect 54290 1702 54340 1744
rect 54128 1638 54270 1688
rect 54334 1638 54340 1702
rect 54128 1632 54340 1638
rect 55760 1744 56108 1844
rect 55760 1702 55914 1744
rect 55760 1638 55902 1702
rect 55970 1688 56108 1744
rect 55966 1638 56108 1688
rect 55760 1632 56108 1638
rect 57528 1744 57740 1844
rect 57528 1702 57594 1744
rect 57528 1638 57534 1702
rect 57650 1688 57740 1744
rect 57598 1638 57740 1688
rect 57528 1632 57740 1638
rect 59160 1744 59372 1844
rect 59160 1702 59274 1744
rect 59160 1638 59166 1702
rect 59230 1688 59274 1702
rect 59330 1688 59372 1744
rect 59230 1638 59372 1688
rect 59160 1632 59372 1638
rect 60928 1744 61140 1844
rect 60928 1702 60954 1744
rect 60928 1638 60934 1702
rect 61010 1688 61140 1744
rect 60998 1638 61140 1688
rect 60928 1632 61140 1638
rect 62560 1744 62772 1844
rect 62560 1688 62634 1744
rect 62690 1702 62772 1744
rect 64192 1744 64404 1844
rect 64192 1708 64314 1744
rect 62690 1688 62702 1702
rect 62560 1638 62702 1688
rect 62766 1638 62772 1702
rect 62560 1632 62772 1638
rect 64056 1702 64314 1708
rect 64056 1638 64062 1702
rect 64126 1688 64314 1702
rect 64370 1688 64404 1744
rect 64126 1638 64404 1688
rect 64056 1632 64404 1638
rect 65960 1744 66172 1844
rect 65960 1702 65994 1744
rect 65960 1638 65966 1702
rect 66050 1688 66172 1744
rect 66030 1638 66172 1688
rect 65960 1632 66172 1638
rect 67592 1744 67804 1844
rect 67592 1688 67674 1744
rect 67730 1702 67804 1744
rect 67730 1688 67734 1702
rect 67592 1638 67734 1688
rect 67798 1638 67804 1702
rect 67592 1632 67804 1638
rect 69224 1744 69436 1844
rect 69224 1702 69354 1744
rect 69224 1638 69230 1702
rect 69294 1688 69354 1702
rect 69410 1688 69436 1744
rect 69294 1638 69436 1688
rect 69224 1632 69436 1638
rect 70992 1744 71204 1844
rect 70992 1702 71034 1744
rect 70992 1638 70998 1702
rect 71090 1688 71204 1744
rect 71062 1638 71204 1688
rect 70992 1632 71204 1638
rect 72624 1744 72836 1844
rect 72624 1702 72714 1744
rect 72624 1638 72630 1702
rect 72694 1688 72714 1702
rect 72770 1688 72836 1744
rect 72694 1638 72836 1688
rect 72624 1632 72836 1638
rect 74256 1744 74604 1844
rect 74256 1702 74394 1744
rect 74256 1638 74262 1702
rect 74326 1688 74394 1702
rect 74450 1688 74604 1744
rect 74326 1638 74604 1688
rect 74256 1632 74604 1638
rect 76024 1744 76236 1844
rect 76024 1688 76074 1744
rect 76130 1702 76236 1744
rect 76130 1688 76166 1702
rect 76024 1638 76166 1688
rect 76230 1638 76236 1702
rect 76024 1632 76236 1638
rect 77656 1744 77868 1844
rect 77656 1702 77754 1744
rect 77656 1638 77662 1702
rect 77726 1688 77754 1702
rect 77810 1688 77868 1744
rect 77726 1638 77868 1688
rect 77656 1632 77868 1638
rect 79288 1744 79636 1844
rect 79288 1702 79434 1744
rect 79490 1702 79636 1744
rect 79288 1638 79430 1702
rect 79494 1638 79636 1702
rect 79288 1632 79636 1638
rect 81056 1744 81268 1844
rect 81056 1688 81114 1744
rect 81170 1702 81268 1744
rect 82688 1744 82900 1844
rect 82688 1708 82794 1744
rect 81170 1688 81198 1702
rect 81056 1638 81198 1688
rect 81262 1638 81268 1702
rect 81056 1632 81268 1638
rect 82552 1702 82794 1708
rect 82552 1638 82558 1702
rect 82622 1688 82794 1702
rect 82850 1688 82900 1744
rect 82622 1638 82900 1688
rect 82552 1632 82900 1638
rect 84320 1744 84668 1844
rect 84320 1702 84474 1744
rect 84320 1638 84462 1702
rect 84530 1688 84668 1744
rect 84526 1638 84668 1688
rect 84320 1632 84668 1638
rect 86088 1744 86300 1844
rect 86088 1688 86154 1744
rect 86210 1702 86300 1744
rect 86210 1688 86230 1702
rect 86088 1638 86230 1688
rect 86294 1638 86300 1702
rect 86088 1632 86300 1638
rect 87720 1744 87932 1844
rect 87720 1702 87834 1744
rect 87720 1638 87726 1702
rect 87790 1688 87834 1702
rect 87890 1688 87932 1744
rect 87790 1638 87932 1688
rect 87720 1632 87932 1638
rect 89488 1744 89700 1844
rect 89488 1702 89514 1744
rect 89488 1638 89494 1702
rect 89570 1688 89700 1744
rect 89558 1638 89700 1688
rect 89488 1632 89700 1638
rect 91120 1744 91332 1844
rect 91120 1702 91194 1744
rect 91120 1638 91126 1702
rect 91190 1688 91194 1702
rect 91250 1688 91332 1744
rect 91190 1638 91332 1688
rect 91120 1632 91332 1638
rect 92752 1744 92964 1844
rect 92752 1702 92874 1744
rect 92752 1638 92758 1702
rect 92822 1688 92874 1702
rect 92930 1688 92964 1744
rect 92822 1638 92964 1688
rect 92752 1632 92964 1638
rect 952 1294 95004 1300
rect 952 1230 958 1294
rect 1022 1230 1094 1294
rect 1158 1230 1230 1294
rect 1294 1230 2182 1294
rect 2246 1230 3950 1294
rect 4014 1230 5446 1294
rect 5510 1230 7214 1294
rect 7278 1230 8982 1294
rect 9046 1230 10478 1294
rect 10542 1230 12246 1294
rect 12310 1230 14014 1294
rect 14078 1230 15782 1294
rect 15846 1230 17414 1294
rect 17478 1230 18910 1294
rect 18974 1230 20678 1294
rect 20742 1230 22446 1294
rect 22510 1230 23942 1294
rect 24006 1230 25710 1294
rect 25774 1230 27478 1294
rect 27542 1230 28974 1294
rect 29038 1230 30606 1294
rect 30670 1230 32374 1294
rect 32438 1230 34006 1294
rect 34070 1230 35774 1294
rect 35838 1230 37406 1294
rect 37470 1230 39174 1294
rect 39238 1230 40534 1294
rect 40598 1230 42302 1294
rect 42366 1230 44206 1294
rect 44270 1230 45838 1294
rect 45902 1230 47470 1294
rect 47534 1230 48966 1294
rect 49030 1230 51006 1294
rect 51070 1230 52638 1294
rect 52702 1230 54270 1294
rect 54334 1230 55902 1294
rect 55966 1230 57534 1294
rect 57598 1230 59166 1294
rect 59230 1230 60934 1294
rect 60998 1230 62702 1294
rect 62766 1230 64062 1294
rect 64126 1230 65966 1294
rect 66030 1230 67734 1294
rect 67798 1230 69230 1294
rect 69294 1230 70998 1294
rect 71062 1230 72630 1294
rect 72694 1230 74262 1294
rect 74326 1230 76166 1294
rect 76230 1230 77662 1294
rect 77726 1230 79430 1294
rect 79494 1230 81198 1294
rect 81262 1230 82558 1294
rect 82622 1230 84462 1294
rect 84526 1230 86230 1294
rect 86294 1230 87726 1294
rect 87790 1230 89494 1294
rect 89558 1230 91126 1294
rect 91190 1230 92758 1294
rect 92822 1230 94662 1294
rect 94726 1230 94798 1294
rect 94862 1230 94934 1294
rect 94998 1230 95004 1294
rect 952 1158 95004 1230
rect 952 1094 958 1158
rect 1022 1094 1094 1158
rect 1158 1094 1230 1158
rect 1294 1094 94662 1158
rect 94726 1094 94798 1158
rect 94862 1094 94934 1158
rect 94998 1094 95004 1158
rect 952 1022 95004 1094
rect 952 958 958 1022
rect 1022 958 1094 1022
rect 1158 958 1230 1022
rect 1294 958 94662 1022
rect 94726 958 94798 1022
rect 94862 958 94934 1022
rect 94998 958 95004 1022
rect 952 952 95004 958
rect 272 614 95684 620
rect 272 550 278 614
rect 342 550 414 614
rect 478 550 550 614
rect 614 550 26662 614
rect 26726 550 95342 614
rect 95406 550 95478 614
rect 95542 550 95614 614
rect 95678 550 95684 614
rect 272 478 95684 550
rect 272 414 278 478
rect 342 414 414 478
rect 478 414 550 478
rect 614 414 95342 478
rect 95406 414 95478 478
rect 95542 414 95614 478
rect 95678 414 95684 478
rect 272 342 95684 414
rect 272 278 278 342
rect 342 278 414 342
rect 478 278 550 342
rect 614 278 95342 342
rect 95406 278 95478 342
rect 95542 278 95614 342
rect 95678 278 95684 342
rect 272 272 95684 278
<< via3 >>
rect 278 79158 342 79222
rect 414 79158 478 79222
rect 550 79158 614 79222
rect 95342 79158 95406 79222
rect 95478 79158 95542 79222
rect 95614 79158 95678 79222
rect 278 79022 342 79086
rect 414 79022 478 79086
rect 550 79022 614 79086
rect 95342 79022 95406 79086
rect 95478 79022 95542 79086
rect 95614 79022 95678 79086
rect 278 78886 342 78950
rect 414 78886 478 78950
rect 550 78886 614 78950
rect 78886 78886 78950 78950
rect 82150 78886 82214 78950
rect 95342 78886 95406 78950
rect 95478 78886 95542 78950
rect 95614 78886 95678 78950
rect 958 78478 1022 78542
rect 1094 78478 1158 78542
rect 1230 78478 1294 78542
rect 94662 78478 94726 78542
rect 94798 78478 94862 78542
rect 94934 78478 94998 78542
rect 958 78342 1022 78406
rect 1094 78342 1158 78406
rect 1230 78342 1294 78406
rect 94662 78342 94726 78406
rect 94798 78342 94862 78406
rect 94934 78342 94998 78406
rect 958 78206 1022 78270
rect 1094 78206 1158 78270
rect 1230 78206 1294 78270
rect 2182 78206 2246 78270
rect 3950 78206 4014 78270
rect 5446 78206 5510 78270
rect 7214 78206 7278 78270
rect 8982 78206 9046 78270
rect 10478 78206 10542 78270
rect 12246 78206 12310 78270
rect 14014 78206 14078 78270
rect 15646 78206 15710 78270
rect 17414 78206 17478 78270
rect 18910 78206 18974 78270
rect 20678 78206 20742 78270
rect 22174 78206 22238 78270
rect 23942 78206 24006 78270
rect 25710 78206 25774 78270
rect 27478 78206 27542 78270
rect 28974 78206 29038 78270
rect 30878 78206 30942 78270
rect 32510 78206 32574 78270
rect 34142 78206 34206 78270
rect 35502 78206 35566 78270
rect 37406 78206 37470 78270
rect 39174 78206 39238 78270
rect 40534 78206 40598 78270
rect 42438 78206 42502 78270
rect 44206 78206 44270 78270
rect 45838 78206 45902 78270
rect 47470 78206 47534 78270
rect 49238 78206 49302 78270
rect 50734 78206 50798 78270
rect 52638 78206 52702 78270
rect 54134 78206 54198 78270
rect 55902 78206 55966 78270
rect 57670 78206 57734 78270
rect 59166 78206 59230 78270
rect 60934 78206 60998 78270
rect 62702 78206 62766 78270
rect 64062 78206 64126 78270
rect 65966 78206 66030 78270
rect 67734 78206 67798 78270
rect 69230 78206 69294 78270
rect 71134 78206 71198 78270
rect 72766 78206 72830 78270
rect 74398 78206 74462 78270
rect 76166 78206 76230 78270
rect 77662 78206 77726 78270
rect 79294 78206 79358 78270
rect 81198 78206 81262 78270
rect 82694 78206 82758 78270
rect 84462 78206 84526 78270
rect 86230 78206 86294 78270
rect 87726 78206 87790 78270
rect 89630 78206 89694 78270
rect 91262 78206 91326 78270
rect 92894 78206 92958 78270
rect 94662 78206 94726 78270
rect 94798 78206 94862 78270
rect 94934 78206 94998 78270
rect 2182 77808 2246 77862
rect 2182 77798 2210 77808
rect 2210 77798 2246 77808
rect 3950 77798 4014 77862
rect 5446 77798 5510 77862
rect 7214 77808 7278 77862
rect 7214 77798 7250 77808
rect 7250 77798 7278 77808
rect 8982 77798 9046 77862
rect 10478 77798 10542 77862
rect 12246 77808 12310 77862
rect 12246 77798 12290 77808
rect 12290 77798 12310 77808
rect 14014 77798 14078 77862
rect 15646 77808 15710 77862
rect 15646 77798 15650 77808
rect 15650 77798 15710 77808
rect 17414 77798 17478 77862
rect 18910 77808 18974 77862
rect 18910 77798 18954 77808
rect 18954 77798 18974 77808
rect 20678 77808 20742 77862
rect 20678 77798 20690 77808
rect 20690 77798 20742 77808
rect 22174 77798 22238 77862
rect 23942 77808 24006 77862
rect 23942 77798 23994 77808
rect 23994 77798 24006 77808
rect 25710 77808 25774 77862
rect 25710 77798 25730 77808
rect 25730 77798 25774 77808
rect 27478 77798 27542 77862
rect 28974 77808 29038 77862
rect 28974 77798 29034 77808
rect 29034 77798 29038 77808
rect 30878 77798 30942 77862
rect 29790 77662 29854 77726
rect 32510 77798 32574 77862
rect 34142 77798 34206 77862
rect 35502 77798 35566 77862
rect 37406 77808 37470 77862
rect 37406 77798 37434 77808
rect 37434 77798 37470 77808
rect 39174 77798 39238 77862
rect 40534 77798 40598 77862
rect 42438 77808 42502 77862
rect 42438 77798 42474 77808
rect 42474 77798 42502 77808
rect 44206 77808 44270 77862
rect 44206 77798 44210 77808
rect 44210 77798 44270 77808
rect 45838 77808 45902 77862
rect 45838 77798 45890 77808
rect 45890 77798 45902 77808
rect 47470 77808 47534 77862
rect 47470 77798 47514 77808
rect 47514 77798 47534 77808
rect 49238 77808 49302 77862
rect 49238 77798 49250 77808
rect 49250 77798 49302 77808
rect 50734 77798 50798 77862
rect 52638 77798 52702 77862
rect 54134 77798 54198 77862
rect 55902 77808 55966 77862
rect 55902 77798 55914 77808
rect 55914 77798 55966 77808
rect 57670 77798 57734 77862
rect 59166 77798 59230 77862
rect 60934 77808 60998 77862
rect 60934 77798 60954 77808
rect 60954 77798 60998 77808
rect 62702 77798 62766 77862
rect 64062 77798 64126 77862
rect 65966 77808 66030 77862
rect 65966 77798 65994 77808
rect 65994 77798 66030 77808
rect 67734 77798 67798 77862
rect 69230 77798 69294 77862
rect 71134 77798 71198 77862
rect 72766 77808 72830 77862
rect 72766 77798 72770 77808
rect 72770 77798 72830 77808
rect 74398 77808 74462 77862
rect 74398 77798 74450 77808
rect 74450 77798 74462 77808
rect 76166 77798 76230 77862
rect 77662 77798 77726 77862
rect 79294 77798 79358 77862
rect 79294 77662 79358 77726
rect 81198 77798 81262 77862
rect 82694 77798 82758 77862
rect 81878 77662 81942 77726
rect 84462 77808 84526 77862
rect 84462 77798 84474 77808
rect 84474 77798 84526 77808
rect 86230 77798 86294 77862
rect 87726 77798 87790 77862
rect 89630 77798 89694 77862
rect 91262 77798 91326 77862
rect 92894 77808 92958 77862
rect 92894 77798 92930 77808
rect 92930 77798 92958 77808
rect 82150 77118 82214 77182
rect 82014 76982 82078 77046
rect 95342 77118 95406 77182
rect 78886 76438 78950 76502
rect 90038 76467 90102 76502
rect 90038 76438 90079 76467
rect 90079 76438 90102 76467
rect 1230 75894 1294 75958
rect 79430 75894 79494 75958
rect 94662 75894 94726 75958
rect 81878 75758 81942 75822
rect 81878 75622 81942 75686
rect 79294 75078 79358 75142
rect 1230 74398 1294 74462
rect 82014 74262 82078 74326
rect 28158 74126 28222 74190
rect 29518 74126 29582 74190
rect 30606 74126 30670 74190
rect 31966 74126 32030 74190
rect 31150 73990 31214 74054
rect 33190 74126 33254 74190
rect 34550 74126 34614 74190
rect 35774 74126 35838 74190
rect 36862 74126 36926 74190
rect 38222 74126 38286 74190
rect 39310 74126 39374 74190
rect 40670 74126 40734 74190
rect 41894 74126 41958 74190
rect 43254 74126 43318 74190
rect 44342 74126 44406 74190
rect 45566 74126 45630 74190
rect 46926 74126 46990 74190
rect 48150 74126 48214 74190
rect 49510 74126 49574 74190
rect 50598 74126 50662 74190
rect 51958 74126 52022 74190
rect 53046 74126 53110 74190
rect 54270 74126 54334 74190
rect 55630 74126 55694 74190
rect 56854 74126 56918 74190
rect 58214 74126 58278 74190
rect 59302 74126 59366 74190
rect 60662 74126 60726 74190
rect 61886 74126 61950 74190
rect 63246 74126 63310 74190
rect 64334 74126 64398 74190
rect 65558 74126 65622 74190
rect 66918 74126 66982 74190
rect 82014 74126 82078 74190
rect 94662 74262 94726 74326
rect 29790 73854 29854 73918
rect 28566 73718 28630 73782
rect 29790 73718 29854 73782
rect 31014 73718 31078 73782
rect 32102 73718 32166 73782
rect 33462 73718 33526 73782
rect 34686 73718 34750 73782
rect 36046 73718 36110 73782
rect 37270 73718 37334 73782
rect 38494 73718 38558 73782
rect 39718 73718 39782 73782
rect 40806 73718 40870 73782
rect 42030 73718 42094 73782
rect 42302 73718 42366 73782
rect 43390 73718 43454 73782
rect 44750 73718 44814 73782
rect 45974 73718 46038 73782
rect 47198 73718 47262 73782
rect 48558 73718 48622 73782
rect 49782 73718 49846 73782
rect 51006 73718 51070 73782
rect 52094 73718 52158 73782
rect 53454 73718 53518 73782
rect 54678 73718 54742 73782
rect 56038 73718 56102 73782
rect 57262 73718 57326 73782
rect 58486 73718 58550 73782
rect 59710 73718 59774 73782
rect 60798 73718 60862 73782
rect 62158 73718 62222 73782
rect 63518 73718 63582 73782
rect 64742 73718 64806 73782
rect 65966 73718 66030 73782
rect 67190 73718 67254 73782
rect 28566 73038 28630 73102
rect 29790 73038 29854 73102
rect 31014 73038 31078 73102
rect 30878 72766 30942 72830
rect 32102 73038 32166 73102
rect 33462 73038 33526 73102
rect 34686 73038 34750 73102
rect 36046 73038 36110 73102
rect 37270 73038 37334 73102
rect 38494 73038 38558 73102
rect 39718 73038 39782 73102
rect 40806 73038 40870 73102
rect 42030 73038 42094 73102
rect 42302 73038 42366 73102
rect 43390 73038 43454 73102
rect 44750 73038 44814 73102
rect 45974 73038 46038 73102
rect 47198 73038 47262 73102
rect 48558 73038 48622 73102
rect 49782 73038 49846 73102
rect 51006 73038 51070 73102
rect 52094 73038 52158 73102
rect 53454 73038 53518 73102
rect 54678 73038 54742 73102
rect 56038 73038 56102 73102
rect 57262 73038 57326 73102
rect 58486 73038 58550 73102
rect 59710 73038 59774 73102
rect 60798 73038 60862 73102
rect 62158 73038 62222 73102
rect 63518 73038 63582 73102
rect 64742 73038 64806 73102
rect 65966 73038 66030 73102
rect 67190 73038 67254 73102
rect 74806 72902 74870 72966
rect 81878 72902 81942 72966
rect 82150 72766 82214 72830
rect 1230 72494 1294 72558
rect 94662 72494 94726 72558
rect 28566 72222 28630 72286
rect 31150 72222 31214 72286
rect 74670 71542 74734 71606
rect 82014 71542 82078 71606
rect 82014 71406 82078 71470
rect 94118 71406 94182 71470
rect 1230 70862 1294 70926
rect 94118 70998 94182 71062
rect 94662 70862 94726 70926
rect 28566 70454 28630 70518
rect 27614 70318 27678 70382
rect 68958 70318 69022 70382
rect 74806 70318 74870 70382
rect 74534 70182 74598 70246
rect 82150 70046 82214 70110
rect 92486 69910 92550 69974
rect 93425 69598 93489 69662
rect 1230 69094 1294 69158
rect 94662 69230 94726 69294
rect 94118 69094 94182 69158
rect 28294 68686 28358 68750
rect 29246 68686 29310 68750
rect 30878 68958 30942 69022
rect 30334 68686 30398 68750
rect 30606 68686 30670 68750
rect 31558 68686 31622 68750
rect 31694 68686 31758 68750
rect 32782 68686 32846 68750
rect 33326 68686 33390 68750
rect 34142 68686 34206 68750
rect 35230 68686 35294 68750
rect 35774 68686 35838 68750
rect 36590 68686 36654 68750
rect 37814 68686 37878 68750
rect 38358 68686 38422 68750
rect 39038 68686 39102 68750
rect 39310 68686 39374 68750
rect 40262 68686 40326 68750
rect 41894 68686 41958 68750
rect 42846 68686 42910 68750
rect 43390 68686 43454 68750
rect 44070 68686 44134 68750
rect 45838 68686 45902 68750
rect 46518 68686 46582 68750
rect 47062 68686 47126 68750
rect 47742 68686 47806 68750
rect 48966 68686 49030 68750
rect 50598 68686 50662 68750
rect 51550 68686 51614 68750
rect 52094 68686 52158 68750
rect 52774 68686 52838 68750
rect 53046 68686 53110 68750
rect 53998 68686 54062 68750
rect 55222 68686 55286 68750
rect 55766 68686 55830 68750
rect 56854 68686 56918 68750
rect 57806 68686 57870 68750
rect 57942 68686 58006 68750
rect 59030 68686 59094 68750
rect 59574 68686 59638 68750
rect 60254 68686 60318 68750
rect 60798 68686 60862 68750
rect 61478 68686 61542 68750
rect 62702 68686 62766 68750
rect 64062 68686 64126 68750
rect 65286 68686 65350 68750
rect 66510 68686 66574 68750
rect 67054 68686 67118 68750
rect 67734 68686 67798 68750
rect 68278 68686 68342 68750
rect 82014 68686 82078 68750
rect 94118 68686 94182 68750
rect 28294 68278 28358 68342
rect 30334 68278 30398 68342
rect 30606 68278 30670 68342
rect 27614 68142 27678 68206
rect 29246 68142 29310 68206
rect 31558 68278 31622 68342
rect 31694 68278 31758 68342
rect 32782 68278 32846 68342
rect 33326 68278 33390 68342
rect 34142 68278 34206 68342
rect 35230 68278 35294 68342
rect 35774 68278 35838 68342
rect 36590 68278 36654 68342
rect 37814 68278 37878 68342
rect 38358 68278 38422 68342
rect 39038 68278 39102 68342
rect 39310 68278 39374 68342
rect 40262 68278 40326 68342
rect 41894 68278 41958 68342
rect 42846 68278 42910 68342
rect 43390 68278 43454 68342
rect 44070 68278 44134 68342
rect 45838 68278 45902 68342
rect 46518 68278 46582 68342
rect 47062 68278 47126 68342
rect 47742 68278 47806 68342
rect 48966 68278 49030 68342
rect 50598 68278 50662 68342
rect 51550 68278 51614 68342
rect 52094 68278 52158 68342
rect 52774 68278 52838 68342
rect 53046 68278 53110 68342
rect 53998 68278 54062 68342
rect 55222 68278 55286 68342
rect 55766 68278 55830 68342
rect 56854 68278 56918 68342
rect 57806 68278 57870 68342
rect 57942 68278 58006 68342
rect 59030 68278 59094 68342
rect 59574 68278 59638 68342
rect 60254 68278 60318 68342
rect 60798 68278 60862 68342
rect 61478 68278 61542 68342
rect 62702 68278 62766 68342
rect 64062 68278 64126 68342
rect 65286 68278 65350 68342
rect 66510 68278 66574 68342
rect 67054 68278 67118 68342
rect 67734 68278 67798 68342
rect 68278 68278 68342 68342
rect 70318 68278 70382 68342
rect 26934 68006 26998 68070
rect 69366 68006 69430 68070
rect 70318 68006 70382 68070
rect 74670 68006 74734 68070
rect 26934 67734 26998 67798
rect 1230 67598 1294 67662
rect 68958 67734 69022 67798
rect 69366 67734 69430 67798
rect 73854 67734 73918 67798
rect 20950 67190 21014 67254
rect 21086 67190 21150 67254
rect 21358 67190 21422 67254
rect 21766 67190 21830 67254
rect 94662 67598 94726 67662
rect 73854 67326 73918 67390
rect 22038 67190 22102 67254
rect 27206 67054 27270 67118
rect 20406 66918 20470 66982
rect 20950 66918 21014 66982
rect 21086 66918 21150 66982
rect 21358 66918 21422 66982
rect 21766 66918 21830 66982
rect 21630 66782 21694 66846
rect 22038 66918 22102 66982
rect 22038 66782 22102 66846
rect 27206 66782 27270 66846
rect 20406 66646 20470 66710
rect 21630 66510 21694 66574
rect 22038 66510 22102 66574
rect 20542 66102 20606 66166
rect 1230 65966 1294 66030
rect 20542 65830 20606 65894
rect 20406 65694 20470 65758
rect 20814 65694 20878 65758
rect 73990 67190 74054 67254
rect 74534 67326 74598 67390
rect 74398 67190 74462 67254
rect 74670 67190 74734 67254
rect 69094 67054 69158 67118
rect 92486 67190 92550 67254
rect 95342 67190 95406 67254
rect 69094 66782 69158 66846
rect 73990 66918 74054 66982
rect 73990 66782 74054 66846
rect 74398 66918 74462 66982
rect 74262 66782 74326 66846
rect 74670 66918 74734 66982
rect 92622 67054 92686 67118
rect 75622 66918 75686 66982
rect 69094 66510 69158 66574
rect 73990 66510 74054 66574
rect 26934 65830 26998 65894
rect 68958 66238 69022 66302
rect 69094 66238 69158 66302
rect 68958 65966 69022 66030
rect 68958 65830 69022 65894
rect 74262 66510 74326 66574
rect 75078 66374 75142 66438
rect 75622 66646 75686 66710
rect 26934 65558 26998 65622
rect 20406 65422 20470 65486
rect 20406 65286 20470 65350
rect 20814 65422 20878 65486
rect 21766 65286 21830 65350
rect 22038 65286 22102 65350
rect 27206 65422 27270 65486
rect 68958 65558 69022 65622
rect 75078 66102 75142 66166
rect 75486 66102 75550 66166
rect 94662 65966 94726 66030
rect 74670 65694 74734 65758
rect 74942 65694 75006 65758
rect 75486 65830 75550 65894
rect 75486 65694 75550 65758
rect 73854 65286 73918 65350
rect 74262 65286 74326 65350
rect 74670 65422 74734 65486
rect 74942 65422 75006 65486
rect 75486 65422 75550 65486
rect 75622 65286 75686 65350
rect 27206 65150 27270 65214
rect 20406 65014 20470 65078
rect 20406 64878 20470 64942
rect 21494 64878 21558 64942
rect 21766 65014 21830 65078
rect 21766 64878 21830 64942
rect 22038 65014 22102 65078
rect 22038 64878 22102 64942
rect 73854 65014 73918 65078
rect 73990 64878 74054 64942
rect 74262 65014 74326 65078
rect 74262 64878 74326 64942
rect 75078 64878 75142 64942
rect 75622 65014 75686 65078
rect 75486 64878 75550 64942
rect 20406 64606 20470 64670
rect 20542 64470 20606 64534
rect 20814 64470 20878 64534
rect 21494 64606 21558 64670
rect 21494 64470 21558 64534
rect 21766 64606 21830 64670
rect 21630 64470 21694 64534
rect 22038 64606 22102 64670
rect 22038 64470 22102 64534
rect 73990 64606 74054 64670
rect 73854 64470 73918 64534
rect 74262 64606 74326 64670
rect 74398 64470 74462 64534
rect 75078 64606 75142 64670
rect 74806 64470 74870 64534
rect 75486 64606 75550 64670
rect 75622 64470 75686 64534
rect 92486 64470 92550 64534
rect 1230 64062 1294 64126
rect 20542 64198 20606 64262
rect 20542 64062 20606 64126
rect 20814 64198 20878 64262
rect 21494 64198 21558 64262
rect 20950 64062 21014 64126
rect 21086 64062 21150 64126
rect 21222 64062 21286 64126
rect 21630 64198 21694 64262
rect 21766 64062 21830 64126
rect 22038 64198 22102 64262
rect 22038 64062 22102 64126
rect 20542 63790 20606 63854
rect 20542 63654 20606 63718
rect 20950 63790 21014 63854
rect 21086 63790 21150 63854
rect 21222 63790 21286 63854
rect 20814 63654 20878 63718
rect 21766 63790 21830 63854
rect 21766 63654 21830 63718
rect 22038 63790 22102 63854
rect 22038 63654 22102 63718
rect 73854 64198 73918 64262
rect 73990 64062 74054 64126
rect 74398 64198 74462 64262
rect 74398 64062 74462 64126
rect 74806 64198 74870 64262
rect 75622 64198 75686 64262
rect 75622 64062 75686 64126
rect 94662 64062 94726 64126
rect 73990 63790 74054 63854
rect 73990 63654 74054 63718
rect 74398 63790 74462 63854
rect 74262 63654 74326 63718
rect 74942 63654 75006 63718
rect 75622 63790 75686 63854
rect 75622 63654 75686 63718
rect 20542 63382 20606 63446
rect 20814 63382 20878 63446
rect 20814 63246 20878 63310
rect 21494 63246 21558 63310
rect 21766 63382 21830 63446
rect 21630 63246 21694 63310
rect 22038 63382 22102 63446
rect 22174 63246 22238 63310
rect 27206 63110 27270 63174
rect 73990 63382 74054 63446
rect 73854 63246 73918 63310
rect 74262 63382 74326 63446
rect 74398 63246 74462 63310
rect 74942 63382 75006 63446
rect 74806 63246 74870 63310
rect 75214 63246 75278 63310
rect 75622 63382 75686 63446
rect 20814 62974 20878 63038
rect 21494 62974 21558 63038
rect 21630 62974 21694 63038
rect 21766 62838 21830 62902
rect 22174 62974 22238 63038
rect 22174 62838 22238 62902
rect 27070 62838 27134 62902
rect 27206 62838 27270 62902
rect 1230 62430 1294 62494
rect 20814 62430 20878 62494
rect 21766 62566 21830 62630
rect 22174 62566 22238 62630
rect 20542 62158 20606 62222
rect 20814 62158 20878 62222
rect 26934 62294 26998 62358
rect 27070 62294 27134 62358
rect 26934 62022 26998 62086
rect 20542 61886 20606 61950
rect 20406 61750 20470 61814
rect 20950 61750 21014 61814
rect 21086 61750 21150 61814
rect 26934 61886 26998 61950
rect 73854 62974 73918 63038
rect 73990 62838 74054 62902
rect 74398 62974 74462 63038
rect 74398 62838 74462 62902
rect 74806 62974 74870 63038
rect 75214 62974 75278 63038
rect 94118 62838 94182 62902
rect 73990 62566 74054 62630
rect 74398 62566 74462 62630
rect 74942 62430 75006 62494
rect 94118 62566 94182 62630
rect 94662 62430 94726 62494
rect 68958 61886 69022 61950
rect 74942 62158 75006 62222
rect 75622 62158 75686 62222
rect 20406 61478 20470 61542
rect 20542 61342 20606 61406
rect 20950 61478 21014 61542
rect 21086 61478 21150 61542
rect 21630 61342 21694 61406
rect 22038 61342 22102 61406
rect 26934 61614 26998 61678
rect 27206 61478 27270 61542
rect 27206 61206 27270 61270
rect 20542 61070 20606 61134
rect 20406 60934 20470 60998
rect 21086 60934 21150 60998
rect 21358 60934 21422 60998
rect 21630 61070 21694 61134
rect 21630 60934 21694 60998
rect 22038 61070 22102 61134
rect 68958 61614 69022 61678
rect 74670 61750 74734 61814
rect 75078 61750 75142 61814
rect 75622 61886 75686 61950
rect 75486 61750 75550 61814
rect 95342 61614 95406 61678
rect 73990 61342 74054 61406
rect 74262 61342 74326 61406
rect 74670 61478 74734 61542
rect 75078 61478 75142 61542
rect 75486 61478 75550 61542
rect 91942 61478 92006 61542
rect 75622 61342 75686 61406
rect 22038 60934 22102 60998
rect 1230 60798 1294 60862
rect 20406 60662 20470 60726
rect 20542 60526 20606 60590
rect 21086 60662 21150 60726
rect 21358 60662 21422 60726
rect 20950 60526 21014 60590
rect 21086 60526 21150 60590
rect 21630 60662 21694 60726
rect 21766 60526 21830 60590
rect 22038 60662 22102 60726
rect 22038 60526 22102 60590
rect 73990 61070 74054 61134
rect 73990 60934 74054 60998
rect 74262 61070 74326 61134
rect 74262 60934 74326 60998
rect 75078 60934 75142 60998
rect 75622 61070 75686 61134
rect 75622 60934 75686 60998
rect 94118 60824 94176 60862
rect 94176 60824 94182 60862
rect 94118 60798 94182 60824
rect 94662 60798 94726 60862
rect 73990 60662 74054 60726
rect 73990 60526 74054 60590
rect 74262 60662 74326 60726
rect 74398 60526 74462 60590
rect 75078 60662 75142 60726
rect 74670 60526 74734 60590
rect 74942 60526 75006 60590
rect 75622 60662 75686 60726
rect 75486 60526 75550 60590
rect 20542 60254 20606 60318
rect 20542 60118 20606 60182
rect 20950 60254 21014 60318
rect 21086 60254 21150 60318
rect 21358 60118 21422 60182
rect 21766 60254 21830 60318
rect 21630 60118 21694 60182
rect 22038 60254 22102 60318
rect 22174 60118 22238 60182
rect 73990 60254 74054 60318
rect 73854 60118 73918 60182
rect 74398 60254 74462 60318
rect 74262 60118 74326 60182
rect 74670 60254 74734 60318
rect 74942 60254 75006 60318
rect 74806 60118 74870 60182
rect 75486 60254 75550 60318
rect 75622 60118 75686 60182
rect 94118 60254 94182 60318
rect 20542 59846 20606 59910
rect 20542 59710 20606 59774
rect 21358 59846 21422 59910
rect 20814 59710 20878 59774
rect 21086 59710 21150 59774
rect 21494 59710 21558 59774
rect 21630 59846 21694 59910
rect 21630 59710 21694 59774
rect 22174 59846 22238 59910
rect 22038 59710 22102 59774
rect 73854 59846 73918 59910
rect 73854 59710 73918 59774
rect 74262 59846 74326 59910
rect 74398 59710 74462 59774
rect 74806 59846 74870 59910
rect 74670 59710 74734 59774
rect 75622 59846 75686 59910
rect 75622 59710 75686 59774
rect 20542 59438 20606 59502
rect 20814 59438 20878 59502
rect 21086 59438 21150 59502
rect 21494 59438 21558 59502
rect 20950 59302 21014 59366
rect 21086 59302 21150 59366
rect 21630 59438 21694 59502
rect 21630 59302 21694 59366
rect 22038 59438 22102 59502
rect 22038 59302 22102 59366
rect 1230 59166 1294 59230
rect 73854 59438 73918 59502
rect 73854 59302 73918 59366
rect 74398 59438 74462 59502
rect 74398 59302 74462 59366
rect 74670 59438 74734 59502
rect 75078 59302 75142 59366
rect 75622 59438 75686 59502
rect 93425 59423 93489 59427
rect 93425 59367 93429 59423
rect 93429 59367 93485 59423
rect 93485 59367 93489 59423
rect 93425 59363 93489 59367
rect 20950 59030 21014 59094
rect 21086 59030 21150 59094
rect 21630 59030 21694 59094
rect 21630 58894 21694 58958
rect 22038 59030 22102 59094
rect 22174 58894 22238 58958
rect 20814 58486 20878 58550
rect 21086 58486 21150 58550
rect 21630 58622 21694 58686
rect 21766 58486 21830 58550
rect 22174 58622 22238 58686
rect 73854 59030 73918 59094
rect 73854 58894 73918 58958
rect 74398 59030 74462 59094
rect 74262 58894 74326 58958
rect 75078 59030 75142 59094
rect 94662 59030 94726 59094
rect 73854 58622 73918 58686
rect 22174 58486 22238 58550
rect 26934 58350 26998 58414
rect 20406 58214 20470 58278
rect 20814 58214 20878 58278
rect 21086 58214 21150 58278
rect 21766 58214 21830 58278
rect 22174 58214 22238 58278
rect 20406 57942 20470 58006
rect 20542 57806 20606 57870
rect 20814 57806 20878 57870
rect 26934 58078 26998 58142
rect 27206 58078 27270 58142
rect 73990 58486 74054 58550
rect 74262 58622 74326 58686
rect 74398 58486 74462 58550
rect 74670 58486 74734 58550
rect 91942 58758 92006 58822
rect 68958 58350 69022 58414
rect 68958 58078 69022 58142
rect 73990 58214 74054 58278
rect 74398 58214 74462 58278
rect 74670 58214 74734 58278
rect 75622 58214 75686 58278
rect 74942 58078 75006 58142
rect 69094 57942 69158 58006
rect 27206 57670 27270 57734
rect 1230 57398 1294 57462
rect 20542 57534 20606 57598
rect 20542 57398 20606 57462
rect 20814 57534 20878 57598
rect 20542 57126 20606 57190
rect 20542 56990 20606 57054
rect 21494 56990 21558 57054
rect 21630 56990 21694 57054
rect 22174 56990 22238 57054
rect 69094 57670 69158 57734
rect 74942 57806 75006 57870
rect 75214 57806 75278 57870
rect 75622 57942 75686 58006
rect 75622 57806 75686 57870
rect 20542 56718 20606 56782
rect 20406 56582 20470 56646
rect 20950 56582 21014 56646
rect 21494 56718 21558 56782
rect 21630 56718 21694 56782
rect 21630 56582 21694 56646
rect 22174 56718 22238 56782
rect 22038 56582 22102 56646
rect 27206 56718 27270 56782
rect 73854 56990 73918 57054
rect 74262 56990 74326 57054
rect 75214 57534 75278 57598
rect 75622 57534 75686 57598
rect 75486 57398 75550 57462
rect 94662 57398 94726 57462
rect 74806 56990 74870 57054
rect 74942 56990 75006 57054
rect 75486 57126 75550 57190
rect 75486 56990 75550 57054
rect 73854 56718 73918 56782
rect 73854 56582 73918 56646
rect 74262 56718 74326 56782
rect 74398 56582 74462 56646
rect 74806 56718 74870 56782
rect 74942 56718 75006 56782
rect 75214 56582 75278 56646
rect 75486 56718 75550 56782
rect 75622 56582 75686 56646
rect 27206 56446 27270 56510
rect 20406 56310 20470 56374
rect 20406 56174 20470 56238
rect 20950 56310 21014 56374
rect 20950 56174 21014 56238
rect 21086 56174 21150 56238
rect 21630 56310 21694 56374
rect 21766 56174 21830 56238
rect 22038 56310 22102 56374
rect 73854 56310 73918 56374
rect 22038 56174 22102 56238
rect 73990 56174 74054 56238
rect 74398 56310 74462 56374
rect 74398 56174 74462 56238
rect 74670 56174 74734 56238
rect 75214 56310 75278 56374
rect 75078 56174 75142 56238
rect 75622 56310 75686 56374
rect 75486 56174 75550 56238
rect 1230 55902 1294 55966
rect 20406 55902 20470 55966
rect 20406 55766 20470 55830
rect 20950 55902 21014 55966
rect 21086 55902 21150 55966
rect 20814 55766 20878 55830
rect 21766 55902 21830 55966
rect 21630 55766 21694 55830
rect 22038 55902 22102 55966
rect 22038 55766 22102 55830
rect 73990 55902 74054 55966
rect 73854 55766 73918 55830
rect 74398 55902 74462 55966
rect 74262 55766 74326 55830
rect 74670 55902 74734 55966
rect 75078 55902 75142 55966
rect 75486 55902 75550 55966
rect 75622 55766 75686 55830
rect 94662 55902 94726 55966
rect 20406 55494 20470 55558
rect 20814 55494 20878 55558
rect 20814 55358 20878 55422
rect 21086 55358 21150 55422
rect 21494 55358 21558 55422
rect 21630 55494 21694 55558
rect 21630 55358 21694 55422
rect 22038 55494 22102 55558
rect 22174 55358 22238 55422
rect 20406 54950 20470 55014
rect 20814 55086 20878 55150
rect 21086 55086 21150 55150
rect 21494 55086 21558 55150
rect 20950 54950 21014 55014
rect 21086 54950 21150 55014
rect 21630 55086 21694 55150
rect 21630 54950 21694 55014
rect 22174 55086 22238 55150
rect 22038 54950 22102 55014
rect 20406 54678 20470 54742
rect 20950 54678 21014 54742
rect 21086 54678 21150 54742
rect 21494 54542 21558 54606
rect 21630 54678 21694 54742
rect 21630 54542 21694 54606
rect 22038 54678 22102 54742
rect 73854 55494 73918 55558
rect 73990 55358 74054 55422
rect 74262 55494 74326 55558
rect 74398 55358 74462 55422
rect 75214 55358 75278 55422
rect 75622 55494 75686 55558
rect 73990 55086 74054 55150
rect 73854 54950 73918 55014
rect 74398 55086 74462 55150
rect 74262 54950 74326 55014
rect 74670 54950 74734 55014
rect 75214 55086 75278 55150
rect 75622 54950 75686 55014
rect 22038 54542 22102 54606
rect 73854 54678 73918 54742
rect 73854 54542 73918 54606
rect 74262 54678 74326 54742
rect 74262 54542 74326 54606
rect 74670 54678 74734 54742
rect 75214 54542 75278 54606
rect 75622 54678 75686 54742
rect 20406 54270 20470 54334
rect 21494 54270 21558 54334
rect 21630 54270 21694 54334
rect 22038 54270 22102 54334
rect 1230 53998 1294 54062
rect 20406 53998 20470 54062
rect 20542 53862 20606 53926
rect 21494 53862 21558 53926
rect 20542 53590 20606 53654
rect 20542 53454 20606 53518
rect 21494 53590 21558 53654
rect 27070 53998 27134 54062
rect 27206 53998 27270 54062
rect 73854 54270 73918 54334
rect 74262 54270 74326 54334
rect 68958 53998 69022 54062
rect 27206 53726 27270 53790
rect 20542 53182 20606 53246
rect 20406 53046 20470 53110
rect 20950 53046 21014 53110
rect 21086 53046 21150 53110
rect 21766 53046 21830 53110
rect 22038 53046 22102 53110
rect 26934 53590 26998 53654
rect 27070 53590 27134 53654
rect 26934 53318 26998 53382
rect 68958 53726 69022 53790
rect 75214 54270 75278 54334
rect 75486 54270 75550 54334
rect 74670 53862 74734 53926
rect 75078 53862 75142 53926
rect 75486 53998 75550 54062
rect 94662 53998 94726 54062
rect 75486 53862 75550 53926
rect 69094 53590 69158 53654
rect 69094 53318 69158 53382
rect 20406 52774 20470 52838
rect 20542 52638 20606 52702
rect 20950 52774 21014 52838
rect 21086 52774 21150 52838
rect 21766 52774 21830 52838
rect 21630 52638 21694 52702
rect 22038 52774 22102 52838
rect 22038 52638 22102 52702
rect 27206 52774 27270 52838
rect 73990 53046 74054 53110
rect 74670 53590 74734 53654
rect 75078 53590 75142 53654
rect 74942 53454 75006 53518
rect 75486 53590 75550 53654
rect 75622 53454 75686 53518
rect 74262 53046 74326 53110
rect 74942 53182 75006 53246
rect 74670 53046 74734 53110
rect 75622 53182 75686 53246
rect 75486 53046 75550 53110
rect 69094 52774 69158 52838
rect 73990 52774 74054 52838
rect 73854 52638 73918 52702
rect 74262 52774 74326 52838
rect 74398 52638 74462 52702
rect 74670 52774 74734 52838
rect 74806 52638 74870 52702
rect 75486 52774 75550 52838
rect 75486 52638 75550 52702
rect 1230 52366 1294 52430
rect 27206 52502 27270 52566
rect 20542 52366 20606 52430
rect 20542 52230 20606 52294
rect 20950 52230 21014 52294
rect 21086 52230 21150 52294
rect 21222 52230 21286 52294
rect 21630 52366 21694 52430
rect 21630 52230 21694 52294
rect 22038 52366 22102 52430
rect 22038 52230 22102 52294
rect 69094 52502 69158 52566
rect 20542 51958 20606 52022
rect 20542 51822 20606 51886
rect 20950 51958 21014 52022
rect 21086 51958 21150 52022
rect 21222 51958 21286 52022
rect 21494 51822 21558 51886
rect 21630 51958 21694 52022
rect 21766 51822 21830 51886
rect 22038 51958 22102 52022
rect 22174 51822 22238 51886
rect 20542 51550 20606 51614
rect 20814 51414 20878 51478
rect 21494 51550 21558 51614
rect 21358 51414 21422 51478
rect 21766 51550 21830 51614
rect 21630 51414 21694 51478
rect 22174 51550 22238 51614
rect 73854 52366 73918 52430
rect 73990 52230 74054 52294
rect 74398 52366 74462 52430
rect 74262 52230 74326 52294
rect 74806 52366 74870 52430
rect 74670 52230 74734 52294
rect 75486 52366 75550 52430
rect 94662 52366 94726 52430
rect 75486 52230 75550 52294
rect 73990 51958 74054 52022
rect 73990 51822 74054 51886
rect 74262 51958 74326 52022
rect 74398 51822 74462 51886
rect 74670 51958 74734 52022
rect 74942 51822 75006 51886
rect 75486 51958 75550 52022
rect 75486 51822 75550 51886
rect 22038 51414 22102 51478
rect 73990 51550 74054 51614
rect 73854 51414 73918 51478
rect 74398 51550 74462 51614
rect 74398 51414 74462 51478
rect 74942 51550 75006 51614
rect 74806 51414 74870 51478
rect 75486 51550 75550 51614
rect 20406 51006 20470 51070
rect 20814 51142 20878 51206
rect 21358 51142 21422 51206
rect 20814 51006 20878 51070
rect 21086 51006 21150 51070
rect 21630 51142 21694 51206
rect 21630 51006 21694 51070
rect 22038 51142 22102 51206
rect 22038 51006 22102 51070
rect 73854 51142 73918 51206
rect 73854 51006 73918 51070
rect 74398 51142 74462 51206
rect 74398 51006 74462 51070
rect 74806 51142 74870 51206
rect 75214 51006 75278 51070
rect 75622 51006 75686 51070
rect 1230 50734 1294 50798
rect 20406 50734 20470 50798
rect 20814 50734 20878 50798
rect 21086 50734 21150 50798
rect 21222 50598 21286 50662
rect 21630 50734 21694 50798
rect 21766 50598 21830 50662
rect 22038 50734 22102 50798
rect 22174 50598 22238 50662
rect 73854 50734 73918 50798
rect 73854 50598 73918 50662
rect 74398 50734 74462 50798
rect 74262 50598 74326 50662
rect 74806 50598 74870 50662
rect 75214 50734 75278 50798
rect 75078 50598 75142 50662
rect 75622 50734 75686 50798
rect 94662 50598 94726 50662
rect 20406 50326 20470 50390
rect 21222 50326 21286 50390
rect 21766 50326 21830 50390
rect 21630 50190 21694 50254
rect 22174 50326 22238 50390
rect 22174 50190 22238 50254
rect 20406 50054 20470 50118
rect 21358 49782 21422 49846
rect 21630 49918 21694 49982
rect 22174 49918 22238 49982
rect 73854 50326 73918 50390
rect 73854 50190 73918 50254
rect 74262 50326 74326 50390
rect 74262 50190 74326 50254
rect 74806 50326 74870 50390
rect 75078 50326 75142 50390
rect 75622 50326 75686 50390
rect 69094 49918 69158 49982
rect 73854 49918 73918 49982
rect 20406 49510 20470 49574
rect 21358 49510 21422 49574
rect 20406 49238 20470 49302
rect 1230 49102 1294 49166
rect 20542 49102 20606 49166
rect 27206 49646 27270 49710
rect 27206 49374 27270 49438
rect 21222 49102 21286 49166
rect 74262 49918 74326 49982
rect 75078 49782 75142 49846
rect 75622 50054 75686 50118
rect 68958 49646 69022 49710
rect 69094 49646 69158 49710
rect 68958 49374 69022 49438
rect 20542 48830 20606 48894
rect 20542 48694 20606 48758
rect 21222 48830 21286 48894
rect 21766 48694 21830 48758
rect 22038 48694 22102 48758
rect 69094 48830 69158 48894
rect 75078 49510 75142 49574
rect 75622 49510 75686 49574
rect 75214 49102 75278 49166
rect 75622 49238 75686 49302
rect 75622 49102 75686 49166
rect 94662 49102 94726 49166
rect 73990 48694 74054 48758
rect 74398 48694 74462 48758
rect 20542 48422 20606 48486
rect 20542 48286 20606 48350
rect 20814 48286 20878 48350
rect 21494 48286 21558 48350
rect 21766 48422 21830 48486
rect 21766 48286 21830 48350
rect 22038 48422 22102 48486
rect 22038 48286 22102 48350
rect 69094 48558 69158 48622
rect 75214 48830 75278 48894
rect 75622 48830 75686 48894
rect 75486 48694 75550 48758
rect 73990 48422 74054 48486
rect 73854 48286 73918 48350
rect 74398 48422 74462 48486
rect 74398 48286 74462 48350
rect 74806 48286 74870 48350
rect 75486 48422 75550 48486
rect 75622 48286 75686 48350
rect 20542 48014 20606 48078
rect 20406 47878 20470 47942
rect 20814 48014 20878 48078
rect 21494 48014 21558 48078
rect 21086 47878 21150 47942
rect 21358 47878 21422 47942
rect 21766 48014 21830 48078
rect 21766 47878 21830 47942
rect 22038 48014 22102 48078
rect 22038 47878 22102 47942
rect 73854 48014 73918 48078
rect 73990 47878 74054 47942
rect 74398 48014 74462 48078
rect 74398 47878 74462 47942
rect 74806 48014 74870 48078
rect 75078 47878 75142 47942
rect 75622 48014 75686 48078
rect 75622 47878 75686 47942
rect 20406 47606 20470 47670
rect 1230 47470 1294 47534
rect 20542 47470 20606 47534
rect 21086 47606 21150 47670
rect 21358 47606 21422 47670
rect 21086 47470 21150 47534
rect 21766 47606 21830 47670
rect 21766 47470 21830 47534
rect 22038 47606 22102 47670
rect 22174 47470 22238 47534
rect 73990 47606 74054 47670
rect 73990 47470 74054 47534
rect 74398 47606 74462 47670
rect 74398 47470 74462 47534
rect 75078 47606 75142 47670
rect 74670 47470 74734 47534
rect 75622 47606 75686 47670
rect 75486 47470 75550 47534
rect 94662 47470 94726 47534
rect 20542 47198 20606 47262
rect 20406 47062 20470 47126
rect 21086 47198 21150 47262
rect 20814 47062 20878 47126
rect 21494 47062 21558 47126
rect 21766 47198 21830 47262
rect 21630 47062 21694 47126
rect 22174 47198 22238 47262
rect 22038 47062 22102 47126
rect 73990 47198 74054 47262
rect 73854 47062 73918 47126
rect 74398 47198 74462 47262
rect 74262 47062 74326 47126
rect 74670 47198 74734 47262
rect 74806 47062 74870 47126
rect 74942 47062 75006 47126
rect 75486 47198 75550 47262
rect 75622 47062 75686 47126
rect 20406 46790 20470 46854
rect 20814 46790 20878 46854
rect 20814 46654 20878 46718
rect 21494 46790 21558 46854
rect 21630 46790 21694 46854
rect 21766 46654 21830 46718
rect 22038 46790 22102 46854
rect 22174 46654 22238 46718
rect 20814 46382 20878 46446
rect 1230 45838 1294 45902
rect 21766 46382 21830 46446
rect 21766 46246 21830 46310
rect 22174 46382 22238 46446
rect 22038 46246 22102 46310
rect 21494 45838 21558 45902
rect 21766 45974 21830 46038
rect 22038 45974 22102 46038
rect 73854 46790 73918 46854
rect 73990 46654 74054 46718
rect 74262 46790 74326 46854
rect 74262 46654 74326 46718
rect 74806 46790 74870 46854
rect 74942 46790 75006 46854
rect 74670 46654 74734 46718
rect 75622 46790 75686 46854
rect 68958 46518 69022 46582
rect 68958 46246 69022 46310
rect 73990 46382 74054 46446
rect 73990 46246 74054 46310
rect 74262 46382 74326 46446
rect 74262 46246 74326 46310
rect 74670 46382 74734 46446
rect 68958 45974 69022 46038
rect 73990 45974 74054 46038
rect 20542 45566 20606 45630
rect 21494 45566 21558 45630
rect 21086 45430 21150 45494
rect 20542 45294 20606 45358
rect 20542 45158 20606 45222
rect 21086 45158 21150 45222
rect 21358 45158 21422 45222
rect 27206 45294 27270 45358
rect 68958 45702 69022 45766
rect 69094 45702 69158 45766
rect 69094 45430 69158 45494
rect 74262 45974 74326 46038
rect 74806 45838 74870 45902
rect 74942 45838 75006 45902
rect 74806 45566 74870 45630
rect 74942 45566 75006 45630
rect 74534 45430 74598 45494
rect 75486 45566 75550 45630
rect 94662 45838 94726 45902
rect 68958 45294 69022 45358
rect 27206 45022 27270 45086
rect 20542 44886 20606 44950
rect 20406 44750 20470 44814
rect 21358 44886 21422 44950
rect 21630 44750 21694 44814
rect 22174 44750 22238 44814
rect 68958 45022 69022 45086
rect 69094 44886 69158 44950
rect 75078 45158 75142 45222
rect 75486 45294 75550 45358
rect 75486 45158 75550 45222
rect 74534 45022 74598 45086
rect 73854 44750 73918 44814
rect 74262 44750 74326 44814
rect 75078 44886 75142 44950
rect 74942 44750 75006 44814
rect 20406 44478 20470 44542
rect 20542 44342 20606 44406
rect 21630 44478 21694 44542
rect 21766 44342 21830 44406
rect 22174 44478 22238 44542
rect 22038 44342 22102 44406
rect 1230 43934 1294 43998
rect 20542 44070 20606 44134
rect 20406 43934 20470 43998
rect 21086 43934 21150 43998
rect 21766 44070 21830 44134
rect 21766 43934 21830 43998
rect 22038 44070 22102 44134
rect 22038 43934 22102 43998
rect 69094 44614 69158 44678
rect 75486 44886 75550 44950
rect 75622 44750 75686 44814
rect 73854 44478 73918 44542
rect 73990 44342 74054 44406
rect 74262 44478 74326 44542
rect 74398 44342 74462 44406
rect 74942 44478 75006 44542
rect 74670 44342 74734 44406
rect 75622 44478 75686 44542
rect 75486 44342 75550 44406
rect 69094 44070 69158 44134
rect 73990 44070 74054 44134
rect 73990 43934 74054 43998
rect 74398 44070 74462 44134
rect 74398 43934 74462 43998
rect 74670 44070 74734 44134
rect 74806 43934 74870 43998
rect 75486 44070 75550 44134
rect 75622 43934 75686 43998
rect 94662 43934 94726 43998
rect 20406 43662 20470 43726
rect 20406 43526 20470 43590
rect 21086 43662 21150 43726
rect 20950 43526 21014 43590
rect 21086 43526 21150 43590
rect 21766 43662 21830 43726
rect 21766 43526 21830 43590
rect 22038 43662 22102 43726
rect 69094 43798 69158 43862
rect 22038 43526 22102 43590
rect 20406 43254 20470 43318
rect 20542 43118 20606 43182
rect 20950 43254 21014 43318
rect 21086 43254 21150 43318
rect 21222 43118 21286 43182
rect 21766 43254 21830 43318
rect 21766 43118 21830 43182
rect 22038 43254 22102 43318
rect 22174 43118 22238 43182
rect 73990 43662 74054 43726
rect 73990 43526 74054 43590
rect 74398 43662 74462 43726
rect 74262 43526 74326 43590
rect 74806 43662 74870 43726
rect 74670 43526 74734 43590
rect 75622 43662 75686 43726
rect 75622 43526 75686 43590
rect 73990 43254 74054 43318
rect 73990 43118 74054 43182
rect 74262 43254 74326 43318
rect 74262 43118 74326 43182
rect 74670 43254 74734 43318
rect 74670 43118 74734 43182
rect 75078 43118 75142 43182
rect 75622 43254 75686 43318
rect 75486 43118 75550 43182
rect 20542 42846 20606 42910
rect 20814 42710 20878 42774
rect 21222 42846 21286 42910
rect 21358 42710 21422 42774
rect 21766 42846 21830 42910
rect 22174 42846 22238 42910
rect 25438 42846 25502 42910
rect 21630 42710 21694 42774
rect 73990 42846 74054 42910
rect 22038 42710 22102 42774
rect 1230 42302 1294 42366
rect 73310 42710 73374 42774
rect 73854 42710 73918 42774
rect 74262 42846 74326 42910
rect 74262 42710 74326 42774
rect 74670 42846 74734 42910
rect 75078 42846 75142 42910
rect 74942 42710 75006 42774
rect 75486 42846 75550 42910
rect 69094 42574 69158 42638
rect 20814 42438 20878 42502
rect 21358 42438 21422 42502
rect 21630 42438 21694 42502
rect 21766 42302 21830 42366
rect 22038 42438 22102 42502
rect 22174 42302 22238 42366
rect 25438 42438 25502 42502
rect 21086 41894 21150 41958
rect 21766 42030 21830 42094
rect 21766 41894 21830 41958
rect 22174 42030 22238 42094
rect 22038 41894 22102 41958
rect 69094 42302 69158 42366
rect 73310 42438 73374 42502
rect 73854 42438 73918 42502
rect 73854 42302 73918 42366
rect 74262 42438 74326 42502
rect 74262 42302 74326 42366
rect 74942 42438 75006 42502
rect 74806 42302 74870 42366
rect 75078 42302 75142 42366
rect 94662 42302 94726 42366
rect 73854 42030 73918 42094
rect 73854 41894 73918 41958
rect 74262 42030 74326 42094
rect 74262 41894 74326 41958
rect 74942 41894 75006 41958
rect 20542 41622 20606 41686
rect 21086 41622 21150 41686
rect 20542 41350 20606 41414
rect 20542 41214 20606 41278
rect 21494 41214 21558 41278
rect 21766 41622 21830 41686
rect 22038 41622 22102 41686
rect 20542 40942 20606 41006
rect 20406 40806 20470 40870
rect 21494 40942 21558 41006
rect 21766 40806 21830 40870
rect 27070 41350 27134 41414
rect 69094 41350 69158 41414
rect 73854 41622 73918 41686
rect 74262 41622 74326 41686
rect 74942 41622 75006 41686
rect 75622 41622 75686 41686
rect 27070 41078 27134 41142
rect 22174 40806 22238 40870
rect 27206 40942 27270 41006
rect 27206 40670 27270 40734
rect 1230 40534 1294 40598
rect 20406 40534 20470 40598
rect 20542 40398 20606 40462
rect 21222 40398 21286 40462
rect 21766 40534 21830 40598
rect 21630 40398 21694 40462
rect 22174 40534 22238 40598
rect 69094 41078 69158 41142
rect 68958 40942 69022 41006
rect 73854 40806 73918 40870
rect 75214 41214 75278 41278
rect 75622 41350 75686 41414
rect 75622 41214 75686 41278
rect 74262 40806 74326 40870
rect 68958 40670 69022 40734
rect 75214 40942 75278 41006
rect 75622 40942 75686 41006
rect 75622 40806 75686 40870
rect 94662 40670 94726 40734
rect 22174 40398 22238 40462
rect 20542 40126 20606 40190
rect 20542 39990 20606 40054
rect 21222 40126 21286 40190
rect 20950 39990 21014 40054
rect 21630 40126 21694 40190
rect 21766 39990 21830 40054
rect 22174 40126 22238 40190
rect 22038 39990 22102 40054
rect 20542 39718 20606 39782
rect 20542 39582 20606 39646
rect 20950 39718 21014 39782
rect 20814 39582 20878 39646
rect 21766 39718 21830 39782
rect 21766 39582 21830 39646
rect 22038 39718 22102 39782
rect 22174 39582 22238 39646
rect 73854 40534 73918 40598
rect 73854 40398 73918 40462
rect 74262 40534 74326 40598
rect 74262 40398 74326 40462
rect 75214 40398 75278 40462
rect 75622 40534 75686 40598
rect 75622 40398 75686 40462
rect 69094 40126 69158 40190
rect 73854 40126 73918 40190
rect 73990 39990 74054 40054
rect 74262 40126 74326 40190
rect 74262 39990 74326 40054
rect 74670 39990 74734 40054
rect 75214 40126 75278 40190
rect 75214 39990 75278 40054
rect 75622 40126 75686 40190
rect 75486 39990 75550 40054
rect 69094 39854 69158 39918
rect 73990 39718 74054 39782
rect 73990 39582 74054 39646
rect 74262 39718 74326 39782
rect 74262 39582 74326 39646
rect 74670 39718 74734 39782
rect 75214 39718 75278 39782
rect 74670 39582 74734 39646
rect 74942 39582 75006 39646
rect 75214 39582 75278 39646
rect 75486 39718 75550 39782
rect 75622 39582 75686 39646
rect 20542 39310 20606 39374
rect 20406 39174 20470 39238
rect 20814 39310 20878 39374
rect 20814 39174 20878 39238
rect 21086 39174 21150 39238
rect 21766 39310 21830 39374
rect 21630 39174 21694 39238
rect 22174 39310 22238 39374
rect 22038 39174 22102 39238
rect 73990 39310 74054 39374
rect 73990 39174 74054 39238
rect 74262 39310 74326 39374
rect 74262 39174 74326 39238
rect 74670 39310 74734 39374
rect 74942 39310 75006 39374
rect 75214 39310 75278 39374
rect 75078 39174 75142 39238
rect 75622 39310 75686 39374
rect 75622 39174 75686 39238
rect 1230 38902 1294 38966
rect 20406 38902 20470 38966
rect 20814 38902 20878 38966
rect 21086 38902 21150 38966
rect 21494 38766 21558 38830
rect 21630 38902 21694 38966
rect 21766 38766 21830 38830
rect 22038 38902 22102 38966
rect 22174 38766 22238 38830
rect 73990 38902 74054 38966
rect 73990 38766 74054 38830
rect 74262 38902 74326 38966
rect 74398 38766 74462 38830
rect 74670 38766 74734 38830
rect 75078 38902 75142 38966
rect 75078 38766 75142 38830
rect 75622 38902 75686 38966
rect 94662 38902 94726 38966
rect 21494 38494 21558 38558
rect 21766 38494 21830 38558
rect 21630 38358 21694 38422
rect 22174 38494 22238 38558
rect 22174 38358 22238 38422
rect 21086 37950 21150 38014
rect 21630 38086 21694 38150
rect 21630 37950 21694 38014
rect 22174 38086 22238 38150
rect 73990 38494 74054 38558
rect 73854 38358 73918 38422
rect 74398 38494 74462 38558
rect 74262 38358 74326 38422
rect 74670 38494 74734 38558
rect 75078 38494 75142 38558
rect 22174 37950 22238 38014
rect 26934 37814 26998 37878
rect 20542 37678 20606 37742
rect 21086 37678 21150 37742
rect 21630 37678 21694 37742
rect 22174 37678 22238 37742
rect 1230 37406 1294 37470
rect 20542 37406 20606 37470
rect 20406 37270 20470 37334
rect 20814 37270 20878 37334
rect 26934 37542 26998 37606
rect 27070 37406 27134 37470
rect 73854 38086 73918 38150
rect 73990 37950 74054 38014
rect 74262 38086 74326 38150
rect 74398 37950 74462 38014
rect 74670 37950 74734 38014
rect 73990 37678 74054 37742
rect 74398 37678 74462 37742
rect 68958 37406 69022 37470
rect 20406 36998 20470 37062
rect 20542 36862 20606 36926
rect 20814 36998 20878 37062
rect 20542 36590 20606 36654
rect 20406 36454 20470 36518
rect 21358 36454 21422 36518
rect 21630 36454 21694 36518
rect 27070 37134 27134 37198
rect 22038 36454 22102 36518
rect 20406 36182 20470 36246
rect 20406 36046 20470 36110
rect 20814 36046 20878 36110
rect 21358 36182 21422 36246
rect 21222 36046 21286 36110
rect 21630 36182 21694 36246
rect 21630 36046 21694 36110
rect 22038 36182 22102 36246
rect 22174 36046 22238 36110
rect 68958 37134 69022 37198
rect 68958 36998 69022 37062
rect 68958 36726 69022 36790
rect 74670 37678 74734 37742
rect 75486 37678 75550 37742
rect 74670 37270 74734 37334
rect 74942 37270 75006 37334
rect 75486 37406 75550 37470
rect 75622 37270 75686 37334
rect 94662 37406 94726 37470
rect 73854 36454 73918 36518
rect 74670 36998 74734 37062
rect 74942 36998 75006 37062
rect 75622 36998 75686 37062
rect 75622 36862 75686 36926
rect 74262 36454 74326 36518
rect 74942 36454 75006 36518
rect 75078 36454 75142 36518
rect 75622 36590 75686 36654
rect 75622 36454 75686 36518
rect 69094 36182 69158 36246
rect 73854 36182 73918 36246
rect 73854 36046 73918 36110
rect 74262 36182 74326 36246
rect 74398 36046 74462 36110
rect 74942 36182 75006 36246
rect 75078 36182 75142 36246
rect 75078 36046 75142 36110
rect 75622 36182 75686 36246
rect 75622 36046 75686 36110
rect 20406 35774 20470 35838
rect 20542 35638 20606 35702
rect 20814 35774 20878 35838
rect 21222 35774 21286 35838
rect 20950 35638 21014 35702
rect 21630 35774 21694 35838
rect 21766 35638 21830 35702
rect 22174 35774 22238 35838
rect 69094 35910 69158 35974
rect 22038 35638 22102 35702
rect 1230 35502 1294 35566
rect 73854 35774 73918 35838
rect 73990 35638 74054 35702
rect 74398 35774 74462 35838
rect 74262 35638 74326 35702
rect 74670 35638 74734 35702
rect 75078 35774 75142 35838
rect 75078 35638 75142 35702
rect 75622 35774 75686 35838
rect 75486 35638 75550 35702
rect 94662 35502 94726 35566
rect 20542 35366 20606 35430
rect 20406 35230 20470 35294
rect 20950 35366 21014 35430
rect 20814 35230 20878 35294
rect 21766 35366 21830 35430
rect 21766 35230 21830 35294
rect 22038 35366 22102 35430
rect 22038 35230 22102 35294
rect 13742 34822 13806 34886
rect 20406 34958 20470 35022
rect 20814 34958 20878 35022
rect 20950 34822 21014 34886
rect 21086 34822 21150 34886
rect 21766 34958 21830 35022
rect 21766 34822 21830 34886
rect 22038 34958 22102 35022
rect 73990 35366 74054 35430
rect 73990 35230 74054 35294
rect 74262 35366 74326 35430
rect 74262 35230 74326 35294
rect 74670 35366 74734 35430
rect 75078 35366 75142 35430
rect 74806 35230 74870 35294
rect 74942 35230 75006 35294
rect 75486 35366 75550 35430
rect 75622 35230 75686 35294
rect 22038 34822 22102 34886
rect 20542 34414 20606 34478
rect 20950 34550 21014 34614
rect 21086 34550 21150 34614
rect 21494 34414 21558 34478
rect 21766 34550 21830 34614
rect 21766 34414 21830 34478
rect 22038 34550 22102 34614
rect 22038 34414 22102 34478
rect 73990 34958 74054 35022
rect 73990 34822 74054 34886
rect 74262 34958 74326 35022
rect 74262 34822 74326 34886
rect 74806 34958 74870 35022
rect 74942 34958 75006 35022
rect 75078 34822 75142 34886
rect 75622 34958 75686 35022
rect 73990 34550 74054 34614
rect 73990 34414 74054 34478
rect 74262 34550 74326 34614
rect 74398 34414 74462 34478
rect 74670 34414 74734 34478
rect 75078 34550 75142 34614
rect 75214 34414 75278 34478
rect 75486 34414 75550 34478
rect 20542 34142 20606 34206
rect 21494 34142 21558 34206
rect 21358 34006 21422 34070
rect 21766 34142 21830 34206
rect 21630 34006 21694 34070
rect 22038 34142 22102 34206
rect 73990 34142 74054 34206
rect 22174 34006 22238 34070
rect 1230 33870 1294 33934
rect 73854 34006 73918 34070
rect 74398 34142 74462 34206
rect 74262 34006 74326 34070
rect 74670 34142 74734 34206
rect 75214 34142 75278 34206
rect 74806 34006 74870 34070
rect 74942 34006 75006 34070
rect 75486 34142 75550 34206
rect 20406 33734 20470 33798
rect 21358 33734 21422 33798
rect 21630 33734 21694 33798
rect 21766 33598 21830 33662
rect 22174 33734 22238 33798
rect 22174 33598 22238 33662
rect 13606 33462 13670 33526
rect 20406 33462 20470 33526
rect 21766 33326 21830 33390
rect 22174 33326 22238 33390
rect 20542 32918 20606 32982
rect 20542 32646 20606 32710
rect 20542 32510 20606 32574
rect 20814 32510 20878 32574
rect 21630 32510 21694 32574
rect 27206 33054 27270 33118
rect 27206 32782 27270 32846
rect 73854 33734 73918 33798
rect 73854 33598 73918 33662
rect 74262 33734 74326 33798
rect 74262 33598 74326 33662
rect 74806 33734 74870 33798
rect 74942 33734 75006 33798
rect 94662 33870 94726 33934
rect 75486 33734 75550 33798
rect 73854 33326 73918 33390
rect 74262 33326 74326 33390
rect 74806 33190 74870 33254
rect 74942 33190 75006 33254
rect 75486 33462 75550 33526
rect 68958 33054 69022 33118
rect 68958 32782 69022 32846
rect 22174 32510 22238 32574
rect 1230 32238 1294 32302
rect 20542 32238 20606 32302
rect 13742 32102 13806 32166
rect 20406 32102 20470 32166
rect 20814 32238 20878 32302
rect 20950 32102 21014 32166
rect 21494 32102 21558 32166
rect 21630 32238 21694 32302
rect 21630 32102 21694 32166
rect 22174 32238 22238 32302
rect 22038 32102 22102 32166
rect 27206 32238 27270 32302
rect 13742 31966 13806 32030
rect 27206 31966 27270 32030
rect 20406 31830 20470 31894
rect 20542 31694 20606 31758
rect 20950 31830 21014 31894
rect 21494 31830 21558 31894
rect 21222 31694 21286 31758
rect 21630 31830 21694 31894
rect 21630 31694 21694 31758
rect 22038 31830 22102 31894
rect 74806 32918 74870 32982
rect 74942 32918 75006 32982
rect 75622 32918 75686 32982
rect 73990 32510 74054 32574
rect 74398 32510 74462 32574
rect 74670 32510 74734 32574
rect 75622 32646 75686 32710
rect 75486 32510 75550 32574
rect 73990 32238 74054 32302
rect 73990 32102 74054 32166
rect 74398 32238 74462 32302
rect 74262 32102 74326 32166
rect 74670 32238 74734 32302
rect 74806 32102 74870 32166
rect 75486 32238 75550 32302
rect 94662 32238 94726 32302
rect 75486 32102 75550 32166
rect 22174 31694 22238 31758
rect 73990 31830 74054 31894
rect 73854 31694 73918 31758
rect 74262 31830 74326 31894
rect 74398 31694 74462 31758
rect 74806 31830 74870 31894
rect 74806 31694 74870 31758
rect 75214 31694 75278 31758
rect 75486 31830 75550 31894
rect 75622 31694 75686 31758
rect 20542 31422 20606 31486
rect 20406 31286 20470 31350
rect 21222 31422 21286 31486
rect 20950 31286 21014 31350
rect 21086 31286 21150 31350
rect 21630 31422 21694 31486
rect 21766 31286 21830 31350
rect 22174 31422 22238 31486
rect 22038 31286 22102 31350
rect 20406 31014 20470 31078
rect 20406 30878 20470 30942
rect 20950 31014 21014 31078
rect 21086 31014 21150 31078
rect 20814 30878 20878 30942
rect 21494 30878 21558 30942
rect 21766 31014 21830 31078
rect 21766 30878 21830 30942
rect 22038 31014 22102 31078
rect 22174 30878 22238 30942
rect 73854 31422 73918 31486
rect 73990 31286 74054 31350
rect 74398 31422 74462 31486
rect 74398 31286 74462 31350
rect 74806 31422 74870 31486
rect 75214 31422 75278 31486
rect 75078 31286 75142 31350
rect 75622 31422 75686 31486
rect 75486 31286 75550 31350
rect 73990 31014 74054 31078
rect 13606 30742 13670 30806
rect 73854 30878 73918 30942
rect 74398 31014 74462 31078
rect 74398 30878 74462 30942
rect 74670 30878 74734 30942
rect 75078 31014 75142 31078
rect 75486 31014 75550 31078
rect 75622 30878 75686 30942
rect 1230 30606 1294 30670
rect 13470 30606 13534 30670
rect 20406 30606 20470 30670
rect 20406 30470 20470 30534
rect 20814 30606 20878 30670
rect 21494 30606 21558 30670
rect 21766 30606 21830 30670
rect 21766 30470 21830 30534
rect 22174 30606 22238 30670
rect 22038 30470 22102 30534
rect 73854 30606 73918 30670
rect 73854 30470 73918 30534
rect 74398 30606 74462 30670
rect 74262 30470 74326 30534
rect 74670 30606 74734 30670
rect 74806 30470 74870 30534
rect 75622 30606 75686 30670
rect 75486 30470 75550 30534
rect 94662 30606 94726 30670
rect 20406 30198 20470 30262
rect 21222 30062 21286 30126
rect 21766 30198 21830 30262
rect 21766 30062 21830 30126
rect 22038 30198 22102 30262
rect 22038 30062 22102 30126
rect 73854 30198 73918 30262
rect 73990 30062 74054 30126
rect 74262 30198 74326 30262
rect 74262 30062 74326 30126
rect 74806 30198 74870 30262
rect 74670 30062 74734 30126
rect 74942 30062 75006 30126
rect 75486 30198 75550 30262
rect 20542 29790 20606 29854
rect 20542 29518 20606 29582
rect 13742 29382 13806 29446
rect 13606 29246 13670 29310
rect 21222 29790 21286 29854
rect 21766 29790 21830 29854
rect 21630 29654 21694 29718
rect 22038 29790 22102 29854
rect 22174 29654 22238 29718
rect 21086 29246 21150 29310
rect 21630 29382 21694 29446
rect 22174 29382 22238 29446
rect 73990 29790 74054 29854
rect 73854 29654 73918 29718
rect 74262 29790 74326 29854
rect 74398 29654 74462 29718
rect 74670 29790 74734 29854
rect 74942 29790 75006 29854
rect 75622 29790 75686 29854
rect 1230 28974 1294 29038
rect 20406 28974 20470 29038
rect 21086 28974 21150 29038
rect 20950 28838 21014 28902
rect 20406 28702 20470 28766
rect 20542 28566 20606 28630
rect 21086 28702 21150 28766
rect 20814 28566 20878 28630
rect 27206 29110 27270 29174
rect 27206 28838 27270 28902
rect 27070 28702 27134 28766
rect 68958 29110 69022 29174
rect 68958 28838 69022 28902
rect 73854 29382 73918 29446
rect 74398 29382 74462 29446
rect 74670 29246 74734 29310
rect 75622 29518 75686 29582
rect 68958 28702 69022 28766
rect 69094 28702 69158 28766
rect 20542 28294 20606 28358
rect 20542 28158 20606 28222
rect 20814 28294 20878 28358
rect 21766 28158 21830 28222
rect 22038 28158 22102 28222
rect 27070 28430 27134 28494
rect 68958 28430 69022 28494
rect 74670 28974 74734 29038
rect 75486 28974 75550 29038
rect 94662 28974 94726 29038
rect 74942 28566 75006 28630
rect 75486 28702 75550 28766
rect 75622 28566 75686 28630
rect 69094 28294 69158 28358
rect 73990 28158 74054 28222
rect 74262 28158 74326 28222
rect 74942 28294 75006 28358
rect 75622 28294 75686 28358
rect 75622 28158 75686 28222
rect 13470 27886 13534 27950
rect 13742 27750 13806 27814
rect 20542 27886 20606 27950
rect 20406 27750 20470 27814
rect 21494 27750 21558 27814
rect 21766 27886 21830 27950
rect 21630 27750 21694 27814
rect 22038 27886 22102 27950
rect 22038 27750 22102 27814
rect 73990 27886 74054 27950
rect 20406 27478 20470 27542
rect 1230 27342 1294 27406
rect 20542 27342 20606 27406
rect 21494 27478 21558 27542
rect 20814 27342 20878 27406
rect 21086 27342 21150 27406
rect 21630 27478 21694 27542
rect 21630 27342 21694 27406
rect 22038 27478 22102 27542
rect 22038 27342 22102 27406
rect 27070 27478 27134 27542
rect 73990 27750 74054 27814
rect 74262 27886 74326 27950
rect 74262 27750 74326 27814
rect 74670 27750 74734 27814
rect 75622 27886 75686 27950
rect 75486 27750 75550 27814
rect 69094 27478 69158 27542
rect 73990 27478 74054 27542
rect 73854 27342 73918 27406
rect 74262 27478 74326 27542
rect 74262 27342 74326 27406
rect 74670 27478 74734 27542
rect 75214 27342 75278 27406
rect 75486 27478 75550 27542
rect 75622 27342 75686 27406
rect 94662 27342 94726 27406
rect 27070 27206 27134 27270
rect 20542 27070 20606 27134
rect 20814 27070 20878 27134
rect 21086 27070 21150 27134
rect 20406 26934 20470 26998
rect 20950 26934 21014 26998
rect 21086 26934 21150 26998
rect 21630 27070 21694 27134
rect 21766 26934 21830 26998
rect 22038 27070 22102 27134
rect 22038 26934 22102 26998
rect 69094 27206 69158 27270
rect 73854 27070 73918 27134
rect 73990 26934 74054 26998
rect 74262 27070 74326 27134
rect 74262 26934 74326 26998
rect 74670 26934 74734 26998
rect 75214 27070 75278 27134
rect 75078 26934 75142 26998
rect 75622 27070 75686 27134
rect 75486 26934 75550 26998
rect 20406 26662 20470 26726
rect 13606 26526 13670 26590
rect 20542 26526 20606 26590
rect 20950 26662 21014 26726
rect 21086 26662 21150 26726
rect 20814 26526 20878 26590
rect 21494 26526 21558 26590
rect 21766 26662 21830 26726
rect 21766 26526 21830 26590
rect 22038 26662 22102 26726
rect 22038 26526 22102 26590
rect 73990 26662 74054 26726
rect 73854 26526 73918 26590
rect 74262 26662 74326 26726
rect 74262 26526 74326 26590
rect 74670 26662 74734 26726
rect 75078 26662 75142 26726
rect 74670 26526 74734 26590
rect 74942 26526 75006 26590
rect 75486 26662 75550 26726
rect 75622 26526 75686 26590
rect 17414 26390 17478 26454
rect 20542 26254 20606 26318
rect 20814 26254 20878 26318
rect 21494 26254 21558 26318
rect 21766 26254 21830 26318
rect 21766 26118 21830 26182
rect 22038 26254 22102 26318
rect 22174 26118 22238 26182
rect 27206 25982 27270 26046
rect 21766 25846 21830 25910
rect 21766 25710 21830 25774
rect 22174 25846 22238 25910
rect 22174 25710 22238 25774
rect 27206 25710 27270 25774
rect 1230 25438 1294 25502
rect 20814 25302 20878 25366
rect 21358 25302 21422 25366
rect 21766 25438 21830 25502
rect 21630 25302 21694 25366
rect 22174 25438 22238 25502
rect 22038 25302 22102 25366
rect 73854 26254 73918 26318
rect 73854 26118 73918 26182
rect 74262 26254 74326 26318
rect 74262 26118 74326 26182
rect 74670 26254 74734 26318
rect 74942 26254 75006 26318
rect 75078 26118 75142 26182
rect 75622 26254 75686 26318
rect 73854 25846 73918 25910
rect 73990 25710 74054 25774
rect 74262 25846 74326 25910
rect 74262 25710 74326 25774
rect 75078 25846 75142 25910
rect 73990 25438 74054 25502
rect 13742 25030 13806 25094
rect 73854 25302 73918 25366
rect 74262 25438 74326 25502
rect 74398 25302 74462 25366
rect 74806 25302 74870 25366
rect 74942 25302 75006 25366
rect 94662 25438 94726 25502
rect 20406 25030 20470 25094
rect 15510 24894 15574 24958
rect 21358 25030 21422 25094
rect 21630 25030 21694 25094
rect 22038 25030 22102 25094
rect 17142 24622 17206 24686
rect 17414 24758 17478 24822
rect 17958 24622 18022 24686
rect 18366 24486 18430 24550
rect 20406 24758 20470 24822
rect 20542 24622 20606 24686
rect 21494 24622 21558 24686
rect 18638 24486 18702 24550
rect 20814 24486 20878 24550
rect 20542 24350 20606 24414
rect 17278 24214 17342 24278
rect 18230 24214 18294 24278
rect 20406 24214 20470 24278
rect 21494 24350 21558 24414
rect 21630 24214 21694 24278
rect 26934 24758 26998 24822
rect 68958 24758 69022 24822
rect 73854 25030 73918 25094
rect 74398 25030 74462 25094
rect 74806 25030 74870 25094
rect 74942 25030 75006 25094
rect 26934 24486 26998 24550
rect 22174 24214 22238 24278
rect 68958 24486 69022 24550
rect 68958 24350 69022 24414
rect 73854 24214 73918 24278
rect 75622 25030 75686 25094
rect 74670 24622 74734 24686
rect 75622 24758 75686 24822
rect 75486 24622 75550 24686
rect 77254 24486 77318 24550
rect 78070 24622 78134 24686
rect 79022 24622 79086 24686
rect 77798 24486 77862 24550
rect 74398 24214 74462 24278
rect 74670 24350 74734 24414
rect 1230 23806 1294 23870
rect 17142 23942 17206 24006
rect 17278 23942 17342 24006
rect 17142 23806 17206 23870
rect 17958 23942 18022 24006
rect 18230 23942 18294 24006
rect 18366 23942 18430 24006
rect 18366 23806 18430 23870
rect 18638 23942 18702 24006
rect 20406 23942 20470 24006
rect 20542 23806 20606 23870
rect 20814 23806 20878 23870
rect 21630 23942 21694 24006
rect 21766 23806 21830 23870
rect 22174 23942 22238 24006
rect 27070 23942 27134 24006
rect 68958 24078 69022 24142
rect 75486 24350 75550 24414
rect 75622 24214 75686 24278
rect 74942 24078 75006 24142
rect 22038 23806 22102 23870
rect 17822 23670 17886 23734
rect 20542 23534 20606 23598
rect 550 23398 614 23462
rect 20406 23398 20470 23462
rect 20814 23534 20878 23598
rect 20950 23398 21014 23462
rect 21494 23398 21558 23462
rect 21766 23534 21830 23598
rect 21766 23398 21830 23462
rect 22038 23534 22102 23598
rect 22038 23398 22102 23462
rect 27070 23534 27134 23598
rect 17142 23126 17206 23190
rect 17006 22990 17070 23054
rect 17822 23126 17886 23190
rect 18366 23126 18430 23190
rect 17686 22990 17750 23054
rect 18366 22990 18430 23054
rect 18774 22990 18838 23054
rect 20406 23126 20470 23190
rect 20542 22990 20606 23054
rect 20950 23126 21014 23190
rect 20814 22990 20878 23054
rect 21494 23126 21558 23190
rect 21766 23126 21830 23190
rect 21630 22990 21694 23054
rect 22038 23126 22102 23190
rect 73854 23942 73918 24006
rect 73990 23806 74054 23870
rect 74398 23942 74462 24006
rect 74398 23806 74462 23870
rect 74942 23806 75006 23870
rect 75214 23806 75278 23870
rect 75622 23942 75686 24006
rect 75486 23806 75550 23870
rect 77254 23942 77318 24006
rect 77798 23942 77862 24006
rect 78070 23942 78134 24006
rect 77662 23806 77726 23870
rect 77798 23806 77862 23870
rect 78342 23806 78406 23870
rect 79022 23942 79086 24006
rect 79022 23806 79086 23870
rect 94662 23806 94726 23870
rect 68958 23534 69022 23598
rect 73990 23534 74054 23598
rect 74398 23534 74462 23598
rect 73990 23398 74054 23462
rect 74262 23398 74326 23462
rect 74806 23398 74870 23462
rect 75214 23534 75278 23598
rect 75486 23534 75550 23598
rect 75486 23398 75550 23462
rect 68958 23262 69022 23326
rect 77662 23262 77726 23326
rect 22038 22990 22102 23054
rect 73990 23126 74054 23190
rect 73854 22990 73918 23054
rect 74262 23126 74326 23190
rect 74398 22990 74462 23054
rect 74806 23126 74870 23190
rect 75214 22990 75278 23054
rect 75486 23126 75550 23190
rect 75622 22990 75686 23054
rect 77798 23126 77862 23190
rect 77254 22990 77318 23054
rect 77798 22990 77862 23054
rect 78342 23126 78406 23190
rect 78614 22990 78678 23054
rect 79022 23126 79086 23190
rect 78886 22990 78950 23054
rect 20542 22718 20606 22782
rect 2561 22665 2625 22669
rect 2561 22609 2565 22665
rect 2565 22609 2621 22665
rect 2621 22609 2625 22665
rect 2561 22605 2625 22609
rect 20406 22582 20470 22646
rect 20814 22718 20878 22782
rect 21630 22718 21694 22782
rect 21766 22582 21830 22646
rect 22038 22718 22102 22782
rect 22038 22582 22102 22646
rect 73854 22718 73918 22782
rect 73990 22582 74054 22646
rect 74398 22718 74462 22782
rect 74262 22582 74326 22646
rect 74670 22582 74734 22646
rect 75214 22718 75278 22782
rect 75078 22582 75142 22646
rect 75622 22718 75686 22782
rect 75486 22582 75550 22646
rect 1230 22174 1294 22238
rect 15510 22310 15574 22374
rect 17006 22310 17070 22374
rect 17686 22310 17750 22374
rect 17278 22174 17342 22238
rect 18366 22310 18430 22374
rect 18774 22310 18838 22374
rect 18502 22174 18566 22238
rect 18638 22174 18702 22238
rect 20406 22310 20470 22374
rect 20814 22174 20878 22238
rect 21494 22174 21558 22238
rect 21766 22310 21830 22374
rect 21766 22174 21830 22238
rect 22038 22310 22102 22374
rect 22174 22174 22238 22238
rect 73990 22310 74054 22374
rect 26934 22038 26998 22102
rect 73854 22174 73918 22238
rect 74262 22310 74326 22374
rect 74262 22174 74326 22238
rect 74670 22310 74734 22374
rect 75078 22310 75142 22374
rect 74806 22174 74870 22238
rect 74942 22174 75006 22238
rect 75214 22174 75278 22238
rect 75486 22310 75550 22374
rect 77254 22310 77318 22374
rect 77390 22174 77454 22238
rect 77798 22310 77862 22374
rect 78614 22310 78678 22374
rect 78886 22310 78950 22374
rect 94662 22310 94726 22374
rect 20814 21902 20878 21966
rect 21494 21902 21558 21966
rect 21766 21902 21830 21966
rect 21766 21766 21830 21830
rect 22174 21902 22238 21966
rect 22038 21766 22102 21830
rect 26934 21766 26998 21830
rect 18502 21630 18566 21694
rect 21086 21358 21150 21422
rect 21766 21494 21830 21558
rect 21766 21358 21830 21422
rect 22038 21494 22102 21558
rect 69094 21766 69158 21830
rect 73854 21902 73918 21966
rect 73854 21766 73918 21830
rect 74262 21902 74326 21966
rect 74398 21766 74462 21830
rect 74806 21902 74870 21966
rect 74942 21902 75006 21966
rect 75214 21902 75278 21966
rect 68958 21494 69022 21558
rect 73854 21494 73918 21558
rect 22038 21358 22102 21422
rect 69094 21358 69158 21422
rect 73990 21358 74054 21422
rect 74398 21494 74462 21558
rect 74398 21358 74462 21422
rect 75078 21358 75142 21422
rect 78478 22038 78542 22102
rect 20542 21086 20606 21150
rect 21086 21086 21150 21150
rect 21766 21086 21830 21150
rect 22038 21086 22102 21150
rect 17278 20814 17342 20878
rect 1230 20406 1294 20470
rect 16462 20542 16526 20606
rect 17414 20542 17478 20606
rect 17822 20542 17886 20606
rect 18366 20542 18430 20606
rect 18638 20814 18702 20878
rect 20542 20814 20606 20878
rect 20406 20678 20470 20742
rect 21494 20678 21558 20742
rect 18774 20542 18838 20606
rect 27206 20814 27270 20878
rect 68958 21086 69022 21150
rect 69094 20814 69158 20878
rect 73990 21086 74054 21150
rect 74398 21086 74462 21150
rect 75078 21086 75142 21150
rect 75486 21086 75550 21150
rect 3814 20406 3878 20470
rect 20406 20406 20470 20470
rect 20406 20270 20470 20334
rect 21494 20406 21558 20470
rect 16462 19998 16526 20062
rect 17414 19998 17478 20062
rect 17822 19998 17886 20062
rect 18366 19998 18430 20062
rect 18230 19862 18294 19926
rect 18774 19998 18838 20062
rect 18638 19862 18702 19926
rect 20406 19998 20470 20062
rect 20406 19862 20470 19926
rect 20814 19862 20878 19926
rect 21494 19862 21558 19926
rect 21630 19862 21694 19926
rect 22038 19862 22102 19926
rect 26934 20406 26998 20470
rect 27206 20406 27270 20470
rect 26934 20134 26998 20198
rect 27070 20134 27134 20198
rect 69094 20542 69158 20606
rect 69094 19998 69158 20062
rect 74670 20678 74734 20742
rect 75486 20814 75550 20878
rect 75486 20678 75550 20742
rect 77390 20814 77454 20878
rect 77662 20542 77726 20606
rect 78478 20814 78542 20878
rect 78206 20542 78270 20606
rect 78614 20542 78678 20606
rect 74670 20406 74734 20470
rect 75486 20406 75550 20470
rect 79430 20406 79494 20470
rect 94662 20406 94726 20470
rect 75486 20270 75550 20334
rect 27070 19862 27134 19926
rect 20406 19590 20470 19654
rect 20406 19454 20470 19518
rect 20814 19590 20878 19654
rect 20950 19454 21014 19518
rect 21494 19590 21558 19654
rect 21630 19590 21694 19654
rect 21630 19454 21694 19518
rect 22038 19590 22102 19654
rect 22174 19454 22238 19518
rect 73854 19862 73918 19926
rect 74262 19862 74326 19926
rect 75486 19998 75550 20062
rect 75622 19862 75686 19926
rect 77662 19998 77726 20062
rect 78206 19998 78270 20062
rect 78206 19862 78270 19926
rect 78614 19998 78678 20062
rect 79430 19998 79494 20062
rect 78614 19862 78678 19926
rect 69094 19590 69158 19654
rect 73854 19590 73918 19654
rect 73854 19454 73918 19518
rect 74262 19590 74326 19654
rect 74262 19454 74326 19518
rect 75622 19590 75686 19654
rect 75214 19454 75278 19518
rect 75486 19454 75550 19518
rect 20406 19182 20470 19246
rect 20406 19046 20470 19110
rect 20950 19182 21014 19246
rect 21358 19046 21422 19110
rect 21630 19182 21694 19246
rect 21630 19046 21694 19110
rect 22174 19182 22238 19246
rect 22038 19046 22102 19110
rect 1230 18910 1294 18974
rect 20406 18774 20470 18838
rect 20406 18638 20470 18702
rect 20814 18638 20878 18702
rect 21358 18774 21422 18838
rect 21222 18638 21286 18702
rect 21630 18774 21694 18838
rect 21630 18638 21694 18702
rect 22038 18774 22102 18838
rect 22038 18638 22102 18702
rect 73854 19182 73918 19246
rect 73854 19046 73918 19110
rect 74262 19182 74326 19246
rect 74262 19046 74326 19110
rect 74806 19046 74870 19110
rect 75214 19182 75278 19246
rect 75486 19182 75550 19246
rect 75486 19046 75550 19110
rect 73854 18774 73918 18838
rect 73854 18638 73918 18702
rect 74262 18774 74326 18838
rect 74262 18638 74326 18702
rect 74806 18774 74870 18838
rect 75078 18638 75142 18702
rect 75486 18774 75550 18838
rect 94662 18774 94726 18838
rect 75622 18638 75686 18702
rect 77934 18638 77998 18702
rect 78478 18638 78542 18702
rect 17550 18230 17614 18294
rect 18230 18366 18294 18430
rect 18230 18230 18294 18294
rect 18638 18366 18702 18430
rect 18774 18230 18838 18294
rect 20406 18366 20470 18430
rect 20814 18366 20878 18430
rect 21222 18366 21286 18430
rect 20950 18230 21014 18294
rect 21630 18366 21694 18430
rect 21766 18230 21830 18294
rect 22038 18366 22102 18430
rect 22174 18230 22238 18294
rect 73854 18366 73918 18430
rect 73990 18230 74054 18294
rect 74262 18366 74326 18430
rect 74398 18230 74462 18294
rect 74670 18230 74734 18294
rect 75078 18366 75142 18430
rect 75078 18230 75142 18294
rect 75622 18366 75686 18430
rect 77934 18366 77998 18430
rect 78206 18366 78270 18430
rect 77390 18230 77454 18294
rect 78478 18366 78542 18430
rect 78614 18366 78678 18430
rect 78614 18230 78678 18294
rect 20542 17822 20606 17886
rect 20950 17958 21014 18022
rect 21766 17958 21830 18022
rect 21630 17822 21694 17886
rect 22174 17958 22238 18022
rect 22174 17822 22238 17886
rect 3814 17686 3878 17750
rect 3814 17550 3878 17614
rect 16190 17414 16254 17478
rect 17550 17550 17614 17614
rect 16598 17414 16662 17478
rect 18230 17550 18294 17614
rect 18774 17550 18838 17614
rect 20542 17550 20606 17614
rect 20678 17414 20742 17478
rect 21630 17550 21694 17614
rect 22174 17550 22238 17614
rect 73990 17958 74054 18022
rect 73854 17822 73918 17886
rect 74398 17958 74462 18022
rect 74262 17822 74326 17886
rect 74670 17958 74734 18022
rect 75078 17958 75142 18022
rect 74806 17822 74870 17886
rect 74942 17822 75006 17886
rect 79430 18094 79494 18158
rect 75622 17822 75686 17886
rect 22038 17414 22102 17478
rect 22854 17414 22918 17478
rect 1230 17278 1294 17342
rect 73854 17550 73918 17614
rect 74262 17550 74326 17614
rect 74806 17550 74870 17614
rect 74942 17550 75006 17614
rect 75622 17550 75686 17614
rect 77390 17550 77454 17614
rect 78614 17550 78678 17614
rect 79430 17550 79494 17614
rect 79702 17414 79766 17478
rect 82422 17414 82486 17478
rect 82422 17142 82486 17206
rect 22038 17006 22102 17070
rect 22038 16870 22102 16934
rect 22854 17006 22918 17070
rect 28566 17006 28630 17070
rect 82422 17006 82486 17070
rect 94662 17006 94726 17070
rect 26526 16870 26590 16934
rect 26526 16598 26590 16662
rect 30470 16598 30534 16662
rect 28294 16462 28358 16526
rect 29246 16462 29310 16526
rect 31558 16462 31622 16526
rect 32102 16462 32166 16526
rect 32782 16462 32846 16526
rect 33326 16462 33390 16526
rect 34142 16462 34206 16526
rect 34550 16462 34614 16526
rect 35774 16462 35838 16526
rect 36590 16462 36654 16526
rect 38358 16462 38422 16526
rect 39038 16462 39102 16526
rect 39582 16462 39646 16526
rect 40262 16462 40326 16526
rect 40806 16462 40870 16526
rect 42030 16462 42094 16526
rect 42846 16462 42910 16526
rect 44614 16462 44678 16526
rect 45294 16462 45358 16526
rect 45838 16462 45902 16526
rect 46518 16462 46582 16526
rect 47062 16462 47126 16526
rect 47742 16462 47806 16526
rect 48286 16462 48350 16526
rect 49374 16462 49438 16526
rect 50326 16462 50390 16526
rect 50734 16462 50798 16526
rect 51550 16462 51614 16526
rect 51958 16462 52022 16526
rect 53318 16462 53382 16526
rect 53998 16462 54062 16526
rect 54542 16462 54606 16526
rect 55358 16462 55422 16526
rect 55766 16462 55830 16526
rect 56446 16462 56510 16526
rect 56990 16462 57054 16526
rect 57806 16462 57870 16526
rect 57942 16462 58006 16526
rect 59030 16462 59094 16526
rect 59574 16462 59638 16526
rect 60254 16462 60318 16526
rect 60798 16462 60862 16526
rect 64198 16598 64262 16662
rect 62022 16462 62086 16526
rect 63246 16462 63310 16526
rect 65286 16462 65350 16526
rect 65694 16462 65758 16526
rect 66510 16462 66574 16526
rect 67054 16462 67118 16526
rect 67734 16462 67798 16526
rect 68278 16462 68342 16526
rect 2318 16190 2382 16254
rect 16190 16326 16254 16390
rect 14286 16190 14350 16254
rect 28294 16054 28358 16118
rect 29246 16054 29310 16118
rect 30470 16054 30534 16118
rect 31558 16054 31622 16118
rect 32102 16054 32166 16118
rect 32782 16054 32846 16118
rect 33326 16054 33390 16118
rect 34142 16054 34206 16118
rect 34550 16054 34614 16118
rect 35774 16054 35838 16118
rect 36590 16054 36654 16118
rect 38358 16054 38422 16118
rect 39038 16054 39102 16118
rect 39582 16054 39646 16118
rect 40262 16054 40326 16118
rect 40806 16054 40870 16118
rect 42030 16054 42094 16118
rect 42846 16054 42910 16118
rect 44614 16054 44678 16118
rect 45294 16054 45358 16118
rect 45838 16054 45902 16118
rect 46518 16054 46582 16118
rect 47062 16054 47126 16118
rect 47742 16054 47806 16118
rect 48286 16054 48350 16118
rect 49374 16054 49438 16118
rect 50326 16054 50390 16118
rect 50734 16054 50798 16118
rect 51550 16054 51614 16118
rect 51958 16054 52022 16118
rect 53318 16054 53382 16118
rect 53998 16054 54062 16118
rect 54542 16054 54606 16118
rect 55358 16054 55422 16118
rect 55766 16054 55830 16118
rect 56446 16054 56510 16118
rect 56990 16054 57054 16118
rect 57806 16054 57870 16118
rect 57942 16054 58006 16118
rect 58078 15918 58142 15982
rect 59030 16054 59094 16118
rect 59574 16054 59638 16118
rect 60254 16054 60318 16118
rect 60798 16054 60862 16118
rect 62022 16054 62086 16118
rect 63246 16054 63310 16118
rect 64198 16054 64262 16118
rect 65286 16054 65350 16118
rect 65694 16054 65758 16118
rect 66510 16054 66574 16118
rect 67054 16054 67118 16118
rect 67734 16054 67798 16118
rect 68278 16054 68342 16118
rect 79702 15782 79766 15846
rect 82558 15646 82622 15710
rect 2318 15510 2382 15574
rect 1230 15374 1294 15438
rect 94662 15374 94726 15438
rect 2561 15198 2625 15262
rect 3814 14694 3878 14758
rect 3950 14694 4014 14758
rect 16598 14830 16662 14894
rect 14150 14694 14214 14758
rect 20678 14694 20742 14758
rect 21086 14558 21150 14622
rect 28566 14558 28630 14622
rect 31150 14286 31214 14350
rect 82422 14422 82486 14486
rect 82286 14150 82350 14214
rect 94662 13878 94726 13942
rect 1230 13742 1294 13806
rect 3134 13742 3198 13806
rect 3134 13470 3198 13534
rect 14286 13470 14350 13534
rect 14014 13334 14078 13398
rect 22038 13198 22102 13262
rect 82558 12926 82622 12990
rect 82422 12790 82486 12854
rect 31150 12654 31214 12718
rect 64606 12654 64670 12718
rect 94662 12246 94726 12310
rect 1230 11974 1294 12038
rect 3814 11974 3878 12038
rect 550 11838 614 11902
rect 14150 11974 14214 12038
rect 14286 11838 14350 11902
rect 21086 11838 21150 11902
rect 28430 11838 28494 11902
rect 29790 11838 29854 11902
rect 31014 11838 31078 11902
rect 32102 11838 32166 11902
rect 33462 11838 33526 11902
rect 34686 11838 34750 11902
rect 36046 11838 36110 11902
rect 37134 11838 37198 11902
rect 38494 11838 38558 11902
rect 39718 11838 39782 11902
rect 40806 11838 40870 11902
rect 42166 11838 42230 11902
rect 43390 11838 43454 11902
rect 44750 11838 44814 11902
rect 45838 11838 45902 11902
rect 47198 11838 47262 11902
rect 48422 11838 48486 11902
rect 49782 11838 49846 11902
rect 51006 11838 51070 11902
rect 52094 11838 52158 11902
rect 53454 11838 53518 11902
rect 54542 11838 54606 11902
rect 56038 11838 56102 11902
rect 58078 11974 58142 12038
rect 57126 11838 57190 11902
rect 58486 11838 58550 11902
rect 59710 11838 59774 11902
rect 60798 11838 60862 11902
rect 62158 11838 62222 11902
rect 63382 11838 63446 11902
rect 64742 11838 64806 11902
rect 65830 11838 65894 11902
rect 83102 11974 83166 12038
rect 67190 11838 67254 11902
rect 82286 11566 82350 11630
rect 82558 11430 82622 11494
rect 28430 11158 28494 11222
rect 29790 11158 29854 11222
rect 31014 11158 31078 11222
rect 32102 11158 32166 11222
rect 33462 11158 33526 11222
rect 34686 11158 34750 11222
rect 36046 11158 36110 11222
rect 37134 11158 37198 11222
rect 38494 11158 38558 11222
rect 39718 11158 39782 11222
rect 40806 11158 40870 11222
rect 42166 11158 42230 11222
rect 43390 11158 43454 11222
rect 44750 11158 44814 11222
rect 45838 11158 45902 11222
rect 47198 11158 47262 11222
rect 48422 11158 48486 11222
rect 38494 11022 38558 11086
rect 49782 11158 49846 11222
rect 51006 11158 51070 11222
rect 52094 11158 52158 11222
rect 53454 11158 53518 11222
rect 54542 11158 54606 11222
rect 56038 11158 56102 11222
rect 57126 11158 57190 11222
rect 58486 11158 58550 11222
rect 59710 11158 59774 11222
rect 60798 11158 60862 11222
rect 62158 11158 62222 11222
rect 63382 11158 63446 11222
rect 64742 11158 64806 11222
rect 65830 11158 65894 11222
rect 67190 11158 67254 11222
rect 14014 10614 14078 10678
rect 27886 10614 27950 10678
rect 28566 10614 28630 10678
rect 29246 10614 29310 10678
rect 29790 10614 29854 10678
rect 30334 10614 30398 10678
rect 30878 10614 30942 10678
rect 31966 10614 32030 10678
rect 32238 10614 32302 10678
rect 33190 10614 33254 10678
rect 33462 10614 33526 10678
rect 34414 10614 34478 10678
rect 34822 10614 34886 10678
rect 35638 10614 35702 10678
rect 36046 10614 36110 10678
rect 36862 10614 36926 10678
rect 37134 10614 37198 10678
rect 37814 10614 37878 10678
rect 38630 10614 38694 10678
rect 39310 10614 39374 10678
rect 39718 10614 39782 10678
rect 40670 10614 40734 10678
rect 40942 10614 41006 10678
rect 41758 10614 41822 10678
rect 41894 10614 41958 10678
rect 42302 10614 42366 10678
rect 43118 10614 43182 10678
rect 43526 10614 43590 10678
rect 44342 10614 44406 10678
rect 44750 10614 44814 10678
rect 45294 10614 45358 10678
rect 45566 10614 45630 10678
rect 45974 10614 46038 10678
rect 46654 10614 46718 10678
rect 47198 10614 47262 10678
rect 47742 10614 47806 10678
rect 47878 10614 47942 10678
rect 48422 10614 48486 10678
rect 48966 10614 49030 10678
rect 49102 10614 49166 10678
rect 49646 10614 49710 10678
rect 49782 10614 49846 10678
rect 50598 10614 50662 10678
rect 51006 10614 51070 10678
rect 51414 10614 51478 10678
rect 52230 10614 52294 10678
rect 53182 10614 53246 10678
rect 53454 10614 53518 10678
rect 54406 10614 54470 10678
rect 54678 10614 54742 10678
rect 55630 10614 55694 10678
rect 55902 10614 55966 10678
rect 56854 10614 56918 10678
rect 57262 10614 57326 10678
rect 57806 10614 57870 10678
rect 58486 10614 58550 10678
rect 59166 10614 59230 10678
rect 59302 10614 59366 10678
rect 59710 10614 59774 10678
rect 60526 10614 60590 10678
rect 60934 10614 60998 10678
rect 61750 10614 61814 10678
rect 61886 10614 61950 10678
rect 62158 10614 62222 10678
rect 62974 10614 63038 10678
rect 63110 10614 63174 10678
rect 63518 10614 63582 10678
rect 64742 10750 64806 10814
rect 64334 10614 64398 10678
rect 64742 10614 64806 10678
rect 65422 10614 65486 10678
rect 65558 10614 65622 10678
rect 65966 10614 66030 10678
rect 82694 10886 82758 10950
rect 66782 10614 66846 10678
rect 67054 10614 67118 10678
rect 1230 10478 1294 10542
rect 14014 10478 14078 10542
rect 94662 10478 94726 10542
rect 48966 10342 49030 10406
rect 49646 10342 49710 10406
rect 28566 10070 28630 10134
rect 29790 10070 29854 10134
rect 30878 10070 30942 10134
rect 28430 9798 28494 9862
rect 29790 9798 29854 9862
rect 30878 9798 30942 9862
rect 32238 10070 32302 10134
rect 33462 10070 33526 10134
rect 34822 10070 34886 10134
rect 36046 10070 36110 10134
rect 37134 10070 37198 10134
rect 38630 10070 38694 10134
rect 39718 10070 39782 10134
rect 32374 9798 32438 9862
rect 33598 9798 33662 9862
rect 34822 9798 34886 9862
rect 36046 9798 36110 9862
rect 37270 9798 37334 9862
rect 38222 9798 38286 9862
rect 39718 9798 39782 9862
rect 40942 10070 41006 10134
rect 41758 10070 41822 10134
rect 42302 10070 42366 10134
rect 43526 10070 43590 10134
rect 44750 10070 44814 10134
rect 45294 10070 45358 10134
rect 45974 10070 46038 10134
rect 47198 10070 47262 10134
rect 47742 10070 47806 10134
rect 48422 10070 48486 10134
rect 41078 9798 41142 9862
rect 42302 9798 42366 9862
rect 43526 9798 43590 9862
rect 44750 9798 44814 9862
rect 45974 9798 46038 9862
rect 47198 9798 47262 9862
rect 48422 9798 48486 9862
rect 49782 10070 49846 10134
rect 51006 10070 51070 10134
rect 52230 10070 52294 10134
rect 53454 10070 53518 10134
rect 54678 10070 54742 10134
rect 49782 9798 49846 9862
rect 50870 9798 50934 9862
rect 52094 9798 52158 9862
rect 53590 9798 53654 9862
rect 54678 9798 54742 9862
rect 55902 10070 55966 10134
rect 57262 10070 57326 10134
rect 58486 10070 58550 10134
rect 59166 10070 59230 10134
rect 59710 10070 59774 10134
rect 60934 10070 60998 10134
rect 61750 10070 61814 10134
rect 62158 10070 62222 10134
rect 62974 10070 63038 10134
rect 63518 10070 63582 10134
rect 56038 9798 56102 9862
rect 56718 9798 56782 9862
rect 57126 9798 57190 9862
rect 58486 9798 58550 9862
rect 59710 9798 59774 9862
rect 64742 10070 64806 10134
rect 65422 10070 65486 10134
rect 65966 10070 66030 10134
rect 67054 10070 67118 10134
rect 60934 9798 60998 9862
rect 62294 9798 62358 9862
rect 63518 9798 63582 9862
rect 64742 9798 64806 9862
rect 65830 9798 65894 9862
rect 82422 10070 82486 10134
rect 82422 9934 82486 9998
rect 67190 9798 67254 9862
rect 28294 9390 28358 9454
rect 29654 9390 29718 9454
rect 30742 9390 30806 9454
rect 32238 9390 32302 9454
rect 33462 9390 33526 9454
rect 34686 9390 34750 9454
rect 35910 9390 35974 9454
rect 37134 9390 37198 9454
rect 38494 9526 38558 9590
rect 38358 9390 38422 9454
rect 39582 9390 39646 9454
rect 40942 9390 41006 9454
rect 42166 9390 42230 9454
rect 43390 9390 43454 9454
rect 44614 9390 44678 9454
rect 45838 9390 45902 9454
rect 47062 9390 47126 9454
rect 48286 9390 48350 9454
rect 49646 9390 49710 9454
rect 50734 9390 50798 9454
rect 51958 9390 52022 9454
rect 53454 9390 53518 9454
rect 54542 9390 54606 9454
rect 55902 9390 55966 9454
rect 56990 9390 57054 9454
rect 58350 9390 58414 9454
rect 59574 9390 59638 9454
rect 60798 9390 60862 9454
rect 62158 9390 62222 9454
rect 63382 9390 63446 9454
rect 64606 9390 64670 9454
rect 65694 9390 65758 9454
rect 67054 9390 67118 9454
rect 14286 9254 14350 9318
rect 14150 9118 14214 9182
rect 28430 9254 28494 9318
rect 29790 9254 29854 9318
rect 30878 9254 30942 9318
rect 32374 9254 32438 9318
rect 33598 9254 33662 9318
rect 34822 9254 34886 9318
rect 1230 8846 1294 8910
rect 27750 8846 27814 8910
rect 36046 9254 36110 9318
rect 37270 9254 37334 9318
rect 38222 9254 38286 9318
rect 39718 9254 39782 9318
rect 41078 9254 41142 9318
rect 42302 9254 42366 9318
rect 44750 9254 44814 9318
rect 45974 9254 46038 9318
rect 47198 9254 47262 9318
rect 48422 9254 48486 9318
rect 49782 9254 49846 9318
rect 50870 9254 50934 9318
rect 53590 9254 53654 9318
rect 54678 9254 54742 9318
rect 56038 9254 56102 9318
rect 56718 9254 56782 9318
rect 57126 9254 57190 9318
rect 43526 8982 43590 9046
rect 52094 8982 52158 9046
rect 58486 9254 58550 9318
rect 59710 9254 59774 9318
rect 60934 9254 60998 9318
rect 62294 9254 62358 9318
rect 63518 9254 63582 9318
rect 65830 9254 65894 9318
rect 67190 9254 67254 9318
rect 64742 8982 64806 9046
rect 82830 9118 82894 9182
rect 68006 8846 68070 8910
rect 94662 8846 94726 8910
rect 82558 8710 82622 8774
rect 28158 8574 28222 8638
rect 28294 8574 28358 8638
rect 29654 8574 29718 8638
rect 30742 8574 30806 8638
rect 32238 8574 32302 8638
rect 33462 8574 33526 8638
rect 34686 8574 34750 8638
rect 35910 8574 35974 8638
rect 37134 8574 37198 8638
rect 38358 8574 38422 8638
rect 39582 8574 39646 8638
rect 40942 8574 41006 8638
rect 42166 8574 42230 8638
rect 43390 8574 43454 8638
rect 44614 8574 44678 8638
rect 45838 8574 45902 8638
rect 47062 8574 47126 8638
rect 48286 8574 48350 8638
rect 49646 8574 49710 8638
rect 50734 8574 50798 8638
rect 51958 8574 52022 8638
rect 53454 8574 53518 8638
rect 54542 8574 54606 8638
rect 55902 8574 55966 8638
rect 56990 8574 57054 8638
rect 58350 8574 58414 8638
rect 59574 8574 59638 8638
rect 60798 8574 60862 8638
rect 62158 8574 62222 8638
rect 63382 8574 63446 8638
rect 64606 8574 64670 8638
rect 65694 8574 65758 8638
rect 67054 8574 67118 8638
rect 67870 8574 67934 8638
rect 28158 8166 28222 8230
rect 67870 8166 67934 8230
rect 82966 8074 82982 8094
rect 82982 8074 83030 8094
rect 82966 8030 83030 8074
rect 14014 7758 14078 7822
rect 550 7622 614 7686
rect 14286 7622 14350 7686
rect 82422 7350 82486 7414
rect 27750 7078 27814 7142
rect 68006 7078 68070 7142
rect 1230 6942 1294 7006
rect 2590 6942 2654 7006
rect 94662 6942 94726 7006
rect 2590 6398 2654 6462
rect 14150 6398 14214 6462
rect 15918 6262 15982 6326
rect 1230 5310 1294 5374
rect 5854 5446 5918 5510
rect 94662 5310 94726 5374
rect 550 5038 614 5102
rect 14286 5038 14350 5102
rect 16054 4766 16118 4830
rect 1230 3678 1294 3742
rect 15918 3814 15982 3878
rect 17278 3678 17342 3742
rect 94662 3678 94726 3742
rect 15510 2862 15574 2926
rect 16734 2924 16764 2926
rect 16764 2924 16798 2926
rect 16734 2862 16798 2924
rect 17822 2862 17886 2926
rect 19182 2862 19246 2926
rect 20134 2862 20198 2926
rect 21358 2862 21422 2926
rect 22582 2924 22604 2926
rect 22604 2924 22646 2926
rect 22582 2862 22646 2924
rect 23670 2862 23734 2926
rect 25030 2862 25094 2926
rect 26118 2924 26164 2926
rect 26164 2924 26182 2926
rect 26118 2862 26182 2924
rect 27206 2862 27270 2926
rect 28294 2862 28358 2926
rect 29654 2924 29668 2926
rect 29668 2924 29718 2926
rect 29654 2862 29718 2924
rect 30742 2924 30780 2926
rect 30780 2924 30806 2926
rect 30742 2862 30806 2924
rect 31830 2862 31894 2926
rect 33054 2924 33116 2926
rect 33116 2924 33118 2926
rect 33054 2862 33118 2924
rect 34142 2862 34206 2926
rect 35502 2924 35508 2926
rect 35508 2924 35566 2926
rect 35502 2862 35566 2924
rect 36590 2924 36620 2926
rect 36620 2924 36654 2926
rect 36590 2862 36654 2924
rect 37678 2862 37742 2926
rect 38902 2924 38956 2926
rect 38956 2924 38966 2926
rect 38902 2862 38966 2924
rect 40262 2862 40326 2926
rect 41350 2862 41414 2926
rect 42438 2924 42460 2926
rect 42460 2924 42502 2926
rect 42438 2862 42502 2924
rect 43526 2862 43590 2926
rect 44886 2862 44950 2926
rect 45974 2924 46020 2926
rect 46020 2924 46038 2926
rect 45974 2862 46038 2924
rect 47062 2862 47126 2926
rect 48286 2924 48300 2926
rect 48300 2924 48350 2926
rect 48286 2862 48350 2924
rect 49374 2862 49438 2926
rect 50734 2862 50798 2926
rect 51822 2924 51860 2926
rect 51860 2924 51886 2926
rect 51822 2862 51886 2924
rect 52910 2924 52972 2926
rect 52972 2924 52974 2926
rect 52910 2862 52974 2924
rect 53998 2862 54062 2926
rect 55222 2862 55286 2926
rect 56582 2862 56646 2926
rect 57670 2924 57700 2926
rect 57700 2924 57734 2926
rect 57670 2862 57734 2924
rect 16054 2454 16118 2518
rect 26662 2318 26726 2382
rect 94662 1910 94726 1974
rect 2182 1688 2210 1702
rect 2210 1688 2246 1702
rect 2182 1638 2246 1688
rect 3950 1638 4014 1702
rect 5446 1638 5510 1702
rect 7214 1688 7250 1702
rect 7250 1688 7278 1702
rect 7214 1638 7278 1688
rect 8982 1638 9046 1702
rect 10478 1638 10542 1702
rect 12246 1688 12290 1702
rect 12290 1688 12310 1702
rect 12246 1638 12310 1688
rect 14014 1638 14078 1702
rect 17278 1774 17342 1838
rect 15782 1638 15846 1702
rect 17414 1638 17478 1702
rect 18910 1688 18954 1702
rect 18954 1688 18974 1702
rect 18910 1638 18974 1688
rect 20678 1688 20690 1702
rect 20690 1688 20742 1702
rect 20678 1638 20742 1688
rect 22446 1638 22510 1702
rect 23942 1688 23994 1702
rect 23994 1688 24006 1702
rect 23942 1638 24006 1688
rect 25710 1688 25730 1702
rect 25730 1688 25774 1702
rect 25710 1638 25774 1688
rect 27478 1638 27542 1702
rect 28974 1688 29034 1702
rect 29034 1688 29038 1702
rect 28974 1638 29038 1688
rect 30606 1638 30670 1702
rect 32374 1688 32394 1702
rect 32394 1688 32438 1702
rect 32374 1638 32438 1688
rect 34006 1638 34070 1702
rect 35774 1688 35810 1702
rect 35810 1688 35838 1702
rect 35774 1638 35838 1688
rect 37406 1688 37434 1702
rect 37434 1688 37470 1702
rect 37406 1638 37470 1688
rect 39174 1638 39238 1702
rect 40534 1638 40598 1702
rect 42302 1638 42366 1702
rect 44206 1688 44210 1702
rect 44210 1688 44270 1702
rect 44206 1638 44270 1688
rect 45838 1688 45890 1702
rect 45890 1688 45902 1702
rect 45838 1638 45902 1688
rect 47470 1688 47514 1702
rect 47514 1688 47534 1702
rect 47470 1638 47534 1688
rect 48966 1638 49030 1702
rect 51006 1638 51070 1702
rect 52638 1638 52702 1702
rect 54270 1688 54290 1702
rect 54290 1688 54334 1702
rect 54270 1638 54334 1688
rect 55902 1688 55914 1702
rect 55914 1688 55966 1702
rect 55902 1638 55966 1688
rect 57534 1688 57594 1702
rect 57594 1688 57598 1702
rect 57534 1638 57598 1688
rect 59166 1638 59230 1702
rect 60934 1688 60954 1702
rect 60954 1688 60998 1702
rect 60934 1638 60998 1688
rect 62702 1638 62766 1702
rect 64062 1638 64126 1702
rect 65966 1688 65994 1702
rect 65994 1688 66030 1702
rect 65966 1638 66030 1688
rect 67734 1638 67798 1702
rect 69230 1638 69294 1702
rect 70998 1688 71034 1702
rect 71034 1688 71062 1702
rect 70998 1638 71062 1688
rect 72630 1638 72694 1702
rect 74262 1638 74326 1702
rect 76166 1638 76230 1702
rect 77662 1638 77726 1702
rect 79430 1688 79434 1702
rect 79434 1688 79490 1702
rect 79490 1688 79494 1702
rect 79430 1638 79494 1688
rect 81198 1638 81262 1702
rect 82558 1638 82622 1702
rect 84462 1688 84474 1702
rect 84474 1688 84526 1702
rect 84462 1638 84526 1688
rect 86230 1638 86294 1702
rect 87726 1638 87790 1702
rect 89494 1688 89514 1702
rect 89514 1688 89558 1702
rect 89494 1638 89558 1688
rect 91126 1638 91190 1702
rect 92758 1638 92822 1702
rect 958 1230 1022 1294
rect 1094 1230 1158 1294
rect 1230 1230 1294 1294
rect 2182 1230 2246 1294
rect 3950 1230 4014 1294
rect 5446 1230 5510 1294
rect 7214 1230 7278 1294
rect 8982 1230 9046 1294
rect 10478 1230 10542 1294
rect 12246 1230 12310 1294
rect 14014 1230 14078 1294
rect 15782 1230 15846 1294
rect 17414 1230 17478 1294
rect 18910 1230 18974 1294
rect 20678 1230 20742 1294
rect 22446 1230 22510 1294
rect 23942 1230 24006 1294
rect 25710 1230 25774 1294
rect 27478 1230 27542 1294
rect 28974 1230 29038 1294
rect 30606 1230 30670 1294
rect 32374 1230 32438 1294
rect 34006 1230 34070 1294
rect 35774 1230 35838 1294
rect 37406 1230 37470 1294
rect 39174 1230 39238 1294
rect 40534 1230 40598 1294
rect 42302 1230 42366 1294
rect 44206 1230 44270 1294
rect 45838 1230 45902 1294
rect 47470 1230 47534 1294
rect 48966 1230 49030 1294
rect 51006 1230 51070 1294
rect 52638 1230 52702 1294
rect 54270 1230 54334 1294
rect 55902 1230 55966 1294
rect 57534 1230 57598 1294
rect 59166 1230 59230 1294
rect 60934 1230 60998 1294
rect 62702 1230 62766 1294
rect 64062 1230 64126 1294
rect 65966 1230 66030 1294
rect 67734 1230 67798 1294
rect 69230 1230 69294 1294
rect 70998 1230 71062 1294
rect 72630 1230 72694 1294
rect 74262 1230 74326 1294
rect 76166 1230 76230 1294
rect 77662 1230 77726 1294
rect 79430 1230 79494 1294
rect 81198 1230 81262 1294
rect 82558 1230 82622 1294
rect 84462 1230 84526 1294
rect 86230 1230 86294 1294
rect 87726 1230 87790 1294
rect 89494 1230 89558 1294
rect 91126 1230 91190 1294
rect 92758 1230 92822 1294
rect 94662 1230 94726 1294
rect 94798 1230 94862 1294
rect 94934 1230 94998 1294
rect 958 1094 1022 1158
rect 1094 1094 1158 1158
rect 1230 1094 1294 1158
rect 94662 1094 94726 1158
rect 94798 1094 94862 1158
rect 94934 1094 94998 1158
rect 958 958 1022 1022
rect 1094 958 1158 1022
rect 1230 958 1294 1022
rect 94662 958 94726 1022
rect 94798 958 94862 1022
rect 94934 958 94998 1022
rect 278 550 342 614
rect 414 550 478 614
rect 550 550 614 614
rect 26662 550 26726 614
rect 95342 550 95406 614
rect 95478 550 95542 614
rect 95614 550 95678 614
rect 278 414 342 478
rect 414 414 478 478
rect 550 414 614 478
rect 95342 414 95406 478
rect 95478 414 95542 478
rect 95614 414 95678 478
rect 278 278 342 342
rect 414 278 478 342
rect 550 278 614 342
rect 95342 278 95406 342
rect 95478 278 95542 342
rect 95614 278 95678 342
<< metal4 >>
rect 272 79222 620 79228
rect 272 79158 278 79222
rect 342 79158 414 79222
rect 478 79158 550 79222
rect 614 79158 620 79222
rect 272 79086 620 79158
rect 272 79022 278 79086
rect 342 79022 414 79086
rect 478 79022 550 79086
rect 614 79022 620 79086
rect 272 78950 620 79022
rect 272 78886 278 78950
rect 342 78886 414 78950
rect 478 78886 550 78950
rect 614 78886 620 78950
rect 272 23462 620 78886
rect 272 23398 550 23462
rect 614 23398 620 23462
rect 272 11902 620 23398
rect 272 11838 550 11902
rect 614 11838 620 11902
rect 272 7686 620 11838
rect 272 7622 550 7686
rect 614 7622 620 7686
rect 272 5102 620 7622
rect 272 5038 550 5102
rect 614 5038 620 5102
rect 272 614 620 5038
rect 952 78542 1300 78548
rect 952 78478 958 78542
rect 1022 78478 1094 78542
rect 1158 78478 1230 78542
rect 1294 78478 1300 78542
rect 952 78406 1300 78478
rect 952 78342 958 78406
rect 1022 78342 1094 78406
rect 1158 78342 1230 78406
rect 1294 78342 1300 78406
rect 952 78270 1300 78342
rect 952 78206 958 78270
rect 1022 78206 1094 78270
rect 1158 78206 1230 78270
rect 1294 78206 1300 78270
rect 952 75958 1300 78206
rect 2176 78270 2252 78276
rect 2176 78206 2182 78270
rect 2246 78206 2252 78270
rect 2176 77862 2252 78206
rect 2176 77830 2182 77862
rect 2181 77798 2182 77830
rect 2246 77830 2252 77862
rect 3944 78270 4020 78276
rect 3944 78206 3950 78270
rect 4014 78206 4020 78270
rect 3944 77862 4020 78206
rect 3944 77830 3950 77862
rect 2246 77798 2247 77830
rect 2181 77797 2247 77798
rect 3949 77798 3950 77830
rect 4014 77830 4020 77862
rect 5440 78270 5516 78276
rect 5440 78206 5446 78270
rect 5510 78206 5516 78270
rect 5440 77862 5516 78206
rect 5440 77830 5446 77862
rect 4014 77798 4015 77830
rect 3949 77797 4015 77798
rect 5445 77798 5446 77830
rect 5510 77830 5516 77862
rect 7208 78270 7284 78276
rect 7208 78206 7214 78270
rect 7278 78206 7284 78270
rect 7208 77862 7284 78206
rect 7208 77830 7214 77862
rect 5510 77798 5511 77830
rect 5445 77797 5511 77798
rect 7213 77798 7214 77830
rect 7278 77830 7284 77862
rect 8976 78270 9052 78276
rect 8976 78206 8982 78270
rect 9046 78206 9052 78270
rect 8976 77862 9052 78206
rect 8976 77830 8982 77862
rect 7278 77798 7279 77830
rect 7213 77797 7279 77798
rect 8981 77798 8982 77830
rect 9046 77830 9052 77862
rect 10472 78270 10548 78276
rect 10472 78206 10478 78270
rect 10542 78206 10548 78270
rect 10472 77862 10548 78206
rect 10472 77830 10478 77862
rect 9046 77798 9047 77830
rect 8981 77797 9047 77798
rect 10477 77798 10478 77830
rect 10542 77830 10548 77862
rect 12240 78270 12316 78276
rect 12240 78206 12246 78270
rect 12310 78206 12316 78270
rect 12240 77862 12316 78206
rect 12240 77830 12246 77862
rect 10542 77798 10543 77830
rect 10477 77797 10543 77798
rect 12245 77798 12246 77830
rect 12310 77830 12316 77862
rect 14008 78270 14084 78276
rect 14008 78206 14014 78270
rect 14078 78206 14084 78270
rect 14008 77862 14084 78206
rect 14008 77830 14014 77862
rect 12310 77798 12311 77830
rect 12245 77797 12311 77798
rect 14013 77798 14014 77830
rect 14078 77830 14084 77862
rect 15640 78270 15716 78276
rect 15640 78206 15646 78270
rect 15710 78206 15716 78270
rect 15640 77862 15716 78206
rect 15640 77830 15646 77862
rect 14078 77798 14079 77830
rect 14013 77797 14079 77798
rect 15645 77798 15646 77830
rect 15710 77830 15716 77862
rect 17408 78270 17484 78276
rect 17408 78206 17414 78270
rect 17478 78206 17484 78270
rect 17408 77862 17484 78206
rect 17408 77830 17414 77862
rect 15710 77798 15711 77830
rect 15645 77797 15711 77798
rect 17413 77798 17414 77830
rect 17478 77830 17484 77862
rect 18904 78270 18980 78276
rect 18904 78206 18910 78270
rect 18974 78206 18980 78270
rect 18904 77862 18980 78206
rect 18904 77830 18910 77862
rect 17478 77798 17479 77830
rect 17413 77797 17479 77798
rect 18909 77798 18910 77830
rect 18974 77830 18980 77862
rect 20672 78270 20748 78276
rect 20672 78206 20678 78270
rect 20742 78206 20748 78270
rect 20672 77862 20748 78206
rect 20672 77830 20678 77862
rect 18974 77798 18975 77830
rect 18909 77797 18975 77798
rect 20677 77798 20678 77830
rect 20742 77830 20748 77862
rect 22168 78270 22244 78276
rect 22168 78206 22174 78270
rect 22238 78206 22244 78270
rect 22168 77862 22244 78206
rect 22168 77830 22174 77862
rect 20742 77798 20743 77830
rect 20677 77797 20743 77798
rect 22173 77798 22174 77830
rect 22238 77830 22244 77862
rect 23936 78270 24012 78276
rect 23936 78206 23942 78270
rect 24006 78206 24012 78270
rect 23936 77862 24012 78206
rect 23936 77830 23942 77862
rect 22238 77798 22239 77830
rect 22173 77797 22239 77798
rect 23941 77798 23942 77830
rect 24006 77830 24012 77862
rect 25704 78270 25780 78276
rect 25704 78206 25710 78270
rect 25774 78206 25780 78270
rect 25704 77862 25780 78206
rect 25704 77830 25710 77862
rect 24006 77798 24007 77830
rect 23941 77797 24007 77798
rect 25709 77798 25710 77830
rect 25774 77830 25780 77862
rect 27472 78270 27548 78276
rect 27472 78206 27478 78270
rect 27542 78206 27548 78270
rect 27472 77862 27548 78206
rect 27472 77830 27478 77862
rect 25774 77798 25775 77830
rect 25709 77797 25775 77798
rect 27477 77798 27478 77830
rect 27542 77830 27548 77862
rect 27542 77798 27543 77830
rect 27477 77797 27543 77798
rect 952 75894 1230 75958
rect 1294 75894 1300 75958
rect 952 74462 1300 75894
rect 952 74398 1230 74462
rect 1294 74398 1300 74462
rect 952 72558 1300 74398
rect 28152 74190 28228 79500
rect 28968 78270 29044 78276
rect 28968 78206 28974 78270
rect 29038 78206 29044 78270
rect 28968 77862 29044 78206
rect 28968 77830 28974 77862
rect 28973 77798 28974 77830
rect 29038 77830 29044 77862
rect 29038 77798 29039 77830
rect 28973 77797 29039 77798
rect 28152 74158 28158 74190
rect 28157 74126 28158 74158
rect 28222 74158 28228 74190
rect 29512 74190 29588 79500
rect 29789 77726 29855 77727
rect 29789 77694 29790 77726
rect 29512 74158 29518 74190
rect 28222 74126 28223 74158
rect 28157 74125 28223 74126
rect 29517 74126 29518 74158
rect 29582 74158 29588 74190
rect 29784 77662 29790 77694
rect 29854 77694 29855 77726
rect 29854 77662 29860 77694
rect 29582 74126 29583 74158
rect 29517 74125 29583 74126
rect 29784 73918 29860 77662
rect 30600 74190 30676 79500
rect 30872 78270 30948 78276
rect 30872 78206 30878 78270
rect 30942 78206 30948 78270
rect 30872 77862 30948 78206
rect 30872 77830 30878 77862
rect 30877 77798 30878 77830
rect 30942 77830 30948 77862
rect 30942 77798 30943 77830
rect 30877 77797 30943 77798
rect 30600 74158 30606 74190
rect 30605 74126 30606 74158
rect 30670 74158 30676 74190
rect 31960 74190 32036 79500
rect 32504 78270 32580 78276
rect 32504 78206 32510 78270
rect 32574 78206 32580 78270
rect 32504 77862 32580 78206
rect 32504 77830 32510 77862
rect 32509 77798 32510 77830
rect 32574 77830 32580 77862
rect 32574 77798 32575 77830
rect 32509 77797 32575 77798
rect 31960 74158 31966 74190
rect 30670 74126 30671 74158
rect 30605 74125 30671 74126
rect 31965 74126 31966 74158
rect 32030 74158 32036 74190
rect 33184 74190 33260 79500
rect 34136 78270 34212 78276
rect 34136 78206 34142 78270
rect 34206 78206 34212 78270
rect 34136 77862 34212 78206
rect 34136 77830 34142 77862
rect 34141 77798 34142 77830
rect 34206 77830 34212 77862
rect 34206 77798 34207 77830
rect 34141 77797 34207 77798
rect 33184 74158 33190 74190
rect 32030 74126 32031 74158
rect 31965 74125 32031 74126
rect 33189 74126 33190 74158
rect 33254 74158 33260 74190
rect 34544 74190 34620 79500
rect 35496 78270 35572 78276
rect 35496 78206 35502 78270
rect 35566 78206 35572 78270
rect 35496 77862 35572 78206
rect 35496 77830 35502 77862
rect 35501 77798 35502 77830
rect 35566 77830 35572 77862
rect 35566 77798 35567 77830
rect 35501 77797 35567 77798
rect 34544 74158 34550 74190
rect 33254 74126 33255 74158
rect 33189 74125 33255 74126
rect 34549 74126 34550 74158
rect 34614 74158 34620 74190
rect 35768 74190 35844 79500
rect 35768 74158 35774 74190
rect 34614 74126 34615 74158
rect 34549 74125 34615 74126
rect 35773 74126 35774 74158
rect 35838 74158 35844 74190
rect 36856 74190 36932 79500
rect 37400 78270 37476 78276
rect 37400 78206 37406 78270
rect 37470 78206 37476 78270
rect 37400 77862 37476 78206
rect 37400 77830 37406 77862
rect 37405 77798 37406 77830
rect 37470 77830 37476 77862
rect 37470 77798 37471 77830
rect 37405 77797 37471 77798
rect 36856 74158 36862 74190
rect 35838 74126 35839 74158
rect 35773 74125 35839 74126
rect 36861 74126 36862 74158
rect 36926 74158 36932 74190
rect 38216 74190 38292 79500
rect 39168 78270 39244 78276
rect 39168 78206 39174 78270
rect 39238 78206 39244 78270
rect 39168 77862 39244 78206
rect 39168 77830 39174 77862
rect 39173 77798 39174 77830
rect 39238 77830 39244 77862
rect 39238 77798 39239 77830
rect 39173 77797 39239 77798
rect 38216 74158 38222 74190
rect 36926 74126 36927 74158
rect 36861 74125 36927 74126
rect 38221 74126 38222 74158
rect 38286 74158 38292 74190
rect 39304 74190 39380 79500
rect 40528 78270 40604 78276
rect 40528 78206 40534 78270
rect 40598 78206 40604 78270
rect 40528 77862 40604 78206
rect 40528 77830 40534 77862
rect 40533 77798 40534 77830
rect 40598 77830 40604 77862
rect 40598 77798 40599 77830
rect 40533 77797 40599 77798
rect 39304 74158 39310 74190
rect 38286 74126 38287 74158
rect 38221 74125 38287 74126
rect 39309 74126 39310 74158
rect 39374 74158 39380 74190
rect 40664 74190 40740 79500
rect 40664 74158 40670 74190
rect 39374 74126 39375 74158
rect 39309 74125 39375 74126
rect 40669 74126 40670 74158
rect 40734 74158 40740 74190
rect 41888 74190 41964 79500
rect 42432 78270 42508 78276
rect 42432 78206 42438 78270
rect 42502 78206 42508 78270
rect 42432 77862 42508 78206
rect 42432 77830 42438 77862
rect 42437 77798 42438 77830
rect 42502 77830 42508 77862
rect 42502 77798 42503 77830
rect 42437 77797 42503 77798
rect 41888 74158 41894 74190
rect 40734 74126 40735 74158
rect 40669 74125 40735 74126
rect 41893 74126 41894 74158
rect 41958 74158 41964 74190
rect 43248 74190 43324 79500
rect 44200 78270 44276 78276
rect 44200 78206 44206 78270
rect 44270 78206 44276 78270
rect 44200 77862 44276 78206
rect 44200 77830 44206 77862
rect 44205 77798 44206 77830
rect 44270 77830 44276 77862
rect 44270 77798 44271 77830
rect 44205 77797 44271 77798
rect 43248 74158 43254 74190
rect 41958 74126 41959 74158
rect 41893 74125 41959 74126
rect 43253 74126 43254 74158
rect 43318 74158 43324 74190
rect 44336 74190 44412 79500
rect 44336 74158 44342 74190
rect 43318 74126 43319 74158
rect 43253 74125 43319 74126
rect 44341 74126 44342 74158
rect 44406 74158 44412 74190
rect 45560 74190 45636 79500
rect 45832 78270 45908 78276
rect 45832 78206 45838 78270
rect 45902 78206 45908 78270
rect 45832 77862 45908 78206
rect 45832 77830 45838 77862
rect 45837 77798 45838 77830
rect 45902 77830 45908 77862
rect 45902 77798 45903 77830
rect 45837 77797 45903 77798
rect 45560 74158 45566 74190
rect 44406 74126 44407 74158
rect 44341 74125 44407 74126
rect 45565 74126 45566 74158
rect 45630 74158 45636 74190
rect 46920 74190 46996 79500
rect 47464 78270 47540 78276
rect 47464 78206 47470 78270
rect 47534 78206 47540 78270
rect 47464 77862 47540 78206
rect 47464 77830 47470 77862
rect 47469 77798 47470 77830
rect 47534 77830 47540 77862
rect 47534 77798 47535 77830
rect 47469 77797 47535 77798
rect 46920 74158 46926 74190
rect 45630 74126 45631 74158
rect 45565 74125 45631 74126
rect 46925 74126 46926 74158
rect 46990 74158 46996 74190
rect 48144 74190 48220 79500
rect 49232 78270 49308 78276
rect 49232 78206 49238 78270
rect 49302 78206 49308 78270
rect 49232 77862 49308 78206
rect 49232 77830 49238 77862
rect 49237 77798 49238 77830
rect 49302 77830 49308 77862
rect 49302 77798 49303 77830
rect 49237 77797 49303 77798
rect 48144 74158 48150 74190
rect 46990 74126 46991 74158
rect 46925 74125 46991 74126
rect 48149 74126 48150 74158
rect 48214 74158 48220 74190
rect 49504 74190 49580 79500
rect 49504 74158 49510 74190
rect 48214 74126 48215 74158
rect 48149 74125 48215 74126
rect 49509 74126 49510 74158
rect 49574 74158 49580 74190
rect 50592 74190 50668 79500
rect 50728 78270 50804 78276
rect 50728 78206 50734 78270
rect 50798 78206 50804 78270
rect 50728 77862 50804 78206
rect 50728 77830 50734 77862
rect 50733 77798 50734 77830
rect 50798 77830 50804 77862
rect 50798 77798 50799 77830
rect 50733 77797 50799 77798
rect 50592 74158 50598 74190
rect 49574 74126 49575 74158
rect 49509 74125 49575 74126
rect 50597 74126 50598 74158
rect 50662 74158 50668 74190
rect 51952 74190 52028 79500
rect 52632 78270 52708 78276
rect 52632 78206 52638 78270
rect 52702 78206 52708 78270
rect 52632 77862 52708 78206
rect 52632 77830 52638 77862
rect 52637 77798 52638 77830
rect 52702 77830 52708 77862
rect 52702 77798 52703 77830
rect 52637 77797 52703 77798
rect 51952 74158 51958 74190
rect 50662 74126 50663 74158
rect 50597 74125 50663 74126
rect 51957 74126 51958 74158
rect 52022 74158 52028 74190
rect 53040 74190 53116 79500
rect 54128 78270 54204 78276
rect 54128 78206 54134 78270
rect 54198 78206 54204 78270
rect 54128 77862 54204 78206
rect 54128 77830 54134 77862
rect 54133 77798 54134 77830
rect 54198 77830 54204 77862
rect 54198 77798 54199 77830
rect 54133 77797 54199 77798
rect 53040 74158 53046 74190
rect 52022 74126 52023 74158
rect 51957 74125 52023 74126
rect 53045 74126 53046 74158
rect 53110 74158 53116 74190
rect 54264 74190 54340 79500
rect 54264 74158 54270 74190
rect 53110 74126 53111 74158
rect 53045 74125 53111 74126
rect 54269 74126 54270 74158
rect 54334 74158 54340 74190
rect 55624 74190 55700 79500
rect 55896 78270 55972 78276
rect 55896 78206 55902 78270
rect 55966 78206 55972 78270
rect 55896 77862 55972 78206
rect 55896 77830 55902 77862
rect 55901 77798 55902 77830
rect 55966 77830 55972 77862
rect 55966 77798 55967 77830
rect 55901 77797 55967 77798
rect 55624 74158 55630 74190
rect 54334 74126 54335 74158
rect 54269 74125 54335 74126
rect 55629 74126 55630 74158
rect 55694 74158 55700 74190
rect 56848 74190 56924 79500
rect 57664 78270 57740 78276
rect 57664 78206 57670 78270
rect 57734 78206 57740 78270
rect 57664 77862 57740 78206
rect 57664 77830 57670 77862
rect 57669 77798 57670 77830
rect 57734 77830 57740 77862
rect 57734 77798 57735 77830
rect 57669 77797 57735 77798
rect 56848 74158 56854 74190
rect 55694 74126 55695 74158
rect 55629 74125 55695 74126
rect 56853 74126 56854 74158
rect 56918 74158 56924 74190
rect 58208 74190 58284 79500
rect 59160 78270 59236 78276
rect 59160 78206 59166 78270
rect 59230 78206 59236 78270
rect 59160 77862 59236 78206
rect 59160 77830 59166 77862
rect 59165 77798 59166 77830
rect 59230 77830 59236 77862
rect 59230 77798 59231 77830
rect 59165 77797 59231 77798
rect 58208 74158 58214 74190
rect 56918 74126 56919 74158
rect 56853 74125 56919 74126
rect 58213 74126 58214 74158
rect 58278 74158 58284 74190
rect 59296 74190 59372 79500
rect 59296 74158 59302 74190
rect 58278 74126 58279 74158
rect 58213 74125 58279 74126
rect 59301 74126 59302 74158
rect 59366 74158 59372 74190
rect 60656 74190 60732 79500
rect 60928 78270 61004 78276
rect 60928 78206 60934 78270
rect 60998 78206 61004 78270
rect 60928 77862 61004 78206
rect 60928 77830 60934 77862
rect 60933 77798 60934 77830
rect 60998 77830 61004 77862
rect 60998 77798 60999 77830
rect 60933 77797 60999 77798
rect 60656 74158 60662 74190
rect 59366 74126 59367 74158
rect 59301 74125 59367 74126
rect 60661 74126 60662 74158
rect 60726 74158 60732 74190
rect 61880 74190 61956 79500
rect 62696 78270 62772 78276
rect 62696 78206 62702 78270
rect 62766 78206 62772 78270
rect 62696 77862 62772 78206
rect 62696 77830 62702 77862
rect 62701 77798 62702 77830
rect 62766 77830 62772 77862
rect 62766 77798 62767 77830
rect 62701 77797 62767 77798
rect 61880 74158 61886 74190
rect 60726 74126 60727 74158
rect 60661 74125 60727 74126
rect 61885 74126 61886 74158
rect 61950 74158 61956 74190
rect 63240 74190 63316 79500
rect 64056 78270 64132 78276
rect 64056 78206 64062 78270
rect 64126 78206 64132 78270
rect 64056 77862 64132 78206
rect 64056 77830 64062 77862
rect 64061 77798 64062 77830
rect 64126 77830 64132 77862
rect 64126 77798 64127 77830
rect 64061 77797 64127 77798
rect 63240 74158 63246 74190
rect 61950 74126 61951 74158
rect 61885 74125 61951 74126
rect 63245 74126 63246 74158
rect 63310 74158 63316 74190
rect 64328 74190 64404 79500
rect 64328 74158 64334 74190
rect 63310 74126 63311 74158
rect 63245 74125 63311 74126
rect 64333 74126 64334 74158
rect 64398 74158 64404 74190
rect 65552 74190 65628 79500
rect 65960 78270 66036 78276
rect 65960 78206 65966 78270
rect 66030 78206 66036 78270
rect 65960 77862 66036 78206
rect 65960 77830 65966 77862
rect 65965 77798 65966 77830
rect 66030 77830 66036 77862
rect 66030 77798 66031 77830
rect 65965 77797 66031 77798
rect 65552 74158 65558 74190
rect 64398 74126 64399 74158
rect 64333 74125 64399 74126
rect 65557 74126 65558 74158
rect 65622 74158 65628 74190
rect 66912 74190 66988 79500
rect 78880 78950 78956 78956
rect 78880 78886 78886 78950
rect 78950 78886 78956 78950
rect 67728 78270 67804 78276
rect 67728 78206 67734 78270
rect 67798 78206 67804 78270
rect 67728 77862 67804 78206
rect 67728 77830 67734 77862
rect 67733 77798 67734 77830
rect 67798 77830 67804 77862
rect 69224 78270 69300 78276
rect 69224 78206 69230 78270
rect 69294 78206 69300 78270
rect 69224 77862 69300 78206
rect 69224 77830 69230 77862
rect 67798 77798 67799 77830
rect 67733 77797 67799 77798
rect 69229 77798 69230 77830
rect 69294 77830 69300 77862
rect 71128 78270 71204 78276
rect 71128 78206 71134 78270
rect 71198 78206 71204 78270
rect 71128 77862 71204 78206
rect 71128 77830 71134 77862
rect 69294 77798 69295 77830
rect 69229 77797 69295 77798
rect 71133 77798 71134 77830
rect 71198 77830 71204 77862
rect 72760 78270 72836 78276
rect 72760 78206 72766 78270
rect 72830 78206 72836 78270
rect 72760 77862 72836 78206
rect 72760 77830 72766 77862
rect 71198 77798 71199 77830
rect 71133 77797 71199 77798
rect 72765 77798 72766 77830
rect 72830 77830 72836 77862
rect 74392 78270 74468 78276
rect 74392 78206 74398 78270
rect 74462 78206 74468 78270
rect 74392 77862 74468 78206
rect 74392 77830 74398 77862
rect 72830 77798 72831 77830
rect 72765 77797 72831 77798
rect 74397 77798 74398 77830
rect 74462 77830 74468 77862
rect 76160 78270 76236 78276
rect 76160 78206 76166 78270
rect 76230 78206 76236 78270
rect 76160 77862 76236 78206
rect 76160 77830 76166 77862
rect 74462 77798 74463 77830
rect 74397 77797 74463 77798
rect 76165 77798 76166 77830
rect 76230 77830 76236 77862
rect 77656 78270 77732 78276
rect 77656 78206 77662 78270
rect 77726 78206 77732 78270
rect 77656 77862 77732 78206
rect 77656 77830 77662 77862
rect 76230 77798 76231 77830
rect 76165 77797 76231 77798
rect 77661 77798 77662 77830
rect 77726 77830 77732 77862
rect 77726 77798 77727 77830
rect 77661 77797 77727 77798
rect 78880 76502 78956 78886
rect 79288 78270 79364 78276
rect 79288 78206 79294 78270
rect 79358 78206 79364 78270
rect 79288 77862 79364 78206
rect 79288 77830 79294 77862
rect 79293 77798 79294 77830
rect 79358 77830 79364 77862
rect 79358 77798 79359 77830
rect 79293 77797 79359 77798
rect 78880 76470 78886 76502
rect 78885 76438 78886 76470
rect 78950 76470 78956 76502
rect 79288 77726 79364 77732
rect 79288 77662 79294 77726
rect 79358 77662 79364 77726
rect 78950 76438 78951 76470
rect 78885 76437 78951 76438
rect 79288 75142 79364 77662
rect 79424 75958 79500 79500
rect 82144 78950 82220 78956
rect 82144 78886 82150 78950
rect 82214 78886 82220 78950
rect 81192 78270 81268 78276
rect 81192 78206 81198 78270
rect 81262 78206 81268 78270
rect 81192 77862 81268 78206
rect 81192 77830 81198 77862
rect 81197 77798 81198 77830
rect 81262 77830 81268 77862
rect 81262 77798 81263 77830
rect 81197 77797 81263 77798
rect 81877 77726 81943 77727
rect 81877 77694 81878 77726
rect 79424 75926 79430 75958
rect 79429 75894 79430 75926
rect 79494 75926 79500 75958
rect 81872 77662 81878 77694
rect 81942 77694 81943 77726
rect 81942 77662 81948 77694
rect 79494 75894 79495 75926
rect 79429 75893 79495 75894
rect 81872 75822 81948 77662
rect 82144 77182 82220 78886
rect 82688 78270 82764 78276
rect 82688 78206 82694 78270
rect 82758 78206 82764 78270
rect 82688 77862 82764 78206
rect 82688 77830 82694 77862
rect 82693 77798 82694 77830
rect 82758 77830 82764 77862
rect 84456 78270 84532 78276
rect 84456 78206 84462 78270
rect 84526 78206 84532 78270
rect 84456 77862 84532 78206
rect 84456 77830 84462 77862
rect 82758 77798 82759 77830
rect 82693 77797 82759 77798
rect 84461 77798 84462 77830
rect 84526 77830 84532 77862
rect 86224 78270 86300 78276
rect 86224 78206 86230 78270
rect 86294 78206 86300 78270
rect 86224 77862 86300 78206
rect 86224 77830 86230 77862
rect 84526 77798 84527 77830
rect 84461 77797 84527 77798
rect 86229 77798 86230 77830
rect 86294 77830 86300 77862
rect 87720 78270 87796 78276
rect 87720 78206 87726 78270
rect 87790 78206 87796 78270
rect 87720 77862 87796 78206
rect 87720 77830 87726 77862
rect 86294 77798 86295 77830
rect 86229 77797 86295 77798
rect 87725 77798 87726 77830
rect 87790 77830 87796 77862
rect 89624 78270 89700 78276
rect 89624 78206 89630 78270
rect 89694 78206 89700 78270
rect 89624 77862 89700 78206
rect 89624 77830 89630 77862
rect 87790 77798 87791 77830
rect 87725 77797 87791 77798
rect 89629 77798 89630 77830
rect 89694 77830 89700 77862
rect 89694 77798 89695 77830
rect 89629 77797 89695 77798
rect 82144 77150 82150 77182
rect 82149 77118 82150 77150
rect 82214 77150 82220 77182
rect 82214 77118 82215 77150
rect 82149 77117 82215 77118
rect 82013 77046 82079 77047
rect 82013 77014 82014 77046
rect 81872 75758 81878 75822
rect 81942 75758 81948 75822
rect 81872 75752 81948 75758
rect 82008 76982 82014 77014
rect 82078 77014 82079 77046
rect 82078 76982 82084 77014
rect 79288 75110 79294 75142
rect 79293 75078 79294 75110
rect 79358 75110 79364 75142
rect 81872 75686 81948 75692
rect 81872 75622 81878 75686
rect 81942 75622 81948 75686
rect 79358 75078 79359 75110
rect 79293 75077 79359 75078
rect 66912 74158 66918 74190
rect 65622 74126 65623 74158
rect 65557 74125 65623 74126
rect 66917 74126 66918 74158
rect 66982 74158 66988 74190
rect 66982 74126 66983 74158
rect 66917 74125 66983 74126
rect 31149 74054 31215 74055
rect 31149 74022 31150 74054
rect 29784 73854 29790 73918
rect 29854 73854 29860 73918
rect 29784 73848 29860 73854
rect 31144 73990 31150 74022
rect 31214 74022 31215 74054
rect 31214 73990 31220 74022
rect 28560 73782 28636 73788
rect 28560 73718 28566 73782
rect 28630 73718 28636 73782
rect 28560 73102 28636 73718
rect 28560 73070 28566 73102
rect 28565 73038 28566 73070
rect 28630 73070 28636 73102
rect 29784 73782 29860 73788
rect 29784 73718 29790 73782
rect 29854 73718 29860 73782
rect 29784 73102 29860 73718
rect 29784 73070 29790 73102
rect 28630 73038 28631 73070
rect 28565 73037 28631 73038
rect 29789 73038 29790 73070
rect 29854 73070 29860 73102
rect 31008 73782 31084 73788
rect 31008 73718 31014 73782
rect 31078 73718 31084 73782
rect 31008 73102 31084 73718
rect 31008 73070 31014 73102
rect 29854 73038 29855 73070
rect 29789 73037 29855 73038
rect 31013 73038 31014 73070
rect 31078 73070 31084 73102
rect 31078 73038 31079 73070
rect 31013 73037 31079 73038
rect 952 72494 1230 72558
rect 1294 72494 1300 72558
rect 952 70926 1300 72494
rect 30872 72830 30948 72836
rect 30872 72766 30878 72830
rect 30942 72766 30948 72830
rect 28565 72286 28631 72287
rect 28565 72254 28566 72286
rect 952 70862 1230 70926
rect 1294 70862 1300 70926
rect 952 69158 1300 70862
rect 28560 72222 28566 72254
rect 28630 72254 28631 72286
rect 28630 72222 28636 72254
rect 28560 70518 28636 72222
rect 28560 70454 28566 70518
rect 28630 70454 28636 70518
rect 28560 70448 28636 70454
rect 952 69094 1230 69158
rect 1294 69094 1300 69158
rect 952 67662 1300 69094
rect 27608 70382 27684 70388
rect 27608 70318 27614 70382
rect 27678 70318 27684 70382
rect 27608 68206 27684 70318
rect 30872 69022 30948 72766
rect 31144 72286 31220 73990
rect 32096 73782 32172 73788
rect 32096 73718 32102 73782
rect 32166 73718 32172 73782
rect 32096 73102 32172 73718
rect 32096 73070 32102 73102
rect 32101 73038 32102 73070
rect 32166 73070 32172 73102
rect 33456 73782 33532 73788
rect 33456 73718 33462 73782
rect 33526 73718 33532 73782
rect 33456 73102 33532 73718
rect 33456 73070 33462 73102
rect 32166 73038 32167 73070
rect 32101 73037 32167 73038
rect 33461 73038 33462 73070
rect 33526 73070 33532 73102
rect 34680 73782 34756 73788
rect 34680 73718 34686 73782
rect 34750 73718 34756 73782
rect 34680 73102 34756 73718
rect 34680 73070 34686 73102
rect 33526 73038 33527 73070
rect 33461 73037 33527 73038
rect 34685 73038 34686 73070
rect 34750 73070 34756 73102
rect 36040 73782 36116 73788
rect 36040 73718 36046 73782
rect 36110 73718 36116 73782
rect 36040 73102 36116 73718
rect 36040 73070 36046 73102
rect 34750 73038 34751 73070
rect 34685 73037 34751 73038
rect 36045 73038 36046 73070
rect 36110 73070 36116 73102
rect 37264 73782 37340 73788
rect 37264 73718 37270 73782
rect 37334 73718 37340 73782
rect 37264 73102 37340 73718
rect 37264 73070 37270 73102
rect 36110 73038 36111 73070
rect 36045 73037 36111 73038
rect 37269 73038 37270 73070
rect 37334 73070 37340 73102
rect 38488 73782 38564 73788
rect 38488 73718 38494 73782
rect 38558 73718 38564 73782
rect 38488 73102 38564 73718
rect 38488 73070 38494 73102
rect 37334 73038 37335 73070
rect 37269 73037 37335 73038
rect 38493 73038 38494 73070
rect 38558 73070 38564 73102
rect 39712 73782 39788 73788
rect 39712 73718 39718 73782
rect 39782 73718 39788 73782
rect 39712 73102 39788 73718
rect 39712 73070 39718 73102
rect 38558 73038 38559 73070
rect 38493 73037 38559 73038
rect 39717 73038 39718 73070
rect 39782 73070 39788 73102
rect 40800 73782 40876 73788
rect 40800 73718 40806 73782
rect 40870 73718 40876 73782
rect 42029 73782 42095 73783
rect 42029 73750 42030 73782
rect 40800 73102 40876 73718
rect 40800 73070 40806 73102
rect 39782 73038 39783 73070
rect 39717 73037 39783 73038
rect 40805 73038 40806 73070
rect 40870 73070 40876 73102
rect 42024 73718 42030 73750
rect 42094 73750 42095 73782
rect 42296 73782 42372 73788
rect 42094 73718 42100 73750
rect 42024 73102 42100 73718
rect 40870 73038 40871 73070
rect 40805 73037 40871 73038
rect 42024 73038 42030 73102
rect 42094 73038 42100 73102
rect 42296 73718 42302 73782
rect 42366 73718 42372 73782
rect 42296 73102 42372 73718
rect 42296 73070 42302 73102
rect 42024 73032 42100 73038
rect 42301 73038 42302 73070
rect 42366 73070 42372 73102
rect 43384 73782 43460 73788
rect 43384 73718 43390 73782
rect 43454 73718 43460 73782
rect 43384 73102 43460 73718
rect 43384 73070 43390 73102
rect 42366 73038 42367 73070
rect 42301 73037 42367 73038
rect 43389 73038 43390 73070
rect 43454 73070 43460 73102
rect 44744 73782 44820 73788
rect 44744 73718 44750 73782
rect 44814 73718 44820 73782
rect 44744 73102 44820 73718
rect 44744 73070 44750 73102
rect 43454 73038 43455 73070
rect 43389 73037 43455 73038
rect 44749 73038 44750 73070
rect 44814 73070 44820 73102
rect 45968 73782 46044 73788
rect 45968 73718 45974 73782
rect 46038 73718 46044 73782
rect 45968 73102 46044 73718
rect 45968 73070 45974 73102
rect 44814 73038 44815 73070
rect 44749 73037 44815 73038
rect 45973 73038 45974 73070
rect 46038 73070 46044 73102
rect 47192 73782 47268 73788
rect 47192 73718 47198 73782
rect 47262 73718 47268 73782
rect 47192 73102 47268 73718
rect 47192 73070 47198 73102
rect 46038 73038 46039 73070
rect 45973 73037 46039 73038
rect 47197 73038 47198 73070
rect 47262 73070 47268 73102
rect 48552 73782 48628 73788
rect 48552 73718 48558 73782
rect 48622 73718 48628 73782
rect 48552 73102 48628 73718
rect 48552 73070 48558 73102
rect 47262 73038 47263 73070
rect 47197 73037 47263 73038
rect 48557 73038 48558 73070
rect 48622 73070 48628 73102
rect 49776 73782 49852 73788
rect 49776 73718 49782 73782
rect 49846 73718 49852 73782
rect 49776 73102 49852 73718
rect 49776 73070 49782 73102
rect 48622 73038 48623 73070
rect 48557 73037 48623 73038
rect 49781 73038 49782 73070
rect 49846 73070 49852 73102
rect 51000 73782 51076 73788
rect 51000 73718 51006 73782
rect 51070 73718 51076 73782
rect 51000 73102 51076 73718
rect 51000 73070 51006 73102
rect 49846 73038 49847 73070
rect 49781 73037 49847 73038
rect 51005 73038 51006 73070
rect 51070 73070 51076 73102
rect 52088 73782 52164 73788
rect 52088 73718 52094 73782
rect 52158 73718 52164 73782
rect 52088 73102 52164 73718
rect 52088 73070 52094 73102
rect 51070 73038 51071 73070
rect 51005 73037 51071 73038
rect 52093 73038 52094 73070
rect 52158 73070 52164 73102
rect 53448 73782 53524 73788
rect 53448 73718 53454 73782
rect 53518 73718 53524 73782
rect 53448 73102 53524 73718
rect 53448 73070 53454 73102
rect 52158 73038 52159 73070
rect 52093 73037 52159 73038
rect 53453 73038 53454 73070
rect 53518 73070 53524 73102
rect 54672 73782 54748 73788
rect 54672 73718 54678 73782
rect 54742 73718 54748 73782
rect 54672 73102 54748 73718
rect 54672 73070 54678 73102
rect 53518 73038 53519 73070
rect 53453 73037 53519 73038
rect 54677 73038 54678 73070
rect 54742 73070 54748 73102
rect 56032 73782 56108 73788
rect 56032 73718 56038 73782
rect 56102 73718 56108 73782
rect 56032 73102 56108 73718
rect 56032 73070 56038 73102
rect 54742 73038 54743 73070
rect 54677 73037 54743 73038
rect 56037 73038 56038 73070
rect 56102 73070 56108 73102
rect 57256 73782 57332 73788
rect 57256 73718 57262 73782
rect 57326 73718 57332 73782
rect 57256 73102 57332 73718
rect 57256 73070 57262 73102
rect 56102 73038 56103 73070
rect 56037 73037 56103 73038
rect 57261 73038 57262 73070
rect 57326 73070 57332 73102
rect 58480 73782 58556 73788
rect 58480 73718 58486 73782
rect 58550 73718 58556 73782
rect 58480 73102 58556 73718
rect 58480 73070 58486 73102
rect 57326 73038 57327 73070
rect 57261 73037 57327 73038
rect 58485 73038 58486 73070
rect 58550 73070 58556 73102
rect 59704 73782 59780 73788
rect 59704 73718 59710 73782
rect 59774 73718 59780 73782
rect 59704 73102 59780 73718
rect 59704 73070 59710 73102
rect 58550 73038 58551 73070
rect 58485 73037 58551 73038
rect 59709 73038 59710 73070
rect 59774 73070 59780 73102
rect 60792 73782 60868 73788
rect 60792 73718 60798 73782
rect 60862 73718 60868 73782
rect 60792 73102 60868 73718
rect 60792 73070 60798 73102
rect 59774 73038 59775 73070
rect 59709 73037 59775 73038
rect 60797 73038 60798 73070
rect 60862 73070 60868 73102
rect 62152 73782 62228 73788
rect 62152 73718 62158 73782
rect 62222 73718 62228 73782
rect 62152 73102 62228 73718
rect 62152 73070 62158 73102
rect 60862 73038 60863 73070
rect 60797 73037 60863 73038
rect 62157 73038 62158 73070
rect 62222 73070 62228 73102
rect 63512 73782 63588 73788
rect 63512 73718 63518 73782
rect 63582 73718 63588 73782
rect 63512 73102 63588 73718
rect 63512 73070 63518 73102
rect 62222 73038 62223 73070
rect 62157 73037 62223 73038
rect 63517 73038 63518 73070
rect 63582 73070 63588 73102
rect 64736 73782 64812 73788
rect 64736 73718 64742 73782
rect 64806 73718 64812 73782
rect 64736 73102 64812 73718
rect 64736 73070 64742 73102
rect 63582 73038 63583 73070
rect 63517 73037 63583 73038
rect 64741 73038 64742 73070
rect 64806 73070 64812 73102
rect 65960 73782 66036 73788
rect 65960 73718 65966 73782
rect 66030 73718 66036 73782
rect 65960 73102 66036 73718
rect 65960 73070 65966 73102
rect 64806 73038 64807 73070
rect 64741 73037 64807 73038
rect 65965 73038 65966 73070
rect 66030 73070 66036 73102
rect 67184 73782 67260 73788
rect 67184 73718 67190 73782
rect 67254 73718 67260 73782
rect 67184 73102 67260 73718
rect 67184 73070 67190 73102
rect 66030 73038 66031 73070
rect 65965 73037 66031 73038
rect 67189 73038 67190 73070
rect 67254 73070 67260 73102
rect 67254 73038 67255 73070
rect 67189 73037 67255 73038
rect 74805 72966 74871 72967
rect 74805 72934 74806 72966
rect 31144 72222 31150 72286
rect 31214 72222 31220 72286
rect 31144 72216 31220 72222
rect 74800 72902 74806 72934
rect 74870 72934 74871 72966
rect 81872 72966 81948 75622
rect 82008 74326 82084 76982
rect 90032 76502 90108 79500
rect 95336 79222 95684 79228
rect 95336 79158 95342 79222
rect 95406 79158 95478 79222
rect 95542 79158 95614 79222
rect 95678 79158 95684 79222
rect 95336 79086 95684 79158
rect 95336 79022 95342 79086
rect 95406 79022 95478 79086
rect 95542 79022 95614 79086
rect 95678 79022 95684 79086
rect 95336 78950 95684 79022
rect 95336 78886 95342 78950
rect 95406 78886 95478 78950
rect 95542 78886 95614 78950
rect 95678 78886 95684 78950
rect 94656 78542 95004 78548
rect 94656 78478 94662 78542
rect 94726 78478 94798 78542
rect 94862 78478 94934 78542
rect 94998 78478 95004 78542
rect 94656 78406 95004 78478
rect 94656 78342 94662 78406
rect 94726 78342 94798 78406
rect 94862 78342 94934 78406
rect 94998 78342 95004 78406
rect 91256 78270 91332 78276
rect 91256 78206 91262 78270
rect 91326 78206 91332 78270
rect 91256 77862 91332 78206
rect 91256 77830 91262 77862
rect 91261 77798 91262 77830
rect 91326 77830 91332 77862
rect 92888 78270 92964 78276
rect 92888 78206 92894 78270
rect 92958 78206 92964 78270
rect 92888 77862 92964 78206
rect 92888 77830 92894 77862
rect 91326 77798 91327 77830
rect 91261 77797 91327 77798
rect 92893 77798 92894 77830
rect 92958 77830 92964 77862
rect 94656 78270 95004 78342
rect 94656 78206 94662 78270
rect 94726 78206 94798 78270
rect 94862 78206 94934 78270
rect 94998 78206 95004 78270
rect 92958 77798 92959 77830
rect 92893 77797 92959 77798
rect 90032 76470 90038 76502
rect 90037 76438 90038 76470
rect 90102 76470 90108 76502
rect 90102 76438 90103 76470
rect 90037 76437 90103 76438
rect 82008 74262 82014 74326
rect 82078 74262 82084 74326
rect 82008 74256 82084 74262
rect 94656 75958 95004 78206
rect 94656 75894 94662 75958
rect 94726 75894 95004 75958
rect 94656 74326 95004 75894
rect 94656 74262 94662 74326
rect 94726 74262 95004 74326
rect 81872 72934 81878 72966
rect 74870 72902 74876 72934
rect 74664 71606 74740 71612
rect 74664 71542 74670 71606
rect 74734 71542 74740 71606
rect 68957 70382 69023 70383
rect 68957 70350 68958 70382
rect 30872 68990 30878 69022
rect 30877 68958 30878 68990
rect 30942 68990 30948 69022
rect 68952 70318 68958 70350
rect 69022 70350 69023 70382
rect 69022 70318 69028 70350
rect 30942 68958 30943 68990
rect 30877 68957 30943 68958
rect 28293 68750 28359 68751
rect 28293 68718 28294 68750
rect 28288 68686 28294 68718
rect 28358 68718 28359 68750
rect 29245 68750 29311 68751
rect 29245 68718 29246 68750
rect 28358 68686 28364 68718
rect 28288 68342 28364 68686
rect 28288 68278 28294 68342
rect 28358 68278 28364 68342
rect 28288 68272 28364 68278
rect 29240 68686 29246 68718
rect 29310 68718 29311 68750
rect 30328 68750 30404 68756
rect 29310 68686 29316 68718
rect 27608 68174 27614 68206
rect 27613 68142 27614 68174
rect 27678 68174 27684 68206
rect 29240 68206 29316 68686
rect 30328 68686 30334 68750
rect 30398 68686 30404 68750
rect 30605 68750 30671 68751
rect 30605 68718 30606 68750
rect 30328 68342 30404 68686
rect 30328 68310 30334 68342
rect 30333 68278 30334 68310
rect 30398 68310 30404 68342
rect 30600 68686 30606 68718
rect 30670 68718 30671 68750
rect 31552 68750 31628 68756
rect 30670 68686 30676 68718
rect 30600 68342 30676 68686
rect 30398 68278 30399 68310
rect 30333 68277 30399 68278
rect 30600 68278 30606 68342
rect 30670 68278 30676 68342
rect 31552 68686 31558 68750
rect 31622 68686 31628 68750
rect 31693 68750 31759 68751
rect 31693 68718 31694 68750
rect 31552 68342 31628 68686
rect 31552 68310 31558 68342
rect 30600 68272 30676 68278
rect 31557 68278 31558 68310
rect 31622 68310 31628 68342
rect 31688 68686 31694 68718
rect 31758 68718 31759 68750
rect 32776 68750 32852 68756
rect 31758 68686 31764 68718
rect 31688 68342 31764 68686
rect 31622 68278 31623 68310
rect 31557 68277 31623 68278
rect 31688 68278 31694 68342
rect 31758 68278 31764 68342
rect 32776 68686 32782 68750
rect 32846 68686 32852 68750
rect 33325 68750 33391 68751
rect 33325 68718 33326 68750
rect 32776 68342 32852 68686
rect 32776 68310 32782 68342
rect 31688 68272 31764 68278
rect 32781 68278 32782 68310
rect 32846 68310 32852 68342
rect 33320 68686 33326 68718
rect 33390 68718 33391 68750
rect 34136 68750 34212 68756
rect 33390 68686 33396 68718
rect 33320 68342 33396 68686
rect 32846 68278 32847 68310
rect 32781 68277 32847 68278
rect 33320 68278 33326 68342
rect 33390 68278 33396 68342
rect 34136 68686 34142 68750
rect 34206 68686 34212 68750
rect 34136 68342 34212 68686
rect 34136 68310 34142 68342
rect 33320 68272 33396 68278
rect 34141 68278 34142 68310
rect 34206 68310 34212 68342
rect 35224 68750 35300 68756
rect 35224 68686 35230 68750
rect 35294 68686 35300 68750
rect 35773 68750 35839 68751
rect 35773 68718 35774 68750
rect 35224 68342 35300 68686
rect 35224 68310 35230 68342
rect 34206 68278 34207 68310
rect 34141 68277 34207 68278
rect 35229 68278 35230 68310
rect 35294 68310 35300 68342
rect 35768 68686 35774 68718
rect 35838 68718 35839 68750
rect 36584 68750 36660 68756
rect 35838 68686 35844 68718
rect 35768 68342 35844 68686
rect 35294 68278 35295 68310
rect 35229 68277 35295 68278
rect 35768 68278 35774 68342
rect 35838 68278 35844 68342
rect 36584 68686 36590 68750
rect 36654 68686 36660 68750
rect 36584 68342 36660 68686
rect 36584 68310 36590 68342
rect 35768 68272 35844 68278
rect 36589 68278 36590 68310
rect 36654 68310 36660 68342
rect 37808 68750 37884 68756
rect 37808 68686 37814 68750
rect 37878 68686 37884 68750
rect 38357 68750 38423 68751
rect 38357 68718 38358 68750
rect 37808 68342 37884 68686
rect 37808 68310 37814 68342
rect 36654 68278 36655 68310
rect 36589 68277 36655 68278
rect 37813 68278 37814 68310
rect 37878 68310 37884 68342
rect 38352 68686 38358 68718
rect 38422 68718 38423 68750
rect 39032 68750 39108 68756
rect 38422 68686 38428 68718
rect 38352 68342 38428 68686
rect 37878 68278 37879 68310
rect 37813 68277 37879 68278
rect 38352 68278 38358 68342
rect 38422 68278 38428 68342
rect 39032 68686 39038 68750
rect 39102 68686 39108 68750
rect 39309 68750 39375 68751
rect 39309 68718 39310 68750
rect 39032 68342 39108 68686
rect 39032 68310 39038 68342
rect 38352 68272 38428 68278
rect 39037 68278 39038 68310
rect 39102 68310 39108 68342
rect 39304 68686 39310 68718
rect 39374 68718 39375 68750
rect 40256 68750 40332 68756
rect 39374 68686 39380 68718
rect 39304 68342 39380 68686
rect 39102 68278 39103 68310
rect 39037 68277 39103 68278
rect 39304 68278 39310 68342
rect 39374 68278 39380 68342
rect 40256 68686 40262 68750
rect 40326 68686 40332 68750
rect 40256 68342 40332 68686
rect 40256 68310 40262 68342
rect 39304 68272 39380 68278
rect 40261 68278 40262 68310
rect 40326 68310 40332 68342
rect 41888 68750 41964 68756
rect 41888 68686 41894 68750
rect 41958 68686 41964 68750
rect 41888 68342 41964 68686
rect 41888 68310 41894 68342
rect 40326 68278 40327 68310
rect 40261 68277 40327 68278
rect 41893 68278 41894 68310
rect 41958 68310 41964 68342
rect 42840 68750 42916 68756
rect 42840 68686 42846 68750
rect 42910 68686 42916 68750
rect 43389 68750 43455 68751
rect 43389 68718 43390 68750
rect 42840 68342 42916 68686
rect 42840 68310 42846 68342
rect 41958 68278 41959 68310
rect 41893 68277 41959 68278
rect 42845 68278 42846 68310
rect 42910 68310 42916 68342
rect 43384 68686 43390 68718
rect 43454 68718 43455 68750
rect 44064 68750 44140 68756
rect 43454 68686 43460 68718
rect 43384 68342 43460 68686
rect 42910 68278 42911 68310
rect 42845 68277 42911 68278
rect 43384 68278 43390 68342
rect 43454 68278 43460 68342
rect 44064 68686 44070 68750
rect 44134 68686 44140 68750
rect 45837 68750 45903 68751
rect 45837 68718 45838 68750
rect 44064 68342 44140 68686
rect 44064 68310 44070 68342
rect 43384 68272 43460 68278
rect 44069 68278 44070 68310
rect 44134 68310 44140 68342
rect 45832 68686 45838 68718
rect 45902 68718 45903 68750
rect 46512 68750 46588 68756
rect 45902 68686 45908 68718
rect 45832 68342 45908 68686
rect 44134 68278 44135 68310
rect 44069 68277 44135 68278
rect 45832 68278 45838 68342
rect 45902 68278 45908 68342
rect 46512 68686 46518 68750
rect 46582 68686 46588 68750
rect 47061 68750 47127 68751
rect 47061 68718 47062 68750
rect 46512 68342 46588 68686
rect 46512 68310 46518 68342
rect 45832 68272 45908 68278
rect 46517 68278 46518 68310
rect 46582 68310 46588 68342
rect 47056 68686 47062 68718
rect 47126 68718 47127 68750
rect 47736 68750 47812 68756
rect 47126 68686 47132 68718
rect 47056 68342 47132 68686
rect 46582 68278 46583 68310
rect 46517 68277 46583 68278
rect 47056 68278 47062 68342
rect 47126 68278 47132 68342
rect 47736 68686 47742 68750
rect 47806 68686 47812 68750
rect 47736 68342 47812 68686
rect 47736 68310 47742 68342
rect 47056 68272 47132 68278
rect 47741 68278 47742 68310
rect 47806 68310 47812 68342
rect 48960 68750 49036 68756
rect 48960 68686 48966 68750
rect 49030 68686 49036 68750
rect 48960 68342 49036 68686
rect 48960 68310 48966 68342
rect 47806 68278 47807 68310
rect 47741 68277 47807 68278
rect 48965 68278 48966 68310
rect 49030 68310 49036 68342
rect 50592 68750 50668 68756
rect 50592 68686 50598 68750
rect 50662 68686 50668 68750
rect 50592 68342 50668 68686
rect 50592 68310 50598 68342
rect 49030 68278 49031 68310
rect 48965 68277 49031 68278
rect 50597 68278 50598 68310
rect 50662 68310 50668 68342
rect 51544 68750 51620 68756
rect 51544 68686 51550 68750
rect 51614 68686 51620 68750
rect 52093 68750 52159 68751
rect 52093 68718 52094 68750
rect 51544 68342 51620 68686
rect 51544 68310 51550 68342
rect 50662 68278 50663 68310
rect 50597 68277 50663 68278
rect 51549 68278 51550 68310
rect 51614 68310 51620 68342
rect 52088 68686 52094 68718
rect 52158 68718 52159 68750
rect 52768 68750 52844 68756
rect 52158 68686 52164 68718
rect 52088 68342 52164 68686
rect 51614 68278 51615 68310
rect 51549 68277 51615 68278
rect 52088 68278 52094 68342
rect 52158 68278 52164 68342
rect 52768 68686 52774 68750
rect 52838 68686 52844 68750
rect 53045 68750 53111 68751
rect 53045 68718 53046 68750
rect 52768 68342 52844 68686
rect 52768 68310 52774 68342
rect 52088 68272 52164 68278
rect 52773 68278 52774 68310
rect 52838 68310 52844 68342
rect 53040 68686 53046 68718
rect 53110 68718 53111 68750
rect 53992 68750 54068 68756
rect 53110 68686 53116 68718
rect 53040 68342 53116 68686
rect 52838 68278 52839 68310
rect 52773 68277 52839 68278
rect 53040 68278 53046 68342
rect 53110 68278 53116 68342
rect 53992 68686 53998 68750
rect 54062 68686 54068 68750
rect 53992 68342 54068 68686
rect 53992 68310 53998 68342
rect 53040 68272 53116 68278
rect 53997 68278 53998 68310
rect 54062 68310 54068 68342
rect 55216 68750 55292 68756
rect 55216 68686 55222 68750
rect 55286 68686 55292 68750
rect 55765 68750 55831 68751
rect 55765 68718 55766 68750
rect 55216 68342 55292 68686
rect 55216 68310 55222 68342
rect 54062 68278 54063 68310
rect 53997 68277 54063 68278
rect 55221 68278 55222 68310
rect 55286 68310 55292 68342
rect 55760 68686 55766 68718
rect 55830 68718 55831 68750
rect 56848 68750 56924 68756
rect 55830 68686 55836 68718
rect 55760 68342 55836 68686
rect 55286 68278 55287 68310
rect 55221 68277 55287 68278
rect 55760 68278 55766 68342
rect 55830 68278 55836 68342
rect 56848 68686 56854 68750
rect 56918 68686 56924 68750
rect 56848 68342 56924 68686
rect 56848 68310 56854 68342
rect 55760 68272 55836 68278
rect 56853 68278 56854 68310
rect 56918 68310 56924 68342
rect 57800 68750 57876 68756
rect 57800 68686 57806 68750
rect 57870 68686 57876 68750
rect 57941 68750 58007 68751
rect 57941 68718 57942 68750
rect 57800 68342 57876 68686
rect 57800 68310 57806 68342
rect 56918 68278 56919 68310
rect 56853 68277 56919 68278
rect 57805 68278 57806 68310
rect 57870 68310 57876 68342
rect 57936 68686 57942 68718
rect 58006 68718 58007 68750
rect 59024 68750 59100 68756
rect 58006 68686 58012 68718
rect 57936 68342 58012 68686
rect 57870 68278 57871 68310
rect 57805 68277 57871 68278
rect 57936 68278 57942 68342
rect 58006 68278 58012 68342
rect 59024 68686 59030 68750
rect 59094 68686 59100 68750
rect 59573 68750 59639 68751
rect 59573 68718 59574 68750
rect 59024 68342 59100 68686
rect 59024 68310 59030 68342
rect 57936 68272 58012 68278
rect 59029 68278 59030 68310
rect 59094 68310 59100 68342
rect 59568 68686 59574 68718
rect 59638 68718 59639 68750
rect 60248 68750 60324 68756
rect 59638 68686 59644 68718
rect 59568 68342 59644 68686
rect 59094 68278 59095 68310
rect 59029 68277 59095 68278
rect 59568 68278 59574 68342
rect 59638 68278 59644 68342
rect 60248 68686 60254 68750
rect 60318 68686 60324 68750
rect 60797 68750 60863 68751
rect 60797 68718 60798 68750
rect 60248 68342 60324 68686
rect 60248 68310 60254 68342
rect 59568 68272 59644 68278
rect 60253 68278 60254 68310
rect 60318 68310 60324 68342
rect 60792 68686 60798 68718
rect 60862 68718 60863 68750
rect 61472 68750 61548 68756
rect 60862 68686 60868 68718
rect 60792 68342 60868 68686
rect 60318 68278 60319 68310
rect 60253 68277 60319 68278
rect 60792 68278 60798 68342
rect 60862 68278 60868 68342
rect 61472 68686 61478 68750
rect 61542 68686 61548 68750
rect 61472 68342 61548 68686
rect 61472 68310 61478 68342
rect 60792 68272 60868 68278
rect 61477 68278 61478 68310
rect 61542 68310 61548 68342
rect 62696 68750 62772 68756
rect 62696 68686 62702 68750
rect 62766 68686 62772 68750
rect 62696 68342 62772 68686
rect 62696 68310 62702 68342
rect 61542 68278 61543 68310
rect 61477 68277 61543 68278
rect 62701 68278 62702 68310
rect 62766 68310 62772 68342
rect 64056 68750 64132 68756
rect 64056 68686 64062 68750
rect 64126 68686 64132 68750
rect 64056 68342 64132 68686
rect 64056 68310 64062 68342
rect 62766 68278 62767 68310
rect 62701 68277 62767 68278
rect 64061 68278 64062 68310
rect 64126 68310 64132 68342
rect 65280 68750 65356 68756
rect 65280 68686 65286 68750
rect 65350 68686 65356 68750
rect 65280 68342 65356 68686
rect 65280 68310 65286 68342
rect 64126 68278 64127 68310
rect 64061 68277 64127 68278
rect 65285 68278 65286 68310
rect 65350 68310 65356 68342
rect 66504 68750 66580 68756
rect 66504 68686 66510 68750
rect 66574 68686 66580 68750
rect 67053 68750 67119 68751
rect 67053 68718 67054 68750
rect 66504 68342 66580 68686
rect 66504 68310 66510 68342
rect 65350 68278 65351 68310
rect 65285 68277 65351 68278
rect 66509 68278 66510 68310
rect 66574 68310 66580 68342
rect 67048 68686 67054 68718
rect 67118 68718 67119 68750
rect 67728 68750 67804 68756
rect 67118 68686 67124 68718
rect 67048 68342 67124 68686
rect 66574 68278 66575 68310
rect 66509 68277 66575 68278
rect 67048 68278 67054 68342
rect 67118 68278 67124 68342
rect 67728 68686 67734 68750
rect 67798 68686 67804 68750
rect 68277 68750 68343 68751
rect 68277 68718 68278 68750
rect 67728 68342 67804 68686
rect 67728 68310 67734 68342
rect 67048 68272 67124 68278
rect 67733 68278 67734 68310
rect 67798 68310 67804 68342
rect 68272 68686 68278 68718
rect 68342 68718 68343 68750
rect 68342 68686 68348 68718
rect 68272 68342 68348 68686
rect 67798 68278 67799 68310
rect 67733 68277 67799 68278
rect 68272 68278 68278 68342
rect 68342 68278 68348 68342
rect 68272 68272 68348 68278
rect 27678 68142 27679 68174
rect 27613 68141 27679 68142
rect 29240 68142 29246 68206
rect 29310 68142 29316 68206
rect 29240 68136 29316 68142
rect 26933 68070 26999 68071
rect 26933 68038 26934 68070
rect 26928 68006 26934 68038
rect 26998 68038 26999 68070
rect 26998 68006 27004 68038
rect 26928 67798 27004 68006
rect 26928 67734 26934 67798
rect 26998 67734 27004 67798
rect 26928 67728 27004 67734
rect 68952 67798 69028 70318
rect 74528 70246 74604 70252
rect 74528 70182 74534 70246
rect 74598 70182 74604 70246
rect 70317 68342 70383 68343
rect 70317 68310 70318 68342
rect 70312 68278 70318 68310
rect 70382 68310 70383 68342
rect 70382 68278 70388 68310
rect 68952 67734 68958 67798
rect 69022 67734 69028 67798
rect 69360 68070 69436 68076
rect 69360 68006 69366 68070
rect 69430 68006 69436 68070
rect 69360 67798 69436 68006
rect 70312 68070 70388 68278
rect 70312 68006 70318 68070
rect 70382 68006 70388 68070
rect 70312 68000 70388 68006
rect 69360 67766 69366 67798
rect 68952 67728 69028 67734
rect 69365 67734 69366 67766
rect 69430 67766 69436 67798
rect 73853 67798 73919 67799
rect 73853 67766 73854 67798
rect 69430 67734 69431 67766
rect 69365 67733 69431 67734
rect 73848 67734 73854 67766
rect 73918 67766 73919 67798
rect 73918 67734 73924 67766
rect 952 67598 1230 67662
rect 1294 67598 1300 67662
rect 952 66030 1300 67598
rect 73848 67390 73924 67734
rect 73848 67326 73854 67390
rect 73918 67326 73924 67390
rect 74528 67390 74604 70182
rect 74664 68070 74740 71542
rect 74800 70382 74876 72902
rect 81877 72902 81878 72934
rect 81942 72934 81948 72966
rect 82008 74190 82084 74196
rect 82008 74126 82014 74190
rect 82078 74126 82084 74190
rect 81942 72902 81943 72934
rect 81877 72901 81943 72902
rect 82008 71606 82084 74126
rect 82149 72830 82215 72831
rect 82149 72798 82150 72830
rect 82008 71574 82014 71606
rect 82013 71542 82014 71574
rect 82078 71574 82084 71606
rect 82144 72766 82150 72798
rect 82214 72798 82215 72830
rect 82214 72766 82220 72798
rect 82078 71542 82079 71574
rect 82013 71541 82079 71542
rect 82013 71470 82079 71471
rect 82013 71438 82014 71470
rect 74800 70318 74806 70382
rect 74870 70318 74876 70382
rect 74800 70312 74876 70318
rect 82008 71406 82014 71438
rect 82078 71438 82079 71470
rect 82078 71406 82084 71438
rect 82008 68750 82084 71406
rect 82144 70110 82220 72766
rect 94656 72558 95004 74262
rect 94656 72494 94662 72558
rect 94726 72494 95004 72558
rect 94117 71470 94183 71471
rect 94117 71438 94118 71470
rect 94112 71406 94118 71438
rect 94182 71438 94183 71470
rect 94182 71406 94188 71438
rect 94112 71062 94188 71406
rect 94112 70998 94118 71062
rect 94182 70998 94188 71062
rect 94112 70992 94188 70998
rect 82144 70046 82150 70110
rect 82214 70046 82220 70110
rect 82144 70040 82220 70046
rect 94656 70926 95004 72494
rect 94656 70862 94662 70926
rect 94726 70862 95004 70926
rect 92485 69974 92551 69975
rect 92485 69942 92486 69974
rect 82008 68686 82014 68750
rect 82078 68686 82084 68750
rect 82008 68680 82084 68686
rect 92480 69910 92486 69942
rect 92550 69942 92551 69974
rect 92550 69910 92556 69942
rect 74664 68038 74670 68070
rect 74669 68006 74670 68038
rect 74734 68038 74740 68070
rect 74734 68006 74735 68038
rect 74669 68005 74735 68006
rect 74528 67358 74534 67390
rect 73848 67320 73924 67326
rect 74533 67326 74534 67358
rect 74598 67358 74604 67390
rect 74598 67326 74599 67358
rect 74533 67325 74599 67326
rect 20944 67254 21020 67260
rect 20944 67190 20950 67254
rect 21014 67190 21020 67254
rect 20400 66982 20476 66988
rect 20400 66918 20406 66982
rect 20470 66918 20476 66982
rect 20944 66982 21020 67190
rect 20944 66950 20950 66982
rect 20400 66710 20476 66918
rect 20949 66918 20950 66950
rect 21014 66950 21020 66982
rect 21080 67254 21156 67260
rect 21080 67190 21086 67254
rect 21150 67190 21156 67254
rect 21357 67254 21423 67255
rect 21357 67222 21358 67254
rect 21080 66982 21156 67190
rect 21080 66950 21086 66982
rect 21014 66918 21015 66950
rect 20949 66917 21015 66918
rect 21085 66918 21086 66950
rect 21150 66950 21156 66982
rect 21352 67190 21358 67222
rect 21422 67222 21423 67254
rect 21765 67254 21831 67255
rect 21765 67222 21766 67254
rect 21422 67190 21428 67222
rect 21352 66982 21428 67190
rect 21150 66918 21151 66950
rect 21085 66917 21151 66918
rect 21352 66918 21358 66982
rect 21422 66918 21428 66982
rect 21352 66912 21428 66918
rect 21760 67190 21766 67222
rect 21830 67222 21831 67254
rect 22037 67254 22103 67255
rect 22037 67222 22038 67254
rect 21830 67190 21836 67222
rect 21760 66982 21836 67190
rect 21760 66918 21766 66982
rect 21830 66918 21836 66982
rect 21760 66912 21836 66918
rect 22032 67190 22038 67222
rect 22102 67222 22103 67254
rect 73989 67254 74055 67255
rect 73989 67222 73990 67254
rect 22102 67190 22108 67222
rect 22032 66982 22108 67190
rect 73984 67190 73990 67222
rect 74054 67222 74055 67254
rect 74392 67254 74468 67260
rect 74054 67190 74060 67222
rect 22032 66918 22038 66982
rect 22102 66918 22108 66982
rect 22032 66912 22108 66918
rect 27200 67118 27276 67124
rect 27200 67054 27206 67118
rect 27270 67054 27276 67118
rect 20400 66678 20406 66710
rect 20405 66646 20406 66678
rect 20470 66678 20476 66710
rect 21624 66846 21700 66852
rect 21624 66782 21630 66846
rect 21694 66782 21700 66846
rect 20470 66646 20471 66678
rect 20405 66645 20471 66646
rect 21624 66574 21700 66782
rect 21624 66542 21630 66574
rect 21629 66510 21630 66542
rect 21694 66542 21700 66574
rect 22032 66846 22108 66852
rect 22032 66782 22038 66846
rect 22102 66782 22108 66846
rect 27200 66846 27276 67054
rect 27200 66814 27206 66846
rect 22032 66574 22108 66782
rect 27205 66782 27206 66814
rect 27270 66814 27276 66846
rect 69088 67118 69164 67124
rect 69088 67054 69094 67118
rect 69158 67054 69164 67118
rect 69088 66846 69164 67054
rect 73984 66982 74060 67190
rect 73984 66918 73990 66982
rect 74054 66918 74060 66982
rect 74392 67190 74398 67254
rect 74462 67190 74468 67254
rect 74669 67254 74735 67255
rect 74669 67222 74670 67254
rect 74392 66982 74468 67190
rect 74392 66950 74398 66982
rect 73984 66912 74060 66918
rect 74397 66918 74398 66950
rect 74462 66950 74468 66982
rect 74664 67190 74670 67222
rect 74734 67222 74735 67254
rect 92480 67254 92556 69910
rect 93424 69662 93490 69663
rect 93424 69598 93425 69662
rect 93489 69598 93490 69662
rect 93424 69597 93490 69598
rect 74734 67190 74740 67222
rect 74664 66982 74740 67190
rect 92480 67190 92486 67254
rect 92550 67190 92556 67254
rect 92480 67184 92556 67190
rect 92480 67118 92692 67124
rect 92480 67054 92622 67118
rect 92686 67054 92692 67118
rect 92480 67048 92692 67054
rect 74462 66918 74463 66950
rect 74397 66917 74463 66918
rect 74664 66918 74670 66982
rect 74734 66918 74740 66982
rect 74664 66912 74740 66918
rect 75616 66982 75692 66988
rect 75616 66918 75622 66982
rect 75686 66918 75692 66982
rect 69088 66814 69094 66846
rect 27270 66782 27271 66814
rect 27205 66781 27271 66782
rect 69093 66782 69094 66814
rect 69158 66814 69164 66846
rect 73989 66846 74055 66847
rect 73989 66814 73990 66846
rect 69158 66782 69159 66814
rect 69093 66781 69159 66782
rect 73984 66782 73990 66814
rect 74054 66814 74055 66846
rect 74256 66846 74332 66852
rect 74054 66782 74060 66814
rect 22032 66542 22038 66574
rect 21694 66510 21695 66542
rect 21629 66509 21695 66510
rect 22037 66510 22038 66542
rect 22102 66542 22108 66574
rect 69088 66574 69164 66580
rect 22102 66510 22103 66542
rect 22037 66509 22103 66510
rect 69088 66510 69094 66574
rect 69158 66510 69164 66574
rect 68952 66302 69028 66308
rect 68952 66238 68958 66302
rect 69022 66238 69028 66302
rect 69088 66302 69164 66510
rect 73984 66574 74060 66782
rect 73984 66510 73990 66574
rect 74054 66510 74060 66574
rect 74256 66782 74262 66846
rect 74326 66782 74332 66846
rect 74256 66574 74332 66782
rect 75616 66710 75692 66918
rect 75616 66678 75622 66710
rect 75621 66646 75622 66678
rect 75686 66678 75692 66710
rect 75686 66646 75687 66678
rect 75621 66645 75687 66646
rect 74256 66542 74262 66574
rect 73984 66504 74060 66510
rect 74261 66510 74262 66542
rect 74326 66542 74332 66574
rect 74326 66510 74327 66542
rect 74261 66509 74327 66510
rect 69088 66270 69094 66302
rect 952 65966 1230 66030
rect 1294 65966 1300 66030
rect 952 64126 1300 65966
rect 20536 66166 20612 66172
rect 20536 66102 20542 66166
rect 20606 66102 20612 66166
rect 20536 65894 20612 66102
rect 68952 66030 69028 66238
rect 69093 66238 69094 66270
rect 69158 66270 69164 66302
rect 75072 66438 75148 66444
rect 75072 66374 75078 66438
rect 75142 66374 75148 66438
rect 69158 66238 69159 66270
rect 69093 66237 69159 66238
rect 75072 66166 75148 66374
rect 75072 66134 75078 66166
rect 75077 66102 75078 66134
rect 75142 66134 75148 66166
rect 75480 66166 75556 66172
rect 75142 66102 75143 66134
rect 75077 66101 75143 66102
rect 75480 66102 75486 66166
rect 75550 66102 75556 66166
rect 68952 65998 68958 66030
rect 68957 65966 68958 65998
rect 69022 65998 69028 66030
rect 69022 65966 69023 65998
rect 68957 65965 69023 65966
rect 20536 65862 20542 65894
rect 20541 65830 20542 65862
rect 20606 65862 20612 65894
rect 26933 65894 26999 65895
rect 26933 65862 26934 65894
rect 20606 65830 20607 65862
rect 20541 65829 20607 65830
rect 26928 65830 26934 65862
rect 26998 65862 26999 65894
rect 68957 65894 69023 65895
rect 68957 65862 68958 65894
rect 26998 65830 27004 65862
rect 20400 65758 20476 65764
rect 20400 65694 20406 65758
rect 20470 65694 20476 65758
rect 20400 65486 20476 65694
rect 20400 65454 20406 65486
rect 20405 65422 20406 65454
rect 20470 65454 20476 65486
rect 20808 65758 20884 65764
rect 20808 65694 20814 65758
rect 20878 65694 20884 65758
rect 20808 65486 20884 65694
rect 26928 65622 27004 65830
rect 26928 65558 26934 65622
rect 26998 65558 27004 65622
rect 26928 65552 27004 65558
rect 68952 65830 68958 65862
rect 69022 65862 69023 65894
rect 75480 65894 75556 66102
rect 75480 65862 75486 65894
rect 69022 65830 69028 65862
rect 68952 65622 69028 65830
rect 75485 65830 75486 65862
rect 75550 65862 75556 65894
rect 75550 65830 75551 65862
rect 75485 65829 75551 65830
rect 74669 65758 74735 65759
rect 74669 65726 74670 65758
rect 68952 65558 68958 65622
rect 69022 65558 69028 65622
rect 68952 65552 69028 65558
rect 74664 65694 74670 65726
rect 74734 65726 74735 65758
rect 74936 65758 75012 65764
rect 74734 65694 74740 65726
rect 20808 65454 20814 65486
rect 20470 65422 20471 65454
rect 20405 65421 20471 65422
rect 20813 65422 20814 65454
rect 20878 65454 20884 65486
rect 27200 65486 27276 65492
rect 20878 65422 20879 65454
rect 20813 65421 20879 65422
rect 27200 65422 27206 65486
rect 27270 65422 27276 65486
rect 20400 65350 20476 65356
rect 20400 65286 20406 65350
rect 20470 65286 20476 65350
rect 20400 65078 20476 65286
rect 20400 65046 20406 65078
rect 20405 65014 20406 65046
rect 20470 65046 20476 65078
rect 21760 65350 21836 65356
rect 21760 65286 21766 65350
rect 21830 65286 21836 65350
rect 21760 65078 21836 65286
rect 21760 65046 21766 65078
rect 20470 65014 20471 65046
rect 20405 65013 20471 65014
rect 21765 65014 21766 65046
rect 21830 65046 21836 65078
rect 22032 65350 22108 65356
rect 22032 65286 22038 65350
rect 22102 65286 22108 65350
rect 22032 65078 22108 65286
rect 27200 65214 27276 65422
rect 74664 65486 74740 65694
rect 74664 65422 74670 65486
rect 74734 65422 74740 65486
rect 74936 65694 74942 65758
rect 75006 65694 75012 65758
rect 75485 65758 75551 65759
rect 75485 65726 75486 65758
rect 74936 65486 75012 65694
rect 74936 65454 74942 65486
rect 74664 65416 74740 65422
rect 74941 65422 74942 65454
rect 75006 65454 75012 65486
rect 75480 65694 75486 65726
rect 75550 65726 75551 65758
rect 75550 65694 75556 65726
rect 75480 65486 75556 65694
rect 75006 65422 75007 65454
rect 74941 65421 75007 65422
rect 75480 65422 75486 65486
rect 75550 65422 75556 65486
rect 75480 65416 75556 65422
rect 73853 65350 73919 65351
rect 73853 65318 73854 65350
rect 27200 65182 27206 65214
rect 27205 65150 27206 65182
rect 27270 65182 27276 65214
rect 73848 65286 73854 65318
rect 73918 65318 73919 65350
rect 74256 65350 74332 65356
rect 73918 65286 73924 65318
rect 27270 65150 27271 65182
rect 27205 65149 27271 65150
rect 22032 65046 22038 65078
rect 21830 65014 21831 65046
rect 21765 65013 21831 65014
rect 22037 65014 22038 65046
rect 22102 65046 22108 65078
rect 73848 65078 73924 65286
rect 22102 65014 22103 65046
rect 22037 65013 22103 65014
rect 73848 65014 73854 65078
rect 73918 65014 73924 65078
rect 74256 65286 74262 65350
rect 74326 65286 74332 65350
rect 75621 65350 75687 65351
rect 75621 65318 75622 65350
rect 74256 65078 74332 65286
rect 74256 65046 74262 65078
rect 73848 65008 73924 65014
rect 74261 65014 74262 65046
rect 74326 65046 74332 65078
rect 75616 65286 75622 65318
rect 75686 65318 75687 65350
rect 75686 65286 75692 65318
rect 75616 65078 75692 65286
rect 74326 65014 74327 65046
rect 74261 65013 74327 65014
rect 75616 65014 75622 65078
rect 75686 65014 75692 65078
rect 75616 65008 75692 65014
rect 20405 64942 20471 64943
rect 20405 64910 20406 64942
rect 20400 64878 20406 64910
rect 20470 64910 20471 64942
rect 21488 64942 21564 64948
rect 20470 64878 20476 64910
rect 20400 64670 20476 64878
rect 20400 64606 20406 64670
rect 20470 64606 20476 64670
rect 21488 64878 21494 64942
rect 21558 64878 21564 64942
rect 21765 64942 21831 64943
rect 21765 64910 21766 64942
rect 21488 64670 21564 64878
rect 21488 64638 21494 64670
rect 20400 64600 20476 64606
rect 21493 64606 21494 64638
rect 21558 64638 21564 64670
rect 21760 64878 21766 64910
rect 21830 64910 21831 64942
rect 22037 64942 22103 64943
rect 22037 64910 22038 64942
rect 21830 64878 21836 64910
rect 21760 64670 21836 64878
rect 21558 64606 21559 64638
rect 21493 64605 21559 64606
rect 21760 64606 21766 64670
rect 21830 64606 21836 64670
rect 21760 64600 21836 64606
rect 22032 64878 22038 64910
rect 22102 64910 22103 64942
rect 73984 64942 74060 64948
rect 22102 64878 22108 64910
rect 22032 64670 22108 64878
rect 22032 64606 22038 64670
rect 22102 64606 22108 64670
rect 73984 64878 73990 64942
rect 74054 64878 74060 64942
rect 74261 64942 74327 64943
rect 74261 64910 74262 64942
rect 73984 64670 74060 64878
rect 73984 64638 73990 64670
rect 22032 64600 22108 64606
rect 73989 64606 73990 64638
rect 74054 64638 74060 64670
rect 74256 64878 74262 64910
rect 74326 64910 74327 64942
rect 75077 64942 75143 64943
rect 75077 64910 75078 64942
rect 74326 64878 74332 64910
rect 74256 64670 74332 64878
rect 74054 64606 74055 64638
rect 73989 64605 74055 64606
rect 74256 64606 74262 64670
rect 74326 64606 74332 64670
rect 74256 64600 74332 64606
rect 75072 64878 75078 64910
rect 75142 64910 75143 64942
rect 75485 64942 75551 64943
rect 75485 64910 75486 64942
rect 75142 64878 75148 64910
rect 75072 64670 75148 64878
rect 75072 64606 75078 64670
rect 75142 64606 75148 64670
rect 75072 64600 75148 64606
rect 75480 64878 75486 64910
rect 75550 64910 75551 64942
rect 75550 64878 75556 64910
rect 75480 64670 75556 64878
rect 75480 64606 75486 64670
rect 75550 64606 75556 64670
rect 75480 64600 75556 64606
rect 20536 64534 20612 64540
rect 20536 64470 20542 64534
rect 20606 64470 20612 64534
rect 20813 64534 20879 64535
rect 20813 64502 20814 64534
rect 20536 64262 20612 64470
rect 20536 64230 20542 64262
rect 20541 64198 20542 64230
rect 20606 64230 20612 64262
rect 20808 64470 20814 64502
rect 20878 64502 20879 64534
rect 21488 64534 21564 64540
rect 20878 64470 20884 64502
rect 20808 64262 20884 64470
rect 20606 64198 20607 64230
rect 20541 64197 20607 64198
rect 20808 64198 20814 64262
rect 20878 64198 20884 64262
rect 21488 64470 21494 64534
rect 21558 64470 21564 64534
rect 21488 64262 21564 64470
rect 21488 64230 21494 64262
rect 20808 64192 20884 64198
rect 21493 64198 21494 64230
rect 21558 64230 21564 64262
rect 21624 64534 21700 64540
rect 21624 64470 21630 64534
rect 21694 64470 21700 64534
rect 22037 64534 22103 64535
rect 22037 64502 22038 64534
rect 21624 64262 21700 64470
rect 21624 64230 21630 64262
rect 21558 64198 21559 64230
rect 21493 64197 21559 64198
rect 21629 64198 21630 64230
rect 21694 64230 21700 64262
rect 22032 64470 22038 64502
rect 22102 64502 22103 64534
rect 73853 64534 73919 64535
rect 73853 64502 73854 64534
rect 22102 64470 22108 64502
rect 22032 64262 22108 64470
rect 21694 64198 21695 64230
rect 21629 64197 21695 64198
rect 22032 64198 22038 64262
rect 22102 64198 22108 64262
rect 22032 64192 22108 64198
rect 73848 64470 73854 64502
rect 73918 64502 73919 64534
rect 74392 64534 74468 64540
rect 73918 64470 73924 64502
rect 73848 64262 73924 64470
rect 73848 64198 73854 64262
rect 73918 64198 73924 64262
rect 74392 64470 74398 64534
rect 74462 64470 74468 64534
rect 74392 64262 74468 64470
rect 74392 64230 74398 64262
rect 73848 64192 73924 64198
rect 74397 64198 74398 64230
rect 74462 64230 74468 64262
rect 74800 64534 74876 64540
rect 74800 64470 74806 64534
rect 74870 64470 74876 64534
rect 74800 64262 74876 64470
rect 74800 64230 74806 64262
rect 74462 64198 74463 64230
rect 74397 64197 74463 64198
rect 74805 64198 74806 64230
rect 74870 64230 74876 64262
rect 75616 64534 75692 64540
rect 75616 64470 75622 64534
rect 75686 64470 75692 64534
rect 92480 64534 92556 67048
rect 92480 64502 92486 64534
rect 75616 64262 75692 64470
rect 92485 64470 92486 64502
rect 92550 64502 92556 64534
rect 92550 64470 92551 64502
rect 92485 64469 92551 64470
rect 75616 64230 75622 64262
rect 74870 64198 74871 64230
rect 74805 64197 74871 64198
rect 75621 64198 75622 64230
rect 75686 64230 75692 64262
rect 75686 64198 75687 64230
rect 75621 64197 75687 64198
rect 952 64062 1230 64126
rect 1294 64062 1300 64126
rect 952 62494 1300 64062
rect 20536 64126 20612 64132
rect 20536 64062 20542 64126
rect 20606 64062 20612 64126
rect 20536 63854 20612 64062
rect 20536 63822 20542 63854
rect 20541 63790 20542 63822
rect 20606 63822 20612 63854
rect 20944 64126 21020 64132
rect 20944 64062 20950 64126
rect 21014 64062 21020 64126
rect 20944 63854 21020 64062
rect 20944 63822 20950 63854
rect 20606 63790 20607 63822
rect 20541 63789 20607 63790
rect 20949 63790 20950 63822
rect 21014 63822 21020 63854
rect 21080 64126 21156 64132
rect 21080 64062 21086 64126
rect 21150 64062 21156 64126
rect 21221 64126 21287 64127
rect 21221 64094 21222 64126
rect 21080 63854 21156 64062
rect 21080 63822 21086 63854
rect 21014 63790 21015 63822
rect 20949 63789 21015 63790
rect 21085 63790 21086 63822
rect 21150 63822 21156 63854
rect 21216 64062 21222 64094
rect 21286 64094 21287 64126
rect 21760 64126 21836 64132
rect 21286 64062 21292 64094
rect 21216 63854 21292 64062
rect 21150 63790 21151 63822
rect 21085 63789 21151 63790
rect 21216 63790 21222 63854
rect 21286 63790 21292 63854
rect 21760 64062 21766 64126
rect 21830 64062 21836 64126
rect 21760 63854 21836 64062
rect 21760 63822 21766 63854
rect 21216 63784 21292 63790
rect 21765 63790 21766 63822
rect 21830 63822 21836 63854
rect 22032 64126 22108 64132
rect 22032 64062 22038 64126
rect 22102 64062 22108 64126
rect 22032 63854 22108 64062
rect 22032 63822 22038 63854
rect 21830 63790 21831 63822
rect 21765 63789 21831 63790
rect 22037 63790 22038 63822
rect 22102 63822 22108 63854
rect 73984 64126 74060 64132
rect 73984 64062 73990 64126
rect 74054 64062 74060 64126
rect 74397 64126 74463 64127
rect 74397 64094 74398 64126
rect 73984 63854 74060 64062
rect 73984 63822 73990 63854
rect 22102 63790 22103 63822
rect 22037 63789 22103 63790
rect 73989 63790 73990 63822
rect 74054 63822 74060 63854
rect 74392 64062 74398 64094
rect 74462 64094 74463 64126
rect 75621 64126 75687 64127
rect 75621 64094 75622 64126
rect 74462 64062 74468 64094
rect 74392 63854 74468 64062
rect 74054 63790 74055 63822
rect 73989 63789 74055 63790
rect 74392 63790 74398 63854
rect 74462 63790 74468 63854
rect 74392 63784 74468 63790
rect 75616 64062 75622 64094
rect 75686 64094 75687 64126
rect 75686 64062 75692 64094
rect 75616 63854 75692 64062
rect 75616 63790 75622 63854
rect 75686 63790 75692 63854
rect 75616 63784 75692 63790
rect 20541 63718 20607 63719
rect 20541 63686 20542 63718
rect 20536 63654 20542 63686
rect 20606 63686 20607 63718
rect 20808 63718 20884 63724
rect 20606 63654 20612 63686
rect 20536 63446 20612 63654
rect 20536 63382 20542 63446
rect 20606 63382 20612 63446
rect 20808 63654 20814 63718
rect 20878 63654 20884 63718
rect 21765 63718 21831 63719
rect 21765 63686 21766 63718
rect 20808 63446 20884 63654
rect 20808 63414 20814 63446
rect 20536 63376 20612 63382
rect 20813 63382 20814 63414
rect 20878 63414 20884 63446
rect 21760 63654 21766 63686
rect 21830 63686 21831 63718
rect 22037 63718 22103 63719
rect 22037 63686 22038 63718
rect 21830 63654 21836 63686
rect 21760 63446 21836 63654
rect 20878 63382 20879 63414
rect 20813 63381 20879 63382
rect 21760 63382 21766 63446
rect 21830 63382 21836 63446
rect 21760 63376 21836 63382
rect 22032 63654 22038 63686
rect 22102 63686 22103 63718
rect 73989 63718 74055 63719
rect 73989 63686 73990 63718
rect 22102 63654 22108 63686
rect 22032 63446 22108 63654
rect 22032 63382 22038 63446
rect 22102 63382 22108 63446
rect 22032 63376 22108 63382
rect 73984 63654 73990 63686
rect 74054 63686 74055 63718
rect 74261 63718 74327 63719
rect 74261 63686 74262 63718
rect 74054 63654 74060 63686
rect 73984 63446 74060 63654
rect 73984 63382 73990 63446
rect 74054 63382 74060 63446
rect 73984 63376 74060 63382
rect 74256 63654 74262 63686
rect 74326 63686 74327 63718
rect 74936 63718 75012 63724
rect 74326 63654 74332 63686
rect 74256 63446 74332 63654
rect 74256 63382 74262 63446
rect 74326 63382 74332 63446
rect 74936 63654 74942 63718
rect 75006 63654 75012 63718
rect 74936 63446 75012 63654
rect 74936 63414 74942 63446
rect 74256 63376 74332 63382
rect 74941 63382 74942 63414
rect 75006 63414 75012 63446
rect 75616 63718 75692 63724
rect 75616 63654 75622 63718
rect 75686 63654 75692 63718
rect 75616 63446 75692 63654
rect 75616 63414 75622 63446
rect 75006 63382 75007 63414
rect 74941 63381 75007 63382
rect 75621 63382 75622 63414
rect 75686 63414 75692 63446
rect 75686 63382 75687 63414
rect 75621 63381 75687 63382
rect 20813 63310 20879 63311
rect 20813 63278 20814 63310
rect 20808 63246 20814 63278
rect 20878 63278 20879 63310
rect 21493 63310 21559 63311
rect 21493 63278 21494 63310
rect 20878 63246 20884 63278
rect 20808 63038 20884 63246
rect 20808 62974 20814 63038
rect 20878 62974 20884 63038
rect 20808 62968 20884 62974
rect 21488 63246 21494 63278
rect 21558 63278 21559 63310
rect 21624 63310 21700 63316
rect 21558 63246 21564 63278
rect 21488 63038 21564 63246
rect 21488 62974 21494 63038
rect 21558 62974 21564 63038
rect 21624 63246 21630 63310
rect 21694 63246 21700 63310
rect 21624 63038 21700 63246
rect 21624 63006 21630 63038
rect 21488 62968 21564 62974
rect 21629 62974 21630 63006
rect 21694 63006 21700 63038
rect 22168 63310 22244 63316
rect 22168 63246 22174 63310
rect 22238 63246 22244 63310
rect 73853 63310 73919 63311
rect 73853 63278 73854 63310
rect 22168 63038 22244 63246
rect 73848 63246 73854 63278
rect 73918 63278 73919 63310
rect 74392 63310 74468 63316
rect 73918 63246 73924 63278
rect 27205 63174 27271 63175
rect 27205 63142 27206 63174
rect 22168 63006 22174 63038
rect 21694 62974 21695 63006
rect 21629 62973 21695 62974
rect 22173 62974 22174 63006
rect 22238 63006 22244 63038
rect 27200 63110 27206 63142
rect 27270 63142 27271 63174
rect 27270 63110 27276 63142
rect 22238 62974 22239 63006
rect 22173 62973 22239 62974
rect 21765 62902 21831 62903
rect 21765 62870 21766 62902
rect 21760 62838 21766 62870
rect 21830 62870 21831 62902
rect 22168 62902 22244 62908
rect 21830 62838 21836 62870
rect 21760 62630 21836 62838
rect 21760 62566 21766 62630
rect 21830 62566 21836 62630
rect 22168 62838 22174 62902
rect 22238 62838 22244 62902
rect 22168 62630 22244 62838
rect 22168 62598 22174 62630
rect 21760 62560 21836 62566
rect 22173 62566 22174 62598
rect 22238 62598 22244 62630
rect 27064 62902 27140 62908
rect 27064 62838 27070 62902
rect 27134 62838 27140 62902
rect 22238 62566 22239 62598
rect 22173 62565 22239 62566
rect 952 62430 1230 62494
rect 1294 62430 1300 62494
rect 952 60862 1300 62430
rect 20808 62494 20884 62500
rect 20808 62430 20814 62494
rect 20878 62430 20884 62494
rect 20536 62222 20612 62228
rect 20536 62158 20542 62222
rect 20606 62158 20612 62222
rect 20808 62222 20884 62430
rect 20808 62190 20814 62222
rect 20536 61950 20612 62158
rect 20813 62158 20814 62190
rect 20878 62190 20884 62222
rect 26928 62358 27004 62364
rect 26928 62294 26934 62358
rect 26998 62294 27004 62358
rect 27064 62358 27140 62838
rect 27200 62902 27276 63110
rect 73848 63038 73924 63246
rect 73848 62974 73854 63038
rect 73918 62974 73924 63038
rect 74392 63246 74398 63310
rect 74462 63246 74468 63310
rect 74392 63038 74468 63246
rect 74392 63006 74398 63038
rect 73848 62968 73924 62974
rect 74397 62974 74398 63006
rect 74462 63006 74468 63038
rect 74800 63310 74876 63316
rect 74800 63246 74806 63310
rect 74870 63246 74876 63310
rect 74800 63038 74876 63246
rect 74800 63006 74806 63038
rect 74462 62974 74463 63006
rect 74397 62973 74463 62974
rect 74805 62974 74806 63006
rect 74870 63006 74876 63038
rect 75208 63310 75284 63316
rect 75208 63246 75214 63310
rect 75278 63246 75284 63310
rect 75208 63038 75284 63246
rect 75208 63006 75214 63038
rect 74870 62974 74871 63006
rect 74805 62973 74871 62974
rect 75213 62974 75214 63006
rect 75278 63006 75284 63038
rect 75278 62974 75279 63006
rect 75213 62973 75279 62974
rect 27200 62838 27206 62902
rect 27270 62838 27276 62902
rect 27200 62832 27276 62838
rect 73984 62902 74060 62908
rect 73984 62838 73990 62902
rect 74054 62838 74060 62902
rect 73984 62630 74060 62838
rect 73984 62598 73990 62630
rect 73989 62566 73990 62598
rect 74054 62598 74060 62630
rect 74392 62902 74468 62908
rect 74392 62838 74398 62902
rect 74462 62838 74468 62902
rect 74392 62630 74468 62838
rect 74392 62598 74398 62630
rect 74054 62566 74055 62598
rect 73989 62565 74055 62566
rect 74397 62566 74398 62598
rect 74462 62598 74468 62630
rect 74462 62566 74463 62598
rect 74397 62565 74463 62566
rect 27064 62326 27070 62358
rect 20878 62158 20879 62190
rect 20813 62157 20879 62158
rect 26928 62086 27004 62294
rect 27069 62294 27070 62326
rect 27134 62326 27140 62358
rect 74936 62494 75012 62500
rect 74936 62430 74942 62494
rect 75006 62430 75012 62494
rect 27134 62294 27135 62326
rect 27069 62293 27135 62294
rect 74936 62222 75012 62430
rect 74936 62190 74942 62222
rect 74941 62158 74942 62190
rect 75006 62190 75012 62222
rect 75621 62222 75687 62223
rect 75621 62190 75622 62222
rect 75006 62158 75007 62190
rect 74941 62157 75007 62158
rect 75616 62158 75622 62190
rect 75686 62190 75687 62222
rect 75686 62158 75692 62190
rect 26928 62054 26934 62086
rect 26933 62022 26934 62054
rect 26998 62054 27004 62086
rect 26998 62022 26999 62054
rect 26933 62021 26999 62022
rect 20536 61918 20542 61950
rect 20541 61886 20542 61918
rect 20606 61918 20612 61950
rect 26933 61950 26999 61951
rect 26933 61918 26934 61950
rect 20606 61886 20607 61918
rect 20541 61885 20607 61886
rect 26928 61886 26934 61918
rect 26998 61918 26999 61950
rect 68952 61950 69028 61956
rect 26998 61886 27004 61918
rect 20405 61814 20471 61815
rect 20405 61782 20406 61814
rect 20400 61750 20406 61782
rect 20470 61782 20471 61814
rect 20949 61814 21015 61815
rect 20949 61782 20950 61814
rect 20470 61750 20476 61782
rect 20400 61542 20476 61750
rect 20400 61478 20406 61542
rect 20470 61478 20476 61542
rect 20400 61472 20476 61478
rect 20944 61750 20950 61782
rect 21014 61782 21015 61814
rect 21085 61814 21151 61815
rect 21085 61782 21086 61814
rect 21014 61750 21020 61782
rect 20944 61542 21020 61750
rect 20944 61478 20950 61542
rect 21014 61478 21020 61542
rect 20944 61472 21020 61478
rect 21080 61750 21086 61782
rect 21150 61782 21151 61814
rect 21150 61750 21156 61782
rect 21080 61542 21156 61750
rect 26928 61678 27004 61886
rect 26928 61614 26934 61678
rect 26998 61614 27004 61678
rect 68952 61886 68958 61950
rect 69022 61886 69028 61950
rect 68952 61678 69028 61886
rect 75616 61950 75692 62158
rect 75616 61886 75622 61950
rect 75686 61886 75692 61950
rect 75616 61880 75692 61886
rect 74669 61814 74735 61815
rect 74669 61782 74670 61814
rect 68952 61646 68958 61678
rect 26928 61608 27004 61614
rect 68957 61614 68958 61646
rect 69022 61646 69028 61678
rect 74664 61750 74670 61782
rect 74734 61782 74735 61814
rect 75072 61814 75148 61820
rect 74734 61750 74740 61782
rect 69022 61614 69023 61646
rect 68957 61613 69023 61614
rect 21080 61478 21086 61542
rect 21150 61478 21156 61542
rect 21080 61472 21156 61478
rect 27200 61542 27276 61548
rect 27200 61478 27206 61542
rect 27270 61478 27276 61542
rect 20541 61406 20607 61407
rect 20541 61374 20542 61406
rect 20536 61342 20542 61374
rect 20606 61374 20607 61406
rect 21624 61406 21700 61412
rect 20606 61342 20612 61374
rect 20536 61134 20612 61342
rect 20536 61070 20542 61134
rect 20606 61070 20612 61134
rect 21624 61342 21630 61406
rect 21694 61342 21700 61406
rect 21624 61134 21700 61342
rect 21624 61102 21630 61134
rect 20536 61064 20612 61070
rect 21629 61070 21630 61102
rect 21694 61102 21700 61134
rect 22032 61406 22108 61412
rect 22032 61342 22038 61406
rect 22102 61342 22108 61406
rect 22032 61134 22108 61342
rect 27200 61270 27276 61478
rect 74664 61542 74740 61750
rect 74664 61478 74670 61542
rect 74734 61478 74740 61542
rect 75072 61750 75078 61814
rect 75142 61750 75148 61814
rect 75072 61542 75148 61750
rect 75072 61510 75078 61542
rect 74664 61472 74740 61478
rect 75077 61478 75078 61510
rect 75142 61510 75148 61542
rect 75480 61814 75556 61820
rect 75480 61750 75486 61814
rect 75550 61750 75556 61814
rect 75480 61542 75556 61750
rect 75480 61510 75486 61542
rect 75142 61478 75143 61510
rect 75077 61477 75143 61478
rect 75485 61478 75486 61510
rect 75550 61510 75556 61542
rect 91936 61542 92012 61548
rect 75550 61478 75551 61510
rect 75485 61477 75551 61478
rect 91936 61478 91942 61542
rect 92006 61478 92012 61542
rect 73989 61406 74055 61407
rect 73989 61374 73990 61406
rect 27200 61238 27206 61270
rect 27205 61206 27206 61238
rect 27270 61238 27276 61270
rect 73984 61342 73990 61374
rect 74054 61374 74055 61406
rect 74256 61406 74332 61412
rect 74054 61342 74060 61374
rect 27270 61206 27271 61238
rect 27205 61205 27271 61206
rect 22032 61102 22038 61134
rect 21694 61070 21695 61102
rect 21629 61069 21695 61070
rect 22037 61070 22038 61102
rect 22102 61102 22108 61134
rect 73984 61134 74060 61342
rect 22102 61070 22103 61102
rect 22037 61069 22103 61070
rect 73984 61070 73990 61134
rect 74054 61070 74060 61134
rect 74256 61342 74262 61406
rect 74326 61342 74332 61406
rect 74256 61134 74332 61342
rect 74256 61102 74262 61134
rect 73984 61064 74060 61070
rect 74261 61070 74262 61102
rect 74326 61102 74332 61134
rect 75616 61406 75692 61412
rect 75616 61342 75622 61406
rect 75686 61342 75692 61406
rect 75616 61134 75692 61342
rect 75616 61102 75622 61134
rect 74326 61070 74327 61102
rect 74261 61069 74327 61070
rect 75621 61070 75622 61102
rect 75686 61102 75692 61134
rect 75686 61070 75687 61102
rect 75621 61069 75687 61070
rect 20405 60998 20471 60999
rect 20405 60966 20406 60998
rect 952 60798 1230 60862
rect 1294 60798 1300 60862
rect 952 59230 1300 60798
rect 20400 60934 20406 60966
rect 20470 60966 20471 60998
rect 21080 60998 21156 61004
rect 20470 60934 20476 60966
rect 20400 60726 20476 60934
rect 20400 60662 20406 60726
rect 20470 60662 20476 60726
rect 21080 60934 21086 60998
rect 21150 60934 21156 60998
rect 21080 60726 21156 60934
rect 21080 60694 21086 60726
rect 20400 60656 20476 60662
rect 21085 60662 21086 60694
rect 21150 60694 21156 60726
rect 21352 60998 21428 61004
rect 21352 60934 21358 60998
rect 21422 60934 21428 60998
rect 21629 60998 21695 60999
rect 21629 60966 21630 60998
rect 21352 60726 21428 60934
rect 21352 60694 21358 60726
rect 21150 60662 21151 60694
rect 21085 60661 21151 60662
rect 21357 60662 21358 60694
rect 21422 60694 21428 60726
rect 21624 60934 21630 60966
rect 21694 60966 21695 60998
rect 22032 60998 22108 61004
rect 21694 60934 21700 60966
rect 21624 60726 21700 60934
rect 21422 60662 21423 60694
rect 21357 60661 21423 60662
rect 21624 60662 21630 60726
rect 21694 60662 21700 60726
rect 22032 60934 22038 60998
rect 22102 60934 22108 60998
rect 22032 60726 22108 60934
rect 22032 60694 22038 60726
rect 21624 60656 21700 60662
rect 22037 60662 22038 60694
rect 22102 60694 22108 60726
rect 73984 60998 74060 61004
rect 73984 60934 73990 60998
rect 74054 60934 74060 60998
rect 74261 60998 74327 60999
rect 74261 60966 74262 60998
rect 73984 60726 74060 60934
rect 73984 60694 73990 60726
rect 22102 60662 22103 60694
rect 22037 60661 22103 60662
rect 73989 60662 73990 60694
rect 74054 60694 74060 60726
rect 74256 60934 74262 60966
rect 74326 60966 74327 60998
rect 75072 60998 75148 61004
rect 74326 60934 74332 60966
rect 74256 60726 74332 60934
rect 74054 60662 74055 60694
rect 73989 60661 74055 60662
rect 74256 60662 74262 60726
rect 74326 60662 74332 60726
rect 75072 60934 75078 60998
rect 75142 60934 75148 60998
rect 75621 60998 75687 60999
rect 75621 60966 75622 60998
rect 75072 60726 75148 60934
rect 75072 60694 75078 60726
rect 74256 60656 74332 60662
rect 75077 60662 75078 60694
rect 75142 60694 75148 60726
rect 75616 60934 75622 60966
rect 75686 60966 75687 60998
rect 75686 60934 75692 60966
rect 75616 60726 75692 60934
rect 75142 60662 75143 60694
rect 75077 60661 75143 60662
rect 75616 60662 75622 60726
rect 75686 60662 75692 60726
rect 75616 60656 75692 60662
rect 20536 60590 20612 60596
rect 20536 60526 20542 60590
rect 20606 60526 20612 60590
rect 20949 60590 21015 60591
rect 20949 60558 20950 60590
rect 20536 60318 20612 60526
rect 20536 60286 20542 60318
rect 20541 60254 20542 60286
rect 20606 60286 20612 60318
rect 20944 60526 20950 60558
rect 21014 60558 21015 60590
rect 21085 60590 21151 60591
rect 21085 60558 21086 60590
rect 21014 60526 21020 60558
rect 20944 60318 21020 60526
rect 20606 60254 20607 60286
rect 20541 60253 20607 60254
rect 20944 60254 20950 60318
rect 21014 60254 21020 60318
rect 20944 60248 21020 60254
rect 21080 60526 21086 60558
rect 21150 60558 21151 60590
rect 21760 60590 21836 60596
rect 21150 60526 21156 60558
rect 21080 60318 21156 60526
rect 21080 60254 21086 60318
rect 21150 60254 21156 60318
rect 21760 60526 21766 60590
rect 21830 60526 21836 60590
rect 22037 60590 22103 60591
rect 22037 60558 22038 60590
rect 21760 60318 21836 60526
rect 21760 60286 21766 60318
rect 21080 60248 21156 60254
rect 21765 60254 21766 60286
rect 21830 60286 21836 60318
rect 22032 60526 22038 60558
rect 22102 60558 22103 60590
rect 73989 60590 74055 60591
rect 73989 60558 73990 60590
rect 22102 60526 22108 60558
rect 22032 60318 22108 60526
rect 21830 60254 21831 60286
rect 21765 60253 21831 60254
rect 22032 60254 22038 60318
rect 22102 60254 22108 60318
rect 22032 60248 22108 60254
rect 73984 60526 73990 60558
rect 74054 60558 74055 60590
rect 74392 60590 74468 60596
rect 74054 60526 74060 60558
rect 73984 60318 74060 60526
rect 73984 60254 73990 60318
rect 74054 60254 74060 60318
rect 74392 60526 74398 60590
rect 74462 60526 74468 60590
rect 74669 60590 74735 60591
rect 74669 60558 74670 60590
rect 74392 60318 74468 60526
rect 74392 60286 74398 60318
rect 73984 60248 74060 60254
rect 74397 60254 74398 60286
rect 74462 60286 74468 60318
rect 74664 60526 74670 60558
rect 74734 60558 74735 60590
rect 74936 60590 75012 60596
rect 74734 60526 74740 60558
rect 74664 60318 74740 60526
rect 74462 60254 74463 60286
rect 74397 60253 74463 60254
rect 74664 60254 74670 60318
rect 74734 60254 74740 60318
rect 74936 60526 74942 60590
rect 75006 60526 75012 60590
rect 74936 60318 75012 60526
rect 74936 60286 74942 60318
rect 74664 60248 74740 60254
rect 74941 60254 74942 60286
rect 75006 60286 75012 60318
rect 75480 60590 75556 60596
rect 75480 60526 75486 60590
rect 75550 60526 75556 60590
rect 75480 60318 75556 60526
rect 75480 60286 75486 60318
rect 75006 60254 75007 60286
rect 74941 60253 75007 60254
rect 75485 60254 75486 60286
rect 75550 60286 75556 60318
rect 75550 60254 75551 60286
rect 75485 60253 75551 60254
rect 20536 60182 20612 60188
rect 20536 60118 20542 60182
rect 20606 60118 20612 60182
rect 21357 60182 21423 60183
rect 21357 60150 21358 60182
rect 20536 59910 20612 60118
rect 20536 59878 20542 59910
rect 20541 59846 20542 59878
rect 20606 59878 20612 59910
rect 21352 60118 21358 60150
rect 21422 60150 21423 60182
rect 21624 60182 21700 60188
rect 21422 60118 21428 60150
rect 21352 59910 21428 60118
rect 20606 59846 20607 59878
rect 20541 59845 20607 59846
rect 21352 59846 21358 59910
rect 21422 59846 21428 59910
rect 21624 60118 21630 60182
rect 21694 60118 21700 60182
rect 21624 59910 21700 60118
rect 21624 59878 21630 59910
rect 21352 59840 21428 59846
rect 21629 59846 21630 59878
rect 21694 59878 21700 59910
rect 22168 60182 22244 60188
rect 22168 60118 22174 60182
rect 22238 60118 22244 60182
rect 22168 59910 22244 60118
rect 22168 59878 22174 59910
rect 21694 59846 21695 59878
rect 21629 59845 21695 59846
rect 22173 59846 22174 59878
rect 22238 59878 22244 59910
rect 73848 60182 73924 60188
rect 73848 60118 73854 60182
rect 73918 60118 73924 60182
rect 74261 60182 74327 60183
rect 74261 60150 74262 60182
rect 73848 59910 73924 60118
rect 73848 59878 73854 59910
rect 22238 59846 22239 59878
rect 22173 59845 22239 59846
rect 73853 59846 73854 59878
rect 73918 59878 73924 59910
rect 74256 60118 74262 60150
rect 74326 60150 74327 60182
rect 74805 60182 74871 60183
rect 74805 60150 74806 60182
rect 74326 60118 74332 60150
rect 74256 59910 74332 60118
rect 73918 59846 73919 59878
rect 73853 59845 73919 59846
rect 74256 59846 74262 59910
rect 74326 59846 74332 59910
rect 74256 59840 74332 59846
rect 74800 60118 74806 60150
rect 74870 60150 74871 60182
rect 75616 60182 75692 60188
rect 74870 60118 74876 60150
rect 74800 59910 74876 60118
rect 74800 59846 74806 59910
rect 74870 59846 74876 59910
rect 75616 60118 75622 60182
rect 75686 60118 75692 60182
rect 75616 59910 75692 60118
rect 75616 59878 75622 59910
rect 74800 59840 74876 59846
rect 75621 59846 75622 59878
rect 75686 59878 75692 59910
rect 75686 59846 75687 59878
rect 75621 59845 75687 59846
rect 20536 59774 20612 59780
rect 20536 59710 20542 59774
rect 20606 59710 20612 59774
rect 20813 59774 20879 59775
rect 20813 59742 20814 59774
rect 20536 59502 20612 59710
rect 20536 59470 20542 59502
rect 20541 59438 20542 59470
rect 20606 59470 20612 59502
rect 20808 59710 20814 59742
rect 20878 59742 20879 59774
rect 21080 59774 21156 59780
rect 20878 59710 20884 59742
rect 20808 59502 20884 59710
rect 20606 59438 20607 59470
rect 20541 59437 20607 59438
rect 20808 59438 20814 59502
rect 20878 59438 20884 59502
rect 21080 59710 21086 59774
rect 21150 59710 21156 59774
rect 21080 59502 21156 59710
rect 21080 59470 21086 59502
rect 20808 59432 20884 59438
rect 21085 59438 21086 59470
rect 21150 59470 21156 59502
rect 21488 59774 21564 59780
rect 21488 59710 21494 59774
rect 21558 59710 21564 59774
rect 21629 59774 21695 59775
rect 21629 59742 21630 59774
rect 21488 59502 21564 59710
rect 21488 59470 21494 59502
rect 21150 59438 21151 59470
rect 21085 59437 21151 59438
rect 21493 59438 21494 59470
rect 21558 59470 21564 59502
rect 21624 59710 21630 59742
rect 21694 59742 21695 59774
rect 22032 59774 22108 59780
rect 21694 59710 21700 59742
rect 21624 59502 21700 59710
rect 21558 59438 21559 59470
rect 21493 59437 21559 59438
rect 21624 59438 21630 59502
rect 21694 59438 21700 59502
rect 22032 59710 22038 59774
rect 22102 59710 22108 59774
rect 73853 59774 73919 59775
rect 73853 59742 73854 59774
rect 22032 59502 22108 59710
rect 22032 59470 22038 59502
rect 21624 59432 21700 59438
rect 22037 59438 22038 59470
rect 22102 59470 22108 59502
rect 73848 59710 73854 59742
rect 73918 59742 73919 59774
rect 74392 59774 74468 59780
rect 73918 59710 73924 59742
rect 73848 59502 73924 59710
rect 22102 59438 22103 59470
rect 22037 59437 22103 59438
rect 73848 59438 73854 59502
rect 73918 59438 73924 59502
rect 74392 59710 74398 59774
rect 74462 59710 74468 59774
rect 74392 59502 74468 59710
rect 74392 59470 74398 59502
rect 73848 59432 73924 59438
rect 74397 59438 74398 59470
rect 74462 59470 74468 59502
rect 74664 59774 74740 59780
rect 74664 59710 74670 59774
rect 74734 59710 74740 59774
rect 75621 59774 75687 59775
rect 75621 59742 75622 59774
rect 74664 59502 74740 59710
rect 74664 59470 74670 59502
rect 74462 59438 74463 59470
rect 74397 59437 74463 59438
rect 74669 59438 74670 59470
rect 74734 59470 74740 59502
rect 75616 59710 75622 59742
rect 75686 59742 75687 59774
rect 75686 59710 75692 59742
rect 75616 59502 75692 59710
rect 74734 59438 74735 59470
rect 74669 59437 74735 59438
rect 75616 59438 75622 59502
rect 75686 59438 75692 59502
rect 75616 59432 75692 59438
rect 20949 59366 21015 59367
rect 20949 59334 20950 59366
rect 952 59166 1230 59230
rect 1294 59166 1300 59230
rect 952 57462 1300 59166
rect 20944 59302 20950 59334
rect 21014 59334 21015 59366
rect 21085 59366 21151 59367
rect 21085 59334 21086 59366
rect 21014 59302 21020 59334
rect 20944 59094 21020 59302
rect 20944 59030 20950 59094
rect 21014 59030 21020 59094
rect 20944 59024 21020 59030
rect 21080 59302 21086 59334
rect 21150 59334 21151 59366
rect 21624 59366 21700 59372
rect 21150 59302 21156 59334
rect 21080 59094 21156 59302
rect 21080 59030 21086 59094
rect 21150 59030 21156 59094
rect 21624 59302 21630 59366
rect 21694 59302 21700 59366
rect 22037 59366 22103 59367
rect 22037 59334 22038 59366
rect 21624 59094 21700 59302
rect 21624 59062 21630 59094
rect 21080 59024 21156 59030
rect 21629 59030 21630 59062
rect 21694 59062 21700 59094
rect 22032 59302 22038 59334
rect 22102 59334 22103 59366
rect 73848 59366 73924 59372
rect 22102 59302 22108 59334
rect 22032 59094 22108 59302
rect 21694 59030 21695 59062
rect 21629 59029 21695 59030
rect 22032 59030 22038 59094
rect 22102 59030 22108 59094
rect 73848 59302 73854 59366
rect 73918 59302 73924 59366
rect 74397 59366 74463 59367
rect 74397 59334 74398 59366
rect 73848 59094 73924 59302
rect 73848 59062 73854 59094
rect 22032 59024 22108 59030
rect 73853 59030 73854 59062
rect 73918 59062 73924 59094
rect 74392 59302 74398 59334
rect 74462 59334 74463 59366
rect 75077 59366 75143 59367
rect 75077 59334 75078 59366
rect 74462 59302 74468 59334
rect 74392 59094 74468 59302
rect 73918 59030 73919 59062
rect 73853 59029 73919 59030
rect 74392 59030 74398 59094
rect 74462 59030 74468 59094
rect 74392 59024 74468 59030
rect 75072 59302 75078 59334
rect 75142 59334 75143 59366
rect 75142 59302 75148 59334
rect 75072 59094 75148 59302
rect 75072 59030 75078 59094
rect 75142 59030 75148 59094
rect 75072 59024 75148 59030
rect 21624 58958 21700 58964
rect 21624 58894 21630 58958
rect 21694 58894 21700 58958
rect 21624 58686 21700 58894
rect 21624 58654 21630 58686
rect 21629 58622 21630 58654
rect 21694 58654 21700 58686
rect 22168 58958 22244 58964
rect 22168 58894 22174 58958
rect 22238 58894 22244 58958
rect 73853 58958 73919 58959
rect 73853 58926 73854 58958
rect 22168 58686 22244 58894
rect 22168 58654 22174 58686
rect 21694 58622 21695 58654
rect 21629 58621 21695 58622
rect 22173 58622 22174 58654
rect 22238 58654 22244 58686
rect 73848 58894 73854 58926
rect 73918 58926 73919 58958
rect 74261 58958 74327 58959
rect 74261 58926 74262 58958
rect 73918 58894 73924 58926
rect 73848 58686 73924 58894
rect 22238 58622 22239 58654
rect 22173 58621 22239 58622
rect 73848 58622 73854 58686
rect 73918 58622 73924 58686
rect 73848 58616 73924 58622
rect 74256 58894 74262 58926
rect 74326 58926 74327 58958
rect 74326 58894 74332 58926
rect 74256 58686 74332 58894
rect 91936 58822 92012 61478
rect 93427 59428 93487 69597
rect 94656 69294 95004 70862
rect 94656 69230 94662 69294
rect 94726 69230 95004 69294
rect 94112 69158 94188 69164
rect 94112 69094 94118 69158
rect 94182 69094 94188 69158
rect 94112 68750 94188 69094
rect 94112 68718 94118 68750
rect 94117 68686 94118 68718
rect 94182 68718 94188 68750
rect 94182 68686 94183 68718
rect 94117 68685 94183 68686
rect 94656 67662 95004 69230
rect 94656 67598 94662 67662
rect 94726 67598 95004 67662
rect 94656 66030 95004 67598
rect 94656 65966 94662 66030
rect 94726 65966 95004 66030
rect 94656 64126 95004 65966
rect 94656 64062 94662 64126
rect 94726 64062 95004 64126
rect 94117 62902 94183 62903
rect 94117 62870 94118 62902
rect 94112 62838 94118 62870
rect 94182 62870 94183 62902
rect 94182 62838 94188 62870
rect 94112 62630 94188 62838
rect 94112 62566 94118 62630
rect 94182 62566 94188 62630
rect 94112 62560 94188 62566
rect 94656 62494 95004 64062
rect 94656 62430 94662 62494
rect 94726 62430 95004 62494
rect 94112 60862 94188 60868
rect 94112 60798 94118 60862
rect 94182 60798 94188 60862
rect 94112 60318 94188 60798
rect 94112 60286 94118 60318
rect 94117 60254 94118 60286
rect 94182 60286 94188 60318
rect 94656 60862 95004 62430
rect 94656 60798 94662 60862
rect 94726 60798 95004 60862
rect 94182 60254 94183 60286
rect 94117 60253 94183 60254
rect 93424 59427 93490 59428
rect 93424 59363 93425 59427
rect 93489 59363 93490 59427
rect 93424 59362 93490 59363
rect 91936 58790 91942 58822
rect 91941 58758 91942 58790
rect 92006 58790 92012 58822
rect 94656 59094 95004 60798
rect 94656 59030 94662 59094
rect 94726 59030 95004 59094
rect 92006 58758 92007 58790
rect 91941 58757 92007 58758
rect 74256 58622 74262 58686
rect 74326 58622 74332 58686
rect 74256 58616 74332 58622
rect 20813 58550 20879 58551
rect 20813 58518 20814 58550
rect 20808 58486 20814 58518
rect 20878 58518 20879 58550
rect 21085 58550 21151 58551
rect 21085 58518 21086 58550
rect 20878 58486 20884 58518
rect 20405 58278 20471 58279
rect 20405 58246 20406 58278
rect 20400 58214 20406 58246
rect 20470 58246 20471 58278
rect 20808 58278 20884 58486
rect 20470 58214 20476 58246
rect 20400 58006 20476 58214
rect 20808 58214 20814 58278
rect 20878 58214 20884 58278
rect 20808 58208 20884 58214
rect 21080 58486 21086 58518
rect 21150 58518 21151 58550
rect 21760 58550 21836 58556
rect 21150 58486 21156 58518
rect 21080 58278 21156 58486
rect 21080 58214 21086 58278
rect 21150 58214 21156 58278
rect 21760 58486 21766 58550
rect 21830 58486 21836 58550
rect 21760 58278 21836 58486
rect 21760 58246 21766 58278
rect 21080 58208 21156 58214
rect 21765 58214 21766 58246
rect 21830 58246 21836 58278
rect 22168 58550 22244 58556
rect 22168 58486 22174 58550
rect 22238 58486 22244 58550
rect 22168 58278 22244 58486
rect 73984 58550 74060 58556
rect 73984 58486 73990 58550
rect 74054 58486 74060 58550
rect 22168 58246 22174 58278
rect 21830 58214 21831 58246
rect 21765 58213 21831 58214
rect 22173 58214 22174 58246
rect 22238 58246 22244 58278
rect 26928 58414 27004 58420
rect 26928 58350 26934 58414
rect 26998 58350 27004 58414
rect 68957 58414 69023 58415
rect 68957 58382 68958 58414
rect 22238 58214 22239 58246
rect 22173 58213 22239 58214
rect 26928 58142 27004 58350
rect 68952 58350 68958 58382
rect 69022 58382 69023 58414
rect 69022 58350 69028 58382
rect 26928 58110 26934 58142
rect 26933 58078 26934 58110
rect 26998 58110 27004 58142
rect 27205 58142 27271 58143
rect 27205 58110 27206 58142
rect 26998 58078 26999 58110
rect 26933 58077 26999 58078
rect 27200 58078 27206 58110
rect 27270 58110 27271 58142
rect 68952 58142 69028 58350
rect 73984 58278 74060 58486
rect 73984 58246 73990 58278
rect 73989 58214 73990 58246
rect 74054 58246 74060 58278
rect 74392 58550 74468 58556
rect 74392 58486 74398 58550
rect 74462 58486 74468 58550
rect 74392 58278 74468 58486
rect 74392 58246 74398 58278
rect 74054 58214 74055 58246
rect 73989 58213 74055 58214
rect 74397 58214 74398 58246
rect 74462 58246 74468 58278
rect 74664 58550 74740 58556
rect 74664 58486 74670 58550
rect 74734 58486 74740 58550
rect 74664 58278 74740 58486
rect 74664 58246 74670 58278
rect 74462 58214 74463 58246
rect 74397 58213 74463 58214
rect 74669 58214 74670 58246
rect 74734 58246 74740 58278
rect 75616 58278 75692 58284
rect 74734 58214 74735 58246
rect 74669 58213 74735 58214
rect 75616 58214 75622 58278
rect 75686 58214 75692 58278
rect 27270 58078 27276 58110
rect 20400 57942 20406 58006
rect 20470 57942 20476 58006
rect 20400 57936 20476 57942
rect 20536 57870 20612 57876
rect 20536 57806 20542 57870
rect 20606 57806 20612 57870
rect 20813 57870 20879 57871
rect 20813 57838 20814 57870
rect 20536 57598 20612 57806
rect 20536 57566 20542 57598
rect 20541 57534 20542 57566
rect 20606 57566 20612 57598
rect 20808 57806 20814 57838
rect 20878 57838 20879 57870
rect 20878 57806 20884 57838
rect 20808 57598 20884 57806
rect 27200 57734 27276 58078
rect 68952 58078 68958 58142
rect 69022 58078 69028 58142
rect 68952 58072 69028 58078
rect 74936 58142 75012 58148
rect 74936 58078 74942 58142
rect 75006 58078 75012 58142
rect 27200 57670 27206 57734
rect 27270 57670 27276 57734
rect 69088 58006 69164 58012
rect 69088 57942 69094 58006
rect 69158 57942 69164 58006
rect 69088 57734 69164 57942
rect 74936 57870 75012 58078
rect 75616 58006 75692 58214
rect 75616 57974 75622 58006
rect 75621 57942 75622 57974
rect 75686 57974 75692 58006
rect 75686 57942 75687 57974
rect 75621 57941 75687 57942
rect 74936 57838 74942 57870
rect 74941 57806 74942 57838
rect 75006 57838 75012 57870
rect 75213 57870 75279 57871
rect 75213 57838 75214 57870
rect 75006 57806 75007 57838
rect 74941 57805 75007 57806
rect 75208 57806 75214 57838
rect 75278 57838 75279 57870
rect 75621 57870 75687 57871
rect 75621 57838 75622 57870
rect 75278 57806 75284 57838
rect 69088 57702 69094 57734
rect 27200 57664 27276 57670
rect 69093 57670 69094 57702
rect 69158 57702 69164 57734
rect 69158 57670 69159 57702
rect 69093 57669 69159 57670
rect 20606 57534 20607 57566
rect 20541 57533 20607 57534
rect 20808 57534 20814 57598
rect 20878 57534 20884 57598
rect 20808 57528 20884 57534
rect 75208 57598 75284 57806
rect 75208 57534 75214 57598
rect 75278 57534 75284 57598
rect 75208 57528 75284 57534
rect 75616 57806 75622 57838
rect 75686 57838 75687 57870
rect 75686 57806 75692 57838
rect 75616 57598 75692 57806
rect 75616 57534 75622 57598
rect 75686 57534 75692 57598
rect 75616 57528 75692 57534
rect 952 57398 1230 57462
rect 1294 57398 1300 57462
rect 952 55966 1300 57398
rect 20536 57462 20612 57468
rect 20536 57398 20542 57462
rect 20606 57398 20612 57462
rect 20536 57190 20612 57398
rect 20536 57158 20542 57190
rect 20541 57126 20542 57158
rect 20606 57158 20612 57190
rect 75480 57462 75556 57468
rect 75480 57398 75486 57462
rect 75550 57398 75556 57462
rect 75480 57190 75556 57398
rect 75480 57158 75486 57190
rect 20606 57126 20607 57158
rect 20541 57125 20607 57126
rect 75485 57126 75486 57158
rect 75550 57158 75556 57190
rect 94656 57462 95004 59030
rect 94656 57398 94662 57462
rect 94726 57398 95004 57462
rect 75550 57126 75551 57158
rect 75485 57125 75551 57126
rect 20541 57054 20607 57055
rect 20541 57022 20542 57054
rect 20536 56990 20542 57022
rect 20606 57022 20607 57054
rect 21493 57054 21559 57055
rect 21493 57022 21494 57054
rect 20606 56990 20612 57022
rect 20536 56782 20612 56990
rect 20536 56718 20542 56782
rect 20606 56718 20612 56782
rect 20536 56712 20612 56718
rect 21488 56990 21494 57022
rect 21558 57022 21559 57054
rect 21624 57054 21700 57060
rect 21558 56990 21564 57022
rect 21488 56782 21564 56990
rect 21488 56718 21494 56782
rect 21558 56718 21564 56782
rect 21624 56990 21630 57054
rect 21694 56990 21700 57054
rect 22173 57054 22239 57055
rect 22173 57022 22174 57054
rect 21624 56782 21700 56990
rect 21624 56750 21630 56782
rect 21488 56712 21564 56718
rect 21629 56718 21630 56750
rect 21694 56750 21700 56782
rect 22168 56990 22174 57022
rect 22238 57022 22239 57054
rect 73848 57054 73924 57060
rect 22238 56990 22244 57022
rect 22168 56782 22244 56990
rect 73848 56990 73854 57054
rect 73918 56990 73924 57054
rect 21694 56718 21695 56750
rect 21629 56717 21695 56718
rect 22168 56718 22174 56782
rect 22238 56718 22244 56782
rect 22168 56712 22244 56718
rect 27200 56782 27276 56788
rect 27200 56718 27206 56782
rect 27270 56718 27276 56782
rect 73848 56782 73924 56990
rect 73848 56750 73854 56782
rect 20400 56646 20476 56652
rect 20400 56582 20406 56646
rect 20470 56582 20476 56646
rect 20400 56374 20476 56582
rect 20400 56342 20406 56374
rect 20405 56310 20406 56342
rect 20470 56342 20476 56374
rect 20944 56646 21020 56652
rect 20944 56582 20950 56646
rect 21014 56582 21020 56646
rect 21629 56646 21695 56647
rect 21629 56614 21630 56646
rect 20944 56374 21020 56582
rect 20944 56342 20950 56374
rect 20470 56310 20471 56342
rect 20405 56309 20471 56310
rect 20949 56310 20950 56342
rect 21014 56342 21020 56374
rect 21624 56582 21630 56614
rect 21694 56614 21695 56646
rect 22032 56646 22108 56652
rect 21694 56582 21700 56614
rect 21624 56374 21700 56582
rect 21014 56310 21015 56342
rect 20949 56309 21015 56310
rect 21624 56310 21630 56374
rect 21694 56310 21700 56374
rect 22032 56582 22038 56646
rect 22102 56582 22108 56646
rect 22032 56374 22108 56582
rect 27200 56510 27276 56718
rect 73853 56718 73854 56750
rect 73918 56750 73924 56782
rect 74256 57054 74332 57060
rect 74256 56990 74262 57054
rect 74326 56990 74332 57054
rect 74256 56782 74332 56990
rect 74256 56750 74262 56782
rect 73918 56718 73919 56750
rect 73853 56717 73919 56718
rect 74261 56718 74262 56750
rect 74326 56750 74332 56782
rect 74800 57054 74876 57060
rect 74800 56990 74806 57054
rect 74870 56990 74876 57054
rect 74800 56782 74876 56990
rect 74800 56750 74806 56782
rect 74326 56718 74327 56750
rect 74261 56717 74327 56718
rect 74805 56718 74806 56750
rect 74870 56750 74876 56782
rect 74936 57054 75012 57060
rect 74936 56990 74942 57054
rect 75006 56990 75012 57054
rect 75485 57054 75551 57055
rect 75485 57022 75486 57054
rect 74936 56782 75012 56990
rect 74936 56750 74942 56782
rect 74870 56718 74871 56750
rect 74805 56717 74871 56718
rect 74941 56718 74942 56750
rect 75006 56750 75012 56782
rect 75480 56990 75486 57022
rect 75550 57022 75551 57054
rect 75550 56990 75556 57022
rect 75480 56782 75556 56990
rect 75006 56718 75007 56750
rect 74941 56717 75007 56718
rect 75480 56718 75486 56782
rect 75550 56718 75556 56782
rect 75480 56712 75556 56718
rect 73853 56646 73919 56647
rect 73853 56614 73854 56646
rect 27200 56478 27206 56510
rect 27205 56446 27206 56478
rect 27270 56478 27276 56510
rect 73848 56582 73854 56614
rect 73918 56614 73919 56646
rect 74397 56646 74463 56647
rect 74397 56614 74398 56646
rect 73918 56582 73924 56614
rect 27270 56446 27271 56478
rect 27205 56445 27271 56446
rect 22032 56342 22038 56374
rect 21624 56304 21700 56310
rect 22037 56310 22038 56342
rect 22102 56342 22108 56374
rect 73848 56374 73924 56582
rect 22102 56310 22103 56342
rect 22037 56309 22103 56310
rect 73848 56310 73854 56374
rect 73918 56310 73924 56374
rect 73848 56304 73924 56310
rect 74392 56582 74398 56614
rect 74462 56614 74463 56646
rect 75213 56646 75279 56647
rect 75213 56614 75214 56646
rect 74462 56582 74468 56614
rect 74392 56374 74468 56582
rect 74392 56310 74398 56374
rect 74462 56310 74468 56374
rect 74392 56304 74468 56310
rect 75208 56582 75214 56614
rect 75278 56614 75279 56646
rect 75621 56646 75687 56647
rect 75621 56614 75622 56646
rect 75278 56582 75284 56614
rect 75208 56374 75284 56582
rect 75208 56310 75214 56374
rect 75278 56310 75284 56374
rect 75208 56304 75284 56310
rect 75616 56582 75622 56614
rect 75686 56614 75687 56646
rect 75686 56582 75692 56614
rect 75616 56374 75692 56582
rect 75616 56310 75622 56374
rect 75686 56310 75692 56374
rect 75616 56304 75692 56310
rect 20405 56238 20471 56239
rect 20405 56206 20406 56238
rect 952 55902 1230 55966
rect 1294 55902 1300 55966
rect 952 54062 1300 55902
rect 20400 56174 20406 56206
rect 20470 56206 20471 56238
rect 20949 56238 21015 56239
rect 20949 56206 20950 56238
rect 20470 56174 20476 56206
rect 20400 55966 20476 56174
rect 20400 55902 20406 55966
rect 20470 55902 20476 55966
rect 20400 55896 20476 55902
rect 20944 56174 20950 56206
rect 21014 56206 21015 56238
rect 21085 56238 21151 56239
rect 21085 56206 21086 56238
rect 21014 56174 21020 56206
rect 20944 55966 21020 56174
rect 20944 55902 20950 55966
rect 21014 55902 21020 55966
rect 20944 55896 21020 55902
rect 21080 56174 21086 56206
rect 21150 56206 21151 56238
rect 21765 56238 21831 56239
rect 21765 56206 21766 56238
rect 21150 56174 21156 56206
rect 21080 55966 21156 56174
rect 21080 55902 21086 55966
rect 21150 55902 21156 55966
rect 21080 55896 21156 55902
rect 21760 56174 21766 56206
rect 21830 56206 21831 56238
rect 22037 56238 22103 56239
rect 22037 56206 22038 56238
rect 21830 56174 21836 56206
rect 21760 55966 21836 56174
rect 21760 55902 21766 55966
rect 21830 55902 21836 55966
rect 21760 55896 21836 55902
rect 22032 56174 22038 56206
rect 22102 56206 22103 56238
rect 73984 56238 74060 56244
rect 22102 56174 22108 56206
rect 22032 55966 22108 56174
rect 22032 55902 22038 55966
rect 22102 55902 22108 55966
rect 73984 56174 73990 56238
rect 74054 56174 74060 56238
rect 73984 55966 74060 56174
rect 73984 55934 73990 55966
rect 22032 55896 22108 55902
rect 73989 55902 73990 55934
rect 74054 55934 74060 55966
rect 74392 56238 74468 56244
rect 74392 56174 74398 56238
rect 74462 56174 74468 56238
rect 74669 56238 74735 56239
rect 74669 56206 74670 56238
rect 74392 55966 74468 56174
rect 74392 55934 74398 55966
rect 74054 55902 74055 55934
rect 73989 55901 74055 55902
rect 74397 55902 74398 55934
rect 74462 55934 74468 55966
rect 74664 56174 74670 56206
rect 74734 56206 74735 56238
rect 75072 56238 75148 56244
rect 74734 56174 74740 56206
rect 74664 55966 74740 56174
rect 74462 55902 74463 55934
rect 74397 55901 74463 55902
rect 74664 55902 74670 55966
rect 74734 55902 74740 55966
rect 75072 56174 75078 56238
rect 75142 56174 75148 56238
rect 75072 55966 75148 56174
rect 75072 55934 75078 55966
rect 74664 55896 74740 55902
rect 75077 55902 75078 55934
rect 75142 55934 75148 55966
rect 75480 56238 75556 56244
rect 75480 56174 75486 56238
rect 75550 56174 75556 56238
rect 75480 55966 75556 56174
rect 75480 55934 75486 55966
rect 75142 55902 75143 55934
rect 75077 55901 75143 55902
rect 75485 55902 75486 55934
rect 75550 55934 75556 55966
rect 94656 55966 95004 57398
rect 75550 55902 75551 55934
rect 75485 55901 75551 55902
rect 94656 55902 94662 55966
rect 94726 55902 95004 55966
rect 20405 55830 20471 55831
rect 20405 55798 20406 55830
rect 20400 55766 20406 55798
rect 20470 55798 20471 55830
rect 20808 55830 20884 55836
rect 20470 55766 20476 55798
rect 20400 55558 20476 55766
rect 20400 55494 20406 55558
rect 20470 55494 20476 55558
rect 20808 55766 20814 55830
rect 20878 55766 20884 55830
rect 20808 55558 20884 55766
rect 20808 55526 20814 55558
rect 20400 55488 20476 55494
rect 20813 55494 20814 55526
rect 20878 55526 20884 55558
rect 21624 55830 21700 55836
rect 21624 55766 21630 55830
rect 21694 55766 21700 55830
rect 22037 55830 22103 55831
rect 22037 55798 22038 55830
rect 21624 55558 21700 55766
rect 21624 55526 21630 55558
rect 20878 55494 20879 55526
rect 20813 55493 20879 55494
rect 21629 55494 21630 55526
rect 21694 55526 21700 55558
rect 22032 55766 22038 55798
rect 22102 55798 22103 55830
rect 73853 55830 73919 55831
rect 73853 55798 73854 55830
rect 22102 55766 22108 55798
rect 22032 55558 22108 55766
rect 21694 55494 21695 55526
rect 21629 55493 21695 55494
rect 22032 55494 22038 55558
rect 22102 55494 22108 55558
rect 22032 55488 22108 55494
rect 73848 55766 73854 55798
rect 73918 55798 73919 55830
rect 74261 55830 74327 55831
rect 74261 55798 74262 55830
rect 73918 55766 73924 55798
rect 73848 55558 73924 55766
rect 73848 55494 73854 55558
rect 73918 55494 73924 55558
rect 73848 55488 73924 55494
rect 74256 55766 74262 55798
rect 74326 55798 74327 55830
rect 75616 55830 75692 55836
rect 74326 55766 74332 55798
rect 74256 55558 74332 55766
rect 74256 55494 74262 55558
rect 74326 55494 74332 55558
rect 75616 55766 75622 55830
rect 75686 55766 75692 55830
rect 75616 55558 75692 55766
rect 75616 55526 75622 55558
rect 74256 55488 74332 55494
rect 75621 55494 75622 55526
rect 75686 55526 75692 55558
rect 75686 55494 75687 55526
rect 75621 55493 75687 55494
rect 20813 55422 20879 55423
rect 20813 55390 20814 55422
rect 20808 55358 20814 55390
rect 20878 55390 20879 55422
rect 21080 55422 21156 55428
rect 20878 55358 20884 55390
rect 20808 55150 20884 55358
rect 20808 55086 20814 55150
rect 20878 55086 20884 55150
rect 21080 55358 21086 55422
rect 21150 55358 21156 55422
rect 21080 55150 21156 55358
rect 21080 55118 21086 55150
rect 20808 55080 20884 55086
rect 21085 55086 21086 55118
rect 21150 55118 21156 55150
rect 21488 55422 21564 55428
rect 21488 55358 21494 55422
rect 21558 55358 21564 55422
rect 21629 55422 21695 55423
rect 21629 55390 21630 55422
rect 21488 55150 21564 55358
rect 21488 55118 21494 55150
rect 21150 55086 21151 55118
rect 21085 55085 21151 55086
rect 21493 55086 21494 55118
rect 21558 55118 21564 55150
rect 21624 55358 21630 55390
rect 21694 55390 21695 55422
rect 22173 55422 22239 55423
rect 22173 55390 22174 55422
rect 21694 55358 21700 55390
rect 21624 55150 21700 55358
rect 21558 55086 21559 55118
rect 21493 55085 21559 55086
rect 21624 55086 21630 55150
rect 21694 55086 21700 55150
rect 21624 55080 21700 55086
rect 22168 55358 22174 55390
rect 22238 55390 22239 55422
rect 73984 55422 74060 55428
rect 22238 55358 22244 55390
rect 22168 55150 22244 55358
rect 22168 55086 22174 55150
rect 22238 55086 22244 55150
rect 73984 55358 73990 55422
rect 74054 55358 74060 55422
rect 74397 55422 74463 55423
rect 74397 55390 74398 55422
rect 73984 55150 74060 55358
rect 73984 55118 73990 55150
rect 22168 55080 22244 55086
rect 73989 55086 73990 55118
rect 74054 55118 74060 55150
rect 74392 55358 74398 55390
rect 74462 55390 74463 55422
rect 75213 55422 75279 55423
rect 75213 55390 75214 55422
rect 74462 55358 74468 55390
rect 74392 55150 74468 55358
rect 74054 55086 74055 55118
rect 73989 55085 74055 55086
rect 74392 55086 74398 55150
rect 74462 55086 74468 55150
rect 74392 55080 74468 55086
rect 75208 55358 75214 55390
rect 75278 55390 75279 55422
rect 75278 55358 75284 55390
rect 75208 55150 75284 55358
rect 75208 55086 75214 55150
rect 75278 55086 75284 55150
rect 75208 55080 75284 55086
rect 20400 55014 20476 55020
rect 20400 54950 20406 55014
rect 20470 54950 20476 55014
rect 20949 55014 21015 55015
rect 20949 54982 20950 55014
rect 20400 54742 20476 54950
rect 20400 54710 20406 54742
rect 20405 54678 20406 54710
rect 20470 54710 20476 54742
rect 20944 54950 20950 54982
rect 21014 54982 21015 55014
rect 21085 55014 21151 55015
rect 21085 54982 21086 55014
rect 21014 54950 21020 54982
rect 20944 54742 21020 54950
rect 20470 54678 20471 54710
rect 20405 54677 20471 54678
rect 20944 54678 20950 54742
rect 21014 54678 21020 54742
rect 20944 54672 21020 54678
rect 21080 54950 21086 54982
rect 21150 54982 21151 55014
rect 21624 55014 21700 55020
rect 21150 54950 21156 54982
rect 21080 54742 21156 54950
rect 21080 54678 21086 54742
rect 21150 54678 21156 54742
rect 21624 54950 21630 55014
rect 21694 54950 21700 55014
rect 21624 54742 21700 54950
rect 21624 54710 21630 54742
rect 21080 54672 21156 54678
rect 21629 54678 21630 54710
rect 21694 54710 21700 54742
rect 22032 55014 22108 55020
rect 22032 54950 22038 55014
rect 22102 54950 22108 55014
rect 22032 54742 22108 54950
rect 22032 54710 22038 54742
rect 21694 54678 21695 54710
rect 21629 54677 21695 54678
rect 22037 54678 22038 54710
rect 22102 54710 22108 54742
rect 73848 55014 73924 55020
rect 73848 54950 73854 55014
rect 73918 54950 73924 55014
rect 73848 54742 73924 54950
rect 73848 54710 73854 54742
rect 22102 54678 22103 54710
rect 22037 54677 22103 54678
rect 73853 54678 73854 54710
rect 73918 54710 73924 54742
rect 74256 55014 74332 55020
rect 74256 54950 74262 55014
rect 74326 54950 74332 55014
rect 74669 55014 74735 55015
rect 74669 54982 74670 55014
rect 74256 54742 74332 54950
rect 74256 54710 74262 54742
rect 73918 54678 73919 54710
rect 73853 54677 73919 54678
rect 74261 54678 74262 54710
rect 74326 54710 74332 54742
rect 74664 54950 74670 54982
rect 74734 54982 74735 55014
rect 75616 55014 75692 55020
rect 74734 54950 74740 54982
rect 74664 54742 74740 54950
rect 74326 54678 74327 54710
rect 74261 54677 74327 54678
rect 74664 54678 74670 54742
rect 74734 54678 74740 54742
rect 75616 54950 75622 55014
rect 75686 54950 75692 55014
rect 75616 54742 75692 54950
rect 75616 54710 75622 54742
rect 74664 54672 74740 54678
rect 75621 54678 75622 54710
rect 75686 54710 75692 54742
rect 75686 54678 75687 54710
rect 75621 54677 75687 54678
rect 21493 54606 21559 54607
rect 21493 54574 21494 54606
rect 21488 54542 21494 54574
rect 21558 54574 21559 54606
rect 21629 54606 21695 54607
rect 21629 54574 21630 54606
rect 21558 54542 21564 54574
rect 952 53998 1230 54062
rect 1294 53998 1300 54062
rect 20400 54334 20476 54340
rect 20400 54270 20406 54334
rect 20470 54270 20476 54334
rect 20400 54062 20476 54270
rect 21488 54334 21564 54542
rect 21488 54270 21494 54334
rect 21558 54270 21564 54334
rect 21488 54264 21564 54270
rect 21624 54542 21630 54574
rect 21694 54574 21695 54606
rect 22037 54606 22103 54607
rect 22037 54574 22038 54606
rect 21694 54542 21700 54574
rect 21624 54334 21700 54542
rect 21624 54270 21630 54334
rect 21694 54270 21700 54334
rect 21624 54264 21700 54270
rect 22032 54542 22038 54574
rect 22102 54574 22103 54606
rect 73853 54606 73919 54607
rect 73853 54574 73854 54606
rect 22102 54542 22108 54574
rect 22032 54334 22108 54542
rect 22032 54270 22038 54334
rect 22102 54270 22108 54334
rect 22032 54264 22108 54270
rect 73848 54542 73854 54574
rect 73918 54574 73919 54606
rect 74261 54606 74327 54607
rect 74261 54574 74262 54606
rect 73918 54542 73924 54574
rect 73848 54334 73924 54542
rect 73848 54270 73854 54334
rect 73918 54270 73924 54334
rect 73848 54264 73924 54270
rect 74256 54542 74262 54574
rect 74326 54574 74327 54606
rect 75213 54606 75279 54607
rect 75213 54574 75214 54606
rect 74326 54542 74332 54574
rect 74256 54334 74332 54542
rect 74256 54270 74262 54334
rect 74326 54270 74332 54334
rect 74256 54264 74332 54270
rect 75208 54542 75214 54574
rect 75278 54574 75279 54606
rect 75278 54542 75284 54574
rect 75208 54334 75284 54542
rect 75208 54270 75214 54334
rect 75278 54270 75284 54334
rect 75208 54264 75284 54270
rect 75480 54334 75556 54340
rect 75480 54270 75486 54334
rect 75550 54270 75556 54334
rect 20400 54030 20406 54062
rect 952 52430 1300 53998
rect 20405 53998 20406 54030
rect 20470 54030 20476 54062
rect 27064 54062 27140 54068
rect 20470 53998 20471 54030
rect 20405 53997 20471 53998
rect 27064 53998 27070 54062
rect 27134 53998 27140 54062
rect 27205 54062 27271 54063
rect 27205 54030 27206 54062
rect 20541 53926 20607 53927
rect 20541 53894 20542 53926
rect 20536 53862 20542 53894
rect 20606 53894 20607 53926
rect 21488 53926 21564 53932
rect 20606 53862 20612 53894
rect 20536 53654 20612 53862
rect 20536 53590 20542 53654
rect 20606 53590 20612 53654
rect 21488 53862 21494 53926
rect 21558 53862 21564 53926
rect 21488 53654 21564 53862
rect 21488 53622 21494 53654
rect 20536 53584 20612 53590
rect 21493 53590 21494 53622
rect 21558 53622 21564 53654
rect 26928 53654 27004 53660
rect 21558 53590 21559 53622
rect 21493 53589 21559 53590
rect 26928 53590 26934 53654
rect 26998 53590 27004 53654
rect 27064 53654 27140 53998
rect 27200 53998 27206 54030
rect 27270 54030 27271 54062
rect 68952 54062 69028 54068
rect 27270 53998 27276 54030
rect 27200 53790 27276 53998
rect 27200 53726 27206 53790
rect 27270 53726 27276 53790
rect 68952 53998 68958 54062
rect 69022 53998 69028 54062
rect 75480 54062 75556 54270
rect 75480 54030 75486 54062
rect 68952 53790 69028 53998
rect 75485 53998 75486 54030
rect 75550 54030 75556 54062
rect 94656 54062 95004 55902
rect 75550 53998 75551 54030
rect 75485 53997 75551 53998
rect 94656 53998 94662 54062
rect 94726 53998 95004 54062
rect 68952 53758 68958 53790
rect 27200 53720 27276 53726
rect 68957 53726 68958 53758
rect 69022 53758 69028 53790
rect 74664 53926 74740 53932
rect 74664 53862 74670 53926
rect 74734 53862 74740 53926
rect 75077 53926 75143 53927
rect 75077 53894 75078 53926
rect 69022 53726 69023 53758
rect 68957 53725 69023 53726
rect 27064 53622 27070 53654
rect 20536 53518 20612 53524
rect 20536 53454 20542 53518
rect 20606 53454 20612 53518
rect 20536 53246 20612 53454
rect 26928 53382 27004 53590
rect 27069 53590 27070 53622
rect 27134 53622 27140 53654
rect 69088 53654 69164 53660
rect 27134 53590 27135 53622
rect 27069 53589 27135 53590
rect 69088 53590 69094 53654
rect 69158 53590 69164 53654
rect 74664 53654 74740 53862
rect 74664 53622 74670 53654
rect 26928 53350 26934 53382
rect 26933 53318 26934 53350
rect 26998 53350 27004 53382
rect 69088 53382 69164 53590
rect 74669 53590 74670 53622
rect 74734 53622 74740 53654
rect 75072 53862 75078 53894
rect 75142 53894 75143 53926
rect 75485 53926 75551 53927
rect 75485 53894 75486 53926
rect 75142 53862 75148 53894
rect 75072 53654 75148 53862
rect 74734 53590 74735 53622
rect 74669 53589 74735 53590
rect 75072 53590 75078 53654
rect 75142 53590 75148 53654
rect 75072 53584 75148 53590
rect 75480 53862 75486 53894
rect 75550 53894 75551 53926
rect 75550 53862 75556 53894
rect 75480 53654 75556 53862
rect 75480 53590 75486 53654
rect 75550 53590 75556 53654
rect 75480 53584 75556 53590
rect 74941 53518 75007 53519
rect 74941 53486 74942 53518
rect 69088 53350 69094 53382
rect 26998 53318 26999 53350
rect 26933 53317 26999 53318
rect 69093 53318 69094 53350
rect 69158 53350 69164 53382
rect 74936 53454 74942 53486
rect 75006 53486 75007 53518
rect 75616 53518 75692 53524
rect 75006 53454 75012 53486
rect 69158 53318 69159 53350
rect 69093 53317 69159 53318
rect 20536 53214 20542 53246
rect 20541 53182 20542 53214
rect 20606 53214 20612 53246
rect 74936 53246 75012 53454
rect 20606 53182 20607 53214
rect 20541 53181 20607 53182
rect 74936 53182 74942 53246
rect 75006 53182 75012 53246
rect 75616 53454 75622 53518
rect 75686 53454 75692 53518
rect 75616 53246 75692 53454
rect 75616 53214 75622 53246
rect 74936 53176 75012 53182
rect 75621 53182 75622 53214
rect 75686 53214 75692 53246
rect 75686 53182 75687 53214
rect 75621 53181 75687 53182
rect 20405 53110 20471 53111
rect 20405 53078 20406 53110
rect 20400 53046 20406 53078
rect 20470 53078 20471 53110
rect 20944 53110 21020 53116
rect 20470 53046 20476 53078
rect 20400 52838 20476 53046
rect 20400 52774 20406 52838
rect 20470 52774 20476 52838
rect 20944 53046 20950 53110
rect 21014 53046 21020 53110
rect 20944 52838 21020 53046
rect 20944 52806 20950 52838
rect 20400 52768 20476 52774
rect 20949 52774 20950 52806
rect 21014 52806 21020 52838
rect 21080 53110 21156 53116
rect 21080 53046 21086 53110
rect 21150 53046 21156 53110
rect 21080 52838 21156 53046
rect 21080 52806 21086 52838
rect 21014 52774 21015 52806
rect 20949 52773 21015 52774
rect 21085 52774 21086 52806
rect 21150 52806 21156 52838
rect 21760 53110 21836 53116
rect 21760 53046 21766 53110
rect 21830 53046 21836 53110
rect 22037 53110 22103 53111
rect 22037 53078 22038 53110
rect 21760 52838 21836 53046
rect 21760 52806 21766 52838
rect 21150 52774 21151 52806
rect 21085 52773 21151 52774
rect 21765 52774 21766 52806
rect 21830 52806 21836 52838
rect 22032 53046 22038 53078
rect 22102 53078 22103 53110
rect 73984 53110 74060 53116
rect 22102 53046 22108 53078
rect 22032 52838 22108 53046
rect 73984 53046 73990 53110
rect 74054 53046 74060 53110
rect 74261 53110 74327 53111
rect 74261 53078 74262 53110
rect 21830 52774 21831 52806
rect 21765 52773 21831 52774
rect 22032 52774 22038 52838
rect 22102 52774 22108 52838
rect 22032 52768 22108 52774
rect 27200 52838 27276 52844
rect 27200 52774 27206 52838
rect 27270 52774 27276 52838
rect 952 52366 1230 52430
rect 1294 52366 1300 52430
rect 20536 52702 20612 52708
rect 20536 52638 20542 52702
rect 20606 52638 20612 52702
rect 20536 52430 20612 52638
rect 20536 52398 20542 52430
rect 952 50798 1300 52366
rect 20541 52366 20542 52398
rect 20606 52398 20612 52430
rect 21624 52702 21700 52708
rect 21624 52638 21630 52702
rect 21694 52638 21700 52702
rect 21624 52430 21700 52638
rect 21624 52398 21630 52430
rect 20606 52366 20607 52398
rect 20541 52365 20607 52366
rect 21629 52366 21630 52398
rect 21694 52398 21700 52430
rect 22032 52702 22108 52708
rect 22032 52638 22038 52702
rect 22102 52638 22108 52702
rect 22032 52430 22108 52638
rect 27200 52566 27276 52774
rect 27200 52534 27206 52566
rect 27205 52502 27206 52534
rect 27270 52534 27276 52566
rect 69088 52838 69164 52844
rect 69088 52774 69094 52838
rect 69158 52774 69164 52838
rect 73984 52838 74060 53046
rect 73984 52806 73990 52838
rect 69088 52566 69164 52774
rect 73989 52774 73990 52806
rect 74054 52806 74060 52838
rect 74256 53046 74262 53078
rect 74326 53078 74327 53110
rect 74669 53110 74735 53111
rect 74669 53078 74670 53110
rect 74326 53046 74332 53078
rect 74256 52838 74332 53046
rect 74054 52774 74055 52806
rect 73989 52773 74055 52774
rect 74256 52774 74262 52838
rect 74326 52774 74332 52838
rect 74256 52768 74332 52774
rect 74664 53046 74670 53078
rect 74734 53078 74735 53110
rect 75485 53110 75551 53111
rect 75485 53078 75486 53110
rect 74734 53046 74740 53078
rect 74664 52838 74740 53046
rect 74664 52774 74670 52838
rect 74734 52774 74740 52838
rect 74664 52768 74740 52774
rect 75480 53046 75486 53078
rect 75550 53078 75551 53110
rect 75550 53046 75556 53078
rect 75480 52838 75556 53046
rect 75480 52774 75486 52838
rect 75550 52774 75556 52838
rect 75480 52768 75556 52774
rect 69088 52534 69094 52566
rect 27270 52502 27271 52534
rect 27205 52501 27271 52502
rect 69093 52502 69094 52534
rect 69158 52534 69164 52566
rect 73848 52702 73924 52708
rect 73848 52638 73854 52702
rect 73918 52638 73924 52702
rect 74397 52702 74463 52703
rect 74397 52670 74398 52702
rect 69158 52502 69159 52534
rect 69093 52501 69159 52502
rect 22032 52398 22038 52430
rect 21694 52366 21695 52398
rect 21629 52365 21695 52366
rect 22037 52366 22038 52398
rect 22102 52398 22108 52430
rect 73848 52430 73924 52638
rect 73848 52398 73854 52430
rect 22102 52366 22103 52398
rect 22037 52365 22103 52366
rect 73853 52366 73854 52398
rect 73918 52398 73924 52430
rect 74392 52638 74398 52670
rect 74462 52670 74463 52702
rect 74800 52702 74876 52708
rect 74462 52638 74468 52670
rect 74392 52430 74468 52638
rect 73918 52366 73919 52398
rect 73853 52365 73919 52366
rect 74392 52366 74398 52430
rect 74462 52366 74468 52430
rect 74800 52638 74806 52702
rect 74870 52638 74876 52702
rect 75485 52702 75551 52703
rect 75485 52670 75486 52702
rect 74800 52430 74876 52638
rect 74800 52398 74806 52430
rect 74392 52360 74468 52366
rect 74805 52366 74806 52398
rect 74870 52398 74876 52430
rect 75480 52638 75486 52670
rect 75550 52670 75551 52702
rect 75550 52638 75556 52670
rect 75480 52430 75556 52638
rect 74870 52366 74871 52398
rect 74805 52365 74871 52366
rect 75480 52366 75486 52430
rect 75550 52366 75556 52430
rect 75480 52360 75556 52366
rect 94656 52430 95004 53998
rect 94656 52366 94662 52430
rect 94726 52366 95004 52430
rect 20541 52294 20607 52295
rect 20541 52262 20542 52294
rect 20536 52230 20542 52262
rect 20606 52262 20607 52294
rect 20944 52294 21020 52300
rect 20606 52230 20612 52262
rect 20536 52022 20612 52230
rect 20536 51958 20542 52022
rect 20606 51958 20612 52022
rect 20944 52230 20950 52294
rect 21014 52230 21020 52294
rect 20944 52022 21020 52230
rect 20944 51990 20950 52022
rect 20536 51952 20612 51958
rect 20949 51958 20950 51990
rect 21014 51990 21020 52022
rect 21080 52294 21156 52300
rect 21080 52230 21086 52294
rect 21150 52230 21156 52294
rect 21221 52294 21287 52295
rect 21221 52262 21222 52294
rect 21080 52022 21156 52230
rect 21080 51990 21086 52022
rect 21014 51958 21015 51990
rect 20949 51957 21015 51958
rect 21085 51958 21086 51990
rect 21150 51990 21156 52022
rect 21216 52230 21222 52262
rect 21286 52262 21287 52294
rect 21629 52294 21695 52295
rect 21629 52262 21630 52294
rect 21286 52230 21292 52262
rect 21216 52022 21292 52230
rect 21150 51958 21151 51990
rect 21085 51957 21151 51958
rect 21216 51958 21222 52022
rect 21286 51958 21292 52022
rect 21216 51952 21292 51958
rect 21624 52230 21630 52262
rect 21694 52262 21695 52294
rect 22037 52294 22103 52295
rect 22037 52262 22038 52294
rect 21694 52230 21700 52262
rect 21624 52022 21700 52230
rect 21624 51958 21630 52022
rect 21694 51958 21700 52022
rect 21624 51952 21700 51958
rect 22032 52230 22038 52262
rect 22102 52262 22103 52294
rect 73984 52294 74060 52300
rect 22102 52230 22108 52262
rect 22032 52022 22108 52230
rect 22032 51958 22038 52022
rect 22102 51958 22108 52022
rect 73984 52230 73990 52294
rect 74054 52230 74060 52294
rect 73984 52022 74060 52230
rect 73984 51990 73990 52022
rect 22032 51952 22108 51958
rect 73989 51958 73990 51990
rect 74054 51990 74060 52022
rect 74256 52294 74332 52300
rect 74256 52230 74262 52294
rect 74326 52230 74332 52294
rect 74256 52022 74332 52230
rect 74256 51990 74262 52022
rect 74054 51958 74055 51990
rect 73989 51957 74055 51958
rect 74261 51958 74262 51990
rect 74326 51990 74332 52022
rect 74664 52294 74740 52300
rect 74664 52230 74670 52294
rect 74734 52230 74740 52294
rect 74664 52022 74740 52230
rect 74664 51990 74670 52022
rect 74326 51958 74327 51990
rect 74261 51957 74327 51958
rect 74669 51958 74670 51990
rect 74734 51990 74740 52022
rect 75480 52294 75556 52300
rect 75480 52230 75486 52294
rect 75550 52230 75556 52294
rect 75480 52022 75556 52230
rect 75480 51990 75486 52022
rect 74734 51958 74735 51990
rect 74669 51957 74735 51958
rect 75485 51958 75486 51990
rect 75550 51990 75556 52022
rect 75550 51958 75551 51990
rect 75485 51957 75551 51958
rect 20536 51886 20612 51892
rect 20536 51822 20542 51886
rect 20606 51822 20612 51886
rect 20536 51614 20612 51822
rect 20536 51582 20542 51614
rect 20541 51550 20542 51582
rect 20606 51582 20612 51614
rect 21488 51886 21564 51892
rect 21488 51822 21494 51886
rect 21558 51822 21564 51886
rect 21765 51886 21831 51887
rect 21765 51854 21766 51886
rect 21488 51614 21564 51822
rect 21488 51582 21494 51614
rect 20606 51550 20607 51582
rect 20541 51549 20607 51550
rect 21493 51550 21494 51582
rect 21558 51582 21564 51614
rect 21760 51822 21766 51854
rect 21830 51854 21831 51886
rect 22168 51886 22244 51892
rect 21830 51822 21836 51854
rect 21760 51614 21836 51822
rect 21558 51550 21559 51582
rect 21493 51549 21559 51550
rect 21760 51550 21766 51614
rect 21830 51550 21836 51614
rect 22168 51822 22174 51886
rect 22238 51822 22244 51886
rect 73989 51886 74055 51887
rect 73989 51854 73990 51886
rect 22168 51614 22244 51822
rect 22168 51582 22174 51614
rect 21760 51544 21836 51550
rect 22173 51550 22174 51582
rect 22238 51582 22244 51614
rect 73984 51822 73990 51854
rect 74054 51854 74055 51886
rect 74392 51886 74468 51892
rect 74054 51822 74060 51854
rect 73984 51614 74060 51822
rect 22238 51550 22239 51582
rect 22173 51549 22239 51550
rect 73984 51550 73990 51614
rect 74054 51550 74060 51614
rect 74392 51822 74398 51886
rect 74462 51822 74468 51886
rect 74941 51886 75007 51887
rect 74941 51854 74942 51886
rect 74392 51614 74468 51822
rect 74392 51582 74398 51614
rect 73984 51544 74060 51550
rect 74397 51550 74398 51582
rect 74462 51582 74468 51614
rect 74936 51822 74942 51854
rect 75006 51854 75007 51886
rect 75480 51886 75556 51892
rect 75006 51822 75012 51854
rect 74936 51614 75012 51822
rect 74462 51550 74463 51582
rect 74397 51549 74463 51550
rect 74936 51550 74942 51614
rect 75006 51550 75012 51614
rect 75480 51822 75486 51886
rect 75550 51822 75556 51886
rect 75480 51614 75556 51822
rect 75480 51582 75486 51614
rect 74936 51544 75012 51550
rect 75485 51550 75486 51582
rect 75550 51582 75556 51614
rect 75550 51550 75551 51582
rect 75485 51549 75551 51550
rect 20813 51478 20879 51479
rect 20813 51446 20814 51478
rect 20808 51414 20814 51446
rect 20878 51446 20879 51478
rect 21357 51478 21423 51479
rect 21357 51446 21358 51478
rect 20878 51414 20884 51446
rect 20808 51206 20884 51414
rect 20808 51142 20814 51206
rect 20878 51142 20884 51206
rect 20808 51136 20884 51142
rect 21352 51414 21358 51446
rect 21422 51446 21423 51478
rect 21624 51478 21700 51484
rect 21422 51414 21428 51446
rect 21352 51206 21428 51414
rect 21352 51142 21358 51206
rect 21422 51142 21428 51206
rect 21624 51414 21630 51478
rect 21694 51414 21700 51478
rect 22037 51478 22103 51479
rect 22037 51446 22038 51478
rect 21624 51206 21700 51414
rect 21624 51174 21630 51206
rect 21352 51136 21428 51142
rect 21629 51142 21630 51174
rect 21694 51174 21700 51206
rect 22032 51414 22038 51446
rect 22102 51446 22103 51478
rect 73853 51478 73919 51479
rect 73853 51446 73854 51478
rect 22102 51414 22108 51446
rect 22032 51206 22108 51414
rect 21694 51142 21695 51174
rect 21629 51141 21695 51142
rect 22032 51142 22038 51206
rect 22102 51142 22108 51206
rect 22032 51136 22108 51142
rect 73848 51414 73854 51446
rect 73918 51446 73919 51478
rect 74392 51478 74468 51484
rect 73918 51414 73924 51446
rect 73848 51206 73924 51414
rect 73848 51142 73854 51206
rect 73918 51142 73924 51206
rect 74392 51414 74398 51478
rect 74462 51414 74468 51478
rect 74392 51206 74468 51414
rect 74392 51174 74398 51206
rect 73848 51136 73924 51142
rect 74397 51142 74398 51174
rect 74462 51174 74468 51206
rect 74800 51478 74876 51484
rect 74800 51414 74806 51478
rect 74870 51414 74876 51478
rect 74800 51206 74876 51414
rect 74800 51174 74806 51206
rect 74462 51142 74463 51174
rect 74397 51141 74463 51142
rect 74805 51142 74806 51174
rect 74870 51174 74876 51206
rect 74870 51142 74871 51174
rect 74805 51141 74871 51142
rect 952 50734 1230 50798
rect 1294 50734 1300 50798
rect 20400 51070 20476 51076
rect 20400 51006 20406 51070
rect 20470 51006 20476 51070
rect 20813 51070 20879 51071
rect 20813 51038 20814 51070
rect 20400 50798 20476 51006
rect 20400 50766 20406 50798
rect 952 49166 1300 50734
rect 20405 50734 20406 50766
rect 20470 50766 20476 50798
rect 20808 51006 20814 51038
rect 20878 51038 20879 51070
rect 21080 51070 21156 51076
rect 20878 51006 20884 51038
rect 20808 50798 20884 51006
rect 20470 50734 20471 50766
rect 20405 50733 20471 50734
rect 20808 50734 20814 50798
rect 20878 50734 20884 50798
rect 21080 51006 21086 51070
rect 21150 51006 21156 51070
rect 21629 51070 21695 51071
rect 21629 51038 21630 51070
rect 21080 50798 21156 51006
rect 21080 50766 21086 50798
rect 20808 50728 20884 50734
rect 21085 50734 21086 50766
rect 21150 50766 21156 50798
rect 21624 51006 21630 51038
rect 21694 51038 21695 51070
rect 22032 51070 22108 51076
rect 21694 51006 21700 51038
rect 21624 50798 21700 51006
rect 21150 50734 21151 50766
rect 21085 50733 21151 50734
rect 21624 50734 21630 50798
rect 21694 50734 21700 50798
rect 22032 51006 22038 51070
rect 22102 51006 22108 51070
rect 73853 51070 73919 51071
rect 73853 51038 73854 51070
rect 22032 50798 22108 51006
rect 22032 50766 22038 50798
rect 21624 50728 21700 50734
rect 22037 50734 22038 50766
rect 22102 50766 22108 50798
rect 73848 51006 73854 51038
rect 73918 51038 73919 51070
rect 74397 51070 74463 51071
rect 74397 51038 74398 51070
rect 73918 51006 73924 51038
rect 73848 50798 73924 51006
rect 22102 50734 22103 50766
rect 22037 50733 22103 50734
rect 73848 50734 73854 50798
rect 73918 50734 73924 50798
rect 73848 50728 73924 50734
rect 74392 51006 74398 51038
rect 74462 51038 74463 51070
rect 75213 51070 75279 51071
rect 75213 51038 75214 51070
rect 74462 51006 74468 51038
rect 74392 50798 74468 51006
rect 74392 50734 74398 50798
rect 74462 50734 74468 50798
rect 74392 50728 74468 50734
rect 75208 51006 75214 51038
rect 75278 51038 75279 51070
rect 75621 51070 75687 51071
rect 75621 51038 75622 51070
rect 75278 51006 75284 51038
rect 75208 50798 75284 51006
rect 75208 50734 75214 50798
rect 75278 50734 75284 50798
rect 75208 50728 75284 50734
rect 75616 51006 75622 51038
rect 75686 51038 75687 51070
rect 75686 51006 75692 51038
rect 75616 50798 75692 51006
rect 75616 50734 75622 50798
rect 75686 50734 75692 50798
rect 75616 50728 75692 50734
rect 21221 50662 21287 50663
rect 21221 50630 21222 50662
rect 21216 50598 21222 50630
rect 21286 50630 21287 50662
rect 21765 50662 21831 50663
rect 21765 50630 21766 50662
rect 21286 50598 21292 50630
rect 20405 50390 20471 50391
rect 20405 50358 20406 50390
rect 20400 50326 20406 50358
rect 20470 50358 20471 50390
rect 21216 50390 21292 50598
rect 20470 50326 20476 50358
rect 20400 50118 20476 50326
rect 21216 50326 21222 50390
rect 21286 50326 21292 50390
rect 21216 50320 21292 50326
rect 21760 50598 21766 50630
rect 21830 50630 21831 50662
rect 22173 50662 22239 50663
rect 22173 50630 22174 50662
rect 21830 50598 21836 50630
rect 21760 50390 21836 50598
rect 21760 50326 21766 50390
rect 21830 50326 21836 50390
rect 21760 50320 21836 50326
rect 22168 50598 22174 50630
rect 22238 50630 22239 50662
rect 73848 50662 73924 50668
rect 22238 50598 22244 50630
rect 22168 50390 22244 50598
rect 22168 50326 22174 50390
rect 22238 50326 22244 50390
rect 73848 50598 73854 50662
rect 73918 50598 73924 50662
rect 74261 50662 74327 50663
rect 74261 50630 74262 50662
rect 73848 50390 73924 50598
rect 73848 50358 73854 50390
rect 22168 50320 22244 50326
rect 73853 50326 73854 50358
rect 73918 50358 73924 50390
rect 74256 50598 74262 50630
rect 74326 50630 74327 50662
rect 74800 50662 74876 50668
rect 74326 50598 74332 50630
rect 74256 50390 74332 50598
rect 73918 50326 73919 50358
rect 73853 50325 73919 50326
rect 74256 50326 74262 50390
rect 74326 50326 74332 50390
rect 74800 50598 74806 50662
rect 74870 50598 74876 50662
rect 75077 50662 75143 50663
rect 75077 50630 75078 50662
rect 74800 50390 74876 50598
rect 74800 50358 74806 50390
rect 74256 50320 74332 50326
rect 74805 50326 74806 50358
rect 74870 50358 74876 50390
rect 75072 50598 75078 50630
rect 75142 50630 75143 50662
rect 94656 50662 95004 52366
rect 75142 50598 75148 50630
rect 75072 50390 75148 50598
rect 94656 50598 94662 50662
rect 94726 50598 95004 50662
rect 74870 50326 74871 50358
rect 74805 50325 74871 50326
rect 75072 50326 75078 50390
rect 75142 50326 75148 50390
rect 75621 50390 75687 50391
rect 75621 50358 75622 50390
rect 75072 50320 75148 50326
rect 75616 50326 75622 50358
rect 75686 50358 75687 50390
rect 75686 50326 75692 50358
rect 20400 50054 20406 50118
rect 20470 50054 20476 50118
rect 20400 50048 20476 50054
rect 21624 50254 21700 50260
rect 21624 50190 21630 50254
rect 21694 50190 21700 50254
rect 21624 49982 21700 50190
rect 21624 49950 21630 49982
rect 21629 49918 21630 49950
rect 21694 49950 21700 49982
rect 22168 50254 22244 50260
rect 22168 50190 22174 50254
rect 22238 50190 22244 50254
rect 73853 50254 73919 50255
rect 73853 50222 73854 50254
rect 22168 49982 22244 50190
rect 73848 50190 73854 50222
rect 73918 50222 73919 50254
rect 74261 50254 74327 50255
rect 74261 50222 74262 50254
rect 73918 50190 73924 50222
rect 22168 49950 22174 49982
rect 21694 49918 21695 49950
rect 21629 49917 21695 49918
rect 22173 49918 22174 49950
rect 22238 49950 22244 49982
rect 69088 49982 69164 49988
rect 22238 49918 22239 49950
rect 22173 49917 22239 49918
rect 69088 49918 69094 49982
rect 69158 49918 69164 49982
rect 21352 49846 21428 49852
rect 21352 49782 21358 49846
rect 21422 49782 21428 49846
rect 20405 49574 20471 49575
rect 20405 49542 20406 49574
rect 20400 49510 20406 49542
rect 20470 49542 20471 49574
rect 21352 49574 21428 49782
rect 21352 49542 21358 49574
rect 20470 49510 20476 49542
rect 20400 49302 20476 49510
rect 21357 49510 21358 49542
rect 21422 49542 21428 49574
rect 27200 49710 27276 49716
rect 27200 49646 27206 49710
rect 27270 49646 27276 49710
rect 68957 49710 69023 49711
rect 68957 49678 68958 49710
rect 21422 49510 21423 49542
rect 21357 49509 21423 49510
rect 27200 49438 27276 49646
rect 27200 49406 27206 49438
rect 27205 49374 27206 49406
rect 27270 49406 27276 49438
rect 68952 49646 68958 49678
rect 69022 49678 69023 49710
rect 69088 49710 69164 49918
rect 73848 49982 73924 50190
rect 73848 49918 73854 49982
rect 73918 49918 73924 49982
rect 73848 49912 73924 49918
rect 74256 50190 74262 50222
rect 74326 50222 74327 50254
rect 74326 50190 74332 50222
rect 74256 49982 74332 50190
rect 75616 50118 75692 50326
rect 75616 50054 75622 50118
rect 75686 50054 75692 50118
rect 75616 50048 75692 50054
rect 74256 49918 74262 49982
rect 74326 49918 74332 49982
rect 74256 49912 74332 49918
rect 69088 49678 69094 49710
rect 69022 49646 69028 49678
rect 68952 49438 69028 49646
rect 69093 49646 69094 49678
rect 69158 49678 69164 49710
rect 75072 49846 75148 49852
rect 75072 49782 75078 49846
rect 75142 49782 75148 49846
rect 69158 49646 69159 49678
rect 69093 49645 69159 49646
rect 75072 49574 75148 49782
rect 75072 49542 75078 49574
rect 75077 49510 75078 49542
rect 75142 49542 75148 49574
rect 75616 49574 75692 49580
rect 75142 49510 75143 49542
rect 75077 49509 75143 49510
rect 75616 49510 75622 49574
rect 75686 49510 75692 49574
rect 27270 49374 27271 49406
rect 27205 49373 27271 49374
rect 68952 49374 68958 49438
rect 69022 49374 69028 49438
rect 68952 49368 69028 49374
rect 20400 49238 20406 49302
rect 20470 49238 20476 49302
rect 75616 49302 75692 49510
rect 75616 49270 75622 49302
rect 20400 49232 20476 49238
rect 75621 49238 75622 49270
rect 75686 49270 75692 49302
rect 75686 49238 75687 49270
rect 75621 49237 75687 49238
rect 952 49102 1230 49166
rect 1294 49102 1300 49166
rect 952 47534 1300 49102
rect 20536 49166 20612 49172
rect 20536 49102 20542 49166
rect 20606 49102 20612 49166
rect 21221 49166 21287 49167
rect 21221 49134 21222 49166
rect 20536 48894 20612 49102
rect 20536 48862 20542 48894
rect 20541 48830 20542 48862
rect 20606 48862 20612 48894
rect 21216 49102 21222 49134
rect 21286 49134 21287 49166
rect 75213 49166 75279 49167
rect 75213 49134 75214 49166
rect 21286 49102 21292 49134
rect 21216 48894 21292 49102
rect 75208 49102 75214 49134
rect 75278 49134 75279 49166
rect 75616 49166 75692 49172
rect 75278 49102 75284 49134
rect 20606 48830 20607 48862
rect 20541 48829 20607 48830
rect 21216 48830 21222 48894
rect 21286 48830 21292 48894
rect 69093 48894 69159 48895
rect 69093 48862 69094 48894
rect 21216 48824 21292 48830
rect 69088 48830 69094 48862
rect 69158 48862 69159 48894
rect 75208 48894 75284 49102
rect 69158 48830 69164 48862
rect 20536 48758 20612 48764
rect 20536 48694 20542 48758
rect 20606 48694 20612 48758
rect 21765 48758 21831 48759
rect 21765 48726 21766 48758
rect 20536 48486 20612 48694
rect 20536 48454 20542 48486
rect 20541 48422 20542 48454
rect 20606 48454 20612 48486
rect 21760 48694 21766 48726
rect 21830 48726 21831 48758
rect 22037 48758 22103 48759
rect 22037 48726 22038 48758
rect 21830 48694 21836 48726
rect 21760 48486 21836 48694
rect 20606 48422 20607 48454
rect 20541 48421 20607 48422
rect 21760 48422 21766 48486
rect 21830 48422 21836 48486
rect 21760 48416 21836 48422
rect 22032 48694 22038 48726
rect 22102 48726 22103 48758
rect 22102 48694 22108 48726
rect 22032 48486 22108 48694
rect 69088 48622 69164 48830
rect 75208 48830 75214 48894
rect 75278 48830 75284 48894
rect 75616 49102 75622 49166
rect 75686 49102 75692 49166
rect 75616 48894 75692 49102
rect 75616 48862 75622 48894
rect 75208 48824 75284 48830
rect 75621 48830 75622 48862
rect 75686 48862 75692 48894
rect 94656 49166 95004 50598
rect 94656 49102 94662 49166
rect 94726 49102 95004 49166
rect 75686 48830 75687 48862
rect 75621 48829 75687 48830
rect 69088 48558 69094 48622
rect 69158 48558 69164 48622
rect 69088 48552 69164 48558
rect 73984 48758 74060 48764
rect 73984 48694 73990 48758
rect 74054 48694 74060 48758
rect 22032 48422 22038 48486
rect 22102 48422 22108 48486
rect 73984 48486 74060 48694
rect 73984 48454 73990 48486
rect 22032 48416 22108 48422
rect 73989 48422 73990 48454
rect 74054 48454 74060 48486
rect 74392 48758 74468 48764
rect 74392 48694 74398 48758
rect 74462 48694 74468 48758
rect 74392 48486 74468 48694
rect 74392 48454 74398 48486
rect 74054 48422 74055 48454
rect 73989 48421 74055 48422
rect 74397 48422 74398 48454
rect 74462 48454 74468 48486
rect 75480 48758 75556 48764
rect 75480 48694 75486 48758
rect 75550 48694 75556 48758
rect 75480 48486 75556 48694
rect 75480 48454 75486 48486
rect 74462 48422 74463 48454
rect 74397 48421 74463 48422
rect 75485 48422 75486 48454
rect 75550 48454 75556 48486
rect 75550 48422 75551 48454
rect 75485 48421 75551 48422
rect 20541 48350 20607 48351
rect 20541 48318 20542 48350
rect 20536 48286 20542 48318
rect 20606 48318 20607 48350
rect 20808 48350 20884 48356
rect 20606 48286 20612 48318
rect 20536 48078 20612 48286
rect 20536 48014 20542 48078
rect 20606 48014 20612 48078
rect 20808 48286 20814 48350
rect 20878 48286 20884 48350
rect 21493 48350 21559 48351
rect 21493 48318 21494 48350
rect 20808 48078 20884 48286
rect 20808 48046 20814 48078
rect 20536 48008 20612 48014
rect 20813 48014 20814 48046
rect 20878 48046 20884 48078
rect 21488 48286 21494 48318
rect 21558 48318 21559 48350
rect 21765 48350 21831 48351
rect 21765 48318 21766 48350
rect 21558 48286 21564 48318
rect 21488 48078 21564 48286
rect 20878 48014 20879 48046
rect 20813 48013 20879 48014
rect 21488 48014 21494 48078
rect 21558 48014 21564 48078
rect 21488 48008 21564 48014
rect 21760 48286 21766 48318
rect 21830 48318 21831 48350
rect 22032 48350 22108 48356
rect 21830 48286 21836 48318
rect 21760 48078 21836 48286
rect 21760 48014 21766 48078
rect 21830 48014 21836 48078
rect 22032 48286 22038 48350
rect 22102 48286 22108 48350
rect 22032 48078 22108 48286
rect 22032 48046 22038 48078
rect 21760 48008 21836 48014
rect 22037 48014 22038 48046
rect 22102 48046 22108 48078
rect 73848 48350 73924 48356
rect 73848 48286 73854 48350
rect 73918 48286 73924 48350
rect 74397 48350 74463 48351
rect 74397 48318 74398 48350
rect 73848 48078 73924 48286
rect 73848 48046 73854 48078
rect 22102 48014 22103 48046
rect 22037 48013 22103 48014
rect 73853 48014 73854 48046
rect 73918 48046 73924 48078
rect 74392 48286 74398 48318
rect 74462 48318 74463 48350
rect 74800 48350 74876 48356
rect 74462 48286 74468 48318
rect 74392 48078 74468 48286
rect 73918 48014 73919 48046
rect 73853 48013 73919 48014
rect 74392 48014 74398 48078
rect 74462 48014 74468 48078
rect 74800 48286 74806 48350
rect 74870 48286 74876 48350
rect 74800 48078 74876 48286
rect 74800 48046 74806 48078
rect 74392 48008 74468 48014
rect 74805 48014 74806 48046
rect 74870 48046 74876 48078
rect 75616 48350 75692 48356
rect 75616 48286 75622 48350
rect 75686 48286 75692 48350
rect 75616 48078 75692 48286
rect 75616 48046 75622 48078
rect 74870 48014 74871 48046
rect 74805 48013 74871 48014
rect 75621 48014 75622 48046
rect 75686 48046 75692 48078
rect 75686 48014 75687 48046
rect 75621 48013 75687 48014
rect 20400 47942 20476 47948
rect 20400 47878 20406 47942
rect 20470 47878 20476 47942
rect 20400 47670 20476 47878
rect 20400 47638 20406 47670
rect 20405 47606 20406 47638
rect 20470 47638 20476 47670
rect 21080 47942 21156 47948
rect 21080 47878 21086 47942
rect 21150 47878 21156 47942
rect 21080 47670 21156 47878
rect 21080 47638 21086 47670
rect 20470 47606 20471 47638
rect 20405 47605 20471 47606
rect 21085 47606 21086 47638
rect 21150 47638 21156 47670
rect 21352 47942 21428 47948
rect 21352 47878 21358 47942
rect 21422 47878 21428 47942
rect 21352 47670 21428 47878
rect 21352 47638 21358 47670
rect 21150 47606 21151 47638
rect 21085 47605 21151 47606
rect 21357 47606 21358 47638
rect 21422 47638 21428 47670
rect 21760 47942 21836 47948
rect 21760 47878 21766 47942
rect 21830 47878 21836 47942
rect 21760 47670 21836 47878
rect 21760 47638 21766 47670
rect 21422 47606 21423 47638
rect 21357 47605 21423 47606
rect 21765 47606 21766 47638
rect 21830 47638 21836 47670
rect 22032 47942 22108 47948
rect 22032 47878 22038 47942
rect 22102 47878 22108 47942
rect 22032 47670 22108 47878
rect 22032 47638 22038 47670
rect 21830 47606 21831 47638
rect 21765 47605 21831 47606
rect 22037 47606 22038 47638
rect 22102 47638 22108 47670
rect 73984 47942 74060 47948
rect 73984 47878 73990 47942
rect 74054 47878 74060 47942
rect 74397 47942 74463 47943
rect 74397 47910 74398 47942
rect 73984 47670 74060 47878
rect 73984 47638 73990 47670
rect 22102 47606 22103 47638
rect 22037 47605 22103 47606
rect 73989 47606 73990 47638
rect 74054 47638 74060 47670
rect 74392 47878 74398 47910
rect 74462 47910 74463 47942
rect 75072 47942 75148 47948
rect 74462 47878 74468 47910
rect 74392 47670 74468 47878
rect 74054 47606 74055 47638
rect 73989 47605 74055 47606
rect 74392 47606 74398 47670
rect 74462 47606 74468 47670
rect 75072 47878 75078 47942
rect 75142 47878 75148 47942
rect 75621 47942 75687 47943
rect 75621 47910 75622 47942
rect 75072 47670 75148 47878
rect 75072 47638 75078 47670
rect 74392 47600 74468 47606
rect 75077 47606 75078 47638
rect 75142 47638 75148 47670
rect 75616 47878 75622 47910
rect 75686 47910 75687 47942
rect 75686 47878 75692 47910
rect 75616 47670 75692 47878
rect 75142 47606 75143 47638
rect 75077 47605 75143 47606
rect 75616 47606 75622 47670
rect 75686 47606 75692 47670
rect 75616 47600 75692 47606
rect 952 47470 1230 47534
rect 1294 47470 1300 47534
rect 952 45902 1300 47470
rect 20536 47534 20612 47540
rect 20536 47470 20542 47534
rect 20606 47470 20612 47534
rect 21085 47534 21151 47535
rect 21085 47502 21086 47534
rect 20536 47262 20612 47470
rect 20536 47230 20542 47262
rect 20541 47198 20542 47230
rect 20606 47230 20612 47262
rect 21080 47470 21086 47502
rect 21150 47502 21151 47534
rect 21765 47534 21831 47535
rect 21765 47502 21766 47534
rect 21150 47470 21156 47502
rect 21080 47262 21156 47470
rect 20606 47198 20607 47230
rect 20541 47197 20607 47198
rect 21080 47198 21086 47262
rect 21150 47198 21156 47262
rect 21080 47192 21156 47198
rect 21760 47470 21766 47502
rect 21830 47502 21831 47534
rect 22168 47534 22244 47540
rect 21830 47470 21836 47502
rect 21760 47262 21836 47470
rect 21760 47198 21766 47262
rect 21830 47198 21836 47262
rect 22168 47470 22174 47534
rect 22238 47470 22244 47534
rect 73989 47534 74055 47535
rect 73989 47502 73990 47534
rect 22168 47262 22244 47470
rect 22168 47230 22174 47262
rect 21760 47192 21836 47198
rect 22173 47198 22174 47230
rect 22238 47230 22244 47262
rect 73984 47470 73990 47502
rect 74054 47502 74055 47534
rect 74392 47534 74468 47540
rect 74054 47470 74060 47502
rect 73984 47262 74060 47470
rect 22238 47198 22239 47230
rect 22173 47197 22239 47198
rect 73984 47198 73990 47262
rect 74054 47198 74060 47262
rect 74392 47470 74398 47534
rect 74462 47470 74468 47534
rect 74669 47534 74735 47535
rect 74669 47502 74670 47534
rect 74392 47262 74468 47470
rect 74392 47230 74398 47262
rect 73984 47192 74060 47198
rect 74397 47198 74398 47230
rect 74462 47230 74468 47262
rect 74664 47470 74670 47502
rect 74734 47502 74735 47534
rect 75480 47534 75556 47540
rect 74734 47470 74740 47502
rect 74664 47262 74740 47470
rect 74462 47198 74463 47230
rect 74397 47197 74463 47198
rect 74664 47198 74670 47262
rect 74734 47198 74740 47262
rect 75480 47470 75486 47534
rect 75550 47470 75556 47534
rect 75480 47262 75556 47470
rect 75480 47230 75486 47262
rect 74664 47192 74740 47198
rect 75485 47198 75486 47230
rect 75550 47230 75556 47262
rect 94656 47534 95004 49102
rect 94656 47470 94662 47534
rect 94726 47470 95004 47534
rect 75550 47198 75551 47230
rect 75485 47197 75551 47198
rect 20405 47126 20471 47127
rect 20405 47094 20406 47126
rect 20400 47062 20406 47094
rect 20470 47094 20471 47126
rect 20813 47126 20879 47127
rect 20813 47094 20814 47126
rect 20470 47062 20476 47094
rect 20400 46854 20476 47062
rect 20400 46790 20406 46854
rect 20470 46790 20476 46854
rect 20400 46784 20476 46790
rect 20808 47062 20814 47094
rect 20878 47094 20879 47126
rect 21488 47126 21564 47132
rect 20878 47062 20884 47094
rect 20808 46854 20884 47062
rect 20808 46790 20814 46854
rect 20878 46790 20884 46854
rect 21488 47062 21494 47126
rect 21558 47062 21564 47126
rect 21488 46854 21564 47062
rect 21488 46822 21494 46854
rect 20808 46784 20884 46790
rect 21493 46790 21494 46822
rect 21558 46822 21564 46854
rect 21624 47126 21700 47132
rect 21624 47062 21630 47126
rect 21694 47062 21700 47126
rect 22037 47126 22103 47127
rect 22037 47094 22038 47126
rect 21624 46854 21700 47062
rect 21624 46822 21630 46854
rect 21558 46790 21559 46822
rect 21493 46789 21559 46790
rect 21629 46790 21630 46822
rect 21694 46822 21700 46854
rect 22032 47062 22038 47094
rect 22102 47094 22103 47126
rect 73848 47126 73924 47132
rect 22102 47062 22108 47094
rect 22032 46854 22108 47062
rect 21694 46790 21695 46822
rect 21629 46789 21695 46790
rect 22032 46790 22038 46854
rect 22102 46790 22108 46854
rect 73848 47062 73854 47126
rect 73918 47062 73924 47126
rect 74261 47126 74327 47127
rect 74261 47094 74262 47126
rect 73848 46854 73924 47062
rect 73848 46822 73854 46854
rect 22032 46784 22108 46790
rect 73853 46790 73854 46822
rect 73918 46822 73924 46854
rect 74256 47062 74262 47094
rect 74326 47094 74327 47126
rect 74800 47126 74876 47132
rect 74326 47062 74332 47094
rect 74256 46854 74332 47062
rect 73918 46790 73919 46822
rect 73853 46789 73919 46790
rect 74256 46790 74262 46854
rect 74326 46790 74332 46854
rect 74800 47062 74806 47126
rect 74870 47062 74876 47126
rect 74800 46854 74876 47062
rect 74800 46822 74806 46854
rect 74256 46784 74332 46790
rect 74805 46790 74806 46822
rect 74870 46822 74876 46854
rect 74936 47126 75012 47132
rect 74936 47062 74942 47126
rect 75006 47062 75012 47126
rect 75621 47126 75687 47127
rect 75621 47094 75622 47126
rect 74936 46854 75012 47062
rect 74936 46822 74942 46854
rect 74870 46790 74871 46822
rect 74805 46789 74871 46790
rect 74941 46790 74942 46822
rect 75006 46822 75012 46854
rect 75616 47062 75622 47094
rect 75686 47094 75687 47126
rect 75686 47062 75692 47094
rect 75616 46854 75692 47062
rect 75006 46790 75007 46822
rect 74941 46789 75007 46790
rect 75616 46790 75622 46854
rect 75686 46790 75692 46854
rect 75616 46784 75692 46790
rect 20813 46718 20879 46719
rect 20813 46686 20814 46718
rect 20808 46654 20814 46686
rect 20878 46686 20879 46718
rect 21760 46718 21836 46724
rect 20878 46654 20884 46686
rect 20808 46446 20884 46654
rect 20808 46382 20814 46446
rect 20878 46382 20884 46446
rect 21760 46654 21766 46718
rect 21830 46654 21836 46718
rect 22173 46718 22239 46719
rect 22173 46686 22174 46718
rect 21760 46446 21836 46654
rect 21760 46414 21766 46446
rect 20808 46376 20884 46382
rect 21765 46382 21766 46414
rect 21830 46414 21836 46446
rect 22168 46654 22174 46686
rect 22238 46686 22239 46718
rect 73984 46718 74060 46724
rect 22238 46654 22244 46686
rect 22168 46446 22244 46654
rect 73984 46654 73990 46718
rect 74054 46654 74060 46718
rect 68957 46582 69023 46583
rect 68957 46550 68958 46582
rect 21830 46382 21831 46414
rect 21765 46381 21831 46382
rect 22168 46382 22174 46446
rect 22238 46382 22244 46446
rect 22168 46376 22244 46382
rect 68952 46518 68958 46550
rect 69022 46550 69023 46582
rect 69022 46518 69028 46550
rect 21765 46310 21831 46311
rect 21765 46278 21766 46310
rect 21760 46246 21766 46278
rect 21830 46278 21831 46310
rect 22032 46310 22108 46316
rect 21830 46246 21836 46278
rect 21760 46038 21836 46246
rect 21760 45974 21766 46038
rect 21830 45974 21836 46038
rect 22032 46246 22038 46310
rect 22102 46246 22108 46310
rect 22032 46038 22108 46246
rect 68952 46310 69028 46518
rect 73984 46446 74060 46654
rect 73984 46414 73990 46446
rect 73989 46382 73990 46414
rect 74054 46414 74060 46446
rect 74256 46718 74332 46724
rect 74256 46654 74262 46718
rect 74326 46654 74332 46718
rect 74256 46446 74332 46654
rect 74256 46414 74262 46446
rect 74054 46382 74055 46414
rect 73989 46381 74055 46382
rect 74261 46382 74262 46414
rect 74326 46414 74332 46446
rect 74664 46718 74740 46724
rect 74664 46654 74670 46718
rect 74734 46654 74740 46718
rect 74664 46446 74740 46654
rect 74664 46414 74670 46446
rect 74326 46382 74327 46414
rect 74261 46381 74327 46382
rect 74669 46382 74670 46414
rect 74734 46414 74740 46446
rect 74734 46382 74735 46414
rect 74669 46381 74735 46382
rect 68952 46246 68958 46310
rect 69022 46246 69028 46310
rect 73989 46310 74055 46311
rect 73989 46278 73990 46310
rect 68952 46240 69028 46246
rect 73984 46246 73990 46278
rect 74054 46278 74055 46310
rect 74261 46310 74327 46311
rect 74261 46278 74262 46310
rect 74054 46246 74060 46278
rect 22032 46006 22038 46038
rect 21760 45968 21836 45974
rect 22037 45974 22038 46006
rect 22102 46006 22108 46038
rect 68952 46038 69028 46044
rect 22102 45974 22103 46006
rect 22037 45973 22103 45974
rect 68952 45974 68958 46038
rect 69022 45974 69028 46038
rect 952 45838 1230 45902
rect 1294 45838 1300 45902
rect 952 43998 1300 45838
rect 21488 45902 21564 45908
rect 21488 45838 21494 45902
rect 21558 45838 21564 45902
rect 20541 45630 20607 45631
rect 20541 45598 20542 45630
rect 20536 45566 20542 45598
rect 20606 45598 20607 45630
rect 21488 45630 21564 45838
rect 68952 45766 69028 45974
rect 73984 46038 74060 46246
rect 73984 45974 73990 46038
rect 74054 45974 74060 46038
rect 73984 45968 74060 45974
rect 74256 46246 74262 46278
rect 74326 46278 74327 46310
rect 74326 46246 74332 46278
rect 74256 46038 74332 46246
rect 74256 45974 74262 46038
rect 74326 45974 74332 46038
rect 74256 45968 74332 45974
rect 74805 45902 74871 45903
rect 74805 45870 74806 45902
rect 74800 45838 74806 45870
rect 74870 45870 74871 45902
rect 74941 45902 75007 45903
rect 74941 45870 74942 45902
rect 74870 45838 74876 45870
rect 68952 45734 68958 45766
rect 68957 45702 68958 45734
rect 69022 45734 69028 45766
rect 69093 45766 69159 45767
rect 69093 45734 69094 45766
rect 69022 45702 69023 45734
rect 68957 45701 69023 45702
rect 69088 45702 69094 45734
rect 69158 45734 69159 45766
rect 69158 45702 69164 45734
rect 21488 45598 21494 45630
rect 20606 45566 20612 45598
rect 20536 45358 20612 45566
rect 21493 45566 21494 45598
rect 21558 45598 21564 45630
rect 21558 45566 21559 45598
rect 21493 45565 21559 45566
rect 20536 45294 20542 45358
rect 20606 45294 20612 45358
rect 20536 45288 20612 45294
rect 21080 45494 21156 45500
rect 21080 45430 21086 45494
rect 21150 45430 21156 45494
rect 20541 45222 20607 45223
rect 20541 45190 20542 45222
rect 20536 45158 20542 45190
rect 20606 45190 20607 45222
rect 21080 45222 21156 45430
rect 69088 45494 69164 45702
rect 74800 45630 74876 45838
rect 74800 45566 74806 45630
rect 74870 45566 74876 45630
rect 74800 45560 74876 45566
rect 74936 45838 74942 45870
rect 75006 45870 75007 45902
rect 94656 45902 95004 47470
rect 75006 45838 75012 45870
rect 74936 45630 75012 45838
rect 94656 45838 94662 45902
rect 94726 45838 95004 45902
rect 74936 45566 74942 45630
rect 75006 45566 75012 45630
rect 74936 45560 75012 45566
rect 75480 45630 75556 45636
rect 75480 45566 75486 45630
rect 75550 45566 75556 45630
rect 69088 45430 69094 45494
rect 69158 45430 69164 45494
rect 74533 45494 74599 45495
rect 74533 45462 74534 45494
rect 69088 45424 69164 45430
rect 74528 45430 74534 45462
rect 74598 45462 74599 45494
rect 74598 45430 74604 45462
rect 27200 45358 27276 45364
rect 27200 45294 27206 45358
rect 27270 45294 27276 45358
rect 68957 45358 69023 45359
rect 68957 45326 68958 45358
rect 21080 45190 21086 45222
rect 20606 45158 20612 45190
rect 20536 44950 20612 45158
rect 21085 45158 21086 45190
rect 21150 45190 21156 45222
rect 21357 45222 21423 45223
rect 21357 45190 21358 45222
rect 21150 45158 21151 45190
rect 21085 45157 21151 45158
rect 21352 45158 21358 45190
rect 21422 45190 21423 45222
rect 21422 45158 21428 45190
rect 20536 44886 20542 44950
rect 20606 44886 20612 44950
rect 20536 44880 20612 44886
rect 21352 44950 21428 45158
rect 27200 45086 27276 45294
rect 27200 45054 27206 45086
rect 27205 45022 27206 45054
rect 27270 45054 27276 45086
rect 68952 45294 68958 45326
rect 69022 45326 69023 45358
rect 69022 45294 69028 45326
rect 68952 45086 69028 45294
rect 27270 45022 27271 45054
rect 27205 45021 27271 45022
rect 68952 45022 68958 45086
rect 69022 45022 69028 45086
rect 68952 45016 69028 45022
rect 74528 45086 74604 45430
rect 75480 45358 75556 45566
rect 75480 45326 75486 45358
rect 75485 45294 75486 45326
rect 75550 45326 75556 45358
rect 75550 45294 75551 45326
rect 75485 45293 75551 45294
rect 75077 45222 75143 45223
rect 75077 45190 75078 45222
rect 74528 45022 74534 45086
rect 74598 45022 74604 45086
rect 74528 45016 74604 45022
rect 75072 45158 75078 45190
rect 75142 45190 75143 45222
rect 75485 45222 75551 45223
rect 75485 45190 75486 45222
rect 75142 45158 75148 45190
rect 21352 44886 21358 44950
rect 21422 44886 21428 44950
rect 21352 44880 21428 44886
rect 69088 44950 69164 44956
rect 69088 44886 69094 44950
rect 69158 44886 69164 44950
rect 20405 44814 20471 44815
rect 20405 44782 20406 44814
rect 20400 44750 20406 44782
rect 20470 44782 20471 44814
rect 21624 44814 21700 44820
rect 20470 44750 20476 44782
rect 20400 44542 20476 44750
rect 20400 44478 20406 44542
rect 20470 44478 20476 44542
rect 21624 44750 21630 44814
rect 21694 44750 21700 44814
rect 21624 44542 21700 44750
rect 21624 44510 21630 44542
rect 20400 44472 20476 44478
rect 21629 44478 21630 44510
rect 21694 44510 21700 44542
rect 22168 44814 22244 44820
rect 22168 44750 22174 44814
rect 22238 44750 22244 44814
rect 22168 44542 22244 44750
rect 69088 44678 69164 44886
rect 75072 44950 75148 45158
rect 75072 44886 75078 44950
rect 75142 44886 75148 44950
rect 75072 44880 75148 44886
rect 75480 45158 75486 45190
rect 75550 45190 75551 45222
rect 75550 45158 75556 45190
rect 75480 44950 75556 45158
rect 75480 44886 75486 44950
rect 75550 44886 75556 44950
rect 75480 44880 75556 44886
rect 69088 44646 69094 44678
rect 69093 44614 69094 44646
rect 69158 44646 69164 44678
rect 73848 44814 73924 44820
rect 73848 44750 73854 44814
rect 73918 44750 73924 44814
rect 74261 44814 74327 44815
rect 74261 44782 74262 44814
rect 69158 44614 69159 44646
rect 69093 44613 69159 44614
rect 22168 44510 22174 44542
rect 21694 44478 21695 44510
rect 21629 44477 21695 44478
rect 22173 44478 22174 44510
rect 22238 44510 22244 44542
rect 73848 44542 73924 44750
rect 73848 44510 73854 44542
rect 22238 44478 22239 44510
rect 22173 44477 22239 44478
rect 73853 44478 73854 44510
rect 73918 44510 73924 44542
rect 74256 44750 74262 44782
rect 74326 44782 74327 44814
rect 74941 44814 75007 44815
rect 74941 44782 74942 44814
rect 74326 44750 74332 44782
rect 74256 44542 74332 44750
rect 73918 44478 73919 44510
rect 73853 44477 73919 44478
rect 74256 44478 74262 44542
rect 74326 44478 74332 44542
rect 74256 44472 74332 44478
rect 74936 44750 74942 44782
rect 75006 44782 75007 44814
rect 75616 44814 75692 44820
rect 75006 44750 75012 44782
rect 74936 44542 75012 44750
rect 74936 44478 74942 44542
rect 75006 44478 75012 44542
rect 75616 44750 75622 44814
rect 75686 44750 75692 44814
rect 75616 44542 75692 44750
rect 75616 44510 75622 44542
rect 74936 44472 75012 44478
rect 75621 44478 75622 44510
rect 75686 44510 75692 44542
rect 75686 44478 75687 44510
rect 75621 44477 75687 44478
rect 20536 44406 20612 44412
rect 20536 44342 20542 44406
rect 20606 44342 20612 44406
rect 20536 44134 20612 44342
rect 20536 44102 20542 44134
rect 20541 44070 20542 44102
rect 20606 44102 20612 44134
rect 21760 44406 21836 44412
rect 21760 44342 21766 44406
rect 21830 44342 21836 44406
rect 22037 44406 22103 44407
rect 22037 44374 22038 44406
rect 21760 44134 21836 44342
rect 21760 44102 21766 44134
rect 20606 44070 20607 44102
rect 20541 44069 20607 44070
rect 21765 44070 21766 44102
rect 21830 44102 21836 44134
rect 22032 44342 22038 44374
rect 22102 44374 22103 44406
rect 73989 44406 74055 44407
rect 73989 44374 73990 44406
rect 22102 44342 22108 44374
rect 22032 44134 22108 44342
rect 73984 44342 73990 44374
rect 74054 44374 74055 44406
rect 74392 44406 74468 44412
rect 74054 44342 74060 44374
rect 21830 44070 21831 44102
rect 21765 44069 21831 44070
rect 22032 44070 22038 44134
rect 22102 44070 22108 44134
rect 22032 44064 22108 44070
rect 69088 44134 69164 44140
rect 69088 44070 69094 44134
rect 69158 44070 69164 44134
rect 952 43934 1230 43998
rect 1294 43934 1300 43998
rect 952 42366 1300 43934
rect 20400 43998 20476 44004
rect 20400 43934 20406 43998
rect 20470 43934 20476 43998
rect 21085 43998 21151 43999
rect 21085 43966 21086 43998
rect 20400 43726 20476 43934
rect 20400 43694 20406 43726
rect 20405 43662 20406 43694
rect 20470 43694 20476 43726
rect 21080 43934 21086 43966
rect 21150 43966 21151 43998
rect 21765 43998 21831 43999
rect 21765 43966 21766 43998
rect 21150 43934 21156 43966
rect 21080 43726 21156 43934
rect 20470 43662 20471 43694
rect 20405 43661 20471 43662
rect 21080 43662 21086 43726
rect 21150 43662 21156 43726
rect 21080 43656 21156 43662
rect 21760 43934 21766 43966
rect 21830 43966 21831 43998
rect 22032 43998 22108 44004
rect 21830 43934 21836 43966
rect 21760 43726 21836 43934
rect 21760 43662 21766 43726
rect 21830 43662 21836 43726
rect 22032 43934 22038 43998
rect 22102 43934 22108 43998
rect 22032 43726 22108 43934
rect 69088 43862 69164 44070
rect 73984 44134 74060 44342
rect 73984 44070 73990 44134
rect 74054 44070 74060 44134
rect 74392 44342 74398 44406
rect 74462 44342 74468 44406
rect 74669 44406 74735 44407
rect 74669 44374 74670 44406
rect 74392 44134 74468 44342
rect 74392 44102 74398 44134
rect 73984 44064 74060 44070
rect 74397 44070 74398 44102
rect 74462 44102 74468 44134
rect 74664 44342 74670 44374
rect 74734 44374 74735 44406
rect 75485 44406 75551 44407
rect 75485 44374 75486 44406
rect 74734 44342 74740 44374
rect 74664 44134 74740 44342
rect 74462 44070 74463 44102
rect 74397 44069 74463 44070
rect 74664 44070 74670 44134
rect 74734 44070 74740 44134
rect 74664 44064 74740 44070
rect 75480 44342 75486 44374
rect 75550 44374 75551 44406
rect 75550 44342 75556 44374
rect 75480 44134 75556 44342
rect 75480 44070 75486 44134
rect 75550 44070 75556 44134
rect 75480 44064 75556 44070
rect 73989 43998 74055 43999
rect 73989 43966 73990 43998
rect 69088 43830 69094 43862
rect 69093 43798 69094 43830
rect 69158 43830 69164 43862
rect 73984 43934 73990 43966
rect 74054 43966 74055 43998
rect 74397 43998 74463 43999
rect 74397 43966 74398 43998
rect 74054 43934 74060 43966
rect 69158 43798 69159 43830
rect 69093 43797 69159 43798
rect 22032 43694 22038 43726
rect 21760 43656 21836 43662
rect 22037 43662 22038 43694
rect 22102 43694 22108 43726
rect 73984 43726 74060 43934
rect 22102 43662 22103 43694
rect 22037 43661 22103 43662
rect 73984 43662 73990 43726
rect 74054 43662 74060 43726
rect 73984 43656 74060 43662
rect 74392 43934 74398 43966
rect 74462 43966 74463 43998
rect 74800 43998 74876 44004
rect 74462 43934 74468 43966
rect 74392 43726 74468 43934
rect 74392 43662 74398 43726
rect 74462 43662 74468 43726
rect 74800 43934 74806 43998
rect 74870 43934 74876 43998
rect 74800 43726 74876 43934
rect 74800 43694 74806 43726
rect 74392 43656 74468 43662
rect 74805 43662 74806 43694
rect 74870 43694 74876 43726
rect 75616 43998 75692 44004
rect 75616 43934 75622 43998
rect 75686 43934 75692 43998
rect 75616 43726 75692 43934
rect 75616 43694 75622 43726
rect 74870 43662 74871 43694
rect 74805 43661 74871 43662
rect 75621 43662 75622 43694
rect 75686 43694 75692 43726
rect 94656 43998 95004 45838
rect 94656 43934 94662 43998
rect 94726 43934 95004 43998
rect 75686 43662 75687 43694
rect 75621 43661 75687 43662
rect 20400 43590 20476 43596
rect 20400 43526 20406 43590
rect 20470 43526 20476 43590
rect 20400 43318 20476 43526
rect 20400 43286 20406 43318
rect 20405 43254 20406 43286
rect 20470 43286 20476 43318
rect 20944 43590 21020 43596
rect 20944 43526 20950 43590
rect 21014 43526 21020 43590
rect 20944 43318 21020 43526
rect 20944 43286 20950 43318
rect 20470 43254 20471 43286
rect 20405 43253 20471 43254
rect 20949 43254 20950 43286
rect 21014 43286 21020 43318
rect 21080 43590 21156 43596
rect 21080 43526 21086 43590
rect 21150 43526 21156 43590
rect 21080 43318 21156 43526
rect 21080 43286 21086 43318
rect 21014 43254 21015 43286
rect 20949 43253 21015 43254
rect 21085 43254 21086 43286
rect 21150 43286 21156 43318
rect 21760 43590 21836 43596
rect 21760 43526 21766 43590
rect 21830 43526 21836 43590
rect 22037 43590 22103 43591
rect 22037 43558 22038 43590
rect 21760 43318 21836 43526
rect 21760 43286 21766 43318
rect 21150 43254 21151 43286
rect 21085 43253 21151 43254
rect 21765 43254 21766 43286
rect 21830 43286 21836 43318
rect 22032 43526 22038 43558
rect 22102 43558 22103 43590
rect 73984 43590 74060 43596
rect 22102 43526 22108 43558
rect 22032 43318 22108 43526
rect 21830 43254 21831 43286
rect 21765 43253 21831 43254
rect 22032 43254 22038 43318
rect 22102 43254 22108 43318
rect 73984 43526 73990 43590
rect 74054 43526 74060 43590
rect 73984 43318 74060 43526
rect 73984 43286 73990 43318
rect 22032 43248 22108 43254
rect 73989 43254 73990 43286
rect 74054 43286 74060 43318
rect 74256 43590 74332 43596
rect 74256 43526 74262 43590
rect 74326 43526 74332 43590
rect 74256 43318 74332 43526
rect 74256 43286 74262 43318
rect 74054 43254 74055 43286
rect 73989 43253 74055 43254
rect 74261 43254 74262 43286
rect 74326 43286 74332 43318
rect 74664 43590 74740 43596
rect 74664 43526 74670 43590
rect 74734 43526 74740 43590
rect 75621 43590 75687 43591
rect 75621 43558 75622 43590
rect 74664 43318 74740 43526
rect 74664 43286 74670 43318
rect 74326 43254 74327 43286
rect 74261 43253 74327 43254
rect 74669 43254 74670 43286
rect 74734 43286 74740 43318
rect 75616 43526 75622 43558
rect 75686 43558 75687 43590
rect 75686 43526 75692 43558
rect 75616 43318 75692 43526
rect 74734 43254 74735 43286
rect 74669 43253 74735 43254
rect 75616 43254 75622 43318
rect 75686 43254 75692 43318
rect 75616 43248 75692 43254
rect 20536 43182 20612 43188
rect 20536 43118 20542 43182
rect 20606 43118 20612 43182
rect 21221 43182 21287 43183
rect 21221 43150 21222 43182
rect 20536 42910 20612 43118
rect 20536 42878 20542 42910
rect 20541 42846 20542 42878
rect 20606 42878 20612 42910
rect 21216 43118 21222 43150
rect 21286 43150 21287 43182
rect 21765 43182 21831 43183
rect 21765 43150 21766 43182
rect 21286 43118 21292 43150
rect 21216 42910 21292 43118
rect 20606 42846 20607 42878
rect 20541 42845 20607 42846
rect 21216 42846 21222 42910
rect 21286 42846 21292 42910
rect 21216 42840 21292 42846
rect 21760 43118 21766 43150
rect 21830 43150 21831 43182
rect 22168 43182 22244 43188
rect 21830 43118 21836 43150
rect 21760 42910 21836 43118
rect 21760 42846 21766 42910
rect 21830 42846 21836 42910
rect 22168 43118 22174 43182
rect 22238 43118 22244 43182
rect 73989 43182 74055 43183
rect 73989 43150 73990 43182
rect 22168 42910 22244 43118
rect 73984 43118 73990 43150
rect 74054 43150 74055 43182
rect 74261 43182 74327 43183
rect 74261 43150 74262 43182
rect 74054 43118 74060 43150
rect 22168 42878 22174 42910
rect 21760 42840 21836 42846
rect 22173 42846 22174 42878
rect 22238 42878 22244 42910
rect 25432 42910 25508 42916
rect 22238 42846 22239 42878
rect 22173 42845 22239 42846
rect 25432 42846 25438 42910
rect 25502 42846 25508 42910
rect 20808 42774 20884 42780
rect 20808 42710 20814 42774
rect 20878 42710 20884 42774
rect 21357 42774 21423 42775
rect 21357 42742 21358 42774
rect 20808 42502 20884 42710
rect 20808 42470 20814 42502
rect 20813 42438 20814 42470
rect 20878 42470 20884 42502
rect 21352 42710 21358 42742
rect 21422 42742 21423 42774
rect 21624 42774 21700 42780
rect 21422 42710 21428 42742
rect 21352 42502 21428 42710
rect 20878 42438 20879 42470
rect 20813 42437 20879 42438
rect 21352 42438 21358 42502
rect 21422 42438 21428 42502
rect 21624 42710 21630 42774
rect 21694 42710 21700 42774
rect 22037 42774 22103 42775
rect 22037 42742 22038 42774
rect 21624 42502 21700 42710
rect 21624 42470 21630 42502
rect 21352 42432 21428 42438
rect 21629 42438 21630 42470
rect 21694 42470 21700 42502
rect 22032 42710 22038 42742
rect 22102 42742 22103 42774
rect 22102 42710 22108 42742
rect 22032 42502 22108 42710
rect 21694 42438 21695 42470
rect 21629 42437 21695 42438
rect 22032 42438 22038 42502
rect 22102 42438 22108 42502
rect 25432 42502 25508 42846
rect 73984 42910 74060 43118
rect 73984 42846 73990 42910
rect 74054 42846 74060 42910
rect 73984 42840 74060 42846
rect 74256 43118 74262 43150
rect 74326 43150 74327 43182
rect 74669 43182 74735 43183
rect 74669 43150 74670 43182
rect 74326 43118 74332 43150
rect 74256 42910 74332 43118
rect 74256 42846 74262 42910
rect 74326 42846 74332 42910
rect 74256 42840 74332 42846
rect 74664 43118 74670 43150
rect 74734 43150 74735 43182
rect 75072 43182 75148 43188
rect 74734 43118 74740 43150
rect 74664 42910 74740 43118
rect 74664 42846 74670 42910
rect 74734 42846 74740 42910
rect 75072 43118 75078 43182
rect 75142 43118 75148 43182
rect 75485 43182 75551 43183
rect 75485 43150 75486 43182
rect 75072 42910 75148 43118
rect 75072 42878 75078 42910
rect 74664 42840 74740 42846
rect 75077 42846 75078 42878
rect 75142 42878 75148 42910
rect 75480 43118 75486 43150
rect 75550 43150 75551 43182
rect 75550 43118 75556 43150
rect 75480 42910 75556 43118
rect 75142 42846 75143 42878
rect 75077 42845 75143 42846
rect 75480 42846 75486 42910
rect 75550 42846 75556 42910
rect 75480 42840 75556 42846
rect 73304 42774 73380 42780
rect 73304 42710 73310 42774
rect 73374 42710 73380 42774
rect 25432 42470 25438 42502
rect 22032 42432 22108 42438
rect 25437 42438 25438 42470
rect 25502 42470 25508 42502
rect 69088 42638 69164 42644
rect 69088 42574 69094 42638
rect 69158 42574 69164 42638
rect 25502 42438 25503 42470
rect 25437 42437 25503 42438
rect 952 42302 1230 42366
rect 1294 42302 1300 42366
rect 952 40598 1300 42302
rect 21760 42366 21836 42372
rect 21760 42302 21766 42366
rect 21830 42302 21836 42366
rect 22173 42366 22239 42367
rect 22173 42334 22174 42366
rect 21760 42094 21836 42302
rect 21760 42062 21766 42094
rect 21765 42030 21766 42062
rect 21830 42062 21836 42094
rect 22168 42302 22174 42334
rect 22238 42334 22239 42366
rect 69088 42366 69164 42574
rect 73304 42502 73380 42710
rect 73304 42470 73310 42502
rect 73309 42438 73310 42470
rect 73374 42470 73380 42502
rect 73848 42774 73924 42780
rect 73848 42710 73854 42774
rect 73918 42710 73924 42774
rect 74261 42774 74327 42775
rect 74261 42742 74262 42774
rect 73848 42502 73924 42710
rect 73848 42470 73854 42502
rect 73374 42438 73375 42470
rect 73309 42437 73375 42438
rect 73853 42438 73854 42470
rect 73918 42470 73924 42502
rect 74256 42710 74262 42742
rect 74326 42742 74327 42774
rect 74941 42774 75007 42775
rect 74941 42742 74942 42774
rect 74326 42710 74332 42742
rect 74256 42502 74332 42710
rect 73918 42438 73919 42470
rect 73853 42437 73919 42438
rect 74256 42438 74262 42502
rect 74326 42438 74332 42502
rect 74256 42432 74332 42438
rect 74936 42710 74942 42742
rect 75006 42742 75007 42774
rect 75006 42710 75012 42742
rect 74936 42502 75012 42710
rect 74936 42438 74942 42502
rect 75006 42438 75012 42502
rect 74936 42432 75012 42438
rect 69088 42334 69094 42366
rect 22238 42302 22244 42334
rect 22168 42094 22244 42302
rect 69093 42302 69094 42334
rect 69158 42334 69164 42366
rect 73853 42366 73919 42367
rect 73853 42334 73854 42366
rect 69158 42302 69159 42334
rect 69093 42301 69159 42302
rect 73848 42302 73854 42334
rect 73918 42334 73919 42366
rect 74256 42366 74332 42372
rect 74838 42367 75148 42372
rect 73918 42302 73924 42334
rect 21830 42030 21831 42062
rect 21765 42029 21831 42030
rect 22168 42030 22174 42094
rect 22238 42030 22244 42094
rect 22168 42024 22244 42030
rect 73848 42094 73924 42302
rect 73848 42030 73854 42094
rect 73918 42030 73924 42094
rect 74256 42302 74262 42366
rect 74326 42302 74332 42366
rect 74256 42094 74332 42302
rect 74805 42366 75148 42367
rect 74805 42302 74806 42366
rect 74870 42302 75078 42366
rect 75142 42302 75148 42366
rect 74805 42301 75148 42302
rect 74838 42296 75148 42301
rect 94656 42366 95004 43934
rect 94656 42302 94662 42366
rect 94726 42302 95004 42366
rect 74256 42062 74262 42094
rect 73848 42024 73924 42030
rect 74261 42030 74262 42062
rect 74326 42062 74332 42094
rect 74326 42030 74327 42062
rect 74261 42029 74327 42030
rect 21085 41958 21151 41959
rect 21085 41926 21086 41958
rect 21080 41894 21086 41926
rect 21150 41926 21151 41958
rect 21765 41958 21831 41959
rect 21765 41926 21766 41958
rect 21150 41894 21156 41926
rect 20536 41686 20612 41692
rect 20536 41622 20542 41686
rect 20606 41622 20612 41686
rect 20536 41414 20612 41622
rect 21080 41686 21156 41894
rect 21080 41622 21086 41686
rect 21150 41622 21156 41686
rect 21080 41616 21156 41622
rect 21760 41894 21766 41926
rect 21830 41926 21831 41958
rect 22032 41958 22108 41964
rect 21830 41894 21836 41926
rect 21760 41686 21836 41894
rect 21760 41622 21766 41686
rect 21830 41622 21836 41686
rect 22032 41894 22038 41958
rect 22102 41894 22108 41958
rect 22032 41686 22108 41894
rect 22032 41654 22038 41686
rect 21760 41616 21836 41622
rect 22037 41622 22038 41654
rect 22102 41654 22108 41686
rect 73848 41958 73924 41964
rect 73848 41894 73854 41958
rect 73918 41894 73924 41958
rect 73848 41686 73924 41894
rect 73848 41654 73854 41686
rect 22102 41622 22103 41654
rect 22037 41621 22103 41622
rect 73853 41622 73854 41654
rect 73918 41654 73924 41686
rect 74256 41958 74332 41964
rect 74256 41894 74262 41958
rect 74326 41894 74332 41958
rect 74256 41686 74332 41894
rect 74256 41654 74262 41686
rect 73918 41622 73919 41654
rect 73853 41621 73919 41622
rect 74261 41622 74262 41654
rect 74326 41654 74332 41686
rect 74936 41958 75012 41964
rect 74936 41894 74942 41958
rect 75006 41894 75012 41958
rect 74936 41686 75012 41894
rect 74936 41654 74942 41686
rect 74326 41622 74327 41654
rect 74261 41621 74327 41622
rect 74941 41622 74942 41654
rect 75006 41654 75012 41686
rect 75616 41686 75692 41692
rect 75006 41622 75007 41654
rect 74941 41621 75007 41622
rect 75616 41622 75622 41686
rect 75686 41622 75692 41686
rect 20536 41382 20542 41414
rect 20541 41350 20542 41382
rect 20606 41382 20612 41414
rect 27064 41414 27140 41420
rect 20606 41350 20607 41382
rect 20541 41349 20607 41350
rect 27064 41350 27070 41414
rect 27134 41350 27140 41414
rect 69093 41414 69159 41415
rect 69093 41382 69094 41414
rect 20541 41278 20607 41279
rect 20541 41246 20542 41278
rect 20536 41214 20542 41246
rect 20606 41246 20607 41278
rect 21488 41278 21564 41284
rect 20606 41214 20612 41246
rect 20536 41006 20612 41214
rect 20536 40942 20542 41006
rect 20606 40942 20612 41006
rect 21488 41214 21494 41278
rect 21558 41214 21564 41278
rect 21488 41006 21564 41214
rect 27064 41142 27140 41350
rect 27064 41110 27070 41142
rect 27069 41078 27070 41110
rect 27134 41110 27140 41142
rect 69088 41350 69094 41382
rect 69158 41382 69159 41414
rect 75616 41414 75692 41622
rect 75616 41382 75622 41414
rect 69158 41350 69164 41382
rect 69088 41142 69164 41350
rect 75621 41350 75622 41382
rect 75686 41382 75692 41414
rect 75686 41350 75687 41382
rect 75621 41349 75687 41350
rect 75213 41278 75279 41279
rect 75213 41246 75214 41278
rect 27134 41078 27135 41110
rect 27069 41077 27135 41078
rect 69088 41078 69094 41142
rect 69158 41078 69164 41142
rect 69088 41072 69164 41078
rect 75208 41214 75214 41246
rect 75278 41246 75279 41278
rect 75621 41278 75687 41279
rect 75621 41246 75622 41278
rect 75278 41214 75284 41246
rect 21488 40974 21494 41006
rect 20536 40936 20612 40942
rect 21493 40942 21494 40974
rect 21558 40974 21564 41006
rect 27200 41006 27276 41012
rect 21558 40942 21559 40974
rect 21493 40941 21559 40942
rect 27200 40942 27206 41006
rect 27270 40942 27276 41006
rect 68957 41006 69023 41007
rect 68957 40974 68958 41006
rect 952 40534 1230 40598
rect 1294 40534 1300 40598
rect 20400 40870 20476 40876
rect 20400 40806 20406 40870
rect 20470 40806 20476 40870
rect 21765 40870 21831 40871
rect 21765 40838 21766 40870
rect 20400 40598 20476 40806
rect 20400 40566 20406 40598
rect 952 38966 1300 40534
rect 20405 40534 20406 40566
rect 20470 40566 20476 40598
rect 21760 40806 21766 40838
rect 21830 40838 21831 40870
rect 22173 40870 22239 40871
rect 22173 40838 22174 40870
rect 21830 40806 21836 40838
rect 21760 40598 21836 40806
rect 20470 40534 20471 40566
rect 20405 40533 20471 40534
rect 21760 40534 21766 40598
rect 21830 40534 21836 40598
rect 21760 40528 21836 40534
rect 22168 40806 22174 40838
rect 22238 40838 22239 40870
rect 22238 40806 22244 40838
rect 22168 40598 22244 40806
rect 27200 40734 27276 40942
rect 27200 40702 27206 40734
rect 27205 40670 27206 40702
rect 27270 40702 27276 40734
rect 68952 40942 68958 40974
rect 69022 40974 69023 41006
rect 75208 41006 75284 41214
rect 69022 40942 69028 40974
rect 68952 40734 69028 40942
rect 75208 40942 75214 41006
rect 75278 40942 75284 41006
rect 75208 40936 75284 40942
rect 75616 41214 75622 41246
rect 75686 41246 75687 41278
rect 75686 41214 75692 41246
rect 75616 41006 75692 41214
rect 75616 40942 75622 41006
rect 75686 40942 75692 41006
rect 75616 40936 75692 40942
rect 27270 40670 27271 40702
rect 27205 40669 27271 40670
rect 68952 40670 68958 40734
rect 69022 40670 69028 40734
rect 68952 40664 69028 40670
rect 73848 40870 73924 40876
rect 73848 40806 73854 40870
rect 73918 40806 73924 40870
rect 22168 40534 22174 40598
rect 22238 40534 22244 40598
rect 73848 40598 73924 40806
rect 73848 40566 73854 40598
rect 22168 40528 22244 40534
rect 73853 40534 73854 40566
rect 73918 40566 73924 40598
rect 74256 40870 74332 40876
rect 74256 40806 74262 40870
rect 74326 40806 74332 40870
rect 74256 40598 74332 40806
rect 74256 40566 74262 40598
rect 73918 40534 73919 40566
rect 73853 40533 73919 40534
rect 74261 40534 74262 40566
rect 74326 40566 74332 40598
rect 75616 40870 75692 40876
rect 75616 40806 75622 40870
rect 75686 40806 75692 40870
rect 75616 40598 75692 40806
rect 75616 40566 75622 40598
rect 74326 40534 74327 40566
rect 74261 40533 74327 40534
rect 75621 40534 75622 40566
rect 75686 40566 75692 40598
rect 94656 40734 95004 42302
rect 94656 40670 94662 40734
rect 94726 40670 95004 40734
rect 75686 40534 75687 40566
rect 75621 40533 75687 40534
rect 20536 40462 20612 40468
rect 20536 40398 20542 40462
rect 20606 40398 20612 40462
rect 20536 40190 20612 40398
rect 20536 40158 20542 40190
rect 20541 40126 20542 40158
rect 20606 40158 20612 40190
rect 21216 40462 21292 40468
rect 21216 40398 21222 40462
rect 21286 40398 21292 40462
rect 21216 40190 21292 40398
rect 21216 40158 21222 40190
rect 20606 40126 20607 40158
rect 20541 40125 20607 40126
rect 21221 40126 21222 40158
rect 21286 40158 21292 40190
rect 21624 40462 21700 40468
rect 21624 40398 21630 40462
rect 21694 40398 21700 40462
rect 21624 40190 21700 40398
rect 21624 40158 21630 40190
rect 21286 40126 21287 40158
rect 21221 40125 21287 40126
rect 21629 40126 21630 40158
rect 21694 40158 21700 40190
rect 22168 40462 22244 40468
rect 22168 40398 22174 40462
rect 22238 40398 22244 40462
rect 22168 40190 22244 40398
rect 73848 40462 73924 40468
rect 73848 40398 73854 40462
rect 73918 40398 73924 40462
rect 74261 40462 74327 40463
rect 74261 40430 74262 40462
rect 22168 40158 22174 40190
rect 21694 40126 21695 40158
rect 21629 40125 21695 40126
rect 22173 40126 22174 40158
rect 22238 40158 22244 40190
rect 69093 40190 69159 40191
rect 69093 40158 69094 40190
rect 22238 40126 22239 40158
rect 22173 40125 22239 40126
rect 69088 40126 69094 40158
rect 69158 40158 69159 40190
rect 73848 40190 73924 40398
rect 73848 40158 73854 40190
rect 69158 40126 69164 40158
rect 20536 40054 20612 40060
rect 20536 39990 20542 40054
rect 20606 39990 20612 40054
rect 20949 40054 21015 40055
rect 20949 40022 20950 40054
rect 20536 39782 20612 39990
rect 20536 39750 20542 39782
rect 20541 39718 20542 39750
rect 20606 39750 20612 39782
rect 20944 39990 20950 40022
rect 21014 40022 21015 40054
rect 21765 40054 21831 40055
rect 21765 40022 21766 40054
rect 21014 39990 21020 40022
rect 20944 39782 21020 39990
rect 20606 39718 20607 39750
rect 20541 39717 20607 39718
rect 20944 39718 20950 39782
rect 21014 39718 21020 39782
rect 20944 39712 21020 39718
rect 21760 39990 21766 40022
rect 21830 40022 21831 40054
rect 22037 40054 22103 40055
rect 22037 40022 22038 40054
rect 21830 39990 21836 40022
rect 21760 39782 21836 39990
rect 21760 39718 21766 39782
rect 21830 39718 21836 39782
rect 21760 39712 21836 39718
rect 22032 39990 22038 40022
rect 22102 40022 22103 40054
rect 22102 39990 22108 40022
rect 22032 39782 22108 39990
rect 69088 39918 69164 40126
rect 73853 40126 73854 40158
rect 73918 40158 73924 40190
rect 74256 40398 74262 40430
rect 74326 40430 74327 40462
rect 75213 40462 75279 40463
rect 75213 40430 75214 40462
rect 74326 40398 74332 40430
rect 74256 40190 74332 40398
rect 73918 40126 73919 40158
rect 73853 40125 73919 40126
rect 74256 40126 74262 40190
rect 74326 40126 74332 40190
rect 74256 40120 74332 40126
rect 75208 40398 75214 40430
rect 75278 40430 75279 40462
rect 75621 40462 75687 40463
rect 75621 40430 75622 40462
rect 75278 40398 75284 40430
rect 75208 40190 75284 40398
rect 75208 40126 75214 40190
rect 75278 40126 75284 40190
rect 75208 40120 75284 40126
rect 75616 40398 75622 40430
rect 75686 40430 75687 40462
rect 75686 40398 75692 40430
rect 75616 40190 75692 40398
rect 75616 40126 75622 40190
rect 75686 40126 75692 40190
rect 75616 40120 75692 40126
rect 73989 40054 74055 40055
rect 73989 40022 73990 40054
rect 69088 39854 69094 39918
rect 69158 39854 69164 39918
rect 69088 39848 69164 39854
rect 73984 39990 73990 40022
rect 74054 40022 74055 40054
rect 74261 40054 74327 40055
rect 74261 40022 74262 40054
rect 74054 39990 74060 40022
rect 22032 39718 22038 39782
rect 22102 39718 22108 39782
rect 22032 39712 22108 39718
rect 73984 39782 74060 39990
rect 73984 39718 73990 39782
rect 74054 39718 74060 39782
rect 73984 39712 74060 39718
rect 74256 39990 74262 40022
rect 74326 40022 74327 40054
rect 74669 40054 74735 40055
rect 74669 40022 74670 40054
rect 74326 39990 74332 40022
rect 74256 39782 74332 39990
rect 74256 39718 74262 39782
rect 74326 39718 74332 39782
rect 74256 39712 74332 39718
rect 74664 39990 74670 40022
rect 74734 40022 74735 40054
rect 75213 40054 75279 40055
rect 75213 40022 75214 40054
rect 74734 39990 74740 40022
rect 74664 39782 74740 39990
rect 74664 39718 74670 39782
rect 74734 39718 74740 39782
rect 74664 39712 74740 39718
rect 75208 39990 75214 40022
rect 75278 40022 75279 40054
rect 75485 40054 75551 40055
rect 75485 40022 75486 40054
rect 75278 39990 75284 40022
rect 75208 39782 75284 39990
rect 75208 39718 75214 39782
rect 75278 39718 75284 39782
rect 75208 39712 75284 39718
rect 75480 39990 75486 40022
rect 75550 40022 75551 40054
rect 75550 39990 75556 40022
rect 75480 39782 75556 39990
rect 75480 39718 75486 39782
rect 75550 39718 75556 39782
rect 75480 39712 75556 39718
rect 20541 39646 20607 39647
rect 20541 39614 20542 39646
rect 20536 39582 20542 39614
rect 20606 39614 20607 39646
rect 20808 39646 20884 39652
rect 20606 39582 20612 39614
rect 20536 39374 20612 39582
rect 20536 39310 20542 39374
rect 20606 39310 20612 39374
rect 20808 39582 20814 39646
rect 20878 39582 20884 39646
rect 21765 39646 21831 39647
rect 21765 39614 21766 39646
rect 20808 39374 20884 39582
rect 20808 39342 20814 39374
rect 20536 39304 20612 39310
rect 20813 39310 20814 39342
rect 20878 39342 20884 39374
rect 21760 39582 21766 39614
rect 21830 39614 21831 39646
rect 22173 39646 22239 39647
rect 22173 39614 22174 39646
rect 21830 39582 21836 39614
rect 21760 39374 21836 39582
rect 20878 39310 20879 39342
rect 20813 39309 20879 39310
rect 21760 39310 21766 39374
rect 21830 39310 21836 39374
rect 21760 39304 21836 39310
rect 22168 39582 22174 39614
rect 22238 39614 22239 39646
rect 73989 39646 74055 39647
rect 73989 39614 73990 39646
rect 22238 39582 22244 39614
rect 22168 39374 22244 39582
rect 22168 39310 22174 39374
rect 22238 39310 22244 39374
rect 22168 39304 22244 39310
rect 73984 39582 73990 39614
rect 74054 39614 74055 39646
rect 74256 39646 74332 39652
rect 74054 39582 74060 39614
rect 73984 39374 74060 39582
rect 73984 39310 73990 39374
rect 74054 39310 74060 39374
rect 74256 39582 74262 39646
rect 74326 39582 74332 39646
rect 74669 39646 74735 39647
rect 74669 39614 74670 39646
rect 74256 39374 74332 39582
rect 74256 39342 74262 39374
rect 73984 39304 74060 39310
rect 74261 39310 74262 39342
rect 74326 39342 74332 39374
rect 74664 39582 74670 39614
rect 74734 39614 74735 39646
rect 74936 39646 75012 39652
rect 74734 39582 74740 39614
rect 74664 39374 74740 39582
rect 74326 39310 74327 39342
rect 74261 39309 74327 39310
rect 74664 39310 74670 39374
rect 74734 39310 74740 39374
rect 74936 39582 74942 39646
rect 75006 39582 75012 39646
rect 74936 39374 75012 39582
rect 74936 39342 74942 39374
rect 74664 39304 74740 39310
rect 74941 39310 74942 39342
rect 75006 39342 75012 39374
rect 75208 39646 75284 39652
rect 75208 39582 75214 39646
rect 75278 39582 75284 39646
rect 75208 39374 75284 39582
rect 75208 39342 75214 39374
rect 75006 39310 75007 39342
rect 74941 39309 75007 39310
rect 75213 39310 75214 39342
rect 75278 39342 75284 39374
rect 75616 39646 75692 39652
rect 75616 39582 75622 39646
rect 75686 39582 75692 39646
rect 75616 39374 75692 39582
rect 75616 39342 75622 39374
rect 75278 39310 75279 39342
rect 75213 39309 75279 39310
rect 75621 39310 75622 39342
rect 75686 39342 75692 39374
rect 75686 39310 75687 39342
rect 75621 39309 75687 39310
rect 952 38902 1230 38966
rect 1294 38902 1300 38966
rect 20400 39238 20476 39244
rect 20400 39174 20406 39238
rect 20470 39174 20476 39238
rect 20813 39238 20879 39239
rect 20813 39206 20814 39238
rect 20400 38966 20476 39174
rect 20400 38934 20406 38966
rect 952 37470 1300 38902
rect 20405 38902 20406 38934
rect 20470 38934 20476 38966
rect 20808 39174 20814 39206
rect 20878 39206 20879 39238
rect 21080 39238 21156 39244
rect 20878 39174 20884 39206
rect 20808 38966 20884 39174
rect 20470 38902 20471 38934
rect 20405 38901 20471 38902
rect 20808 38902 20814 38966
rect 20878 38902 20884 38966
rect 21080 39174 21086 39238
rect 21150 39174 21156 39238
rect 21629 39238 21695 39239
rect 21629 39206 21630 39238
rect 21080 38966 21156 39174
rect 21080 38934 21086 38966
rect 20808 38896 20884 38902
rect 21085 38902 21086 38934
rect 21150 38934 21156 38966
rect 21624 39174 21630 39206
rect 21694 39206 21695 39238
rect 22032 39238 22108 39244
rect 21694 39174 21700 39206
rect 21624 38966 21700 39174
rect 21150 38902 21151 38934
rect 21085 38901 21151 38902
rect 21624 38902 21630 38966
rect 21694 38902 21700 38966
rect 22032 39174 22038 39238
rect 22102 39174 22108 39238
rect 22032 38966 22108 39174
rect 22032 38934 22038 38966
rect 21624 38896 21700 38902
rect 22037 38902 22038 38934
rect 22102 38934 22108 38966
rect 73984 39238 74060 39244
rect 73984 39174 73990 39238
rect 74054 39174 74060 39238
rect 73984 38966 74060 39174
rect 73984 38934 73990 38966
rect 22102 38902 22103 38934
rect 22037 38901 22103 38902
rect 73989 38902 73990 38934
rect 74054 38934 74060 38966
rect 74256 39238 74332 39244
rect 74256 39174 74262 39238
rect 74326 39174 74332 39238
rect 74256 38966 74332 39174
rect 74256 38934 74262 38966
rect 74054 38902 74055 38934
rect 73989 38901 74055 38902
rect 74261 38902 74262 38934
rect 74326 38934 74332 38966
rect 75072 39238 75148 39244
rect 75072 39174 75078 39238
rect 75142 39174 75148 39238
rect 75621 39238 75687 39239
rect 75621 39206 75622 39238
rect 75072 38966 75148 39174
rect 75072 38934 75078 38966
rect 74326 38902 74327 38934
rect 74261 38901 74327 38902
rect 75077 38902 75078 38934
rect 75142 38934 75148 38966
rect 75616 39174 75622 39206
rect 75686 39206 75687 39238
rect 75686 39174 75692 39206
rect 75616 38966 75692 39174
rect 75142 38902 75143 38934
rect 75077 38901 75143 38902
rect 75616 38902 75622 38966
rect 75686 38902 75692 38966
rect 75616 38896 75692 38902
rect 94656 38966 95004 40670
rect 94656 38902 94662 38966
rect 94726 38902 95004 38966
rect 21488 38830 21564 38836
rect 21488 38766 21494 38830
rect 21558 38766 21564 38830
rect 21488 38558 21564 38766
rect 21488 38526 21494 38558
rect 21493 38494 21494 38526
rect 21558 38526 21564 38558
rect 21760 38830 21836 38836
rect 21760 38766 21766 38830
rect 21830 38766 21836 38830
rect 21760 38558 21836 38766
rect 21760 38526 21766 38558
rect 21558 38494 21559 38526
rect 21493 38493 21559 38494
rect 21765 38494 21766 38526
rect 21830 38526 21836 38558
rect 22168 38830 22244 38836
rect 22168 38766 22174 38830
rect 22238 38766 22244 38830
rect 22168 38558 22244 38766
rect 22168 38526 22174 38558
rect 21830 38494 21831 38526
rect 21765 38493 21831 38494
rect 22173 38494 22174 38526
rect 22238 38526 22244 38558
rect 73984 38830 74060 38836
rect 73984 38766 73990 38830
rect 74054 38766 74060 38830
rect 73984 38558 74060 38766
rect 73984 38526 73990 38558
rect 22238 38494 22239 38526
rect 22173 38493 22239 38494
rect 73989 38494 73990 38526
rect 74054 38526 74060 38558
rect 74392 38830 74468 38836
rect 74392 38766 74398 38830
rect 74462 38766 74468 38830
rect 74669 38830 74735 38831
rect 74669 38798 74670 38830
rect 74392 38558 74468 38766
rect 74392 38526 74398 38558
rect 74054 38494 74055 38526
rect 73989 38493 74055 38494
rect 74397 38494 74398 38526
rect 74462 38526 74468 38558
rect 74664 38766 74670 38798
rect 74734 38798 74735 38830
rect 75072 38830 75148 38836
rect 74734 38766 74740 38798
rect 74664 38558 74740 38766
rect 74462 38494 74463 38526
rect 74397 38493 74463 38494
rect 74664 38494 74670 38558
rect 74734 38494 74740 38558
rect 75072 38766 75078 38830
rect 75142 38766 75148 38830
rect 75072 38558 75148 38766
rect 75072 38526 75078 38558
rect 74664 38488 74740 38494
rect 75077 38494 75078 38526
rect 75142 38526 75148 38558
rect 75142 38494 75143 38526
rect 75077 38493 75143 38494
rect 21624 38422 21700 38428
rect 21624 38358 21630 38422
rect 21694 38358 21700 38422
rect 21624 38150 21700 38358
rect 21624 38118 21630 38150
rect 21629 38086 21630 38118
rect 21694 38118 21700 38150
rect 22168 38422 22244 38428
rect 22168 38358 22174 38422
rect 22238 38358 22244 38422
rect 22168 38150 22244 38358
rect 22168 38118 22174 38150
rect 21694 38086 21695 38118
rect 21629 38085 21695 38086
rect 22173 38086 22174 38118
rect 22238 38118 22244 38150
rect 73848 38422 73924 38428
rect 73848 38358 73854 38422
rect 73918 38358 73924 38422
rect 74261 38422 74327 38423
rect 74261 38390 74262 38422
rect 73848 38150 73924 38358
rect 73848 38118 73854 38150
rect 22238 38086 22239 38118
rect 22173 38085 22239 38086
rect 73853 38086 73854 38118
rect 73918 38118 73924 38150
rect 74256 38358 74262 38390
rect 74326 38390 74327 38422
rect 74326 38358 74332 38390
rect 74256 38150 74332 38358
rect 73918 38086 73919 38118
rect 73853 38085 73919 38086
rect 74256 38086 74262 38150
rect 74326 38086 74332 38150
rect 74256 38080 74332 38086
rect 21080 38014 21156 38020
rect 21080 37950 21086 38014
rect 21150 37950 21156 38014
rect 21629 38014 21695 38015
rect 21629 37982 21630 38014
rect 952 37406 1230 37470
rect 1294 37406 1300 37470
rect 20536 37742 20612 37748
rect 20536 37678 20542 37742
rect 20606 37678 20612 37742
rect 21080 37742 21156 37950
rect 21080 37710 21086 37742
rect 20536 37470 20612 37678
rect 21085 37678 21086 37710
rect 21150 37710 21156 37742
rect 21624 37950 21630 37982
rect 21694 37982 21695 38014
rect 22173 38014 22239 38015
rect 22173 37982 22174 38014
rect 21694 37950 21700 37982
rect 21624 37742 21700 37950
rect 21150 37678 21151 37710
rect 21085 37677 21151 37678
rect 21624 37678 21630 37742
rect 21694 37678 21700 37742
rect 21624 37672 21700 37678
rect 22168 37950 22174 37982
rect 22238 37982 22239 38014
rect 73984 38014 74060 38020
rect 22238 37950 22244 37982
rect 22168 37742 22244 37950
rect 73984 37950 73990 38014
rect 74054 37950 74060 38014
rect 74397 38014 74463 38015
rect 74397 37982 74398 38014
rect 26933 37878 26999 37879
rect 26933 37846 26934 37878
rect 22168 37678 22174 37742
rect 22238 37678 22244 37742
rect 22168 37672 22244 37678
rect 26928 37814 26934 37846
rect 26998 37846 26999 37878
rect 26998 37814 27004 37846
rect 26928 37606 27004 37814
rect 73984 37742 74060 37950
rect 73984 37710 73990 37742
rect 73989 37678 73990 37710
rect 74054 37710 74060 37742
rect 74392 37950 74398 37982
rect 74462 37982 74463 38014
rect 74664 38014 74740 38020
rect 74462 37950 74468 37982
rect 74392 37742 74468 37950
rect 74054 37678 74055 37710
rect 73989 37677 74055 37678
rect 74392 37678 74398 37742
rect 74462 37678 74468 37742
rect 74664 37950 74670 38014
rect 74734 37950 74740 38014
rect 74664 37742 74740 37950
rect 74664 37710 74670 37742
rect 74392 37672 74468 37678
rect 74669 37678 74670 37710
rect 74734 37710 74740 37742
rect 75480 37742 75556 37748
rect 74734 37678 74735 37710
rect 74669 37677 74735 37678
rect 75480 37678 75486 37742
rect 75550 37678 75556 37742
rect 26928 37542 26934 37606
rect 26998 37542 27004 37606
rect 26928 37536 27004 37542
rect 20536 37438 20542 37470
rect 952 35566 1300 37406
rect 20541 37406 20542 37438
rect 20606 37438 20612 37470
rect 27069 37470 27135 37471
rect 27069 37438 27070 37470
rect 20606 37406 20607 37438
rect 20541 37405 20607 37406
rect 27064 37406 27070 37438
rect 27134 37438 27135 37470
rect 68957 37470 69023 37471
rect 68957 37438 68958 37470
rect 27134 37406 27140 37438
rect 20405 37334 20471 37335
rect 20405 37302 20406 37334
rect 20400 37270 20406 37302
rect 20470 37302 20471 37334
rect 20813 37334 20879 37335
rect 20813 37302 20814 37334
rect 20470 37270 20476 37302
rect 20400 37062 20476 37270
rect 20400 36998 20406 37062
rect 20470 36998 20476 37062
rect 20400 36992 20476 36998
rect 20808 37270 20814 37302
rect 20878 37302 20879 37334
rect 20878 37270 20884 37302
rect 20808 37062 20884 37270
rect 27064 37198 27140 37406
rect 27064 37134 27070 37198
rect 27134 37134 27140 37198
rect 27064 37128 27140 37134
rect 68952 37406 68958 37438
rect 69022 37438 69023 37470
rect 75480 37470 75556 37678
rect 75480 37438 75486 37470
rect 69022 37406 69028 37438
rect 68952 37198 69028 37406
rect 75485 37406 75486 37438
rect 75550 37438 75556 37470
rect 94656 37470 95004 38902
rect 75550 37406 75551 37438
rect 75485 37405 75551 37406
rect 94656 37406 94662 37470
rect 94726 37406 95004 37470
rect 68952 37134 68958 37198
rect 69022 37134 69028 37198
rect 68952 37128 69028 37134
rect 74664 37334 74740 37340
rect 74664 37270 74670 37334
rect 74734 37270 74740 37334
rect 20808 36998 20814 37062
rect 20878 36998 20884 37062
rect 20808 36992 20884 36998
rect 68952 37062 69028 37068
rect 68952 36998 68958 37062
rect 69022 36998 69028 37062
rect 74664 37062 74740 37270
rect 74664 37030 74670 37062
rect 20541 36926 20607 36927
rect 20541 36894 20542 36926
rect 20536 36862 20542 36894
rect 20606 36894 20607 36926
rect 20606 36862 20612 36894
rect 20536 36654 20612 36862
rect 68952 36790 69028 36998
rect 74669 36998 74670 37030
rect 74734 37030 74740 37062
rect 74936 37334 75012 37340
rect 74936 37270 74942 37334
rect 75006 37270 75012 37334
rect 75621 37334 75687 37335
rect 75621 37302 75622 37334
rect 74936 37062 75012 37270
rect 74936 37030 74942 37062
rect 74734 36998 74735 37030
rect 74669 36997 74735 36998
rect 74941 36998 74942 37030
rect 75006 37030 75012 37062
rect 75616 37270 75622 37302
rect 75686 37302 75687 37334
rect 75686 37270 75692 37302
rect 75616 37062 75692 37270
rect 75006 36998 75007 37030
rect 74941 36997 75007 36998
rect 75616 36998 75622 37062
rect 75686 36998 75692 37062
rect 75616 36992 75692 36998
rect 75621 36926 75687 36927
rect 75621 36894 75622 36926
rect 68952 36758 68958 36790
rect 68957 36726 68958 36758
rect 69022 36758 69028 36790
rect 75616 36862 75622 36894
rect 75686 36894 75687 36926
rect 75686 36862 75692 36894
rect 69022 36726 69023 36758
rect 68957 36725 69023 36726
rect 20536 36590 20542 36654
rect 20606 36590 20612 36654
rect 20536 36584 20612 36590
rect 75616 36654 75692 36862
rect 75616 36590 75622 36654
rect 75686 36590 75692 36654
rect 75616 36584 75692 36590
rect 20400 36518 20476 36524
rect 20400 36454 20406 36518
rect 20470 36454 20476 36518
rect 21357 36518 21423 36519
rect 21357 36486 21358 36518
rect 20400 36246 20476 36454
rect 20400 36214 20406 36246
rect 20405 36182 20406 36214
rect 20470 36214 20476 36246
rect 21352 36454 21358 36486
rect 21422 36486 21423 36518
rect 21624 36518 21700 36524
rect 21422 36454 21428 36486
rect 21352 36246 21428 36454
rect 20470 36182 20471 36214
rect 20405 36181 20471 36182
rect 21352 36182 21358 36246
rect 21422 36182 21428 36246
rect 21624 36454 21630 36518
rect 21694 36454 21700 36518
rect 22037 36518 22103 36519
rect 22037 36486 22038 36518
rect 21624 36246 21700 36454
rect 21624 36214 21630 36246
rect 21352 36176 21428 36182
rect 21629 36182 21630 36214
rect 21694 36214 21700 36246
rect 22032 36454 22038 36486
rect 22102 36486 22103 36518
rect 73848 36518 73924 36524
rect 22102 36454 22108 36486
rect 22032 36246 22108 36454
rect 73848 36454 73854 36518
rect 73918 36454 73924 36518
rect 21694 36182 21695 36214
rect 21629 36181 21695 36182
rect 22032 36182 22038 36246
rect 22102 36182 22108 36246
rect 22032 36176 22108 36182
rect 69088 36246 69164 36252
rect 69088 36182 69094 36246
rect 69158 36182 69164 36246
rect 73848 36246 73924 36454
rect 73848 36214 73854 36246
rect 20405 36110 20471 36111
rect 20405 36078 20406 36110
rect 20400 36046 20406 36078
rect 20470 36078 20471 36110
rect 20813 36110 20879 36111
rect 20813 36078 20814 36110
rect 20470 36046 20476 36078
rect 20400 35838 20476 36046
rect 20400 35774 20406 35838
rect 20470 35774 20476 35838
rect 20400 35768 20476 35774
rect 20808 36046 20814 36078
rect 20878 36078 20879 36110
rect 21221 36110 21287 36111
rect 21221 36078 21222 36110
rect 20878 36046 20884 36078
rect 20808 35838 20884 36046
rect 20808 35774 20814 35838
rect 20878 35774 20884 35838
rect 20808 35768 20884 35774
rect 21216 36046 21222 36078
rect 21286 36078 21287 36110
rect 21629 36110 21695 36111
rect 21629 36078 21630 36110
rect 21286 36046 21292 36078
rect 21216 35838 21292 36046
rect 21216 35774 21222 35838
rect 21286 35774 21292 35838
rect 21216 35768 21292 35774
rect 21624 36046 21630 36078
rect 21694 36078 21695 36110
rect 22168 36110 22244 36116
rect 21694 36046 21700 36078
rect 21624 35838 21700 36046
rect 21624 35774 21630 35838
rect 21694 35774 21700 35838
rect 22168 36046 22174 36110
rect 22238 36046 22244 36110
rect 22168 35838 22244 36046
rect 69088 35974 69164 36182
rect 73853 36182 73854 36214
rect 73918 36214 73924 36246
rect 74256 36518 74332 36524
rect 74256 36454 74262 36518
rect 74326 36454 74332 36518
rect 74256 36246 74332 36454
rect 74256 36214 74262 36246
rect 73918 36182 73919 36214
rect 73853 36181 73919 36182
rect 74261 36182 74262 36214
rect 74326 36214 74332 36246
rect 74936 36518 75012 36524
rect 74936 36454 74942 36518
rect 75006 36454 75012 36518
rect 75077 36518 75143 36519
rect 75077 36486 75078 36518
rect 74936 36246 75012 36454
rect 74936 36214 74942 36246
rect 74326 36182 74327 36214
rect 74261 36181 74327 36182
rect 74941 36182 74942 36214
rect 75006 36214 75012 36246
rect 75072 36454 75078 36486
rect 75142 36486 75143 36518
rect 75616 36518 75692 36524
rect 75142 36454 75148 36486
rect 75072 36246 75148 36454
rect 75006 36182 75007 36214
rect 74941 36181 75007 36182
rect 75072 36182 75078 36246
rect 75142 36182 75148 36246
rect 75616 36454 75622 36518
rect 75686 36454 75692 36518
rect 75616 36246 75692 36454
rect 75616 36214 75622 36246
rect 75072 36176 75148 36182
rect 75621 36182 75622 36214
rect 75686 36214 75692 36246
rect 75686 36182 75687 36214
rect 75621 36181 75687 36182
rect 69088 35942 69094 35974
rect 69093 35910 69094 35942
rect 69158 35942 69164 35974
rect 73848 36110 73924 36116
rect 73848 36046 73854 36110
rect 73918 36046 73924 36110
rect 69158 35910 69159 35942
rect 69093 35909 69159 35910
rect 22168 35806 22174 35838
rect 21624 35768 21700 35774
rect 22173 35774 22174 35806
rect 22238 35806 22244 35838
rect 73848 35838 73924 36046
rect 73848 35806 73854 35838
rect 22238 35774 22239 35806
rect 22173 35773 22239 35774
rect 73853 35774 73854 35806
rect 73918 35806 73924 35838
rect 74392 36110 74468 36116
rect 74392 36046 74398 36110
rect 74462 36046 74468 36110
rect 74392 35838 74468 36046
rect 74392 35806 74398 35838
rect 73918 35774 73919 35806
rect 73853 35773 73919 35774
rect 74397 35774 74398 35806
rect 74462 35806 74468 35838
rect 75072 36110 75148 36116
rect 75072 36046 75078 36110
rect 75142 36046 75148 36110
rect 75621 36110 75687 36111
rect 75621 36078 75622 36110
rect 75072 35838 75148 36046
rect 75072 35806 75078 35838
rect 74462 35774 74463 35806
rect 74397 35773 74463 35774
rect 75077 35774 75078 35806
rect 75142 35806 75148 35838
rect 75616 36046 75622 36078
rect 75686 36078 75687 36110
rect 75686 36046 75692 36078
rect 75616 35838 75692 36046
rect 75142 35774 75143 35806
rect 75077 35773 75143 35774
rect 75616 35774 75622 35838
rect 75686 35774 75692 35838
rect 75616 35768 75692 35774
rect 952 35502 1230 35566
rect 1294 35502 1300 35566
rect 952 33934 1300 35502
rect 20536 35702 20612 35708
rect 20536 35638 20542 35702
rect 20606 35638 20612 35702
rect 20949 35702 21015 35703
rect 20949 35670 20950 35702
rect 20536 35430 20612 35638
rect 20536 35398 20542 35430
rect 20541 35366 20542 35398
rect 20606 35398 20612 35430
rect 20944 35638 20950 35670
rect 21014 35670 21015 35702
rect 21760 35702 21836 35708
rect 21014 35638 21020 35670
rect 20944 35430 21020 35638
rect 20606 35366 20607 35398
rect 20541 35365 20607 35366
rect 20944 35366 20950 35430
rect 21014 35366 21020 35430
rect 21760 35638 21766 35702
rect 21830 35638 21836 35702
rect 22037 35702 22103 35703
rect 22037 35670 22038 35702
rect 21760 35430 21836 35638
rect 21760 35398 21766 35430
rect 20944 35360 21020 35366
rect 21765 35366 21766 35398
rect 21830 35398 21836 35430
rect 22032 35638 22038 35670
rect 22102 35670 22103 35702
rect 73984 35702 74060 35708
rect 22102 35638 22108 35670
rect 22032 35430 22108 35638
rect 21830 35366 21831 35398
rect 21765 35365 21831 35366
rect 22032 35366 22038 35430
rect 22102 35366 22108 35430
rect 73984 35638 73990 35702
rect 74054 35638 74060 35702
rect 74261 35702 74327 35703
rect 74261 35670 74262 35702
rect 73984 35430 74060 35638
rect 73984 35398 73990 35430
rect 22032 35360 22108 35366
rect 73989 35366 73990 35398
rect 74054 35398 74060 35430
rect 74256 35638 74262 35670
rect 74326 35670 74327 35702
rect 74669 35702 74735 35703
rect 74669 35670 74670 35702
rect 74326 35638 74332 35670
rect 74256 35430 74332 35638
rect 74054 35366 74055 35398
rect 73989 35365 74055 35366
rect 74256 35366 74262 35430
rect 74326 35366 74332 35430
rect 74256 35360 74332 35366
rect 74664 35638 74670 35670
rect 74734 35670 74735 35702
rect 75072 35702 75148 35708
rect 74734 35638 74740 35670
rect 74664 35430 74740 35638
rect 74664 35366 74670 35430
rect 74734 35366 74740 35430
rect 75072 35638 75078 35702
rect 75142 35638 75148 35702
rect 75485 35702 75551 35703
rect 75485 35670 75486 35702
rect 75072 35430 75148 35638
rect 75072 35398 75078 35430
rect 74664 35360 74740 35366
rect 75077 35366 75078 35398
rect 75142 35398 75148 35430
rect 75480 35638 75486 35670
rect 75550 35670 75551 35702
rect 75550 35638 75556 35670
rect 75480 35430 75556 35638
rect 75142 35366 75143 35398
rect 75077 35365 75143 35366
rect 75480 35366 75486 35430
rect 75550 35366 75556 35430
rect 75480 35360 75556 35366
rect 94656 35566 95004 37406
rect 94656 35502 94662 35566
rect 94726 35502 95004 35566
rect 20400 35294 20476 35300
rect 20400 35230 20406 35294
rect 20470 35230 20476 35294
rect 20400 35022 20476 35230
rect 20400 34990 20406 35022
rect 20405 34958 20406 34990
rect 20470 34990 20476 35022
rect 20808 35294 20884 35300
rect 20808 35230 20814 35294
rect 20878 35230 20884 35294
rect 21765 35294 21831 35295
rect 21765 35262 21766 35294
rect 20808 35022 20884 35230
rect 20808 34990 20814 35022
rect 20470 34958 20471 34990
rect 20405 34957 20471 34958
rect 20813 34958 20814 34990
rect 20878 34990 20884 35022
rect 21760 35230 21766 35262
rect 21830 35262 21831 35294
rect 22032 35294 22108 35300
rect 21830 35230 21836 35262
rect 21760 35022 21836 35230
rect 20878 34958 20879 34990
rect 20813 34957 20879 34958
rect 21760 34958 21766 35022
rect 21830 34958 21836 35022
rect 22032 35230 22038 35294
rect 22102 35230 22108 35294
rect 73989 35294 74055 35295
rect 73989 35262 73990 35294
rect 22032 35022 22108 35230
rect 22032 34990 22038 35022
rect 21760 34952 21836 34958
rect 22037 34958 22038 34990
rect 22102 34990 22108 35022
rect 73984 35230 73990 35262
rect 74054 35262 74055 35294
rect 74256 35294 74332 35300
rect 74054 35230 74060 35262
rect 73984 35022 74060 35230
rect 22102 34958 22103 34990
rect 22037 34957 22103 34958
rect 73984 34958 73990 35022
rect 74054 34958 74060 35022
rect 74256 35230 74262 35294
rect 74326 35230 74332 35294
rect 74256 35022 74332 35230
rect 74256 34990 74262 35022
rect 73984 34952 74060 34958
rect 74261 34958 74262 34990
rect 74326 34990 74332 35022
rect 74800 35294 74876 35300
rect 74800 35230 74806 35294
rect 74870 35230 74876 35294
rect 74800 35022 74876 35230
rect 74800 34990 74806 35022
rect 74326 34958 74327 34990
rect 74261 34957 74327 34958
rect 74805 34958 74806 34990
rect 74870 34990 74876 35022
rect 74936 35294 75012 35300
rect 74936 35230 74942 35294
rect 75006 35230 75012 35294
rect 74936 35022 75012 35230
rect 74936 34990 74942 35022
rect 74870 34958 74871 34990
rect 74805 34957 74871 34958
rect 74941 34958 74942 34990
rect 75006 34990 75012 35022
rect 75616 35294 75692 35300
rect 75616 35230 75622 35294
rect 75686 35230 75692 35294
rect 75616 35022 75692 35230
rect 75616 34990 75622 35022
rect 75006 34958 75007 34990
rect 74941 34957 75007 34958
rect 75621 34958 75622 34990
rect 75686 34990 75692 35022
rect 75686 34958 75687 34990
rect 75621 34957 75687 34958
rect 952 33870 1230 33934
rect 1294 33870 1300 33934
rect 952 32302 1300 33870
rect 13736 34886 13812 34892
rect 13736 34822 13742 34886
rect 13806 34822 13812 34886
rect 13605 33526 13671 33527
rect 13605 33494 13606 33526
rect 952 32238 1230 32302
rect 1294 32238 1300 32302
rect 952 30670 1300 32238
rect 13600 33462 13606 33494
rect 13670 33494 13671 33526
rect 13670 33462 13676 33494
rect 13600 30806 13676 33462
rect 13736 32166 13812 34822
rect 20944 34886 21020 34892
rect 20944 34822 20950 34886
rect 21014 34822 21020 34886
rect 20944 34614 21020 34822
rect 20944 34582 20950 34614
rect 20949 34550 20950 34582
rect 21014 34582 21020 34614
rect 21080 34886 21156 34892
rect 21080 34822 21086 34886
rect 21150 34822 21156 34886
rect 21080 34614 21156 34822
rect 21080 34582 21086 34614
rect 21014 34550 21015 34582
rect 20949 34549 21015 34550
rect 21085 34550 21086 34582
rect 21150 34582 21156 34614
rect 21760 34886 21836 34892
rect 21760 34822 21766 34886
rect 21830 34822 21836 34886
rect 21760 34614 21836 34822
rect 21760 34582 21766 34614
rect 21150 34550 21151 34582
rect 21085 34549 21151 34550
rect 21765 34550 21766 34582
rect 21830 34582 21836 34614
rect 22032 34886 22108 34892
rect 22032 34822 22038 34886
rect 22102 34822 22108 34886
rect 22032 34614 22108 34822
rect 22032 34582 22038 34614
rect 21830 34550 21831 34582
rect 21765 34549 21831 34550
rect 22037 34550 22038 34582
rect 22102 34582 22108 34614
rect 73984 34886 74060 34892
rect 73984 34822 73990 34886
rect 74054 34822 74060 34886
rect 73984 34614 74060 34822
rect 73984 34582 73990 34614
rect 22102 34550 22103 34582
rect 22037 34549 22103 34550
rect 73989 34550 73990 34582
rect 74054 34582 74060 34614
rect 74256 34886 74332 34892
rect 74256 34822 74262 34886
rect 74326 34822 74332 34886
rect 74256 34614 74332 34822
rect 74256 34582 74262 34614
rect 74054 34550 74055 34582
rect 73989 34549 74055 34550
rect 74261 34550 74262 34582
rect 74326 34582 74332 34614
rect 75072 34886 75148 34892
rect 75072 34822 75078 34886
rect 75142 34822 75148 34886
rect 75072 34614 75148 34822
rect 75072 34582 75078 34614
rect 74326 34550 74327 34582
rect 74261 34549 74327 34550
rect 75077 34550 75078 34582
rect 75142 34582 75148 34614
rect 75142 34550 75143 34582
rect 75077 34549 75143 34550
rect 20536 34478 20612 34484
rect 20536 34414 20542 34478
rect 20606 34414 20612 34478
rect 20536 34206 20612 34414
rect 20536 34174 20542 34206
rect 20541 34142 20542 34174
rect 20606 34174 20612 34206
rect 21488 34478 21564 34484
rect 21488 34414 21494 34478
rect 21558 34414 21564 34478
rect 21488 34206 21564 34414
rect 21488 34174 21494 34206
rect 20606 34142 20607 34174
rect 20541 34141 20607 34142
rect 21493 34142 21494 34174
rect 21558 34174 21564 34206
rect 21760 34478 21836 34484
rect 21760 34414 21766 34478
rect 21830 34414 21836 34478
rect 22037 34478 22103 34479
rect 22037 34446 22038 34478
rect 21760 34206 21836 34414
rect 21760 34174 21766 34206
rect 21558 34142 21559 34174
rect 21493 34141 21559 34142
rect 21765 34142 21766 34174
rect 21830 34174 21836 34206
rect 22032 34414 22038 34446
rect 22102 34446 22103 34478
rect 73984 34478 74060 34484
rect 22102 34414 22108 34446
rect 22032 34206 22108 34414
rect 21830 34142 21831 34174
rect 21765 34141 21831 34142
rect 22032 34142 22038 34206
rect 22102 34142 22108 34206
rect 73984 34414 73990 34478
rect 74054 34414 74060 34478
rect 73984 34206 74060 34414
rect 73984 34174 73990 34206
rect 22032 34136 22108 34142
rect 73989 34142 73990 34174
rect 74054 34174 74060 34206
rect 74392 34478 74468 34484
rect 74392 34414 74398 34478
rect 74462 34414 74468 34478
rect 74669 34478 74735 34479
rect 74669 34446 74670 34478
rect 74392 34206 74468 34414
rect 74392 34174 74398 34206
rect 74054 34142 74055 34174
rect 73989 34141 74055 34142
rect 74397 34142 74398 34174
rect 74462 34174 74468 34206
rect 74664 34414 74670 34446
rect 74734 34446 74735 34478
rect 75208 34478 75284 34484
rect 74734 34414 74740 34446
rect 74664 34206 74740 34414
rect 74462 34142 74463 34174
rect 74397 34141 74463 34142
rect 74664 34142 74670 34206
rect 74734 34142 74740 34206
rect 75208 34414 75214 34478
rect 75278 34414 75284 34478
rect 75485 34478 75551 34479
rect 75485 34446 75486 34478
rect 75208 34206 75284 34414
rect 75208 34174 75214 34206
rect 74664 34136 74740 34142
rect 75213 34142 75214 34174
rect 75278 34174 75284 34206
rect 75480 34414 75486 34446
rect 75550 34446 75551 34478
rect 75550 34414 75556 34446
rect 75480 34206 75556 34414
rect 75278 34142 75279 34174
rect 75213 34141 75279 34142
rect 75480 34142 75486 34206
rect 75550 34142 75556 34206
rect 75480 34136 75556 34142
rect 21357 34070 21423 34071
rect 21357 34038 21358 34070
rect 21352 34006 21358 34038
rect 21422 34038 21423 34070
rect 21629 34070 21695 34071
rect 21629 34038 21630 34070
rect 21422 34006 21428 34038
rect 20400 33798 20476 33804
rect 20400 33734 20406 33798
rect 20470 33734 20476 33798
rect 20400 33526 20476 33734
rect 21352 33798 21428 34006
rect 21352 33734 21358 33798
rect 21422 33734 21428 33798
rect 21352 33728 21428 33734
rect 21624 34006 21630 34038
rect 21694 34038 21695 34070
rect 22168 34070 22244 34076
rect 21694 34006 21700 34038
rect 21624 33798 21700 34006
rect 21624 33734 21630 33798
rect 21694 33734 21700 33798
rect 22168 34006 22174 34070
rect 22238 34006 22244 34070
rect 22168 33798 22244 34006
rect 22168 33766 22174 33798
rect 21624 33728 21700 33734
rect 22173 33734 22174 33766
rect 22238 33766 22244 33798
rect 73848 34070 73924 34076
rect 73848 34006 73854 34070
rect 73918 34006 73924 34070
rect 74261 34070 74327 34071
rect 74261 34038 74262 34070
rect 73848 33798 73924 34006
rect 73848 33766 73854 33798
rect 22238 33734 22239 33766
rect 22173 33733 22239 33734
rect 73853 33734 73854 33766
rect 73918 33766 73924 33798
rect 74256 34006 74262 34038
rect 74326 34038 74327 34070
rect 74800 34070 74876 34076
rect 74326 34006 74332 34038
rect 74256 33798 74332 34006
rect 73918 33734 73919 33766
rect 73853 33733 73919 33734
rect 74256 33734 74262 33798
rect 74326 33734 74332 33798
rect 74800 34006 74806 34070
rect 74870 34006 74876 34070
rect 74800 33798 74876 34006
rect 74800 33766 74806 33798
rect 74256 33728 74332 33734
rect 74805 33734 74806 33766
rect 74870 33766 74876 33798
rect 74936 34070 75012 34076
rect 74936 34006 74942 34070
rect 75006 34006 75012 34070
rect 74936 33798 75012 34006
rect 94656 33934 95004 35502
rect 94656 33870 94662 33934
rect 94726 33870 95004 33934
rect 74936 33766 74942 33798
rect 74870 33734 74871 33766
rect 74805 33733 74871 33734
rect 74941 33734 74942 33766
rect 75006 33766 75012 33798
rect 75480 33798 75556 33804
rect 75006 33734 75007 33766
rect 74941 33733 75007 33734
rect 75480 33734 75486 33798
rect 75550 33734 75556 33798
rect 20400 33494 20406 33526
rect 20405 33462 20406 33494
rect 20470 33494 20476 33526
rect 21760 33662 21836 33668
rect 21760 33598 21766 33662
rect 21830 33598 21836 33662
rect 22173 33662 22239 33663
rect 22173 33630 22174 33662
rect 20470 33462 20471 33494
rect 20405 33461 20471 33462
rect 21760 33390 21836 33598
rect 21760 33358 21766 33390
rect 21765 33326 21766 33358
rect 21830 33358 21836 33390
rect 22168 33598 22174 33630
rect 22238 33630 22239 33662
rect 73853 33662 73919 33663
rect 73853 33630 73854 33662
rect 22238 33598 22244 33630
rect 22168 33390 22244 33598
rect 21830 33326 21831 33358
rect 21765 33325 21831 33326
rect 22168 33326 22174 33390
rect 22238 33326 22244 33390
rect 22168 33320 22244 33326
rect 73848 33598 73854 33630
rect 73918 33630 73919 33662
rect 74256 33662 74332 33668
rect 73918 33598 73924 33630
rect 73848 33390 73924 33598
rect 73848 33326 73854 33390
rect 73918 33326 73924 33390
rect 74256 33598 74262 33662
rect 74326 33598 74332 33662
rect 74256 33390 74332 33598
rect 75480 33526 75556 33734
rect 75480 33494 75486 33526
rect 75485 33462 75486 33494
rect 75550 33494 75556 33526
rect 75550 33462 75551 33494
rect 75485 33461 75551 33462
rect 74256 33358 74262 33390
rect 73848 33320 73924 33326
rect 74261 33326 74262 33358
rect 74326 33358 74332 33390
rect 74326 33326 74327 33358
rect 74261 33325 74327 33326
rect 74800 33254 74876 33260
rect 74800 33190 74806 33254
rect 74870 33190 74876 33254
rect 27200 33118 27276 33124
rect 27200 33054 27206 33118
rect 27270 33054 27276 33118
rect 68957 33118 69023 33119
rect 68957 33086 68958 33118
rect 20536 32982 20612 32988
rect 20536 32918 20542 32982
rect 20606 32918 20612 32982
rect 20536 32710 20612 32918
rect 27200 32846 27276 33054
rect 27200 32814 27206 32846
rect 27205 32782 27206 32814
rect 27270 32814 27276 32846
rect 68952 33054 68958 33086
rect 69022 33086 69023 33118
rect 69022 33054 69028 33086
rect 68952 32846 69028 33054
rect 74800 32982 74876 33190
rect 74800 32950 74806 32982
rect 74805 32918 74806 32950
rect 74870 32950 74876 32982
rect 74936 33254 75012 33260
rect 74936 33190 74942 33254
rect 75006 33190 75012 33254
rect 74936 32982 75012 33190
rect 74936 32950 74942 32982
rect 74870 32918 74871 32950
rect 74805 32917 74871 32918
rect 74941 32918 74942 32950
rect 75006 32950 75012 32982
rect 75616 32982 75692 32988
rect 75006 32918 75007 32950
rect 74941 32917 75007 32918
rect 75616 32918 75622 32982
rect 75686 32918 75692 32982
rect 27270 32782 27271 32814
rect 27205 32781 27271 32782
rect 68952 32782 68958 32846
rect 69022 32782 69028 32846
rect 68952 32776 69028 32782
rect 20536 32678 20542 32710
rect 20541 32646 20542 32678
rect 20606 32678 20612 32710
rect 75616 32710 75692 32918
rect 75616 32678 75622 32710
rect 20606 32646 20607 32678
rect 20541 32645 20607 32646
rect 75621 32646 75622 32678
rect 75686 32678 75692 32710
rect 75686 32646 75687 32678
rect 75621 32645 75687 32646
rect 20541 32574 20607 32575
rect 20541 32542 20542 32574
rect 20536 32510 20542 32542
rect 20606 32542 20607 32574
rect 20813 32574 20879 32575
rect 20813 32542 20814 32574
rect 20606 32510 20612 32542
rect 20536 32302 20612 32510
rect 20536 32238 20542 32302
rect 20606 32238 20612 32302
rect 20536 32232 20612 32238
rect 20808 32510 20814 32542
rect 20878 32542 20879 32574
rect 21629 32574 21695 32575
rect 21629 32542 21630 32574
rect 20878 32510 20884 32542
rect 20808 32302 20884 32510
rect 20808 32238 20814 32302
rect 20878 32238 20884 32302
rect 20808 32232 20884 32238
rect 21624 32510 21630 32542
rect 21694 32542 21695 32574
rect 22173 32574 22239 32575
rect 22173 32542 22174 32574
rect 21694 32510 21700 32542
rect 21624 32302 21700 32510
rect 21624 32238 21630 32302
rect 21694 32238 21700 32302
rect 21624 32232 21700 32238
rect 22168 32510 22174 32542
rect 22238 32542 22239 32574
rect 73984 32574 74060 32580
rect 22238 32510 22244 32542
rect 22168 32302 22244 32510
rect 73984 32510 73990 32574
rect 74054 32510 74060 32574
rect 74397 32574 74463 32575
rect 74397 32542 74398 32574
rect 22168 32238 22174 32302
rect 22238 32238 22244 32302
rect 22168 32232 22244 32238
rect 27200 32302 27276 32308
rect 27200 32238 27206 32302
rect 27270 32238 27276 32302
rect 73984 32302 74060 32510
rect 73984 32270 73990 32302
rect 13736 32134 13742 32166
rect 13741 32102 13742 32134
rect 13806 32134 13812 32166
rect 20405 32166 20471 32167
rect 20405 32134 20406 32166
rect 13806 32102 13807 32134
rect 13741 32101 13807 32102
rect 20400 32102 20406 32134
rect 20470 32134 20471 32166
rect 20949 32166 21015 32167
rect 20949 32134 20950 32166
rect 20470 32102 20476 32134
rect 13741 32030 13807 32031
rect 13741 31998 13742 32030
rect 13600 30742 13606 30806
rect 13670 30742 13676 30806
rect 13600 30736 13676 30742
rect 13736 31966 13742 31998
rect 13806 31998 13807 32030
rect 13806 31966 13812 31998
rect 952 30606 1230 30670
rect 1294 30606 1300 30670
rect 13469 30670 13535 30671
rect 13469 30638 13470 30670
rect 952 29038 1300 30606
rect 952 28974 1230 29038
rect 1294 28974 1300 29038
rect 952 27406 1300 28974
rect 13464 30606 13470 30638
rect 13534 30638 13535 30670
rect 13534 30606 13540 30638
rect 13464 27950 13540 30606
rect 13736 29446 13812 31966
rect 20400 31894 20476 32102
rect 20400 31830 20406 31894
rect 20470 31830 20476 31894
rect 20400 31824 20476 31830
rect 20944 32102 20950 32134
rect 21014 32134 21015 32166
rect 21488 32166 21564 32172
rect 21014 32102 21020 32134
rect 20944 31894 21020 32102
rect 20944 31830 20950 31894
rect 21014 31830 21020 31894
rect 21488 32102 21494 32166
rect 21558 32102 21564 32166
rect 21488 31894 21564 32102
rect 21488 31862 21494 31894
rect 20944 31824 21020 31830
rect 21493 31830 21494 31862
rect 21558 31862 21564 31894
rect 21624 32166 21700 32172
rect 21624 32102 21630 32166
rect 21694 32102 21700 32166
rect 21624 31894 21700 32102
rect 21624 31862 21630 31894
rect 21558 31830 21559 31862
rect 21493 31829 21559 31830
rect 21629 31830 21630 31862
rect 21694 31862 21700 31894
rect 22032 32166 22108 32172
rect 22032 32102 22038 32166
rect 22102 32102 22108 32166
rect 22032 31894 22108 32102
rect 27200 32030 27276 32238
rect 73989 32238 73990 32270
rect 74054 32270 74060 32302
rect 74392 32510 74398 32542
rect 74462 32542 74463 32574
rect 74664 32574 74740 32580
rect 74462 32510 74468 32542
rect 74392 32302 74468 32510
rect 74054 32238 74055 32270
rect 73989 32237 74055 32238
rect 74392 32238 74398 32302
rect 74462 32238 74468 32302
rect 74664 32510 74670 32574
rect 74734 32510 74740 32574
rect 74664 32302 74740 32510
rect 74664 32270 74670 32302
rect 74392 32232 74468 32238
rect 74669 32238 74670 32270
rect 74734 32270 74740 32302
rect 75480 32574 75556 32580
rect 75480 32510 75486 32574
rect 75550 32510 75556 32574
rect 75480 32302 75556 32510
rect 75480 32270 75486 32302
rect 74734 32238 74735 32270
rect 74669 32237 74735 32238
rect 75485 32238 75486 32270
rect 75550 32270 75556 32302
rect 94656 32302 95004 33870
rect 75550 32238 75551 32270
rect 75485 32237 75551 32238
rect 94656 32238 94662 32302
rect 94726 32238 95004 32302
rect 73989 32166 74055 32167
rect 73989 32134 73990 32166
rect 27200 31998 27206 32030
rect 27205 31966 27206 31998
rect 27270 31998 27276 32030
rect 73984 32102 73990 32134
rect 74054 32134 74055 32166
rect 74256 32166 74332 32172
rect 74054 32102 74060 32134
rect 27270 31966 27271 31998
rect 27205 31965 27271 31966
rect 22032 31862 22038 31894
rect 21694 31830 21695 31862
rect 21629 31829 21695 31830
rect 22037 31830 22038 31862
rect 22102 31862 22108 31894
rect 73984 31894 74060 32102
rect 22102 31830 22103 31862
rect 22037 31829 22103 31830
rect 73984 31830 73990 31894
rect 74054 31830 74060 31894
rect 74256 32102 74262 32166
rect 74326 32102 74332 32166
rect 74256 31894 74332 32102
rect 74256 31862 74262 31894
rect 73984 31824 74060 31830
rect 74261 31830 74262 31862
rect 74326 31862 74332 31894
rect 74800 32166 74876 32172
rect 74800 32102 74806 32166
rect 74870 32102 74876 32166
rect 75485 32166 75551 32167
rect 75485 32134 75486 32166
rect 74800 31894 74876 32102
rect 74800 31862 74806 31894
rect 74326 31830 74327 31862
rect 74261 31829 74327 31830
rect 74805 31830 74806 31862
rect 74870 31862 74876 31894
rect 75480 32102 75486 32134
rect 75550 32134 75551 32166
rect 75550 32102 75556 32134
rect 75480 31894 75556 32102
rect 74870 31830 74871 31862
rect 74805 31829 74871 31830
rect 75480 31830 75486 31894
rect 75550 31830 75556 31894
rect 75480 31824 75556 31830
rect 20536 31758 20612 31764
rect 20536 31694 20542 31758
rect 20606 31694 20612 31758
rect 21221 31758 21287 31759
rect 21221 31726 21222 31758
rect 20536 31486 20612 31694
rect 20536 31454 20542 31486
rect 20541 31422 20542 31454
rect 20606 31454 20612 31486
rect 21216 31694 21222 31726
rect 21286 31726 21287 31758
rect 21624 31758 21700 31764
rect 21286 31694 21292 31726
rect 21216 31486 21292 31694
rect 20606 31422 20607 31454
rect 20541 31421 20607 31422
rect 21216 31422 21222 31486
rect 21286 31422 21292 31486
rect 21624 31694 21630 31758
rect 21694 31694 21700 31758
rect 21624 31486 21700 31694
rect 21624 31454 21630 31486
rect 21216 31416 21292 31422
rect 21629 31422 21630 31454
rect 21694 31454 21700 31486
rect 22168 31758 22244 31764
rect 22168 31694 22174 31758
rect 22238 31694 22244 31758
rect 22168 31486 22244 31694
rect 22168 31454 22174 31486
rect 21694 31422 21695 31454
rect 21629 31421 21695 31422
rect 22173 31422 22174 31454
rect 22238 31454 22244 31486
rect 73848 31758 73924 31764
rect 73848 31694 73854 31758
rect 73918 31694 73924 31758
rect 73848 31486 73924 31694
rect 73848 31454 73854 31486
rect 22238 31422 22239 31454
rect 22173 31421 22239 31422
rect 73853 31422 73854 31454
rect 73918 31454 73924 31486
rect 74392 31758 74468 31764
rect 74392 31694 74398 31758
rect 74462 31694 74468 31758
rect 74805 31758 74871 31759
rect 74805 31726 74806 31758
rect 74392 31486 74468 31694
rect 74392 31454 74398 31486
rect 73918 31422 73919 31454
rect 73853 31421 73919 31422
rect 74397 31422 74398 31454
rect 74462 31454 74468 31486
rect 74800 31694 74806 31726
rect 74870 31726 74871 31758
rect 75213 31758 75279 31759
rect 75213 31726 75214 31758
rect 74870 31694 74876 31726
rect 74800 31486 74876 31694
rect 74462 31422 74463 31454
rect 74397 31421 74463 31422
rect 74800 31422 74806 31486
rect 74870 31422 74876 31486
rect 74800 31416 74876 31422
rect 75208 31694 75214 31726
rect 75278 31726 75279 31758
rect 75616 31758 75692 31764
rect 75278 31694 75284 31726
rect 75208 31486 75284 31694
rect 75208 31422 75214 31486
rect 75278 31422 75284 31486
rect 75616 31694 75622 31758
rect 75686 31694 75692 31758
rect 75616 31486 75692 31694
rect 75616 31454 75622 31486
rect 75208 31416 75284 31422
rect 75621 31422 75622 31454
rect 75686 31454 75692 31486
rect 75686 31422 75687 31454
rect 75621 31421 75687 31422
rect 20405 31350 20471 31351
rect 20405 31318 20406 31350
rect 20400 31286 20406 31318
rect 20470 31318 20471 31350
rect 20949 31350 21015 31351
rect 20949 31318 20950 31350
rect 20470 31286 20476 31318
rect 20400 31078 20476 31286
rect 20400 31014 20406 31078
rect 20470 31014 20476 31078
rect 20400 31008 20476 31014
rect 20944 31286 20950 31318
rect 21014 31318 21015 31350
rect 21085 31350 21151 31351
rect 21085 31318 21086 31350
rect 21014 31286 21020 31318
rect 20944 31078 21020 31286
rect 20944 31014 20950 31078
rect 21014 31014 21020 31078
rect 20944 31008 21020 31014
rect 21080 31286 21086 31318
rect 21150 31318 21151 31350
rect 21765 31350 21831 31351
rect 21765 31318 21766 31350
rect 21150 31286 21156 31318
rect 21080 31078 21156 31286
rect 21080 31014 21086 31078
rect 21150 31014 21156 31078
rect 21080 31008 21156 31014
rect 21760 31286 21766 31318
rect 21830 31318 21831 31350
rect 22037 31350 22103 31351
rect 22037 31318 22038 31350
rect 21830 31286 21836 31318
rect 21760 31078 21836 31286
rect 21760 31014 21766 31078
rect 21830 31014 21836 31078
rect 21760 31008 21836 31014
rect 22032 31286 22038 31318
rect 22102 31318 22103 31350
rect 73984 31350 74060 31356
rect 22102 31286 22108 31318
rect 22032 31078 22108 31286
rect 22032 31014 22038 31078
rect 22102 31014 22108 31078
rect 73984 31286 73990 31350
rect 74054 31286 74060 31350
rect 73984 31078 74060 31286
rect 73984 31046 73990 31078
rect 22032 31008 22108 31014
rect 73989 31014 73990 31046
rect 74054 31046 74060 31078
rect 74392 31350 74468 31356
rect 74392 31286 74398 31350
rect 74462 31286 74468 31350
rect 74392 31078 74468 31286
rect 74392 31046 74398 31078
rect 74054 31014 74055 31046
rect 73989 31013 74055 31014
rect 74397 31014 74398 31046
rect 74462 31046 74468 31078
rect 75072 31350 75148 31356
rect 75072 31286 75078 31350
rect 75142 31286 75148 31350
rect 75485 31350 75551 31351
rect 75485 31318 75486 31350
rect 75072 31078 75148 31286
rect 75072 31046 75078 31078
rect 74462 31014 74463 31046
rect 74397 31013 74463 31014
rect 75077 31014 75078 31046
rect 75142 31046 75148 31078
rect 75480 31286 75486 31318
rect 75550 31318 75551 31350
rect 75550 31286 75556 31318
rect 75480 31078 75556 31286
rect 75142 31014 75143 31046
rect 75077 31013 75143 31014
rect 75480 31014 75486 31078
rect 75550 31014 75556 31078
rect 75480 31008 75556 31014
rect 20400 30942 20476 30948
rect 20400 30878 20406 30942
rect 20470 30878 20476 30942
rect 20400 30670 20476 30878
rect 20400 30638 20406 30670
rect 20405 30606 20406 30638
rect 20470 30638 20476 30670
rect 20808 30942 20884 30948
rect 20808 30878 20814 30942
rect 20878 30878 20884 30942
rect 21493 30942 21559 30943
rect 21493 30910 21494 30942
rect 20808 30670 20884 30878
rect 20808 30638 20814 30670
rect 20470 30606 20471 30638
rect 20405 30605 20471 30606
rect 20813 30606 20814 30638
rect 20878 30638 20884 30670
rect 21488 30878 21494 30910
rect 21558 30910 21559 30942
rect 21765 30942 21831 30943
rect 21765 30910 21766 30942
rect 21558 30878 21564 30910
rect 21488 30670 21564 30878
rect 20878 30606 20879 30638
rect 20813 30605 20879 30606
rect 21488 30606 21494 30670
rect 21558 30606 21564 30670
rect 21488 30600 21564 30606
rect 21760 30878 21766 30910
rect 21830 30910 21831 30942
rect 22168 30942 22244 30948
rect 21830 30878 21836 30910
rect 21760 30670 21836 30878
rect 21760 30606 21766 30670
rect 21830 30606 21836 30670
rect 22168 30878 22174 30942
rect 22238 30878 22244 30942
rect 22168 30670 22244 30878
rect 22168 30638 22174 30670
rect 21760 30600 21836 30606
rect 22173 30606 22174 30638
rect 22238 30638 22244 30670
rect 73848 30942 73924 30948
rect 73848 30878 73854 30942
rect 73918 30878 73924 30942
rect 74397 30942 74463 30943
rect 74397 30910 74398 30942
rect 73848 30670 73924 30878
rect 73848 30638 73854 30670
rect 22238 30606 22239 30638
rect 22173 30605 22239 30606
rect 73853 30606 73854 30638
rect 73918 30638 73924 30670
rect 74392 30878 74398 30910
rect 74462 30910 74463 30942
rect 74669 30942 74735 30943
rect 74669 30910 74670 30942
rect 74462 30878 74468 30910
rect 74392 30670 74468 30878
rect 73918 30606 73919 30638
rect 73853 30605 73919 30606
rect 74392 30606 74398 30670
rect 74462 30606 74468 30670
rect 74392 30600 74468 30606
rect 74664 30878 74670 30910
rect 74734 30910 74735 30942
rect 75616 30942 75692 30948
rect 74734 30878 74740 30910
rect 74664 30670 74740 30878
rect 74664 30606 74670 30670
rect 74734 30606 74740 30670
rect 75616 30878 75622 30942
rect 75686 30878 75692 30942
rect 75616 30670 75692 30878
rect 75616 30638 75622 30670
rect 74664 30600 74740 30606
rect 75621 30606 75622 30638
rect 75686 30638 75692 30670
rect 94656 30670 95004 32238
rect 75686 30606 75687 30638
rect 75621 30605 75687 30606
rect 94656 30606 94662 30670
rect 94726 30606 95004 30670
rect 20400 30534 20476 30540
rect 20400 30470 20406 30534
rect 20470 30470 20476 30534
rect 20400 30262 20476 30470
rect 20400 30230 20406 30262
rect 20405 30198 20406 30230
rect 20470 30230 20476 30262
rect 21760 30534 21836 30540
rect 21760 30470 21766 30534
rect 21830 30470 21836 30534
rect 22037 30534 22103 30535
rect 22037 30502 22038 30534
rect 21760 30262 21836 30470
rect 21760 30230 21766 30262
rect 20470 30198 20471 30230
rect 20405 30197 20471 30198
rect 21765 30198 21766 30230
rect 21830 30230 21836 30262
rect 22032 30470 22038 30502
rect 22102 30502 22103 30534
rect 73853 30534 73919 30535
rect 73853 30502 73854 30534
rect 22102 30470 22108 30502
rect 22032 30262 22108 30470
rect 21830 30198 21831 30230
rect 21765 30197 21831 30198
rect 22032 30198 22038 30262
rect 22102 30198 22108 30262
rect 22032 30192 22108 30198
rect 73848 30470 73854 30502
rect 73918 30502 73919 30534
rect 74256 30534 74332 30540
rect 73918 30470 73924 30502
rect 73848 30262 73924 30470
rect 73848 30198 73854 30262
rect 73918 30198 73924 30262
rect 74256 30470 74262 30534
rect 74326 30470 74332 30534
rect 74805 30534 74871 30535
rect 74805 30502 74806 30534
rect 74256 30262 74332 30470
rect 74256 30230 74262 30262
rect 73848 30192 73924 30198
rect 74261 30198 74262 30230
rect 74326 30230 74332 30262
rect 74800 30470 74806 30502
rect 74870 30502 74871 30534
rect 75480 30534 75556 30540
rect 74870 30470 74876 30502
rect 74800 30262 74876 30470
rect 74326 30198 74327 30230
rect 74261 30197 74327 30198
rect 74800 30198 74806 30262
rect 74870 30198 74876 30262
rect 75480 30470 75486 30534
rect 75550 30470 75556 30534
rect 75480 30262 75556 30470
rect 75480 30230 75486 30262
rect 74800 30192 74876 30198
rect 75485 30198 75486 30230
rect 75550 30230 75556 30262
rect 75550 30198 75551 30230
rect 75485 30197 75551 30198
rect 21221 30126 21287 30127
rect 21221 30094 21222 30126
rect 21216 30062 21222 30094
rect 21286 30094 21287 30126
rect 21765 30126 21831 30127
rect 21765 30094 21766 30126
rect 21286 30062 21292 30094
rect 20536 29854 20612 29860
rect 20536 29790 20542 29854
rect 20606 29790 20612 29854
rect 20536 29582 20612 29790
rect 21216 29854 21292 30062
rect 21216 29790 21222 29854
rect 21286 29790 21292 29854
rect 21216 29784 21292 29790
rect 21760 30062 21766 30094
rect 21830 30094 21831 30126
rect 22037 30126 22103 30127
rect 22037 30094 22038 30126
rect 21830 30062 21836 30094
rect 21760 29854 21836 30062
rect 21760 29790 21766 29854
rect 21830 29790 21836 29854
rect 21760 29784 21836 29790
rect 22032 30062 22038 30094
rect 22102 30094 22103 30126
rect 73989 30126 74055 30127
rect 73989 30094 73990 30126
rect 22102 30062 22108 30094
rect 22032 29854 22108 30062
rect 22032 29790 22038 29854
rect 22102 29790 22108 29854
rect 22032 29784 22108 29790
rect 73984 30062 73990 30094
rect 74054 30094 74055 30126
rect 74261 30126 74327 30127
rect 74261 30094 74262 30126
rect 74054 30062 74060 30094
rect 73984 29854 74060 30062
rect 73984 29790 73990 29854
rect 74054 29790 74060 29854
rect 73984 29784 74060 29790
rect 74256 30062 74262 30094
rect 74326 30094 74327 30126
rect 74664 30126 74740 30132
rect 74326 30062 74332 30094
rect 74256 29854 74332 30062
rect 74256 29790 74262 29854
rect 74326 29790 74332 29854
rect 74664 30062 74670 30126
rect 74734 30062 74740 30126
rect 74664 29854 74740 30062
rect 74664 29822 74670 29854
rect 74256 29784 74332 29790
rect 74669 29790 74670 29822
rect 74734 29822 74740 29854
rect 74936 30126 75012 30132
rect 74936 30062 74942 30126
rect 75006 30062 75012 30126
rect 74936 29854 75012 30062
rect 74936 29822 74942 29854
rect 74734 29790 74735 29822
rect 74669 29789 74735 29790
rect 74941 29790 74942 29822
rect 75006 29822 75012 29854
rect 75616 29854 75692 29860
rect 75006 29790 75007 29822
rect 74941 29789 75007 29790
rect 75616 29790 75622 29854
rect 75686 29790 75692 29854
rect 21629 29718 21695 29719
rect 21629 29686 21630 29718
rect 20536 29550 20542 29582
rect 20541 29518 20542 29550
rect 20606 29550 20612 29582
rect 21624 29654 21630 29686
rect 21694 29686 21695 29718
rect 22168 29718 22244 29724
rect 21694 29654 21700 29686
rect 20606 29518 20607 29550
rect 20541 29517 20607 29518
rect 13736 29382 13742 29446
rect 13806 29382 13812 29446
rect 13736 29376 13812 29382
rect 21624 29446 21700 29654
rect 21624 29382 21630 29446
rect 21694 29382 21700 29446
rect 22168 29654 22174 29718
rect 22238 29654 22244 29718
rect 22168 29446 22244 29654
rect 22168 29414 22174 29446
rect 21624 29376 21700 29382
rect 22173 29382 22174 29414
rect 22238 29414 22244 29446
rect 73848 29718 73924 29724
rect 73848 29654 73854 29718
rect 73918 29654 73924 29718
rect 73848 29446 73924 29654
rect 73848 29414 73854 29446
rect 22238 29382 22239 29414
rect 22173 29381 22239 29382
rect 73853 29382 73854 29414
rect 73918 29414 73924 29446
rect 74392 29718 74468 29724
rect 74392 29654 74398 29718
rect 74462 29654 74468 29718
rect 74392 29446 74468 29654
rect 75616 29582 75692 29790
rect 75616 29550 75622 29582
rect 75621 29518 75622 29550
rect 75686 29550 75692 29582
rect 75686 29518 75687 29550
rect 75621 29517 75687 29518
rect 74392 29414 74398 29446
rect 73918 29382 73919 29414
rect 73853 29381 73919 29382
rect 74397 29382 74398 29414
rect 74462 29414 74468 29446
rect 74462 29382 74463 29414
rect 74397 29381 74463 29382
rect 13464 27886 13470 27950
rect 13534 27886 13540 27950
rect 13464 27880 13540 27886
rect 13600 29310 13676 29316
rect 13600 29246 13606 29310
rect 13670 29246 13676 29310
rect 952 27342 1230 27406
rect 1294 27342 1300 27406
rect 952 25502 1300 27342
rect 13600 26590 13676 29246
rect 21080 29310 21156 29316
rect 21080 29246 21086 29310
rect 21150 29246 21156 29310
rect 20405 29038 20471 29039
rect 20405 29006 20406 29038
rect 20400 28974 20406 29006
rect 20470 29006 20471 29038
rect 21080 29038 21156 29246
rect 74664 29310 74740 29316
rect 74664 29246 74670 29310
rect 74734 29246 74740 29310
rect 21080 29006 21086 29038
rect 20470 28974 20476 29006
rect 20400 28766 20476 28974
rect 21085 28974 21086 29006
rect 21150 29006 21156 29038
rect 27200 29174 27276 29180
rect 27200 29110 27206 29174
rect 27270 29110 27276 29174
rect 68957 29174 69023 29175
rect 68957 29142 68958 29174
rect 21150 28974 21151 29006
rect 21085 28973 21151 28974
rect 20949 28902 21015 28903
rect 20949 28870 20950 28902
rect 20400 28702 20406 28766
rect 20470 28702 20476 28766
rect 20400 28696 20476 28702
rect 20944 28838 20950 28870
rect 21014 28870 21015 28902
rect 27200 28902 27276 29110
rect 27200 28870 27206 28902
rect 21014 28838 21020 28870
rect 20944 28772 21020 28838
rect 27205 28838 27206 28870
rect 27270 28870 27276 28902
rect 68952 29110 68958 29142
rect 69022 29142 69023 29174
rect 69022 29110 69028 29142
rect 68952 28902 69028 29110
rect 74664 29038 74740 29246
rect 74664 29006 74670 29038
rect 74669 28974 74670 29006
rect 74734 29006 74740 29038
rect 75485 29038 75551 29039
rect 75485 29006 75486 29038
rect 74734 28974 74735 29006
rect 74669 28973 74735 28974
rect 75480 28974 75486 29006
rect 75550 29006 75551 29038
rect 94656 29038 95004 30606
rect 75550 28974 75556 29006
rect 27270 28838 27271 28870
rect 27205 28837 27271 28838
rect 68952 28838 68958 28902
rect 69022 28838 69028 28902
rect 68952 28832 69028 28838
rect 20944 28766 21156 28772
rect 20944 28702 21086 28766
rect 21150 28702 21156 28766
rect 27069 28766 27135 28767
rect 27069 28734 27070 28766
rect 20944 28696 21156 28702
rect 27064 28702 27070 28734
rect 27134 28734 27135 28766
rect 68952 28766 69028 28772
rect 27134 28702 27140 28734
rect 20536 28630 20612 28636
rect 20536 28566 20542 28630
rect 20606 28566 20612 28630
rect 20813 28630 20879 28631
rect 20813 28598 20814 28630
rect 20536 28358 20612 28566
rect 20536 28326 20542 28358
rect 20541 28294 20542 28326
rect 20606 28326 20612 28358
rect 20808 28566 20814 28598
rect 20878 28598 20879 28630
rect 20878 28566 20884 28598
rect 20808 28358 20884 28566
rect 27064 28494 27140 28702
rect 27064 28430 27070 28494
rect 27134 28430 27140 28494
rect 68952 28702 68958 28766
rect 69022 28702 69028 28766
rect 68952 28494 69028 28702
rect 68952 28462 68958 28494
rect 27064 28424 27140 28430
rect 68957 28430 68958 28462
rect 69022 28462 69028 28494
rect 69088 28766 69164 28772
rect 69088 28702 69094 28766
rect 69158 28702 69164 28766
rect 69022 28430 69023 28462
rect 68957 28429 69023 28430
rect 20606 28294 20607 28326
rect 20541 28293 20607 28294
rect 20808 28294 20814 28358
rect 20878 28294 20884 28358
rect 69088 28358 69164 28702
rect 75480 28766 75556 28974
rect 75480 28702 75486 28766
rect 75550 28702 75556 28766
rect 75480 28696 75556 28702
rect 94656 28974 94662 29038
rect 94726 28974 95004 29038
rect 74941 28630 75007 28631
rect 74941 28598 74942 28630
rect 69088 28326 69094 28358
rect 20808 28288 20884 28294
rect 69093 28294 69094 28326
rect 69158 28326 69164 28358
rect 74936 28566 74942 28598
rect 75006 28598 75007 28630
rect 75621 28630 75687 28631
rect 75621 28598 75622 28630
rect 75006 28566 75012 28598
rect 74936 28358 75012 28566
rect 69158 28294 69159 28326
rect 69093 28293 69159 28294
rect 74936 28294 74942 28358
rect 75006 28294 75012 28358
rect 74936 28288 75012 28294
rect 75616 28566 75622 28598
rect 75686 28598 75687 28630
rect 75686 28566 75692 28598
rect 75616 28358 75692 28566
rect 75616 28294 75622 28358
rect 75686 28294 75692 28358
rect 75616 28288 75692 28294
rect 20541 28222 20607 28223
rect 20541 28190 20542 28222
rect 20536 28158 20542 28190
rect 20606 28190 20607 28222
rect 21760 28222 21836 28228
rect 20606 28158 20612 28190
rect 20536 27950 20612 28158
rect 20536 27886 20542 27950
rect 20606 27886 20612 27950
rect 21760 28158 21766 28222
rect 21830 28158 21836 28222
rect 21760 27950 21836 28158
rect 21760 27918 21766 27950
rect 20536 27880 20612 27886
rect 21765 27886 21766 27918
rect 21830 27918 21836 27950
rect 22032 28222 22108 28228
rect 22032 28158 22038 28222
rect 22102 28158 22108 28222
rect 22032 27950 22108 28158
rect 22032 27918 22038 27950
rect 21830 27886 21831 27918
rect 21765 27885 21831 27886
rect 22037 27886 22038 27918
rect 22102 27918 22108 27950
rect 73984 28222 74060 28228
rect 73984 28158 73990 28222
rect 74054 28158 74060 28222
rect 73984 27950 74060 28158
rect 73984 27918 73990 27950
rect 22102 27886 22103 27918
rect 22037 27885 22103 27886
rect 73989 27886 73990 27918
rect 74054 27918 74060 27950
rect 74256 28222 74332 28228
rect 74256 28158 74262 28222
rect 74326 28158 74332 28222
rect 75621 28222 75687 28223
rect 75621 28190 75622 28222
rect 74256 27950 74332 28158
rect 74256 27918 74262 27950
rect 74054 27886 74055 27918
rect 73989 27885 74055 27886
rect 74261 27886 74262 27918
rect 74326 27918 74332 27950
rect 75616 28158 75622 28190
rect 75686 28190 75687 28222
rect 75686 28158 75692 28190
rect 75616 27950 75692 28158
rect 74326 27886 74327 27918
rect 74261 27885 74327 27886
rect 75616 27886 75622 27950
rect 75686 27886 75692 27950
rect 75616 27880 75692 27886
rect 13600 26558 13606 26590
rect 13605 26526 13606 26558
rect 13670 26558 13676 26590
rect 13736 27814 13812 27820
rect 13736 27750 13742 27814
rect 13806 27750 13812 27814
rect 13670 26526 13671 26558
rect 13605 26525 13671 26526
rect 952 25438 1230 25502
rect 1294 25438 1300 25502
rect 952 23870 1300 25438
rect 13736 25094 13812 27750
rect 20400 27814 20476 27820
rect 20400 27750 20406 27814
rect 20470 27750 20476 27814
rect 20400 27542 20476 27750
rect 20400 27510 20406 27542
rect 20405 27478 20406 27510
rect 20470 27510 20476 27542
rect 21488 27814 21564 27820
rect 21488 27750 21494 27814
rect 21558 27750 21564 27814
rect 21488 27542 21564 27750
rect 21488 27510 21494 27542
rect 20470 27478 20471 27510
rect 20405 27477 20471 27478
rect 21493 27478 21494 27510
rect 21558 27510 21564 27542
rect 21624 27814 21700 27820
rect 21624 27750 21630 27814
rect 21694 27750 21700 27814
rect 22037 27814 22103 27815
rect 22037 27782 22038 27814
rect 21624 27542 21700 27750
rect 21624 27510 21630 27542
rect 21558 27478 21559 27510
rect 21493 27477 21559 27478
rect 21629 27478 21630 27510
rect 21694 27510 21700 27542
rect 22032 27750 22038 27782
rect 22102 27782 22103 27814
rect 73989 27814 74055 27815
rect 73989 27782 73990 27814
rect 22102 27750 22108 27782
rect 22032 27542 22108 27750
rect 73984 27750 73990 27782
rect 74054 27782 74055 27814
rect 74256 27814 74332 27820
rect 74054 27750 74060 27782
rect 21694 27478 21695 27510
rect 21629 27477 21695 27478
rect 22032 27478 22038 27542
rect 22102 27478 22108 27542
rect 27069 27542 27135 27543
rect 27069 27510 27070 27542
rect 22032 27472 22108 27478
rect 27064 27478 27070 27510
rect 27134 27510 27135 27542
rect 69088 27542 69164 27548
rect 27134 27478 27140 27510
rect 20536 27406 20612 27412
rect 20536 27342 20542 27406
rect 20606 27342 20612 27406
rect 20813 27406 20879 27407
rect 20813 27374 20814 27406
rect 20536 27134 20612 27342
rect 20536 27102 20542 27134
rect 20541 27070 20542 27102
rect 20606 27102 20612 27134
rect 20808 27342 20814 27374
rect 20878 27374 20879 27406
rect 21080 27406 21156 27412
rect 20878 27342 20884 27374
rect 20808 27134 20884 27342
rect 20606 27070 20607 27102
rect 20541 27069 20607 27070
rect 20808 27070 20814 27134
rect 20878 27070 20884 27134
rect 21080 27342 21086 27406
rect 21150 27342 21156 27406
rect 21629 27406 21695 27407
rect 21629 27374 21630 27406
rect 21080 27134 21156 27342
rect 21080 27102 21086 27134
rect 20808 27064 20884 27070
rect 21085 27070 21086 27102
rect 21150 27102 21156 27134
rect 21624 27342 21630 27374
rect 21694 27374 21695 27406
rect 22037 27406 22103 27407
rect 22037 27374 22038 27406
rect 21694 27342 21700 27374
rect 21624 27134 21700 27342
rect 21150 27070 21151 27102
rect 21085 27069 21151 27070
rect 21624 27070 21630 27134
rect 21694 27070 21700 27134
rect 21624 27064 21700 27070
rect 22032 27342 22038 27374
rect 22102 27374 22103 27406
rect 22102 27342 22108 27374
rect 22032 27134 22108 27342
rect 27064 27270 27140 27478
rect 27064 27206 27070 27270
rect 27134 27206 27140 27270
rect 69088 27478 69094 27542
rect 69158 27478 69164 27542
rect 69088 27270 69164 27478
rect 73984 27542 74060 27750
rect 73984 27478 73990 27542
rect 74054 27478 74060 27542
rect 74256 27750 74262 27814
rect 74326 27750 74332 27814
rect 74669 27814 74735 27815
rect 74669 27782 74670 27814
rect 74256 27542 74332 27750
rect 74256 27510 74262 27542
rect 73984 27472 74060 27478
rect 74261 27478 74262 27510
rect 74326 27510 74332 27542
rect 74664 27750 74670 27782
rect 74734 27782 74735 27814
rect 75485 27814 75551 27815
rect 75485 27782 75486 27814
rect 74734 27750 74740 27782
rect 74664 27542 74740 27750
rect 74326 27478 74327 27510
rect 74261 27477 74327 27478
rect 74664 27478 74670 27542
rect 74734 27478 74740 27542
rect 74664 27472 74740 27478
rect 75480 27750 75486 27782
rect 75550 27782 75551 27814
rect 75550 27750 75556 27782
rect 75480 27542 75556 27750
rect 75480 27478 75486 27542
rect 75550 27478 75556 27542
rect 75480 27472 75556 27478
rect 73853 27406 73919 27407
rect 73853 27374 73854 27406
rect 69088 27238 69094 27270
rect 27064 27200 27140 27206
rect 69093 27206 69094 27238
rect 69158 27238 69164 27270
rect 73848 27342 73854 27374
rect 73918 27374 73919 27406
rect 74261 27406 74327 27407
rect 74261 27374 74262 27406
rect 73918 27342 73924 27374
rect 69158 27206 69159 27238
rect 69093 27205 69159 27206
rect 22032 27070 22038 27134
rect 22102 27070 22108 27134
rect 22032 27064 22108 27070
rect 73848 27134 73924 27342
rect 73848 27070 73854 27134
rect 73918 27070 73924 27134
rect 73848 27064 73924 27070
rect 74256 27342 74262 27374
rect 74326 27374 74327 27406
rect 75213 27406 75279 27407
rect 75213 27374 75214 27406
rect 74326 27342 74332 27374
rect 74256 27134 74332 27342
rect 74256 27070 74262 27134
rect 74326 27070 74332 27134
rect 74256 27064 74332 27070
rect 75208 27342 75214 27374
rect 75278 27374 75279 27406
rect 75616 27406 75692 27412
rect 75278 27342 75284 27374
rect 75208 27134 75284 27342
rect 75208 27070 75214 27134
rect 75278 27070 75284 27134
rect 75616 27342 75622 27406
rect 75686 27342 75692 27406
rect 75616 27134 75692 27342
rect 75616 27102 75622 27134
rect 75208 27064 75284 27070
rect 75621 27070 75622 27102
rect 75686 27102 75692 27134
rect 94656 27406 95004 28974
rect 94656 27342 94662 27406
rect 94726 27342 95004 27406
rect 75686 27070 75687 27102
rect 75621 27069 75687 27070
rect 20405 26998 20471 26999
rect 20405 26966 20406 26998
rect 20400 26934 20406 26966
rect 20470 26966 20471 26998
rect 20944 26998 21020 27004
rect 20470 26934 20476 26966
rect 20400 26726 20476 26934
rect 20400 26662 20406 26726
rect 20470 26662 20476 26726
rect 20944 26934 20950 26998
rect 21014 26934 21020 26998
rect 21085 26998 21151 26999
rect 21085 26966 21086 26998
rect 20944 26726 21020 26934
rect 20944 26694 20950 26726
rect 20400 26656 20476 26662
rect 20949 26662 20950 26694
rect 21014 26694 21020 26726
rect 21080 26934 21086 26966
rect 21150 26966 21151 26998
rect 21760 26998 21836 27004
rect 21150 26934 21156 26966
rect 21080 26726 21156 26934
rect 21014 26662 21015 26694
rect 20949 26661 21015 26662
rect 21080 26662 21086 26726
rect 21150 26662 21156 26726
rect 21760 26934 21766 26998
rect 21830 26934 21836 26998
rect 22037 26998 22103 26999
rect 22037 26966 22038 26998
rect 21760 26726 21836 26934
rect 21760 26694 21766 26726
rect 21080 26656 21156 26662
rect 21765 26662 21766 26694
rect 21830 26694 21836 26726
rect 22032 26934 22038 26966
rect 22102 26966 22103 26998
rect 73989 26998 74055 26999
rect 73989 26966 73990 26998
rect 22102 26934 22108 26966
rect 22032 26726 22108 26934
rect 21830 26662 21831 26694
rect 21765 26661 21831 26662
rect 22032 26662 22038 26726
rect 22102 26662 22108 26726
rect 22032 26656 22108 26662
rect 73984 26934 73990 26966
rect 74054 26966 74055 26998
rect 74261 26998 74327 26999
rect 74261 26966 74262 26998
rect 74054 26934 74060 26966
rect 73984 26726 74060 26934
rect 73984 26662 73990 26726
rect 74054 26662 74060 26726
rect 73984 26656 74060 26662
rect 74256 26934 74262 26966
rect 74326 26966 74327 26998
rect 74669 26998 74735 26999
rect 74669 26966 74670 26998
rect 74326 26934 74332 26966
rect 74256 26726 74332 26934
rect 74256 26662 74262 26726
rect 74326 26662 74332 26726
rect 74256 26656 74332 26662
rect 74664 26934 74670 26966
rect 74734 26966 74735 26998
rect 75072 26998 75148 27004
rect 74734 26934 74740 26966
rect 74664 26726 74740 26934
rect 74664 26662 74670 26726
rect 74734 26662 74740 26726
rect 75072 26934 75078 26998
rect 75142 26934 75148 26998
rect 75485 26998 75551 26999
rect 75485 26966 75486 26998
rect 75072 26726 75148 26934
rect 75072 26694 75078 26726
rect 74664 26656 74740 26662
rect 75077 26662 75078 26694
rect 75142 26694 75148 26726
rect 75480 26934 75486 26966
rect 75550 26966 75551 26998
rect 75550 26934 75556 26966
rect 75480 26726 75556 26934
rect 75142 26662 75143 26694
rect 75077 26661 75143 26662
rect 75480 26662 75486 26726
rect 75550 26662 75556 26726
rect 75480 26656 75556 26662
rect 20541 26590 20607 26591
rect 20541 26558 20542 26590
rect 20536 26526 20542 26558
rect 20606 26558 20607 26590
rect 20808 26590 20884 26596
rect 20606 26526 20612 26558
rect 17413 26454 17479 26455
rect 17413 26422 17414 26454
rect 13736 25062 13742 25094
rect 13741 25030 13742 25062
rect 13806 25062 13812 25094
rect 17408 26390 17414 26422
rect 17478 26422 17479 26454
rect 17478 26390 17484 26422
rect 13806 25030 13807 25062
rect 13741 25029 13807 25030
rect 15509 24958 15575 24959
rect 15509 24926 15510 24958
rect 952 23806 1230 23870
rect 1294 23806 1300 23870
rect 952 22238 1300 23806
rect 15504 24894 15510 24926
rect 15574 24926 15575 24958
rect 15574 24894 15580 24926
rect 2560 22669 2626 22670
rect 2560 22605 2561 22669
rect 2625 22605 2626 22669
rect 2560 22604 2626 22605
rect 952 22174 1230 22238
rect 1294 22174 1300 22238
rect 952 20470 1300 22174
rect 952 20406 1230 20470
rect 1294 20406 1300 20470
rect 952 18974 1300 20406
rect 952 18910 1230 18974
rect 1294 18910 1300 18974
rect 952 17342 1300 18910
rect 952 17278 1230 17342
rect 1294 17278 1300 17342
rect 952 15438 1300 17278
rect 2312 16254 2388 16260
rect 2312 16190 2318 16254
rect 2382 16190 2388 16254
rect 2312 15574 2388 16190
rect 2312 15542 2318 15574
rect 2317 15510 2318 15542
rect 2382 15542 2388 15574
rect 2382 15510 2383 15542
rect 2317 15509 2383 15510
rect 952 15374 1230 15438
rect 1294 15374 1300 15438
rect 952 13806 1300 15374
rect 2563 15263 2623 22604
rect 15504 22374 15580 24894
rect 17408 24822 17484 26390
rect 20536 26318 20612 26526
rect 20536 26254 20542 26318
rect 20606 26254 20612 26318
rect 20808 26526 20814 26590
rect 20878 26526 20884 26590
rect 21493 26590 21559 26591
rect 21493 26558 21494 26590
rect 20808 26318 20884 26526
rect 20808 26286 20814 26318
rect 20536 26248 20612 26254
rect 20813 26254 20814 26286
rect 20878 26286 20884 26318
rect 21488 26526 21494 26558
rect 21558 26558 21559 26590
rect 21765 26590 21831 26591
rect 21765 26558 21766 26590
rect 21558 26526 21564 26558
rect 21488 26318 21564 26526
rect 20878 26254 20879 26286
rect 20813 26253 20879 26254
rect 21488 26254 21494 26318
rect 21558 26254 21564 26318
rect 21488 26248 21564 26254
rect 21760 26526 21766 26558
rect 21830 26558 21831 26590
rect 22032 26590 22108 26596
rect 21830 26526 21836 26558
rect 21760 26318 21836 26526
rect 21760 26254 21766 26318
rect 21830 26254 21836 26318
rect 22032 26526 22038 26590
rect 22102 26526 22108 26590
rect 22032 26318 22108 26526
rect 22032 26286 22038 26318
rect 21760 26248 21836 26254
rect 22037 26254 22038 26286
rect 22102 26286 22108 26318
rect 73848 26590 73924 26596
rect 73848 26526 73854 26590
rect 73918 26526 73924 26590
rect 73848 26318 73924 26526
rect 73848 26286 73854 26318
rect 22102 26254 22103 26286
rect 22037 26253 22103 26254
rect 73853 26254 73854 26286
rect 73918 26286 73924 26318
rect 74256 26590 74332 26596
rect 74256 26526 74262 26590
rect 74326 26526 74332 26590
rect 74669 26590 74735 26591
rect 74669 26558 74670 26590
rect 74256 26318 74332 26526
rect 74256 26286 74262 26318
rect 73918 26254 73919 26286
rect 73853 26253 73919 26254
rect 74261 26254 74262 26286
rect 74326 26286 74332 26318
rect 74664 26526 74670 26558
rect 74734 26558 74735 26590
rect 74936 26590 75012 26596
rect 74734 26526 74740 26558
rect 74664 26318 74740 26526
rect 74326 26254 74327 26286
rect 74261 26253 74327 26254
rect 74664 26254 74670 26318
rect 74734 26254 74740 26318
rect 74936 26526 74942 26590
rect 75006 26526 75012 26590
rect 74936 26318 75012 26526
rect 74936 26286 74942 26318
rect 74664 26248 74740 26254
rect 74941 26254 74942 26286
rect 75006 26286 75012 26318
rect 75616 26590 75692 26596
rect 75616 26526 75622 26590
rect 75686 26526 75692 26590
rect 75616 26318 75692 26526
rect 75616 26286 75622 26318
rect 75006 26254 75007 26286
rect 74941 26253 75007 26254
rect 75621 26254 75622 26286
rect 75686 26286 75692 26318
rect 75686 26254 75687 26286
rect 75621 26253 75687 26254
rect 21760 26182 21836 26188
rect 21760 26118 21766 26182
rect 21830 26118 21836 26182
rect 22173 26182 22239 26183
rect 22173 26150 22174 26182
rect 21760 25910 21836 26118
rect 21760 25878 21766 25910
rect 21765 25846 21766 25878
rect 21830 25878 21836 25910
rect 22168 26118 22174 26150
rect 22238 26150 22239 26182
rect 73853 26182 73919 26183
rect 73853 26150 73854 26182
rect 22238 26118 22244 26150
rect 22168 25910 22244 26118
rect 73848 26118 73854 26150
rect 73918 26150 73919 26182
rect 74256 26182 74332 26188
rect 73918 26118 73924 26150
rect 21830 25846 21831 25878
rect 21765 25845 21831 25846
rect 22168 25846 22174 25910
rect 22238 25846 22244 25910
rect 22168 25840 22244 25846
rect 27200 26046 27276 26052
rect 27200 25982 27206 26046
rect 27270 25982 27276 26046
rect 21765 25774 21831 25775
rect 21765 25742 21766 25774
rect 21760 25710 21766 25742
rect 21830 25742 21831 25774
rect 22168 25774 22244 25780
rect 21830 25710 21836 25742
rect 21760 25502 21836 25710
rect 21760 25438 21766 25502
rect 21830 25438 21836 25502
rect 22168 25710 22174 25774
rect 22238 25710 22244 25774
rect 27200 25774 27276 25982
rect 73848 25910 73924 26118
rect 73848 25846 73854 25910
rect 73918 25846 73924 25910
rect 74256 26118 74262 26182
rect 74326 26118 74332 26182
rect 74256 25910 74332 26118
rect 74256 25878 74262 25910
rect 73848 25840 73924 25846
rect 74261 25846 74262 25878
rect 74326 25878 74332 25910
rect 75072 26182 75148 26188
rect 75072 26118 75078 26182
rect 75142 26118 75148 26182
rect 75072 25910 75148 26118
rect 75072 25878 75078 25910
rect 74326 25846 74327 25878
rect 74261 25845 74327 25846
rect 75077 25846 75078 25878
rect 75142 25878 75148 25910
rect 75142 25846 75143 25878
rect 75077 25845 75143 25846
rect 27200 25742 27206 25774
rect 22168 25502 22244 25710
rect 27205 25710 27206 25742
rect 27270 25742 27276 25774
rect 73989 25774 74055 25775
rect 73989 25742 73990 25774
rect 27270 25710 27271 25742
rect 27205 25709 27271 25710
rect 73984 25710 73990 25742
rect 74054 25742 74055 25774
rect 74261 25774 74327 25775
rect 74261 25742 74262 25774
rect 74054 25710 74060 25742
rect 22168 25470 22174 25502
rect 21760 25432 21836 25438
rect 22173 25438 22174 25470
rect 22238 25470 22244 25502
rect 73984 25502 74060 25710
rect 22238 25438 22239 25470
rect 22173 25437 22239 25438
rect 73984 25438 73990 25502
rect 74054 25438 74060 25502
rect 73984 25432 74060 25438
rect 74256 25710 74262 25742
rect 74326 25742 74327 25774
rect 74326 25710 74332 25742
rect 74256 25502 74332 25710
rect 74256 25438 74262 25502
rect 74326 25438 74332 25502
rect 74256 25432 74332 25438
rect 94656 25502 95004 27342
rect 94656 25438 94662 25502
rect 94726 25438 95004 25502
rect 20808 25366 20884 25372
rect 20808 25302 20814 25366
rect 20878 25302 20884 25366
rect 21357 25366 21423 25367
rect 21357 25334 21358 25366
rect 17408 24758 17414 24822
rect 17478 24758 17484 24822
rect 20400 25094 20476 25100
rect 20400 25030 20406 25094
rect 20470 25030 20476 25094
rect 20400 24822 20476 25030
rect 20400 24790 20406 24822
rect 17408 24752 17484 24758
rect 20405 24758 20406 24790
rect 20470 24790 20476 24822
rect 20470 24758 20471 24790
rect 20405 24757 20471 24758
rect 17136 24686 17212 24692
rect 17136 24622 17142 24686
rect 17206 24622 17212 24686
rect 17136 24006 17212 24622
rect 17952 24686 18028 24692
rect 17952 24622 17958 24686
rect 18022 24622 18028 24686
rect 17136 23974 17142 24006
rect 17141 23942 17142 23974
rect 17206 23974 17212 24006
rect 17272 24278 17348 24284
rect 17272 24214 17278 24278
rect 17342 24214 17348 24278
rect 17272 24006 17348 24214
rect 17272 23974 17278 24006
rect 17206 23942 17207 23974
rect 17141 23941 17207 23942
rect 17277 23942 17278 23974
rect 17342 23974 17348 24006
rect 17952 24006 18028 24622
rect 20536 24686 20612 24692
rect 20536 24622 20542 24686
rect 20606 24622 20612 24686
rect 18365 24550 18431 24551
rect 18365 24518 18366 24550
rect 18360 24486 18366 24518
rect 18430 24518 18431 24550
rect 18637 24550 18703 24551
rect 18637 24518 18638 24550
rect 18430 24486 18436 24518
rect 18229 24278 18295 24279
rect 18229 24246 18230 24278
rect 17952 23974 17958 24006
rect 17342 23942 17343 23974
rect 17277 23941 17343 23942
rect 17957 23942 17958 23974
rect 18022 23974 18028 24006
rect 18224 24214 18230 24246
rect 18294 24246 18295 24278
rect 18294 24214 18300 24246
rect 18224 24006 18300 24214
rect 18022 23942 18023 23974
rect 17957 23941 18023 23942
rect 18224 23942 18230 24006
rect 18294 23942 18300 24006
rect 18224 23936 18300 23942
rect 18360 24006 18436 24486
rect 18360 23942 18366 24006
rect 18430 23942 18436 24006
rect 18360 23936 18436 23942
rect 18632 24486 18638 24518
rect 18702 24518 18703 24550
rect 18702 24486 18708 24518
rect 18632 24006 18708 24486
rect 20536 24414 20612 24622
rect 20808 24550 20884 25302
rect 21352 25302 21358 25334
rect 21422 25334 21423 25366
rect 21629 25366 21695 25367
rect 21629 25334 21630 25366
rect 21422 25302 21428 25334
rect 21352 25094 21428 25302
rect 21352 25030 21358 25094
rect 21422 25030 21428 25094
rect 21352 25024 21428 25030
rect 21624 25302 21630 25334
rect 21694 25334 21695 25366
rect 22037 25366 22103 25367
rect 22037 25334 22038 25366
rect 21694 25302 21700 25334
rect 21624 25094 21700 25302
rect 21624 25030 21630 25094
rect 21694 25030 21700 25094
rect 21624 25024 21700 25030
rect 22032 25302 22038 25334
rect 22102 25334 22103 25366
rect 73853 25366 73919 25367
rect 73853 25334 73854 25366
rect 22102 25302 22108 25334
rect 22032 25094 22108 25302
rect 22032 25030 22038 25094
rect 22102 25030 22108 25094
rect 22032 25024 22108 25030
rect 73848 25302 73854 25334
rect 73918 25334 73919 25366
rect 74392 25366 74468 25372
rect 73918 25302 73924 25334
rect 73848 25094 73924 25302
rect 73848 25030 73854 25094
rect 73918 25030 73924 25094
rect 74392 25302 74398 25366
rect 74462 25302 74468 25366
rect 74392 25094 74468 25302
rect 74392 25062 74398 25094
rect 73848 25024 73924 25030
rect 74397 25030 74398 25062
rect 74462 25062 74468 25094
rect 74800 25366 74876 25372
rect 74800 25302 74806 25366
rect 74870 25302 74876 25366
rect 74800 25094 74876 25302
rect 74800 25062 74806 25094
rect 74462 25030 74463 25062
rect 74397 25029 74463 25030
rect 74805 25030 74806 25062
rect 74870 25062 74876 25094
rect 74936 25366 75012 25372
rect 74936 25302 74942 25366
rect 75006 25302 75012 25366
rect 74936 25094 75012 25302
rect 74936 25062 74942 25094
rect 74870 25030 74871 25062
rect 74805 25029 74871 25030
rect 74941 25030 74942 25062
rect 75006 25062 75012 25094
rect 75621 25094 75687 25095
rect 75621 25062 75622 25094
rect 75006 25030 75007 25062
rect 74941 25029 75007 25030
rect 75616 25030 75622 25062
rect 75686 25062 75687 25094
rect 75686 25030 75692 25062
rect 26933 24822 26999 24823
rect 26933 24790 26934 24822
rect 26928 24758 26934 24790
rect 26998 24790 26999 24822
rect 68957 24822 69023 24823
rect 68957 24790 68958 24822
rect 26998 24758 27004 24790
rect 21493 24686 21559 24687
rect 21493 24654 21494 24686
rect 20808 24518 20814 24550
rect 20813 24486 20814 24518
rect 20878 24518 20884 24550
rect 21488 24622 21494 24654
rect 21558 24654 21559 24686
rect 21558 24622 21564 24654
rect 20878 24486 20879 24518
rect 20813 24485 20879 24486
rect 20536 24382 20542 24414
rect 20541 24350 20542 24382
rect 20606 24382 20612 24414
rect 21488 24414 21564 24622
rect 26928 24550 27004 24758
rect 26928 24486 26934 24550
rect 26998 24486 27004 24550
rect 26928 24480 27004 24486
rect 68952 24758 68958 24790
rect 69022 24790 69023 24822
rect 75616 24822 75692 25030
rect 69022 24758 69028 24790
rect 68952 24550 69028 24758
rect 75616 24758 75622 24822
rect 75686 24758 75692 24822
rect 75616 24752 75692 24758
rect 74669 24686 74735 24687
rect 74669 24654 74670 24686
rect 68952 24486 68958 24550
rect 69022 24486 69028 24550
rect 68952 24480 69028 24486
rect 74664 24622 74670 24654
rect 74734 24654 74735 24686
rect 75480 24686 75556 24692
rect 74734 24622 74740 24654
rect 20606 24350 20607 24382
rect 20541 24349 20607 24350
rect 21488 24350 21494 24414
rect 21558 24350 21564 24414
rect 68957 24414 69023 24415
rect 68957 24382 68958 24414
rect 21488 24344 21564 24350
rect 68952 24350 68958 24382
rect 69022 24382 69023 24414
rect 74664 24414 74740 24622
rect 69022 24350 69028 24382
rect 20405 24278 20471 24279
rect 20405 24246 20406 24278
rect 18632 23942 18638 24006
rect 18702 23942 18708 24006
rect 18632 23936 18708 23942
rect 20400 24214 20406 24246
rect 20470 24246 20471 24278
rect 21629 24278 21695 24279
rect 21629 24246 21630 24278
rect 20470 24214 20476 24246
rect 20400 24006 20476 24214
rect 20400 23942 20406 24006
rect 20470 23942 20476 24006
rect 20400 23936 20476 23942
rect 21624 24214 21630 24246
rect 21694 24246 21695 24278
rect 22168 24278 22244 24284
rect 21694 24214 21700 24246
rect 21624 24006 21700 24214
rect 21624 23942 21630 24006
rect 21694 23942 21700 24006
rect 22168 24214 22174 24278
rect 22238 24214 22244 24278
rect 22168 24006 22244 24214
rect 68952 24142 69028 24350
rect 74664 24350 74670 24414
rect 74734 24350 74740 24414
rect 75480 24622 75486 24686
rect 75550 24622 75556 24686
rect 78069 24686 78135 24687
rect 78069 24654 78070 24686
rect 75480 24414 75556 24622
rect 78064 24622 78070 24654
rect 78134 24654 78135 24686
rect 79016 24686 79092 24692
rect 78134 24622 78140 24654
rect 77253 24550 77319 24551
rect 77253 24518 77254 24550
rect 75480 24382 75486 24414
rect 74664 24344 74740 24350
rect 75485 24350 75486 24382
rect 75550 24382 75556 24414
rect 77248 24486 77254 24518
rect 77318 24518 77319 24550
rect 77792 24550 77868 24556
rect 77318 24486 77324 24518
rect 75550 24350 75551 24382
rect 75485 24349 75551 24350
rect 73853 24278 73919 24279
rect 73853 24246 73854 24278
rect 68952 24078 68958 24142
rect 69022 24078 69028 24142
rect 68952 24072 69028 24078
rect 73848 24214 73854 24246
rect 73918 24246 73919 24278
rect 74392 24278 74468 24284
rect 73918 24214 73924 24246
rect 22168 23974 22174 24006
rect 21624 23936 21700 23942
rect 22173 23942 22174 23974
rect 22238 23974 22244 24006
rect 27064 24006 27140 24012
rect 22238 23942 22239 23974
rect 22173 23941 22239 23942
rect 27064 23942 27070 24006
rect 27134 23942 27140 24006
rect 17141 23870 17207 23871
rect 17141 23838 17142 23870
rect 17136 23806 17142 23838
rect 17206 23838 17207 23870
rect 18365 23870 18431 23871
rect 18365 23838 18366 23870
rect 17206 23806 17212 23838
rect 17136 23190 17212 23806
rect 18360 23806 18366 23838
rect 18430 23838 18431 23870
rect 20541 23870 20607 23871
rect 20541 23838 20542 23870
rect 18430 23806 18436 23838
rect 17821 23734 17887 23735
rect 17821 23702 17822 23734
rect 17136 23126 17142 23190
rect 17206 23126 17212 23190
rect 17136 23120 17212 23126
rect 17816 23670 17822 23702
rect 17886 23702 17887 23734
rect 17886 23670 17892 23702
rect 17816 23190 17892 23670
rect 17816 23126 17822 23190
rect 17886 23126 17892 23190
rect 17816 23120 17892 23126
rect 18360 23190 18436 23806
rect 20536 23806 20542 23838
rect 20606 23838 20607 23870
rect 20813 23870 20879 23871
rect 20813 23838 20814 23870
rect 20606 23806 20612 23838
rect 20536 23598 20612 23806
rect 20536 23534 20542 23598
rect 20606 23534 20612 23598
rect 20536 23528 20612 23534
rect 20808 23806 20814 23838
rect 20878 23838 20879 23870
rect 21760 23870 21836 23876
rect 20878 23806 20884 23838
rect 20808 23598 20884 23806
rect 20808 23534 20814 23598
rect 20878 23534 20884 23598
rect 21760 23806 21766 23870
rect 21830 23806 21836 23870
rect 21760 23598 21836 23806
rect 21760 23566 21766 23598
rect 20808 23528 20884 23534
rect 21765 23534 21766 23566
rect 21830 23566 21836 23598
rect 22032 23870 22108 23876
rect 22032 23806 22038 23870
rect 22102 23806 22108 23870
rect 22032 23598 22108 23806
rect 22032 23566 22038 23598
rect 21830 23534 21831 23566
rect 21765 23533 21831 23534
rect 22037 23534 22038 23566
rect 22102 23566 22108 23598
rect 27064 23598 27140 23942
rect 73848 24006 73924 24214
rect 73848 23942 73854 24006
rect 73918 23942 73924 24006
rect 74392 24214 74398 24278
rect 74462 24214 74468 24278
rect 74392 24006 74468 24214
rect 75616 24278 75692 24284
rect 75616 24214 75622 24278
rect 75686 24214 75692 24278
rect 74392 23974 74398 24006
rect 73848 23936 73924 23942
rect 74397 23942 74398 23974
rect 74462 23974 74468 24006
rect 74936 24142 75012 24148
rect 74936 24078 74942 24142
rect 75006 24078 75012 24142
rect 74462 23942 74463 23974
rect 74397 23941 74463 23942
rect 73984 23870 74060 23876
rect 73984 23806 73990 23870
rect 74054 23806 74060 23870
rect 74397 23870 74463 23871
rect 74397 23838 74398 23870
rect 27064 23566 27070 23598
rect 22102 23534 22103 23566
rect 22037 23533 22103 23534
rect 27069 23534 27070 23566
rect 27134 23566 27140 23598
rect 68957 23598 69023 23599
rect 68957 23566 68958 23598
rect 27134 23534 27135 23566
rect 27069 23533 27135 23534
rect 68952 23534 68958 23566
rect 69022 23566 69023 23598
rect 73984 23598 74060 23806
rect 73984 23566 73990 23598
rect 69022 23534 69028 23566
rect 20405 23462 20471 23463
rect 20405 23430 20406 23462
rect 18360 23126 18366 23190
rect 18430 23126 18436 23190
rect 18360 23120 18436 23126
rect 20400 23398 20406 23430
rect 20470 23430 20471 23462
rect 20949 23462 21015 23463
rect 20949 23430 20950 23462
rect 20470 23398 20476 23430
rect 20400 23190 20476 23398
rect 20400 23126 20406 23190
rect 20470 23126 20476 23190
rect 20400 23120 20476 23126
rect 20944 23398 20950 23430
rect 21014 23430 21015 23462
rect 21488 23462 21564 23468
rect 21014 23398 21020 23430
rect 20944 23190 21020 23398
rect 20944 23126 20950 23190
rect 21014 23126 21020 23190
rect 21488 23398 21494 23462
rect 21558 23398 21564 23462
rect 21765 23462 21831 23463
rect 21765 23430 21766 23462
rect 21488 23190 21564 23398
rect 21488 23158 21494 23190
rect 20944 23120 21020 23126
rect 21493 23126 21494 23158
rect 21558 23158 21564 23190
rect 21760 23398 21766 23430
rect 21830 23430 21831 23462
rect 22032 23462 22108 23468
rect 21830 23398 21836 23430
rect 21760 23190 21836 23398
rect 21558 23126 21559 23158
rect 21493 23125 21559 23126
rect 21760 23126 21766 23190
rect 21830 23126 21836 23190
rect 22032 23398 22038 23462
rect 22102 23398 22108 23462
rect 22032 23190 22108 23398
rect 68952 23326 69028 23534
rect 73989 23534 73990 23566
rect 74054 23566 74060 23598
rect 74392 23806 74398 23838
rect 74462 23838 74463 23870
rect 74936 23870 75012 24078
rect 75616 24006 75692 24214
rect 75616 23974 75622 24006
rect 75621 23942 75622 23974
rect 75686 23974 75692 24006
rect 77248 24006 77324 24486
rect 75686 23942 75687 23974
rect 75621 23941 75687 23942
rect 77248 23942 77254 24006
rect 77318 23942 77324 24006
rect 77792 24486 77798 24550
rect 77862 24486 77868 24550
rect 77792 24006 77868 24486
rect 77792 23974 77798 24006
rect 77248 23936 77324 23942
rect 77797 23942 77798 23974
rect 77862 23974 77868 24006
rect 78064 24006 78140 24622
rect 77862 23942 77863 23974
rect 77797 23941 77863 23942
rect 78064 23942 78070 24006
rect 78134 23942 78140 24006
rect 79016 24622 79022 24686
rect 79086 24622 79092 24686
rect 79016 24006 79092 24622
rect 79016 23974 79022 24006
rect 78064 23936 78140 23942
rect 79021 23942 79022 23974
rect 79086 23974 79092 24006
rect 79086 23942 79087 23974
rect 79021 23941 79087 23942
rect 74936 23838 74942 23870
rect 74462 23806 74468 23838
rect 74392 23598 74468 23806
rect 74941 23806 74942 23838
rect 75006 23838 75012 23870
rect 75213 23870 75279 23871
rect 75213 23838 75214 23870
rect 75006 23806 75007 23838
rect 74941 23805 75007 23806
rect 75208 23806 75214 23838
rect 75278 23838 75279 23870
rect 75480 23870 75556 23876
rect 75278 23806 75284 23838
rect 74054 23534 74055 23566
rect 73989 23533 74055 23534
rect 74392 23534 74398 23598
rect 74462 23534 74468 23598
rect 74392 23528 74468 23534
rect 75208 23598 75284 23806
rect 75208 23534 75214 23598
rect 75278 23534 75284 23598
rect 75480 23806 75486 23870
rect 75550 23806 75556 23870
rect 75480 23598 75556 23806
rect 75480 23566 75486 23598
rect 75208 23528 75284 23534
rect 75485 23534 75486 23566
rect 75550 23566 75556 23598
rect 77656 23870 77732 23876
rect 77656 23806 77662 23870
rect 77726 23806 77732 23870
rect 77797 23870 77863 23871
rect 77797 23838 77798 23870
rect 75550 23534 75551 23566
rect 75485 23533 75551 23534
rect 73989 23462 74055 23463
rect 73989 23430 73990 23462
rect 68952 23262 68958 23326
rect 69022 23262 69028 23326
rect 68952 23256 69028 23262
rect 73984 23398 73990 23430
rect 74054 23430 74055 23462
rect 74261 23462 74327 23463
rect 74261 23430 74262 23462
rect 74054 23398 74060 23430
rect 22032 23158 22038 23190
rect 21760 23120 21836 23126
rect 22037 23126 22038 23158
rect 22102 23158 22108 23190
rect 73984 23190 74060 23398
rect 22102 23126 22103 23158
rect 22037 23125 22103 23126
rect 73984 23126 73990 23190
rect 74054 23126 74060 23190
rect 73984 23120 74060 23126
rect 74256 23398 74262 23430
rect 74326 23430 74327 23462
rect 74800 23462 74876 23468
rect 74326 23398 74332 23430
rect 74256 23190 74332 23398
rect 74256 23126 74262 23190
rect 74326 23126 74332 23190
rect 74800 23398 74806 23462
rect 74870 23398 74876 23462
rect 75485 23462 75551 23463
rect 75485 23430 75486 23462
rect 74800 23190 74876 23398
rect 74800 23158 74806 23190
rect 74256 23120 74332 23126
rect 74805 23126 74806 23158
rect 74870 23158 74876 23190
rect 75480 23398 75486 23430
rect 75550 23430 75551 23462
rect 75550 23398 75556 23430
rect 75480 23190 75556 23398
rect 77656 23326 77732 23806
rect 77656 23294 77662 23326
rect 77661 23262 77662 23294
rect 77726 23294 77732 23326
rect 77792 23806 77798 23838
rect 77862 23838 77863 23870
rect 78341 23870 78407 23871
rect 78341 23838 78342 23870
rect 77862 23806 77868 23838
rect 77726 23262 77727 23294
rect 77661 23261 77727 23262
rect 74870 23126 74871 23158
rect 74805 23125 74871 23126
rect 75480 23126 75486 23190
rect 75550 23126 75556 23190
rect 75480 23120 75556 23126
rect 77792 23190 77868 23806
rect 77792 23126 77798 23190
rect 77862 23126 77868 23190
rect 77792 23120 77868 23126
rect 78336 23806 78342 23838
rect 78406 23838 78407 23870
rect 79016 23870 79092 23876
rect 78406 23806 78412 23838
rect 78336 23190 78412 23806
rect 78336 23126 78342 23190
rect 78406 23126 78412 23190
rect 79016 23806 79022 23870
rect 79086 23806 79092 23870
rect 79016 23190 79092 23806
rect 79016 23158 79022 23190
rect 78336 23120 78412 23126
rect 79021 23126 79022 23158
rect 79086 23158 79092 23190
rect 94656 23870 95004 25438
rect 94656 23806 94662 23870
rect 94726 23806 95004 23870
rect 79086 23126 79087 23158
rect 79021 23125 79087 23126
rect 15504 22310 15510 22374
rect 15574 22310 15580 22374
rect 17000 23054 17076 23060
rect 17000 22990 17006 23054
rect 17070 22990 17076 23054
rect 17000 22374 17076 22990
rect 17000 22342 17006 22374
rect 15504 22304 15580 22310
rect 17005 22310 17006 22342
rect 17070 22342 17076 22374
rect 17680 23054 17756 23060
rect 17680 22990 17686 23054
rect 17750 22990 17756 23054
rect 17680 22374 17756 22990
rect 17680 22342 17686 22374
rect 17070 22310 17071 22342
rect 17005 22309 17071 22310
rect 17685 22310 17686 22342
rect 17750 22342 17756 22374
rect 18360 23054 18436 23060
rect 18360 22990 18366 23054
rect 18430 22990 18436 23054
rect 18360 22374 18436 22990
rect 18360 22342 18366 22374
rect 17750 22310 17751 22342
rect 17685 22309 17751 22310
rect 18365 22310 18366 22342
rect 18430 22342 18436 22374
rect 18768 23054 18844 23060
rect 18768 22990 18774 23054
rect 18838 22990 18844 23054
rect 18768 22374 18844 22990
rect 20536 23054 20612 23060
rect 20536 22990 20542 23054
rect 20606 22990 20612 23054
rect 20536 22782 20612 22990
rect 20536 22750 20542 22782
rect 20541 22718 20542 22750
rect 20606 22750 20612 22782
rect 20808 23054 20884 23060
rect 20808 22990 20814 23054
rect 20878 22990 20884 23054
rect 20808 22782 20884 22990
rect 20808 22750 20814 22782
rect 20606 22718 20607 22750
rect 20541 22717 20607 22718
rect 20813 22718 20814 22750
rect 20878 22750 20884 22782
rect 21624 23054 21700 23060
rect 21624 22990 21630 23054
rect 21694 22990 21700 23054
rect 22037 23054 22103 23055
rect 22037 23022 22038 23054
rect 21624 22782 21700 22990
rect 21624 22750 21630 22782
rect 20878 22718 20879 22750
rect 20813 22717 20879 22718
rect 21629 22718 21630 22750
rect 21694 22750 21700 22782
rect 22032 22990 22038 23022
rect 22102 23022 22103 23054
rect 73848 23054 73924 23060
rect 22102 22990 22108 23022
rect 22032 22782 22108 22990
rect 21694 22718 21695 22750
rect 21629 22717 21695 22718
rect 22032 22718 22038 22782
rect 22102 22718 22108 22782
rect 73848 22990 73854 23054
rect 73918 22990 73924 23054
rect 73848 22782 73924 22990
rect 73848 22750 73854 22782
rect 22032 22712 22108 22718
rect 73853 22718 73854 22750
rect 73918 22750 73924 22782
rect 74392 23054 74468 23060
rect 74392 22990 74398 23054
rect 74462 22990 74468 23054
rect 75213 23054 75279 23055
rect 75213 23022 75214 23054
rect 74392 22782 74468 22990
rect 74392 22750 74398 22782
rect 73918 22718 73919 22750
rect 73853 22717 73919 22718
rect 74397 22718 74398 22750
rect 74462 22750 74468 22782
rect 75208 22990 75214 23022
rect 75278 23022 75279 23054
rect 75621 23054 75687 23055
rect 75621 23022 75622 23054
rect 75278 22990 75284 23022
rect 75208 22782 75284 22990
rect 74462 22718 74463 22750
rect 74397 22717 74463 22718
rect 75208 22718 75214 22782
rect 75278 22718 75284 22782
rect 75208 22712 75284 22718
rect 75616 22990 75622 23022
rect 75686 23022 75687 23054
rect 77248 23054 77324 23060
rect 75686 22990 75692 23022
rect 75616 22782 75692 22990
rect 75616 22718 75622 22782
rect 75686 22718 75692 22782
rect 75616 22712 75692 22718
rect 77248 22990 77254 23054
rect 77318 22990 77324 23054
rect 77797 23054 77863 23055
rect 77797 23022 77798 23054
rect 20405 22646 20471 22647
rect 20405 22614 20406 22646
rect 18768 22342 18774 22374
rect 18430 22310 18431 22342
rect 18365 22309 18431 22310
rect 18773 22310 18774 22342
rect 18838 22342 18844 22374
rect 20400 22582 20406 22614
rect 20470 22614 20471 22646
rect 21760 22646 21836 22652
rect 20470 22582 20476 22614
rect 20400 22374 20476 22582
rect 18838 22310 18839 22342
rect 18773 22309 18839 22310
rect 20400 22310 20406 22374
rect 20470 22310 20476 22374
rect 21760 22582 21766 22646
rect 21830 22582 21836 22646
rect 22037 22646 22103 22647
rect 22037 22614 22038 22646
rect 21760 22374 21836 22582
rect 21760 22342 21766 22374
rect 20400 22304 20476 22310
rect 21765 22310 21766 22342
rect 21830 22342 21836 22374
rect 22032 22582 22038 22614
rect 22102 22614 22103 22646
rect 73984 22646 74060 22652
rect 22102 22582 22108 22614
rect 22032 22374 22108 22582
rect 21830 22310 21831 22342
rect 21765 22309 21831 22310
rect 22032 22310 22038 22374
rect 22102 22310 22108 22374
rect 73984 22582 73990 22646
rect 74054 22582 74060 22646
rect 74261 22646 74327 22647
rect 74261 22614 74262 22646
rect 73984 22374 74060 22582
rect 73984 22342 73990 22374
rect 22032 22304 22108 22310
rect 73989 22310 73990 22342
rect 74054 22342 74060 22374
rect 74256 22582 74262 22614
rect 74326 22614 74327 22646
rect 74669 22646 74735 22647
rect 74669 22614 74670 22646
rect 74326 22582 74332 22614
rect 74256 22374 74332 22582
rect 74054 22310 74055 22342
rect 73989 22309 74055 22310
rect 74256 22310 74262 22374
rect 74326 22310 74332 22374
rect 74256 22304 74332 22310
rect 74664 22582 74670 22614
rect 74734 22614 74735 22646
rect 75072 22646 75148 22652
rect 74734 22582 74740 22614
rect 74664 22374 74740 22582
rect 74664 22310 74670 22374
rect 74734 22310 74740 22374
rect 75072 22582 75078 22646
rect 75142 22582 75148 22646
rect 75072 22374 75148 22582
rect 75072 22342 75078 22374
rect 74664 22304 74740 22310
rect 75077 22310 75078 22342
rect 75142 22342 75148 22374
rect 75480 22646 75556 22652
rect 75480 22582 75486 22646
rect 75550 22582 75556 22646
rect 75480 22374 75556 22582
rect 75480 22342 75486 22374
rect 75142 22310 75143 22342
rect 75077 22309 75143 22310
rect 75485 22310 75486 22342
rect 75550 22342 75556 22374
rect 77248 22374 77324 22990
rect 77248 22342 77254 22374
rect 75550 22310 75551 22342
rect 75485 22309 75551 22310
rect 77253 22310 77254 22342
rect 77318 22342 77324 22374
rect 77792 22990 77798 23022
rect 77862 23022 77863 23054
rect 78608 23054 78684 23060
rect 77862 22990 77868 23022
rect 77792 22374 77868 22990
rect 77318 22310 77319 22342
rect 77253 22309 77319 22310
rect 77792 22310 77798 22374
rect 77862 22310 77868 22374
rect 78608 22990 78614 23054
rect 78678 22990 78684 23054
rect 78885 23054 78951 23055
rect 78885 23022 78886 23054
rect 78608 22374 78684 22990
rect 78608 22342 78614 22374
rect 77792 22304 77868 22310
rect 78613 22310 78614 22342
rect 78678 22342 78684 22374
rect 78880 22990 78886 23022
rect 78950 23022 78951 23054
rect 78950 22990 78956 23022
rect 78880 22374 78956 22990
rect 78678 22310 78679 22342
rect 78613 22309 78679 22310
rect 78880 22310 78886 22374
rect 78950 22310 78956 22374
rect 78880 22304 78956 22310
rect 94656 22374 95004 23806
rect 94656 22310 94662 22374
rect 94726 22310 95004 22374
rect 17277 22238 17343 22239
rect 17277 22206 17278 22238
rect 17272 22174 17278 22206
rect 17342 22206 17343 22238
rect 18501 22238 18567 22239
rect 18501 22206 18502 22238
rect 17342 22174 17348 22206
rect 17272 20878 17348 22174
rect 18496 22174 18502 22206
rect 18566 22206 18567 22238
rect 18632 22238 18708 22244
rect 18566 22174 18572 22206
rect 18496 21694 18572 22174
rect 18496 21630 18502 21694
rect 18566 21630 18572 21694
rect 18496 21624 18572 21630
rect 18632 22174 18638 22238
rect 18702 22174 18708 22238
rect 17272 20814 17278 20878
rect 17342 20814 17348 20878
rect 18632 20878 18708 22174
rect 20808 22238 20884 22244
rect 20808 22174 20814 22238
rect 20878 22174 20884 22238
rect 21493 22238 21559 22239
rect 21493 22206 21494 22238
rect 20808 21966 20884 22174
rect 20808 21934 20814 21966
rect 20813 21902 20814 21934
rect 20878 21934 20884 21966
rect 21488 22174 21494 22206
rect 21558 22206 21559 22238
rect 21765 22238 21831 22239
rect 21765 22206 21766 22238
rect 21558 22174 21564 22206
rect 21488 21966 21564 22174
rect 20878 21902 20879 21934
rect 20813 21901 20879 21902
rect 21488 21902 21494 21966
rect 21558 21902 21564 21966
rect 21488 21896 21564 21902
rect 21760 22174 21766 22206
rect 21830 22206 21831 22238
rect 22173 22238 22239 22239
rect 22173 22206 22174 22238
rect 21830 22174 21836 22206
rect 21760 21966 21836 22174
rect 21760 21902 21766 21966
rect 21830 21902 21836 21966
rect 21760 21896 21836 21902
rect 22168 22174 22174 22206
rect 22238 22206 22239 22238
rect 73848 22238 73924 22244
rect 22238 22174 22244 22206
rect 22168 21966 22244 22174
rect 73848 22174 73854 22238
rect 73918 22174 73924 22238
rect 22168 21902 22174 21966
rect 22238 21902 22244 21966
rect 22168 21896 22244 21902
rect 26928 22102 27004 22108
rect 26928 22038 26934 22102
rect 26998 22038 27004 22102
rect 21760 21830 21836 21836
rect 21760 21766 21766 21830
rect 21830 21766 21836 21830
rect 21760 21558 21836 21766
rect 21760 21526 21766 21558
rect 21765 21494 21766 21526
rect 21830 21526 21836 21558
rect 22032 21830 22108 21836
rect 22032 21766 22038 21830
rect 22102 21766 22108 21830
rect 26928 21830 27004 22038
rect 73848 21966 73924 22174
rect 73848 21934 73854 21966
rect 73853 21902 73854 21934
rect 73918 21934 73924 21966
rect 74256 22238 74332 22244
rect 74256 22174 74262 22238
rect 74326 22174 74332 22238
rect 74256 21966 74332 22174
rect 74256 21934 74262 21966
rect 73918 21902 73919 21934
rect 73853 21901 73919 21902
rect 74261 21902 74262 21934
rect 74326 21934 74332 21966
rect 74800 22238 74876 22244
rect 74800 22174 74806 22238
rect 74870 22174 74876 22238
rect 74800 21966 74876 22174
rect 74800 21934 74806 21966
rect 74326 21902 74327 21934
rect 74261 21901 74327 21902
rect 74805 21902 74806 21934
rect 74870 21934 74876 21966
rect 74936 22238 75012 22244
rect 74936 22174 74942 22238
rect 75006 22174 75012 22238
rect 74936 21966 75012 22174
rect 74936 21934 74942 21966
rect 74870 21902 74871 21934
rect 74805 21901 74871 21902
rect 74941 21902 74942 21934
rect 75006 21934 75012 21966
rect 75208 22238 75284 22244
rect 75208 22174 75214 22238
rect 75278 22174 75284 22238
rect 75208 21966 75284 22174
rect 75208 21934 75214 21966
rect 75006 21902 75007 21934
rect 74941 21901 75007 21902
rect 75213 21902 75214 21934
rect 75278 21934 75284 21966
rect 77384 22238 77460 22244
rect 77384 22174 77390 22238
rect 77454 22174 77460 22238
rect 75278 21902 75279 21934
rect 75213 21901 75279 21902
rect 26928 21798 26934 21830
rect 22032 21558 22108 21766
rect 26933 21766 26934 21798
rect 26998 21798 27004 21830
rect 69093 21830 69159 21831
rect 69093 21798 69094 21830
rect 26998 21766 26999 21798
rect 26933 21765 26999 21766
rect 69088 21766 69094 21798
rect 69158 21798 69159 21830
rect 73853 21830 73919 21831
rect 73853 21798 73854 21830
rect 69158 21766 69164 21798
rect 22032 21526 22038 21558
rect 21830 21494 21831 21526
rect 21765 21493 21831 21494
rect 22037 21494 22038 21526
rect 22102 21526 22108 21558
rect 68952 21558 69028 21564
rect 22102 21494 22103 21526
rect 22037 21493 22103 21494
rect 68952 21494 68958 21558
rect 69022 21494 69028 21558
rect 21085 21422 21151 21423
rect 21085 21390 21086 21422
rect 21080 21358 21086 21390
rect 21150 21390 21151 21422
rect 21760 21422 21836 21428
rect 21150 21358 21156 21390
rect 20541 21150 20607 21151
rect 20541 21118 20542 21150
rect 18632 20846 18638 20878
rect 17272 20808 17348 20814
rect 18637 20814 18638 20846
rect 18702 20846 18708 20878
rect 20536 21086 20542 21118
rect 20606 21118 20607 21150
rect 21080 21150 21156 21358
rect 20606 21086 20612 21118
rect 20536 20878 20612 21086
rect 21080 21086 21086 21150
rect 21150 21086 21156 21150
rect 21760 21358 21766 21422
rect 21830 21358 21836 21422
rect 22037 21422 22103 21423
rect 22037 21390 22038 21422
rect 21760 21150 21836 21358
rect 21760 21118 21766 21150
rect 21080 21080 21156 21086
rect 21765 21086 21766 21118
rect 21830 21118 21836 21150
rect 22032 21358 22038 21390
rect 22102 21390 22103 21422
rect 22102 21358 22108 21390
rect 22032 21150 22108 21358
rect 21830 21086 21831 21118
rect 21765 21085 21831 21086
rect 22032 21086 22038 21150
rect 22102 21086 22108 21150
rect 68952 21150 69028 21494
rect 69088 21422 69164 21766
rect 73848 21766 73854 21798
rect 73918 21798 73919 21830
rect 74397 21830 74463 21831
rect 74397 21798 74398 21830
rect 73918 21766 73924 21798
rect 73848 21558 73924 21766
rect 73848 21494 73854 21558
rect 73918 21494 73924 21558
rect 73848 21488 73924 21494
rect 74392 21766 74398 21798
rect 74462 21798 74463 21830
rect 74462 21766 74468 21798
rect 74392 21558 74468 21766
rect 74392 21494 74398 21558
rect 74462 21494 74468 21558
rect 74392 21488 74468 21494
rect 69088 21358 69094 21422
rect 69158 21358 69164 21422
rect 73989 21422 74055 21423
rect 73989 21390 73990 21422
rect 69088 21352 69164 21358
rect 73984 21358 73990 21390
rect 74054 21390 74055 21422
rect 74392 21422 74468 21428
rect 74054 21358 74060 21390
rect 68952 21118 68958 21150
rect 22032 21080 22108 21086
rect 68957 21086 68958 21118
rect 69022 21118 69028 21150
rect 73984 21150 74060 21358
rect 69022 21086 69023 21118
rect 68957 21085 69023 21086
rect 73984 21086 73990 21150
rect 74054 21086 74060 21150
rect 74392 21358 74398 21422
rect 74462 21358 74468 21422
rect 74392 21150 74468 21358
rect 74392 21118 74398 21150
rect 73984 21080 74060 21086
rect 74397 21086 74398 21118
rect 74462 21118 74468 21150
rect 75072 21422 75148 21428
rect 75072 21358 75078 21422
rect 75142 21358 75148 21422
rect 75072 21150 75148 21358
rect 75072 21118 75078 21150
rect 74462 21086 74463 21118
rect 74397 21085 74463 21086
rect 75077 21086 75078 21118
rect 75142 21118 75148 21150
rect 75485 21150 75551 21151
rect 75485 21118 75486 21150
rect 75142 21086 75143 21118
rect 75077 21085 75143 21086
rect 75480 21086 75486 21118
rect 75550 21118 75551 21150
rect 75550 21086 75556 21118
rect 18702 20814 18703 20846
rect 18637 20813 18703 20814
rect 20536 20814 20542 20878
rect 20606 20814 20612 20878
rect 27205 20878 27271 20879
rect 27205 20846 27206 20878
rect 20536 20808 20612 20814
rect 27200 20814 27206 20846
rect 27270 20846 27271 20878
rect 69093 20878 69159 20879
rect 69093 20846 69094 20878
rect 27270 20814 27276 20846
rect 20400 20742 20476 20748
rect 20400 20678 20406 20742
rect 20470 20678 20476 20742
rect 21493 20742 21559 20743
rect 21493 20710 21494 20742
rect 16456 20606 16532 20612
rect 16456 20542 16462 20606
rect 16526 20542 16532 20606
rect 3808 20470 3884 20476
rect 3808 20406 3814 20470
rect 3878 20406 3884 20470
rect 3808 17750 3884 20406
rect 16456 20062 16532 20542
rect 16456 20030 16462 20062
rect 16461 19998 16462 20030
rect 16526 20030 16532 20062
rect 17408 20606 17484 20612
rect 17408 20542 17414 20606
rect 17478 20542 17484 20606
rect 17408 20062 17484 20542
rect 17408 20030 17414 20062
rect 16526 19998 16527 20030
rect 16461 19997 16527 19998
rect 17413 19998 17414 20030
rect 17478 20030 17484 20062
rect 17816 20606 17892 20612
rect 17816 20542 17822 20606
rect 17886 20542 17892 20606
rect 17816 20062 17892 20542
rect 17816 20030 17822 20062
rect 17478 19998 17479 20030
rect 17413 19997 17479 19998
rect 17821 19998 17822 20030
rect 17886 20030 17892 20062
rect 18360 20606 18436 20612
rect 18360 20542 18366 20606
rect 18430 20542 18436 20606
rect 18360 20062 18436 20542
rect 18360 20030 18366 20062
rect 17886 19998 17887 20030
rect 17821 19997 17887 19998
rect 18365 19998 18366 20030
rect 18430 20030 18436 20062
rect 18768 20606 18844 20612
rect 18768 20542 18774 20606
rect 18838 20542 18844 20606
rect 18768 20062 18844 20542
rect 20400 20470 20476 20678
rect 20400 20438 20406 20470
rect 20405 20406 20406 20438
rect 20470 20438 20476 20470
rect 21488 20678 21494 20710
rect 21558 20710 21559 20742
rect 21558 20678 21564 20710
rect 21488 20470 21564 20678
rect 20470 20406 20471 20438
rect 20405 20405 20471 20406
rect 21488 20406 21494 20470
rect 21558 20406 21564 20470
rect 26933 20470 26999 20471
rect 26933 20438 26934 20470
rect 21488 20400 21564 20406
rect 26928 20406 26934 20438
rect 26998 20438 26999 20470
rect 27200 20470 27276 20814
rect 69088 20814 69094 20846
rect 69158 20846 69159 20878
rect 75480 20878 75556 21086
rect 69158 20814 69164 20846
rect 69088 20606 69164 20814
rect 75480 20814 75486 20878
rect 75550 20814 75556 20878
rect 77384 20878 77460 22174
rect 78477 22102 78543 22103
rect 78477 22070 78478 22102
rect 77384 20846 77390 20878
rect 75480 20808 75556 20814
rect 77389 20814 77390 20846
rect 77454 20846 77460 20878
rect 78472 22038 78478 22070
rect 78542 22070 78543 22102
rect 78542 22038 78548 22070
rect 78472 20878 78548 22038
rect 77454 20814 77455 20846
rect 77389 20813 77455 20814
rect 78472 20814 78478 20878
rect 78542 20814 78548 20878
rect 78472 20808 78548 20814
rect 69088 20542 69094 20606
rect 69158 20542 69164 20606
rect 69088 20536 69164 20542
rect 74664 20742 74740 20748
rect 74664 20678 74670 20742
rect 74734 20678 74740 20742
rect 26998 20406 27004 20438
rect 20405 20334 20471 20335
rect 20405 20302 20406 20334
rect 18768 20030 18774 20062
rect 18430 19998 18431 20030
rect 18365 19997 18431 19998
rect 18773 19998 18774 20030
rect 18838 20030 18844 20062
rect 20400 20270 20406 20302
rect 20470 20302 20471 20334
rect 20470 20270 20476 20302
rect 20400 20062 20476 20270
rect 26928 20198 27004 20406
rect 27200 20406 27206 20470
rect 27270 20406 27276 20470
rect 74664 20470 74740 20678
rect 74664 20438 74670 20470
rect 27200 20400 27276 20406
rect 74669 20406 74670 20438
rect 74734 20438 74740 20470
rect 75480 20742 75556 20748
rect 75480 20678 75486 20742
rect 75550 20678 75556 20742
rect 75480 20470 75556 20678
rect 75480 20438 75486 20470
rect 74734 20406 74735 20438
rect 74669 20405 74735 20406
rect 75485 20406 75486 20438
rect 75550 20438 75556 20470
rect 77656 20606 77732 20612
rect 77656 20542 77662 20606
rect 77726 20542 77732 20606
rect 75550 20406 75551 20438
rect 75485 20405 75551 20406
rect 75485 20334 75551 20335
rect 75485 20302 75486 20334
rect 75480 20270 75486 20302
rect 75550 20302 75551 20334
rect 75550 20270 75556 20302
rect 26928 20134 26934 20198
rect 26998 20134 27004 20198
rect 26928 20128 27004 20134
rect 27064 20198 27140 20204
rect 27064 20134 27070 20198
rect 27134 20134 27140 20198
rect 18838 19998 18839 20030
rect 18773 19997 18839 19998
rect 20400 19998 20406 20062
rect 20470 19998 20476 20062
rect 20400 19992 20476 19998
rect 18229 19926 18295 19927
rect 18229 19894 18230 19926
rect 18224 19862 18230 19894
rect 18294 19894 18295 19926
rect 18637 19926 18703 19927
rect 18637 19894 18638 19926
rect 18294 19862 18300 19894
rect 18224 18430 18300 19862
rect 18224 18366 18230 18430
rect 18294 18366 18300 18430
rect 18224 18360 18300 18366
rect 18632 19862 18638 19894
rect 18702 19894 18703 19926
rect 20405 19926 20471 19927
rect 20405 19894 20406 19926
rect 18702 19862 18708 19894
rect 18632 18430 18708 19862
rect 20400 19862 20406 19894
rect 20470 19894 20471 19926
rect 20813 19926 20879 19927
rect 20813 19894 20814 19926
rect 20470 19862 20476 19894
rect 20400 19654 20476 19862
rect 20400 19590 20406 19654
rect 20470 19590 20476 19654
rect 20400 19584 20476 19590
rect 20808 19862 20814 19894
rect 20878 19894 20879 19926
rect 21488 19926 21564 19932
rect 20878 19862 20884 19894
rect 20808 19654 20884 19862
rect 20808 19590 20814 19654
rect 20878 19590 20884 19654
rect 21488 19862 21494 19926
rect 21558 19862 21564 19926
rect 21488 19654 21564 19862
rect 21488 19622 21494 19654
rect 20808 19584 20884 19590
rect 21493 19590 21494 19622
rect 21558 19622 21564 19654
rect 21624 19926 21700 19932
rect 21624 19862 21630 19926
rect 21694 19862 21700 19926
rect 22037 19926 22103 19927
rect 22037 19894 22038 19926
rect 21624 19654 21700 19862
rect 21624 19622 21630 19654
rect 21558 19590 21559 19622
rect 21493 19589 21559 19590
rect 21629 19590 21630 19622
rect 21694 19622 21700 19654
rect 22032 19862 22038 19894
rect 22102 19894 22103 19926
rect 27064 19926 27140 20134
rect 27064 19894 27070 19926
rect 22102 19862 22108 19894
rect 22032 19654 22108 19862
rect 27069 19862 27070 19894
rect 27134 19894 27140 19926
rect 69088 20062 69164 20068
rect 69088 19998 69094 20062
rect 69158 19998 69164 20062
rect 27134 19862 27135 19894
rect 27069 19861 27135 19862
rect 21694 19590 21695 19622
rect 21629 19589 21695 19590
rect 22032 19590 22038 19654
rect 22102 19590 22108 19654
rect 69088 19654 69164 19998
rect 75480 20062 75556 20270
rect 75480 19998 75486 20062
rect 75550 19998 75556 20062
rect 77656 20062 77732 20542
rect 77656 20030 77662 20062
rect 75480 19992 75556 19998
rect 77661 19998 77662 20030
rect 77726 20030 77732 20062
rect 78200 20606 78276 20612
rect 78200 20542 78206 20606
rect 78270 20542 78276 20606
rect 78200 20062 78276 20542
rect 78200 20030 78206 20062
rect 77726 19998 77727 20030
rect 77661 19997 77727 19998
rect 78205 19998 78206 20030
rect 78270 20030 78276 20062
rect 78608 20606 78684 20612
rect 78608 20542 78614 20606
rect 78678 20542 78684 20606
rect 78608 20062 78684 20542
rect 79429 20470 79495 20471
rect 79429 20438 79430 20470
rect 78608 20030 78614 20062
rect 78270 19998 78271 20030
rect 78205 19997 78271 19998
rect 78613 19998 78614 20030
rect 78678 20030 78684 20062
rect 79424 20406 79430 20438
rect 79494 20438 79495 20470
rect 94656 20470 95004 22310
rect 79494 20406 79500 20438
rect 79424 20062 79500 20406
rect 78678 19998 78679 20030
rect 78613 19997 78679 19998
rect 79424 19998 79430 20062
rect 79494 19998 79500 20062
rect 79424 19992 79500 19998
rect 94656 20406 94662 20470
rect 94726 20406 95004 20470
rect 69088 19622 69094 19654
rect 22032 19584 22108 19590
rect 69093 19590 69094 19622
rect 69158 19622 69164 19654
rect 73848 19926 73924 19932
rect 73848 19862 73854 19926
rect 73918 19862 73924 19926
rect 74261 19926 74327 19927
rect 74261 19894 74262 19926
rect 73848 19654 73924 19862
rect 73848 19622 73854 19654
rect 69158 19590 69159 19622
rect 69093 19589 69159 19590
rect 73853 19590 73854 19622
rect 73918 19622 73924 19654
rect 74256 19862 74262 19894
rect 74326 19894 74327 19926
rect 75621 19926 75687 19927
rect 75621 19894 75622 19926
rect 74326 19862 74332 19894
rect 74256 19654 74332 19862
rect 73918 19590 73919 19622
rect 73853 19589 73919 19590
rect 74256 19590 74262 19654
rect 74326 19590 74332 19654
rect 74256 19584 74332 19590
rect 75616 19862 75622 19894
rect 75686 19894 75687 19926
rect 78200 19926 78276 19932
rect 75686 19862 75692 19894
rect 75616 19654 75692 19862
rect 75616 19590 75622 19654
rect 75686 19590 75692 19654
rect 75616 19584 75692 19590
rect 78200 19862 78206 19926
rect 78270 19862 78276 19926
rect 78613 19926 78679 19927
rect 78613 19894 78614 19926
rect 20400 19518 20476 19524
rect 20400 19454 20406 19518
rect 20470 19454 20476 19518
rect 20400 19246 20476 19454
rect 20400 19214 20406 19246
rect 20405 19182 20406 19214
rect 20470 19214 20476 19246
rect 20944 19518 21020 19524
rect 20944 19454 20950 19518
rect 21014 19454 21020 19518
rect 21629 19518 21695 19519
rect 21629 19486 21630 19518
rect 20944 19246 21020 19454
rect 20944 19214 20950 19246
rect 20470 19182 20471 19214
rect 20405 19181 20471 19182
rect 20949 19182 20950 19214
rect 21014 19214 21020 19246
rect 21624 19454 21630 19486
rect 21694 19486 21695 19518
rect 22173 19518 22239 19519
rect 22173 19486 22174 19518
rect 21694 19454 21700 19486
rect 21624 19246 21700 19454
rect 21014 19182 21015 19214
rect 20949 19181 21015 19182
rect 21624 19182 21630 19246
rect 21694 19182 21700 19246
rect 21624 19176 21700 19182
rect 22168 19454 22174 19486
rect 22238 19486 22239 19518
rect 73853 19518 73919 19519
rect 73853 19486 73854 19518
rect 22238 19454 22244 19486
rect 22168 19246 22244 19454
rect 22168 19182 22174 19246
rect 22238 19182 22244 19246
rect 22168 19176 22244 19182
rect 73848 19454 73854 19486
rect 73918 19486 73919 19518
rect 74256 19518 74332 19524
rect 73918 19454 73924 19486
rect 73848 19246 73924 19454
rect 73848 19182 73854 19246
rect 73918 19182 73924 19246
rect 74256 19454 74262 19518
rect 74326 19454 74332 19518
rect 75213 19518 75279 19519
rect 75213 19486 75214 19518
rect 74256 19246 74332 19454
rect 74256 19214 74262 19246
rect 73848 19176 73924 19182
rect 74261 19182 74262 19214
rect 74326 19214 74332 19246
rect 75208 19454 75214 19486
rect 75278 19486 75279 19518
rect 75480 19518 75556 19524
rect 75278 19454 75284 19486
rect 75208 19246 75284 19454
rect 74326 19182 74327 19214
rect 74261 19181 74327 19182
rect 75208 19182 75214 19246
rect 75278 19182 75284 19246
rect 75480 19454 75486 19518
rect 75550 19454 75556 19518
rect 75480 19246 75556 19454
rect 75480 19214 75486 19246
rect 75208 19176 75284 19182
rect 75485 19182 75486 19214
rect 75550 19214 75556 19246
rect 75550 19182 75551 19214
rect 75485 19181 75551 19182
rect 20405 19110 20471 19111
rect 20405 19078 20406 19110
rect 20400 19046 20406 19078
rect 20470 19078 20471 19110
rect 21357 19110 21423 19111
rect 21357 19078 21358 19110
rect 20470 19046 20476 19078
rect 20400 18838 20476 19046
rect 20400 18774 20406 18838
rect 20470 18774 20476 18838
rect 20400 18768 20476 18774
rect 21352 19046 21358 19078
rect 21422 19078 21423 19110
rect 21624 19110 21700 19116
rect 21422 19046 21428 19078
rect 21352 18838 21428 19046
rect 21352 18774 21358 18838
rect 21422 18774 21428 18838
rect 21624 19046 21630 19110
rect 21694 19046 21700 19110
rect 21624 18838 21700 19046
rect 21624 18806 21630 18838
rect 21352 18768 21428 18774
rect 21629 18774 21630 18806
rect 21694 18806 21700 18838
rect 22032 19110 22108 19116
rect 22032 19046 22038 19110
rect 22102 19046 22108 19110
rect 22032 18838 22108 19046
rect 22032 18806 22038 18838
rect 21694 18774 21695 18806
rect 21629 18773 21695 18774
rect 22037 18774 22038 18806
rect 22102 18806 22108 18838
rect 73848 19110 73924 19116
rect 73848 19046 73854 19110
rect 73918 19046 73924 19110
rect 73848 18838 73924 19046
rect 73848 18806 73854 18838
rect 22102 18774 22103 18806
rect 22037 18773 22103 18774
rect 73853 18774 73854 18806
rect 73918 18806 73924 18838
rect 74256 19110 74332 19116
rect 74256 19046 74262 19110
rect 74326 19046 74332 19110
rect 74256 18838 74332 19046
rect 74256 18806 74262 18838
rect 73918 18774 73919 18806
rect 73853 18773 73919 18774
rect 74261 18774 74262 18806
rect 74326 18806 74332 18838
rect 74800 19110 74876 19116
rect 74800 19046 74806 19110
rect 74870 19046 74876 19110
rect 75485 19110 75551 19111
rect 75485 19078 75486 19110
rect 74800 18838 74876 19046
rect 74800 18806 74806 18838
rect 74326 18774 74327 18806
rect 74261 18773 74327 18774
rect 74805 18774 74806 18806
rect 74870 18806 74876 18838
rect 75480 19046 75486 19078
rect 75550 19078 75551 19110
rect 75550 19046 75556 19078
rect 75480 18838 75556 19046
rect 74870 18774 74871 18806
rect 74805 18773 74871 18774
rect 75480 18774 75486 18838
rect 75550 18774 75556 18838
rect 75480 18768 75556 18774
rect 20405 18702 20471 18703
rect 20405 18670 20406 18702
rect 18632 18366 18638 18430
rect 18702 18366 18708 18430
rect 18632 18360 18708 18366
rect 20400 18638 20406 18670
rect 20470 18670 20471 18702
rect 20813 18702 20879 18703
rect 20813 18670 20814 18702
rect 20470 18638 20476 18670
rect 20400 18430 20476 18638
rect 20400 18366 20406 18430
rect 20470 18366 20476 18430
rect 20400 18360 20476 18366
rect 20808 18638 20814 18670
rect 20878 18670 20879 18702
rect 21221 18702 21287 18703
rect 21221 18670 21222 18702
rect 20878 18638 20884 18670
rect 20808 18430 20884 18638
rect 20808 18366 20814 18430
rect 20878 18366 20884 18430
rect 20808 18360 20884 18366
rect 21216 18638 21222 18670
rect 21286 18670 21287 18702
rect 21624 18702 21700 18708
rect 21286 18638 21292 18670
rect 21216 18430 21292 18638
rect 21216 18366 21222 18430
rect 21286 18366 21292 18430
rect 21624 18638 21630 18702
rect 21694 18638 21700 18702
rect 22037 18702 22103 18703
rect 22037 18670 22038 18702
rect 21624 18430 21700 18638
rect 21624 18398 21630 18430
rect 21216 18360 21292 18366
rect 21629 18366 21630 18398
rect 21694 18398 21700 18430
rect 22032 18638 22038 18670
rect 22102 18670 22103 18702
rect 73853 18702 73919 18703
rect 73853 18670 73854 18702
rect 22102 18638 22108 18670
rect 22032 18430 22108 18638
rect 21694 18366 21695 18398
rect 21629 18365 21695 18366
rect 22032 18366 22038 18430
rect 22102 18366 22108 18430
rect 22032 18360 22108 18366
rect 73848 18638 73854 18670
rect 73918 18670 73919 18702
rect 74261 18702 74327 18703
rect 74261 18670 74262 18702
rect 73918 18638 73924 18670
rect 73848 18430 73924 18638
rect 73848 18366 73854 18430
rect 73918 18366 73924 18430
rect 73848 18360 73924 18366
rect 74256 18638 74262 18670
rect 74326 18670 74327 18702
rect 75072 18702 75148 18708
rect 74326 18638 74332 18670
rect 74256 18430 74332 18638
rect 74256 18366 74262 18430
rect 74326 18366 74332 18430
rect 75072 18638 75078 18702
rect 75142 18638 75148 18702
rect 75072 18430 75148 18638
rect 75072 18398 75078 18430
rect 74256 18360 74332 18366
rect 75077 18366 75078 18398
rect 75142 18398 75148 18430
rect 75616 18702 75692 18708
rect 75616 18638 75622 18702
rect 75686 18638 75692 18702
rect 75616 18430 75692 18638
rect 75616 18398 75622 18430
rect 75142 18366 75143 18398
rect 75077 18365 75143 18366
rect 75621 18366 75622 18398
rect 75686 18398 75692 18430
rect 77928 18702 78004 18708
rect 77928 18638 77934 18702
rect 77998 18638 78004 18702
rect 77928 18430 78004 18638
rect 77928 18398 77934 18430
rect 75686 18366 75687 18398
rect 75621 18365 75687 18366
rect 77933 18366 77934 18398
rect 77998 18398 78004 18430
rect 78200 18430 78276 19862
rect 78608 19862 78614 19894
rect 78678 19894 78679 19926
rect 78678 19862 78684 19894
rect 78477 18702 78543 18703
rect 78477 18670 78478 18702
rect 78200 18398 78206 18430
rect 77998 18366 77999 18398
rect 77933 18365 77999 18366
rect 78205 18366 78206 18398
rect 78270 18398 78276 18430
rect 78472 18638 78478 18670
rect 78542 18670 78543 18702
rect 78542 18638 78548 18670
rect 78472 18430 78548 18638
rect 78270 18366 78271 18398
rect 78205 18365 78271 18366
rect 78472 18366 78478 18430
rect 78542 18366 78548 18430
rect 78472 18360 78548 18366
rect 78608 18430 78684 19862
rect 78608 18366 78614 18430
rect 78678 18366 78684 18430
rect 78608 18360 78684 18366
rect 94656 18838 95004 20406
rect 94656 18774 94662 18838
rect 94726 18774 95004 18838
rect 3808 17718 3814 17750
rect 3813 17686 3814 17718
rect 3878 17718 3884 17750
rect 17544 18294 17620 18300
rect 17544 18230 17550 18294
rect 17614 18230 17620 18294
rect 3878 17686 3879 17718
rect 3813 17685 3879 17686
rect 3808 17614 3884 17620
rect 3808 17550 3814 17614
rect 3878 17550 3884 17614
rect 17544 17614 17620 18230
rect 17544 17582 17550 17614
rect 2560 15262 2626 15263
rect 2560 15198 2561 15262
rect 2625 15198 2626 15262
rect 2560 15197 2626 15198
rect 3808 14758 3884 17550
rect 17549 17550 17550 17582
rect 17614 17582 17620 17614
rect 18224 18294 18300 18300
rect 18224 18230 18230 18294
rect 18294 18230 18300 18294
rect 18773 18294 18839 18295
rect 18773 18262 18774 18294
rect 18224 17614 18300 18230
rect 18224 17582 18230 17614
rect 17614 17550 17615 17582
rect 17549 17549 17615 17550
rect 18229 17550 18230 17582
rect 18294 17582 18300 17614
rect 18768 18230 18774 18262
rect 18838 18262 18839 18294
rect 20944 18294 21020 18300
rect 18838 18230 18844 18262
rect 18768 17614 18844 18230
rect 20944 18230 20950 18294
rect 21014 18230 21020 18294
rect 21765 18294 21831 18295
rect 21765 18262 21766 18294
rect 20944 18022 21020 18230
rect 20944 17990 20950 18022
rect 20949 17958 20950 17990
rect 21014 17990 21020 18022
rect 21760 18230 21766 18262
rect 21830 18262 21831 18294
rect 22168 18294 22244 18300
rect 21830 18230 21836 18262
rect 21760 18022 21836 18230
rect 21014 17958 21015 17990
rect 20949 17957 21015 17958
rect 21760 17958 21766 18022
rect 21830 17958 21836 18022
rect 22168 18230 22174 18294
rect 22238 18230 22244 18294
rect 22168 18022 22244 18230
rect 22168 17990 22174 18022
rect 21760 17952 21836 17958
rect 22173 17958 22174 17990
rect 22238 17990 22244 18022
rect 73984 18294 74060 18300
rect 73984 18230 73990 18294
rect 74054 18230 74060 18294
rect 73984 18022 74060 18230
rect 73984 17990 73990 18022
rect 22238 17958 22239 17990
rect 22173 17957 22239 17958
rect 73989 17958 73990 17990
rect 74054 17990 74060 18022
rect 74392 18294 74468 18300
rect 74392 18230 74398 18294
rect 74462 18230 74468 18294
rect 74669 18294 74735 18295
rect 74669 18262 74670 18294
rect 74392 18022 74468 18230
rect 74392 17990 74398 18022
rect 74054 17958 74055 17990
rect 73989 17957 74055 17958
rect 74397 17958 74398 17990
rect 74462 17990 74468 18022
rect 74664 18230 74670 18262
rect 74734 18262 74735 18294
rect 75077 18294 75143 18295
rect 75077 18262 75078 18294
rect 74734 18230 74740 18262
rect 74664 18022 74740 18230
rect 74462 17958 74463 17990
rect 74397 17957 74463 17958
rect 74664 17958 74670 18022
rect 74734 17958 74740 18022
rect 74664 17952 74740 17958
rect 75072 18230 75078 18262
rect 75142 18262 75143 18294
rect 77384 18294 77460 18300
rect 75142 18230 75148 18262
rect 75072 18022 75148 18230
rect 75072 17958 75078 18022
rect 75142 17958 75148 18022
rect 75072 17952 75148 17958
rect 77384 18230 77390 18294
rect 77454 18230 77460 18294
rect 78613 18294 78679 18295
rect 78613 18262 78614 18294
rect 18294 17550 18295 17582
rect 18229 17549 18295 17550
rect 18768 17550 18774 17614
rect 18838 17550 18844 17614
rect 20536 17886 20612 17892
rect 20536 17822 20542 17886
rect 20606 17822 20612 17886
rect 20536 17614 20612 17822
rect 20536 17582 20542 17614
rect 18768 17544 18844 17550
rect 20541 17550 20542 17582
rect 20606 17582 20612 17614
rect 21624 17886 21700 17892
rect 21624 17822 21630 17886
rect 21694 17822 21700 17886
rect 22173 17886 22239 17887
rect 22173 17854 22174 17886
rect 21624 17614 21700 17822
rect 21624 17582 21630 17614
rect 20606 17550 20607 17582
rect 20541 17549 20607 17550
rect 21629 17550 21630 17582
rect 21694 17582 21700 17614
rect 22168 17822 22174 17854
rect 22238 17854 22239 17886
rect 73848 17886 73924 17892
rect 22238 17822 22244 17854
rect 22168 17614 22244 17822
rect 21694 17550 21695 17582
rect 21629 17549 21695 17550
rect 22168 17550 22174 17614
rect 22238 17550 22244 17614
rect 73848 17822 73854 17886
rect 73918 17822 73924 17886
rect 73848 17614 73924 17822
rect 73848 17582 73854 17614
rect 22168 17544 22244 17550
rect 73853 17550 73854 17582
rect 73918 17582 73924 17614
rect 74256 17886 74332 17892
rect 74256 17822 74262 17886
rect 74326 17822 74332 17886
rect 74256 17614 74332 17822
rect 74256 17582 74262 17614
rect 73918 17550 73919 17582
rect 73853 17549 73919 17550
rect 74261 17550 74262 17582
rect 74326 17582 74332 17614
rect 74800 17886 74876 17892
rect 74800 17822 74806 17886
rect 74870 17822 74876 17886
rect 74800 17614 74876 17822
rect 74800 17582 74806 17614
rect 74326 17550 74327 17582
rect 74261 17549 74327 17550
rect 74805 17550 74806 17582
rect 74870 17582 74876 17614
rect 74936 17886 75012 17892
rect 74936 17822 74942 17886
rect 75006 17822 75012 17886
rect 74936 17614 75012 17822
rect 74936 17582 74942 17614
rect 74870 17550 74871 17582
rect 74805 17549 74871 17550
rect 74941 17550 74942 17582
rect 75006 17582 75012 17614
rect 75616 17886 75692 17892
rect 75616 17822 75622 17886
rect 75686 17822 75692 17886
rect 75616 17614 75692 17822
rect 75616 17582 75622 17614
rect 75006 17550 75007 17582
rect 74941 17549 75007 17550
rect 75621 17550 75622 17582
rect 75686 17582 75692 17614
rect 77384 17614 77460 18230
rect 77384 17582 77390 17614
rect 75686 17550 75687 17582
rect 75621 17549 75687 17550
rect 77389 17550 77390 17582
rect 77454 17582 77460 17614
rect 78608 18230 78614 18262
rect 78678 18262 78679 18294
rect 78678 18230 78684 18262
rect 78608 17614 78684 18230
rect 79429 18158 79495 18159
rect 79429 18126 79430 18158
rect 77454 17550 77455 17582
rect 77389 17549 77455 17550
rect 78608 17550 78614 17614
rect 78678 17550 78684 17614
rect 78608 17544 78684 17550
rect 79424 18094 79430 18126
rect 79494 18126 79495 18158
rect 79494 18094 79500 18126
rect 79424 17614 79500 18094
rect 79424 17550 79430 17614
rect 79494 17550 79500 17614
rect 79424 17544 79500 17550
rect 16184 17478 16260 17484
rect 16184 17414 16190 17478
rect 16254 17414 16260 17478
rect 16184 16390 16260 17414
rect 16184 16358 16190 16390
rect 16189 16326 16190 16358
rect 16254 16358 16260 16390
rect 16592 17478 16668 17484
rect 16592 17414 16598 17478
rect 16662 17414 16668 17478
rect 20677 17478 20743 17479
rect 20677 17446 20678 17478
rect 16254 16326 16255 16358
rect 16189 16325 16255 16326
rect 14280 16254 14356 16260
rect 14280 16190 14286 16254
rect 14350 16190 14356 16254
rect 3808 14726 3814 14758
rect 3813 14694 3814 14726
rect 3878 14726 3884 14758
rect 3944 14758 4020 14764
rect 3878 14694 3879 14726
rect 3813 14693 3879 14694
rect 3944 14694 3950 14758
rect 4014 14694 4020 14758
rect 3944 14628 4020 14694
rect 3808 14552 4020 14628
rect 14144 14758 14220 14764
rect 14144 14694 14150 14758
rect 14214 14694 14220 14758
rect 952 13742 1230 13806
rect 1294 13742 1300 13806
rect 3133 13806 3199 13807
rect 3133 13774 3134 13806
rect 952 12038 1300 13742
rect 3128 13742 3134 13774
rect 3198 13774 3199 13806
rect 3198 13742 3204 13774
rect 3128 13534 3204 13742
rect 3128 13470 3134 13534
rect 3198 13470 3204 13534
rect 3128 13464 3204 13470
rect 952 11974 1230 12038
rect 1294 11974 1300 12038
rect 3808 12038 3884 14552
rect 3808 12006 3814 12038
rect 952 10542 1300 11974
rect 3813 11974 3814 12006
rect 3878 12006 3884 12038
rect 14008 13398 14084 13404
rect 14008 13334 14014 13398
rect 14078 13334 14084 13398
rect 3878 11974 3879 12006
rect 3813 11973 3879 11974
rect 14008 10678 14084 13334
rect 14144 12038 14220 14694
rect 14280 13534 14356 16190
rect 16592 14894 16668 17414
rect 16592 14862 16598 14894
rect 16597 14830 16598 14862
rect 16662 14862 16668 14894
rect 20672 17414 20678 17446
rect 20742 17446 20743 17478
rect 22037 17478 22103 17479
rect 22037 17446 22038 17478
rect 20742 17414 20748 17446
rect 16662 14830 16663 14862
rect 16597 14829 16663 14830
rect 20672 14758 20748 17414
rect 22032 17414 22038 17446
rect 22102 17446 22103 17478
rect 22853 17478 22919 17479
rect 22853 17446 22854 17478
rect 22102 17414 22108 17446
rect 22032 17070 22108 17414
rect 22032 17006 22038 17070
rect 22102 17006 22108 17070
rect 22032 17000 22108 17006
rect 22848 17414 22854 17446
rect 22918 17446 22919 17478
rect 79701 17478 79767 17479
rect 79701 17446 79702 17478
rect 22918 17414 22924 17446
rect 22848 17070 22924 17414
rect 79696 17414 79702 17446
rect 79766 17446 79767 17478
rect 82421 17478 82487 17479
rect 82421 17446 82422 17478
rect 79766 17414 79772 17446
rect 22848 17006 22854 17070
rect 22918 17006 22924 17070
rect 28565 17070 28631 17071
rect 28565 17038 28566 17070
rect 22848 17000 22924 17006
rect 28560 17006 28566 17038
rect 28630 17038 28631 17070
rect 28630 17006 28636 17038
rect 20672 14694 20678 14758
rect 20742 14694 20748 14758
rect 20672 14688 20748 14694
rect 22032 16934 22108 16940
rect 22032 16870 22038 16934
rect 22102 16870 22108 16934
rect 26525 16934 26591 16935
rect 26525 16902 26526 16934
rect 21085 14622 21151 14623
rect 21085 14590 21086 14622
rect 14280 13502 14286 13534
rect 14285 13470 14286 13502
rect 14350 13502 14356 13534
rect 21080 14558 21086 14590
rect 21150 14590 21151 14622
rect 21150 14558 21156 14590
rect 14350 13470 14351 13502
rect 14285 13469 14351 13470
rect 14144 12006 14150 12038
rect 14149 11974 14150 12006
rect 14214 12006 14220 12038
rect 14214 11974 14215 12006
rect 14149 11973 14215 11974
rect 14285 11902 14351 11903
rect 14285 11870 14286 11902
rect 14008 10646 14014 10678
rect 14013 10614 14014 10646
rect 14078 10646 14084 10678
rect 14280 11838 14286 11870
rect 14350 11870 14351 11902
rect 21080 11902 21156 14558
rect 22032 13262 22108 16870
rect 26520 16870 26526 16902
rect 26590 16902 26591 16934
rect 26590 16870 26596 16902
rect 26520 16662 26596 16870
rect 26520 16598 26526 16662
rect 26590 16598 26596 16662
rect 26520 16592 26596 16598
rect 28288 16526 28364 16532
rect 28288 16462 28294 16526
rect 28358 16462 28364 16526
rect 28288 16118 28364 16462
rect 28288 16086 28294 16118
rect 28293 16054 28294 16086
rect 28358 16086 28364 16118
rect 28358 16054 28359 16086
rect 28293 16053 28359 16054
rect 28560 14622 28636 17006
rect 30464 16662 30540 16668
rect 30464 16598 30470 16662
rect 30534 16598 30540 16662
rect 29240 16526 29316 16532
rect 29240 16462 29246 16526
rect 29310 16462 29316 16526
rect 29240 16118 29316 16462
rect 29240 16086 29246 16118
rect 29245 16054 29246 16086
rect 29310 16086 29316 16118
rect 30464 16118 30540 16598
rect 64192 16662 64268 16668
rect 64192 16598 64198 16662
rect 64262 16598 64268 16662
rect 31557 16526 31623 16527
rect 31557 16494 31558 16526
rect 30464 16086 30470 16118
rect 29310 16054 29311 16086
rect 29245 16053 29311 16054
rect 30469 16054 30470 16086
rect 30534 16086 30540 16118
rect 31552 16462 31558 16494
rect 31622 16494 31623 16526
rect 32096 16526 32172 16532
rect 31622 16462 31628 16494
rect 31552 16118 31628 16462
rect 30534 16054 30535 16086
rect 30469 16053 30535 16054
rect 31552 16054 31558 16118
rect 31622 16054 31628 16118
rect 32096 16462 32102 16526
rect 32166 16462 32172 16526
rect 32781 16526 32847 16527
rect 32781 16494 32782 16526
rect 32096 16118 32172 16462
rect 32096 16086 32102 16118
rect 31552 16048 31628 16054
rect 32101 16054 32102 16086
rect 32166 16086 32172 16118
rect 32776 16462 32782 16494
rect 32846 16494 32847 16526
rect 33320 16526 33396 16532
rect 32846 16462 32852 16494
rect 32776 16118 32852 16462
rect 32166 16054 32167 16086
rect 32101 16053 32167 16054
rect 32776 16054 32782 16118
rect 32846 16054 32852 16118
rect 33320 16462 33326 16526
rect 33390 16462 33396 16526
rect 34141 16526 34207 16527
rect 34141 16494 34142 16526
rect 33320 16118 33396 16462
rect 33320 16086 33326 16118
rect 32776 16048 32852 16054
rect 33325 16054 33326 16086
rect 33390 16086 33396 16118
rect 34136 16462 34142 16494
rect 34206 16494 34207 16526
rect 34544 16526 34620 16532
rect 34206 16462 34212 16494
rect 34136 16118 34212 16462
rect 33390 16054 33391 16086
rect 33325 16053 33391 16054
rect 34136 16054 34142 16118
rect 34206 16054 34212 16118
rect 34544 16462 34550 16526
rect 34614 16462 34620 16526
rect 34544 16118 34620 16462
rect 34544 16086 34550 16118
rect 34136 16048 34212 16054
rect 34549 16054 34550 16086
rect 34614 16086 34620 16118
rect 35768 16526 35844 16532
rect 35768 16462 35774 16526
rect 35838 16462 35844 16526
rect 36589 16526 36655 16527
rect 36589 16494 36590 16526
rect 35768 16118 35844 16462
rect 35768 16086 35774 16118
rect 34614 16054 34615 16086
rect 34549 16053 34615 16054
rect 35773 16054 35774 16086
rect 35838 16086 35844 16118
rect 36584 16462 36590 16494
rect 36654 16494 36655 16526
rect 38352 16526 38428 16532
rect 36654 16462 36660 16494
rect 36584 16118 36660 16462
rect 35838 16054 35839 16086
rect 35773 16053 35839 16054
rect 36584 16054 36590 16118
rect 36654 16054 36660 16118
rect 38352 16462 38358 16526
rect 38422 16462 38428 16526
rect 39037 16526 39103 16527
rect 39037 16494 39038 16526
rect 38352 16118 38428 16462
rect 38352 16086 38358 16118
rect 36584 16048 36660 16054
rect 38357 16054 38358 16086
rect 38422 16086 38428 16118
rect 39032 16462 39038 16494
rect 39102 16494 39103 16526
rect 39576 16526 39652 16532
rect 39102 16462 39108 16494
rect 39032 16118 39108 16462
rect 38422 16054 38423 16086
rect 38357 16053 38423 16054
rect 39032 16054 39038 16118
rect 39102 16054 39108 16118
rect 39576 16462 39582 16526
rect 39646 16462 39652 16526
rect 40261 16526 40327 16527
rect 40261 16494 40262 16526
rect 39576 16118 39652 16462
rect 39576 16086 39582 16118
rect 39032 16048 39108 16054
rect 39581 16054 39582 16086
rect 39646 16086 39652 16118
rect 40256 16462 40262 16494
rect 40326 16494 40327 16526
rect 40800 16526 40876 16532
rect 40326 16462 40332 16494
rect 40256 16118 40332 16462
rect 39646 16054 39647 16086
rect 39581 16053 39647 16054
rect 40256 16054 40262 16118
rect 40326 16054 40332 16118
rect 40800 16462 40806 16526
rect 40870 16462 40876 16526
rect 40800 16118 40876 16462
rect 40800 16086 40806 16118
rect 40256 16048 40332 16054
rect 40805 16054 40806 16086
rect 40870 16086 40876 16118
rect 42024 16526 42100 16532
rect 42024 16462 42030 16526
rect 42094 16462 42100 16526
rect 42845 16526 42911 16527
rect 42845 16494 42846 16526
rect 42024 16118 42100 16462
rect 42024 16086 42030 16118
rect 40870 16054 40871 16086
rect 40805 16053 40871 16054
rect 42029 16054 42030 16086
rect 42094 16086 42100 16118
rect 42840 16462 42846 16494
rect 42910 16494 42911 16526
rect 44608 16526 44684 16532
rect 42910 16462 42916 16494
rect 42840 16118 42916 16462
rect 42094 16054 42095 16086
rect 42029 16053 42095 16054
rect 42840 16054 42846 16118
rect 42910 16054 42916 16118
rect 44608 16462 44614 16526
rect 44678 16462 44684 16526
rect 45293 16526 45359 16527
rect 45293 16494 45294 16526
rect 44608 16118 44684 16462
rect 44608 16086 44614 16118
rect 42840 16048 42916 16054
rect 44613 16054 44614 16086
rect 44678 16086 44684 16118
rect 45288 16462 45294 16494
rect 45358 16494 45359 16526
rect 45832 16526 45908 16532
rect 45358 16462 45364 16494
rect 45288 16118 45364 16462
rect 44678 16054 44679 16086
rect 44613 16053 44679 16054
rect 45288 16054 45294 16118
rect 45358 16054 45364 16118
rect 45832 16462 45838 16526
rect 45902 16462 45908 16526
rect 46517 16526 46583 16527
rect 46517 16494 46518 16526
rect 45832 16118 45908 16462
rect 45832 16086 45838 16118
rect 45288 16048 45364 16054
rect 45837 16054 45838 16086
rect 45902 16086 45908 16118
rect 46512 16462 46518 16494
rect 46582 16494 46583 16526
rect 47056 16526 47132 16532
rect 46582 16462 46588 16494
rect 46512 16118 46588 16462
rect 45902 16054 45903 16086
rect 45837 16053 45903 16054
rect 46512 16054 46518 16118
rect 46582 16054 46588 16118
rect 47056 16462 47062 16526
rect 47126 16462 47132 16526
rect 47741 16526 47807 16527
rect 47741 16494 47742 16526
rect 47056 16118 47132 16462
rect 47056 16086 47062 16118
rect 46512 16048 46588 16054
rect 47061 16054 47062 16086
rect 47126 16086 47132 16118
rect 47736 16462 47742 16494
rect 47806 16494 47807 16526
rect 48280 16526 48356 16532
rect 47806 16462 47812 16494
rect 47736 16118 47812 16462
rect 47126 16054 47127 16086
rect 47061 16053 47127 16054
rect 47736 16054 47742 16118
rect 47806 16054 47812 16118
rect 48280 16462 48286 16526
rect 48350 16462 48356 16526
rect 49373 16526 49439 16527
rect 49373 16494 49374 16526
rect 48280 16118 48356 16462
rect 48280 16086 48286 16118
rect 47736 16048 47812 16054
rect 48285 16054 48286 16086
rect 48350 16086 48356 16118
rect 49368 16462 49374 16494
rect 49438 16494 49439 16526
rect 50325 16526 50391 16527
rect 50325 16494 50326 16526
rect 49438 16462 49444 16494
rect 49368 16118 49444 16462
rect 48350 16054 48351 16086
rect 48285 16053 48351 16054
rect 49368 16054 49374 16118
rect 49438 16054 49444 16118
rect 49368 16048 49444 16054
rect 50320 16462 50326 16494
rect 50390 16494 50391 16526
rect 50728 16526 50804 16532
rect 50390 16462 50396 16494
rect 50320 16118 50396 16462
rect 50320 16054 50326 16118
rect 50390 16054 50396 16118
rect 50728 16462 50734 16526
rect 50798 16462 50804 16526
rect 51549 16526 51615 16527
rect 51549 16494 51550 16526
rect 50728 16118 50804 16462
rect 50728 16086 50734 16118
rect 50320 16048 50396 16054
rect 50733 16054 50734 16086
rect 50798 16086 50804 16118
rect 51544 16462 51550 16494
rect 51614 16494 51615 16526
rect 51952 16526 52028 16532
rect 51614 16462 51620 16494
rect 51544 16118 51620 16462
rect 50798 16054 50799 16086
rect 50733 16053 50799 16054
rect 51544 16054 51550 16118
rect 51614 16054 51620 16118
rect 51952 16462 51958 16526
rect 52022 16462 52028 16526
rect 51952 16118 52028 16462
rect 51952 16086 51958 16118
rect 51544 16048 51620 16054
rect 51957 16054 51958 16086
rect 52022 16086 52028 16118
rect 53312 16526 53388 16532
rect 53312 16462 53318 16526
rect 53382 16462 53388 16526
rect 53997 16526 54063 16527
rect 53997 16494 53998 16526
rect 53312 16118 53388 16462
rect 53312 16086 53318 16118
rect 52022 16054 52023 16086
rect 51957 16053 52023 16054
rect 53317 16054 53318 16086
rect 53382 16086 53388 16118
rect 53992 16462 53998 16494
rect 54062 16494 54063 16526
rect 54536 16526 54612 16532
rect 54062 16462 54068 16494
rect 53992 16118 54068 16462
rect 53382 16054 53383 16086
rect 53317 16053 53383 16054
rect 53992 16054 53998 16118
rect 54062 16054 54068 16118
rect 54536 16462 54542 16526
rect 54606 16462 54612 16526
rect 55357 16526 55423 16527
rect 55357 16494 55358 16526
rect 54536 16118 54612 16462
rect 54536 16086 54542 16118
rect 53992 16048 54068 16054
rect 54541 16054 54542 16086
rect 54606 16086 54612 16118
rect 55352 16462 55358 16494
rect 55422 16494 55423 16526
rect 55760 16526 55836 16532
rect 55422 16462 55428 16494
rect 55352 16118 55428 16462
rect 54606 16054 54607 16086
rect 54541 16053 54607 16054
rect 55352 16054 55358 16118
rect 55422 16054 55428 16118
rect 55760 16462 55766 16526
rect 55830 16462 55836 16526
rect 56445 16526 56511 16527
rect 56445 16494 56446 16526
rect 55760 16118 55836 16462
rect 55760 16086 55766 16118
rect 55352 16048 55428 16054
rect 55765 16054 55766 16086
rect 55830 16086 55836 16118
rect 56440 16462 56446 16494
rect 56510 16494 56511 16526
rect 56984 16526 57060 16532
rect 56510 16462 56516 16494
rect 56440 16118 56516 16462
rect 55830 16054 55831 16086
rect 55765 16053 55831 16054
rect 56440 16054 56446 16118
rect 56510 16054 56516 16118
rect 56984 16462 56990 16526
rect 57054 16462 57060 16526
rect 57805 16526 57871 16527
rect 57805 16494 57806 16526
rect 56984 16118 57060 16462
rect 56984 16086 56990 16118
rect 56440 16048 56516 16054
rect 56989 16054 56990 16086
rect 57054 16086 57060 16118
rect 57800 16462 57806 16494
rect 57870 16494 57871 16526
rect 57936 16526 58012 16532
rect 57870 16462 57876 16494
rect 57800 16118 57876 16462
rect 57054 16054 57055 16086
rect 56989 16053 57055 16054
rect 57800 16054 57806 16118
rect 57870 16054 57876 16118
rect 57936 16462 57942 16526
rect 58006 16462 58012 16526
rect 59029 16526 59095 16527
rect 59029 16494 59030 16526
rect 57936 16118 58012 16462
rect 57936 16086 57942 16118
rect 57800 16048 57876 16054
rect 57941 16054 57942 16086
rect 58006 16086 58012 16118
rect 59024 16462 59030 16494
rect 59094 16494 59095 16526
rect 59568 16526 59644 16532
rect 59094 16462 59100 16494
rect 59024 16118 59100 16462
rect 58006 16054 58007 16086
rect 57941 16053 58007 16054
rect 59024 16054 59030 16118
rect 59094 16054 59100 16118
rect 59568 16462 59574 16526
rect 59638 16462 59644 16526
rect 60253 16526 60319 16527
rect 60253 16494 60254 16526
rect 59568 16118 59644 16462
rect 59568 16086 59574 16118
rect 59024 16048 59100 16054
rect 59573 16054 59574 16086
rect 59638 16086 59644 16118
rect 60248 16462 60254 16494
rect 60318 16494 60319 16526
rect 60792 16526 60868 16532
rect 60318 16462 60324 16494
rect 60248 16118 60324 16462
rect 59638 16054 59639 16086
rect 59573 16053 59639 16054
rect 60248 16054 60254 16118
rect 60318 16054 60324 16118
rect 60792 16462 60798 16526
rect 60862 16462 60868 16526
rect 60792 16118 60868 16462
rect 60792 16086 60798 16118
rect 60248 16048 60324 16054
rect 60797 16054 60798 16086
rect 60862 16086 60868 16118
rect 62016 16526 62092 16532
rect 62016 16462 62022 16526
rect 62086 16462 62092 16526
rect 62016 16118 62092 16462
rect 62016 16086 62022 16118
rect 60862 16054 60863 16086
rect 60797 16053 60863 16054
rect 62021 16054 62022 16086
rect 62086 16086 62092 16118
rect 63240 16526 63316 16532
rect 63240 16462 63246 16526
rect 63310 16462 63316 16526
rect 63240 16118 63316 16462
rect 63240 16086 63246 16118
rect 62086 16054 62087 16086
rect 62021 16053 62087 16054
rect 63245 16054 63246 16086
rect 63310 16086 63316 16118
rect 64192 16118 64268 16598
rect 65285 16526 65351 16527
rect 65285 16494 65286 16526
rect 64192 16086 64198 16118
rect 63310 16054 63311 16086
rect 63245 16053 63311 16054
rect 64197 16054 64198 16086
rect 64262 16086 64268 16118
rect 65280 16462 65286 16494
rect 65350 16494 65351 16526
rect 65688 16526 65764 16532
rect 65350 16462 65356 16494
rect 65280 16118 65356 16462
rect 64262 16054 64263 16086
rect 64197 16053 64263 16054
rect 65280 16054 65286 16118
rect 65350 16054 65356 16118
rect 65688 16462 65694 16526
rect 65758 16462 65764 16526
rect 66509 16526 66575 16527
rect 66509 16494 66510 16526
rect 65688 16118 65764 16462
rect 65688 16086 65694 16118
rect 65280 16048 65356 16054
rect 65693 16054 65694 16086
rect 65758 16086 65764 16118
rect 66504 16462 66510 16494
rect 66574 16494 66575 16526
rect 67048 16526 67124 16532
rect 66574 16462 66580 16494
rect 66504 16118 66580 16462
rect 65758 16054 65759 16086
rect 65693 16053 65759 16054
rect 66504 16054 66510 16118
rect 66574 16054 66580 16118
rect 67048 16462 67054 16526
rect 67118 16462 67124 16526
rect 67733 16526 67799 16527
rect 67733 16494 67734 16526
rect 67048 16118 67124 16462
rect 67048 16086 67054 16118
rect 66504 16048 66580 16054
rect 67053 16054 67054 16086
rect 67118 16086 67124 16118
rect 67728 16462 67734 16494
rect 67798 16494 67799 16526
rect 68272 16526 68348 16532
rect 67798 16462 67804 16494
rect 67728 16118 67804 16462
rect 67118 16054 67119 16086
rect 67053 16053 67119 16054
rect 67728 16054 67734 16118
rect 67798 16054 67804 16118
rect 68272 16462 68278 16526
rect 68342 16462 68348 16526
rect 68272 16118 68348 16462
rect 68272 16086 68278 16118
rect 67728 16048 67804 16054
rect 68277 16054 68278 16086
rect 68342 16086 68348 16118
rect 68342 16054 68343 16086
rect 68277 16053 68343 16054
rect 28560 14558 28566 14622
rect 28630 14558 28636 14622
rect 28560 14552 28636 14558
rect 58072 15982 58148 15988
rect 58072 15918 58078 15982
rect 58142 15918 58148 15982
rect 22032 13230 22038 13262
rect 22037 13198 22038 13230
rect 22102 13230 22108 13262
rect 31144 14350 31220 14356
rect 31144 14286 31150 14350
rect 31214 14286 31220 14350
rect 22102 13198 22103 13230
rect 22037 13197 22103 13198
rect 31144 12718 31220 14286
rect 31144 12686 31150 12718
rect 31149 12654 31150 12686
rect 31214 12686 31220 12718
rect 31214 12654 31215 12686
rect 31149 12653 31215 12654
rect 58072 12038 58148 15918
rect 79696 15846 79772 17414
rect 82416 17414 82422 17446
rect 82486 17446 82487 17478
rect 82486 17414 82492 17446
rect 82416 17206 82492 17414
rect 82416 17142 82422 17206
rect 82486 17142 82492 17206
rect 82416 17136 82492 17142
rect 79696 15782 79702 15846
rect 79766 15782 79772 15846
rect 79696 15776 79772 15782
rect 82416 17070 82492 17076
rect 82416 17006 82422 17070
rect 82486 17006 82492 17070
rect 82416 14486 82492 17006
rect 94656 17070 95004 18774
rect 94656 17006 94662 17070
rect 94726 17006 95004 17070
rect 82557 15710 82623 15711
rect 82557 15678 82558 15710
rect 82416 14454 82422 14486
rect 82421 14422 82422 14454
rect 82486 14454 82492 14486
rect 82552 15646 82558 15678
rect 82622 15678 82623 15710
rect 82622 15646 82628 15678
rect 82486 14422 82487 14454
rect 82421 14421 82487 14422
rect 82285 14214 82351 14215
rect 82285 14182 82286 14214
rect 82280 14150 82286 14182
rect 82350 14182 82351 14214
rect 82350 14150 82356 14182
rect 58072 12006 58078 12038
rect 58077 11974 58078 12006
rect 58142 12006 58148 12038
rect 64600 12718 64676 12724
rect 64600 12654 64606 12718
rect 64670 12654 64676 12718
rect 58142 11974 58143 12006
rect 58077 11973 58143 11974
rect 14350 11838 14356 11870
rect 14078 10614 14079 10646
rect 14013 10613 14079 10614
rect 952 10478 1230 10542
rect 1294 10478 1300 10542
rect 14013 10542 14079 10543
rect 14013 10510 14014 10542
rect 952 8910 1300 10478
rect 952 8846 1230 8910
rect 1294 8846 1300 8910
rect 952 7006 1300 8846
rect 14008 10478 14014 10510
rect 14078 10510 14079 10542
rect 14078 10478 14084 10510
rect 14008 7822 14084 10478
rect 14280 9318 14356 11838
rect 21080 11838 21086 11902
rect 21150 11838 21156 11902
rect 28429 11902 28495 11903
rect 28429 11870 28430 11902
rect 21080 11832 21156 11838
rect 28424 11838 28430 11870
rect 28494 11870 28495 11902
rect 29789 11902 29855 11903
rect 29789 11870 29790 11902
rect 28494 11838 28500 11870
rect 28424 11222 28500 11838
rect 28424 11158 28430 11222
rect 28494 11158 28500 11222
rect 28424 11152 28500 11158
rect 29784 11838 29790 11870
rect 29854 11870 29855 11902
rect 31013 11902 31079 11903
rect 31013 11870 31014 11902
rect 29854 11838 29860 11870
rect 29784 11222 29860 11838
rect 29784 11158 29790 11222
rect 29854 11158 29860 11222
rect 29784 11152 29860 11158
rect 31008 11838 31014 11870
rect 31078 11870 31079 11902
rect 32101 11902 32167 11903
rect 32101 11870 32102 11902
rect 31078 11838 31084 11870
rect 31008 11222 31084 11838
rect 31008 11158 31014 11222
rect 31078 11158 31084 11222
rect 31008 11152 31084 11158
rect 32096 11838 32102 11870
rect 32166 11870 32167 11902
rect 33461 11902 33527 11903
rect 33461 11870 33462 11902
rect 32166 11838 32172 11870
rect 32096 11222 32172 11838
rect 32096 11158 32102 11222
rect 32166 11158 32172 11222
rect 32096 11152 32172 11158
rect 33456 11838 33462 11870
rect 33526 11870 33527 11902
rect 34685 11902 34751 11903
rect 34685 11870 34686 11902
rect 33526 11838 33532 11870
rect 33456 11222 33532 11838
rect 33456 11158 33462 11222
rect 33526 11158 33532 11222
rect 33456 11152 33532 11158
rect 34680 11838 34686 11870
rect 34750 11870 34751 11902
rect 36045 11902 36111 11903
rect 36045 11870 36046 11902
rect 34750 11838 34756 11870
rect 34680 11222 34756 11838
rect 34680 11158 34686 11222
rect 34750 11158 34756 11222
rect 34680 11152 34756 11158
rect 36040 11838 36046 11870
rect 36110 11870 36111 11902
rect 37133 11902 37199 11903
rect 37133 11870 37134 11902
rect 36110 11838 36116 11870
rect 36040 11222 36116 11838
rect 36040 11158 36046 11222
rect 36110 11158 36116 11222
rect 36040 11152 36116 11158
rect 37128 11838 37134 11870
rect 37198 11870 37199 11902
rect 38493 11902 38559 11903
rect 38493 11870 38494 11902
rect 37198 11838 37204 11870
rect 37128 11222 37204 11838
rect 37128 11158 37134 11222
rect 37198 11158 37204 11222
rect 37128 11152 37204 11158
rect 38488 11838 38494 11870
rect 38558 11870 38559 11902
rect 39717 11902 39783 11903
rect 39717 11870 39718 11902
rect 38558 11838 38564 11870
rect 38488 11222 38564 11838
rect 38488 11158 38494 11222
rect 38558 11158 38564 11222
rect 38488 11152 38564 11158
rect 39712 11838 39718 11870
rect 39782 11870 39783 11902
rect 40805 11902 40871 11903
rect 40805 11870 40806 11902
rect 39782 11838 39788 11870
rect 39712 11222 39788 11838
rect 39712 11158 39718 11222
rect 39782 11158 39788 11222
rect 39712 11152 39788 11158
rect 40800 11838 40806 11870
rect 40870 11870 40871 11902
rect 42165 11902 42231 11903
rect 42165 11870 42166 11902
rect 40870 11838 40876 11870
rect 40800 11222 40876 11838
rect 40800 11158 40806 11222
rect 40870 11158 40876 11222
rect 40800 11152 40876 11158
rect 42160 11838 42166 11870
rect 42230 11870 42231 11902
rect 43389 11902 43455 11903
rect 43389 11870 43390 11902
rect 42230 11838 42236 11870
rect 42160 11222 42236 11838
rect 42160 11158 42166 11222
rect 42230 11158 42236 11222
rect 42160 11152 42236 11158
rect 43384 11838 43390 11870
rect 43454 11870 43455 11902
rect 44749 11902 44815 11903
rect 44749 11870 44750 11902
rect 43454 11838 43460 11870
rect 43384 11222 43460 11838
rect 43384 11158 43390 11222
rect 43454 11158 43460 11222
rect 43384 11152 43460 11158
rect 44744 11838 44750 11870
rect 44814 11870 44815 11902
rect 45837 11902 45903 11903
rect 45837 11870 45838 11902
rect 44814 11838 44820 11870
rect 44744 11222 44820 11838
rect 44744 11158 44750 11222
rect 44814 11158 44820 11222
rect 44744 11152 44820 11158
rect 45832 11838 45838 11870
rect 45902 11870 45903 11902
rect 47197 11902 47263 11903
rect 47197 11870 47198 11902
rect 45902 11838 45908 11870
rect 45832 11222 45908 11838
rect 45832 11158 45838 11222
rect 45902 11158 45908 11222
rect 45832 11152 45908 11158
rect 47192 11838 47198 11870
rect 47262 11870 47263 11902
rect 48421 11902 48487 11903
rect 48421 11870 48422 11902
rect 47262 11838 47268 11870
rect 47192 11222 47268 11838
rect 47192 11158 47198 11222
rect 47262 11158 47268 11222
rect 47192 11152 47268 11158
rect 48416 11838 48422 11870
rect 48486 11870 48487 11902
rect 49781 11902 49847 11903
rect 49781 11870 49782 11902
rect 48486 11838 48492 11870
rect 48416 11222 48492 11838
rect 48416 11158 48422 11222
rect 48486 11158 48492 11222
rect 48416 11152 48492 11158
rect 49776 11838 49782 11870
rect 49846 11870 49847 11902
rect 51005 11902 51071 11903
rect 51005 11870 51006 11902
rect 49846 11838 49852 11870
rect 49776 11222 49852 11838
rect 49776 11158 49782 11222
rect 49846 11158 49852 11222
rect 49776 11152 49852 11158
rect 51000 11838 51006 11870
rect 51070 11870 51071 11902
rect 52093 11902 52159 11903
rect 52093 11870 52094 11902
rect 51070 11838 51076 11870
rect 51000 11222 51076 11838
rect 51000 11158 51006 11222
rect 51070 11158 51076 11222
rect 51000 11152 51076 11158
rect 52088 11838 52094 11870
rect 52158 11870 52159 11902
rect 53453 11902 53519 11903
rect 53453 11870 53454 11902
rect 52158 11838 52164 11870
rect 52088 11222 52164 11838
rect 52088 11158 52094 11222
rect 52158 11158 52164 11222
rect 52088 11152 52164 11158
rect 53448 11838 53454 11870
rect 53518 11870 53519 11902
rect 54541 11902 54607 11903
rect 54541 11870 54542 11902
rect 53518 11838 53524 11870
rect 53448 11222 53524 11838
rect 53448 11158 53454 11222
rect 53518 11158 53524 11222
rect 53448 11152 53524 11158
rect 54536 11838 54542 11870
rect 54606 11870 54607 11902
rect 56037 11902 56103 11903
rect 56037 11870 56038 11902
rect 54606 11838 54612 11870
rect 54536 11222 54612 11838
rect 54536 11158 54542 11222
rect 54606 11158 54612 11222
rect 54536 11152 54612 11158
rect 56032 11838 56038 11870
rect 56102 11870 56103 11902
rect 57125 11902 57191 11903
rect 57125 11870 57126 11902
rect 56102 11838 56108 11870
rect 56032 11222 56108 11838
rect 56032 11158 56038 11222
rect 56102 11158 56108 11222
rect 56032 11152 56108 11158
rect 57120 11838 57126 11870
rect 57190 11870 57191 11902
rect 58485 11902 58551 11903
rect 58485 11870 58486 11902
rect 57190 11838 57196 11870
rect 57120 11222 57196 11838
rect 57120 11158 57126 11222
rect 57190 11158 57196 11222
rect 57120 11152 57196 11158
rect 58480 11838 58486 11870
rect 58550 11870 58551 11902
rect 59709 11902 59775 11903
rect 59709 11870 59710 11902
rect 58550 11838 58556 11870
rect 58480 11222 58556 11838
rect 58480 11158 58486 11222
rect 58550 11158 58556 11222
rect 58480 11152 58556 11158
rect 59704 11838 59710 11870
rect 59774 11870 59775 11902
rect 60797 11902 60863 11903
rect 60797 11870 60798 11902
rect 59774 11838 59780 11870
rect 59704 11222 59780 11838
rect 59704 11158 59710 11222
rect 59774 11158 59780 11222
rect 59704 11152 59780 11158
rect 60792 11838 60798 11870
rect 60862 11870 60863 11902
rect 62157 11902 62223 11903
rect 62157 11870 62158 11902
rect 60862 11838 60868 11870
rect 60792 11222 60868 11838
rect 60792 11158 60798 11222
rect 60862 11158 60868 11222
rect 60792 11152 60868 11158
rect 62152 11838 62158 11870
rect 62222 11870 62223 11902
rect 63381 11902 63447 11903
rect 63381 11870 63382 11902
rect 62222 11838 62228 11870
rect 62152 11222 62228 11838
rect 62152 11158 62158 11222
rect 62222 11158 62228 11222
rect 62152 11152 62228 11158
rect 63376 11838 63382 11870
rect 63446 11870 63447 11902
rect 63446 11838 63452 11870
rect 63376 11222 63452 11838
rect 63376 11158 63382 11222
rect 63446 11158 63452 11222
rect 63376 11152 63452 11158
rect 64600 11092 64676 12654
rect 64741 11902 64807 11903
rect 64741 11870 64742 11902
rect 64736 11838 64742 11870
rect 64806 11870 64807 11902
rect 65829 11902 65895 11903
rect 65829 11870 65830 11902
rect 64806 11838 64812 11870
rect 64736 11222 64812 11838
rect 64736 11158 64742 11222
rect 64806 11158 64812 11222
rect 64736 11152 64812 11158
rect 65824 11838 65830 11870
rect 65894 11870 65895 11902
rect 67189 11902 67255 11903
rect 67189 11870 67190 11902
rect 65894 11838 65900 11870
rect 65824 11222 65900 11838
rect 65824 11158 65830 11222
rect 65894 11158 65900 11222
rect 65824 11152 65900 11158
rect 67184 11838 67190 11870
rect 67254 11870 67255 11902
rect 67254 11838 67260 11870
rect 67184 11222 67260 11838
rect 82280 11630 82356 14150
rect 82552 12990 82628 15646
rect 82552 12926 82558 12990
rect 82622 12926 82628 12990
rect 82552 12920 82628 12926
rect 94656 15438 95004 17006
rect 94656 15374 94662 15438
rect 94726 15374 95004 15438
rect 94656 13942 95004 15374
rect 94656 13878 94662 13942
rect 94726 13878 95004 13942
rect 82421 12854 82487 12855
rect 82421 12822 82422 12854
rect 82280 11566 82286 11630
rect 82350 11566 82356 11630
rect 82280 11560 82356 11566
rect 82416 12790 82422 12822
rect 82486 12822 82487 12854
rect 82486 12790 82492 12822
rect 67184 11158 67190 11222
rect 67254 11158 67260 11222
rect 67184 11152 67260 11158
rect 38488 11086 38564 11092
rect 38488 11022 38494 11086
rect 38558 11022 38564 11086
rect 27885 10678 27951 10679
rect 27885 10646 27886 10678
rect 14280 9254 14286 9318
rect 14350 9254 14356 9318
rect 14280 9248 14356 9254
rect 27880 10614 27886 10646
rect 27950 10646 27951 10678
rect 28560 10678 28636 10684
rect 27950 10614 27956 10646
rect 14008 7758 14014 7822
rect 14078 7758 14084 7822
rect 14008 7752 14084 7758
rect 14144 9182 14220 9188
rect 14144 9118 14150 9182
rect 14214 9118 14220 9182
rect 952 6942 1230 7006
rect 1294 6942 1300 7006
rect 2589 7006 2655 7007
rect 2589 6974 2590 7006
rect 952 5374 1300 6942
rect 2584 6942 2590 6974
rect 2654 6974 2655 7006
rect 2654 6942 2660 6974
rect 2584 6462 2660 6942
rect 2584 6398 2590 6462
rect 2654 6398 2660 6462
rect 14144 6462 14220 9118
rect 27744 8910 27820 8916
rect 27744 8846 27750 8910
rect 27814 8846 27820 8910
rect 14285 7686 14351 7687
rect 14285 7654 14286 7686
rect 14144 6430 14150 6462
rect 2584 6392 2660 6398
rect 14149 6398 14150 6430
rect 14214 6430 14220 6462
rect 14280 7622 14286 7654
rect 14350 7654 14351 7686
rect 14350 7622 14356 7654
rect 14214 6398 14215 6430
rect 14149 6397 14215 6398
rect 5853 5510 5919 5511
rect 5853 5478 5854 5510
rect 952 5310 1230 5374
rect 1294 5310 1300 5374
rect 952 3742 1300 5310
rect 952 3678 1230 3742
rect 1294 3678 1300 3742
rect 952 1294 1300 3678
rect 5848 5446 5854 5478
rect 5918 5478 5919 5510
rect 5918 5446 5924 5478
rect 2181 1702 2247 1703
rect 2181 1670 2182 1702
rect 952 1230 958 1294
rect 1022 1230 1094 1294
rect 1158 1230 1230 1294
rect 1294 1230 1300 1294
rect 952 1158 1300 1230
rect 2176 1638 2182 1670
rect 2246 1670 2247 1702
rect 3949 1702 4015 1703
rect 3949 1670 3950 1702
rect 2246 1638 2252 1670
rect 2176 1294 2252 1638
rect 2176 1230 2182 1294
rect 2246 1230 2252 1294
rect 2176 1224 2252 1230
rect 3944 1638 3950 1670
rect 4014 1670 4015 1702
rect 5445 1702 5511 1703
rect 5445 1670 5446 1702
rect 4014 1638 4020 1670
rect 3944 1294 4020 1638
rect 3944 1230 3950 1294
rect 4014 1230 4020 1294
rect 3944 1224 4020 1230
rect 5440 1638 5446 1670
rect 5510 1670 5511 1702
rect 5510 1638 5516 1670
rect 5440 1294 5516 1638
rect 5440 1230 5446 1294
rect 5510 1230 5516 1294
rect 5440 1224 5516 1230
rect 952 1094 958 1158
rect 1022 1094 1094 1158
rect 1158 1094 1230 1158
rect 1294 1094 1300 1158
rect 952 1022 1300 1094
rect 952 958 958 1022
rect 1022 958 1094 1022
rect 1158 958 1230 1022
rect 1294 958 1300 1022
rect 952 952 1300 958
rect 272 550 278 614
rect 342 550 414 614
rect 478 550 550 614
rect 614 550 620 614
rect 272 478 620 550
rect 272 414 278 478
rect 342 414 414 478
rect 478 414 550 478
rect 614 414 620 478
rect 272 342 620 414
rect 272 278 278 342
rect 342 278 414 342
rect 478 278 550 342
rect 614 278 620 342
rect 272 272 620 278
rect 5848 0 5924 5446
rect 14280 5102 14356 7622
rect 27744 7142 27820 8846
rect 27744 7110 27750 7142
rect 27749 7078 27750 7110
rect 27814 7110 27820 7142
rect 27814 7078 27815 7110
rect 27749 7077 27815 7078
rect 15917 6326 15983 6327
rect 15917 6294 15918 6326
rect 14280 5038 14286 5102
rect 14350 5038 14356 5102
rect 14280 5032 14356 5038
rect 15912 6262 15918 6294
rect 15982 6294 15983 6326
rect 15982 6262 15988 6294
rect 15912 3878 15988 6262
rect 16053 4830 16119 4831
rect 16053 4798 16054 4830
rect 15912 3814 15918 3878
rect 15982 3814 15988 3878
rect 15912 3808 15988 3814
rect 16048 4766 16054 4798
rect 16118 4798 16119 4830
rect 16118 4766 16124 4798
rect 15509 2926 15575 2927
rect 15509 2894 15510 2926
rect 15504 2862 15510 2894
rect 15574 2894 15575 2926
rect 15574 2862 15580 2894
rect 7213 1702 7279 1703
rect 7213 1670 7214 1702
rect 7208 1638 7214 1670
rect 7278 1670 7279 1702
rect 8981 1702 9047 1703
rect 8981 1670 8982 1702
rect 7278 1638 7284 1670
rect 7208 1294 7284 1638
rect 7208 1230 7214 1294
rect 7278 1230 7284 1294
rect 7208 1224 7284 1230
rect 8976 1638 8982 1670
rect 9046 1670 9047 1702
rect 10477 1702 10543 1703
rect 10477 1670 10478 1702
rect 9046 1638 9052 1670
rect 8976 1294 9052 1638
rect 8976 1230 8982 1294
rect 9046 1230 9052 1294
rect 8976 1224 9052 1230
rect 10472 1638 10478 1670
rect 10542 1670 10543 1702
rect 12245 1702 12311 1703
rect 12245 1670 12246 1702
rect 10542 1638 10548 1670
rect 10472 1294 10548 1638
rect 10472 1230 10478 1294
rect 10542 1230 10548 1294
rect 10472 1224 10548 1230
rect 12240 1638 12246 1670
rect 12310 1670 12311 1702
rect 14013 1702 14079 1703
rect 14013 1670 14014 1702
rect 12310 1638 12316 1670
rect 12240 1294 12316 1638
rect 12240 1230 12246 1294
rect 12310 1230 12316 1294
rect 12240 1224 12316 1230
rect 14008 1638 14014 1670
rect 14078 1670 14079 1702
rect 14078 1638 14084 1670
rect 14008 1294 14084 1638
rect 14008 1230 14014 1294
rect 14078 1230 14084 1294
rect 14008 1224 14084 1230
rect 15504 0 15580 2862
rect 16048 2518 16124 4766
rect 17277 3742 17343 3743
rect 17277 3710 17278 3742
rect 17272 3678 17278 3710
rect 17342 3710 17343 3742
rect 17342 3678 17348 3710
rect 16733 2926 16799 2927
rect 16733 2894 16734 2926
rect 16048 2454 16054 2518
rect 16118 2454 16124 2518
rect 16048 2448 16124 2454
rect 16728 2862 16734 2894
rect 16798 2894 16799 2926
rect 16798 2862 16804 2894
rect 15781 1702 15847 1703
rect 15781 1670 15782 1702
rect 15776 1638 15782 1670
rect 15846 1670 15847 1702
rect 15846 1638 15852 1670
rect 15776 1294 15852 1638
rect 15776 1230 15782 1294
rect 15846 1230 15852 1294
rect 15776 1224 15852 1230
rect 16728 0 16804 2862
rect 17272 1838 17348 3678
rect 17821 2926 17887 2927
rect 17821 2894 17822 2926
rect 17272 1774 17278 1838
rect 17342 1774 17348 1838
rect 17272 1768 17348 1774
rect 17816 2862 17822 2894
rect 17886 2894 17887 2926
rect 19181 2926 19247 2927
rect 19181 2894 19182 2926
rect 17886 2862 17892 2894
rect 17413 1702 17479 1703
rect 17413 1670 17414 1702
rect 17408 1638 17414 1670
rect 17478 1670 17479 1702
rect 17478 1638 17484 1670
rect 17408 1294 17484 1638
rect 17408 1230 17414 1294
rect 17478 1230 17484 1294
rect 17408 1224 17484 1230
rect 17816 0 17892 2862
rect 19176 2862 19182 2894
rect 19246 2894 19247 2926
rect 20133 2926 20199 2927
rect 20133 2894 20134 2926
rect 19246 2862 19252 2894
rect 18909 1702 18975 1703
rect 18909 1670 18910 1702
rect 18904 1638 18910 1670
rect 18974 1670 18975 1702
rect 18974 1638 18980 1670
rect 18904 1294 18980 1638
rect 18904 1230 18910 1294
rect 18974 1230 18980 1294
rect 18904 1224 18980 1230
rect 19176 0 19252 2862
rect 20128 2862 20134 2894
rect 20198 2894 20199 2926
rect 21357 2926 21423 2927
rect 21357 2894 21358 2926
rect 20198 2862 20204 2894
rect 20128 0 20204 2862
rect 21352 2862 21358 2894
rect 21422 2894 21423 2926
rect 22581 2926 22647 2927
rect 22581 2894 22582 2926
rect 21422 2862 21428 2894
rect 20677 1702 20743 1703
rect 20677 1670 20678 1702
rect 20672 1638 20678 1670
rect 20742 1670 20743 1702
rect 20742 1638 20748 1670
rect 20672 1294 20748 1638
rect 20672 1230 20678 1294
rect 20742 1230 20748 1294
rect 20672 1224 20748 1230
rect 21352 0 21428 2862
rect 22576 2862 22582 2894
rect 22646 2894 22647 2926
rect 23669 2926 23735 2927
rect 23669 2894 23670 2926
rect 22646 2862 22652 2894
rect 22445 1702 22511 1703
rect 22445 1670 22446 1702
rect 22440 1638 22446 1670
rect 22510 1670 22511 1702
rect 22510 1638 22516 1670
rect 22440 1294 22516 1638
rect 22440 1230 22446 1294
rect 22510 1230 22516 1294
rect 22440 1224 22516 1230
rect 22576 0 22652 2862
rect 23664 2862 23670 2894
rect 23734 2894 23735 2926
rect 25029 2926 25095 2927
rect 25029 2894 25030 2926
rect 23734 2862 23740 2894
rect 23664 0 23740 2862
rect 25024 2862 25030 2894
rect 25094 2894 25095 2926
rect 26117 2926 26183 2927
rect 26117 2894 26118 2926
rect 25094 2862 25100 2894
rect 23941 1702 24007 1703
rect 23941 1670 23942 1702
rect 23936 1638 23942 1670
rect 24006 1670 24007 1702
rect 24006 1638 24012 1670
rect 23936 1294 24012 1638
rect 23936 1230 23942 1294
rect 24006 1230 24012 1294
rect 23936 1224 24012 1230
rect 25024 0 25100 2862
rect 26112 2862 26118 2894
rect 26182 2894 26183 2926
rect 27205 2926 27271 2927
rect 27205 2894 27206 2926
rect 26182 2862 26188 2894
rect 25709 1702 25775 1703
rect 25709 1670 25710 1702
rect 25704 1638 25710 1670
rect 25774 1670 25775 1702
rect 25774 1638 25780 1670
rect 25704 1294 25780 1638
rect 25704 1230 25710 1294
rect 25774 1230 25780 1294
rect 25704 1224 25780 1230
rect 26112 0 26188 2862
rect 27200 2862 27206 2894
rect 27270 2894 27271 2926
rect 27270 2862 27276 2894
rect 26661 2382 26727 2383
rect 26661 2350 26662 2382
rect 26656 2318 26662 2350
rect 26726 2350 26727 2382
rect 26726 2318 26732 2350
rect 26656 614 26732 2318
rect 26656 550 26662 614
rect 26726 550 26732 614
rect 26656 544 26732 550
rect 27200 0 27276 2862
rect 27477 1702 27543 1703
rect 27477 1670 27478 1702
rect 27472 1638 27478 1670
rect 27542 1670 27543 1702
rect 27542 1638 27548 1670
rect 27472 1294 27548 1638
rect 27472 1230 27478 1294
rect 27542 1230 27548 1294
rect 27472 1224 27548 1230
rect 27880 0 27956 10614
rect 28560 10614 28566 10678
rect 28630 10614 28636 10678
rect 29245 10678 29311 10679
rect 29245 10646 29246 10678
rect 28560 10134 28636 10614
rect 28560 10102 28566 10134
rect 28565 10070 28566 10102
rect 28630 10102 28636 10134
rect 29240 10614 29246 10646
rect 29310 10646 29311 10678
rect 29784 10678 29860 10684
rect 29310 10614 29316 10646
rect 28630 10070 28631 10102
rect 28565 10069 28631 10070
rect 28429 9862 28495 9863
rect 28429 9830 28430 9862
rect 28424 9798 28430 9830
rect 28494 9830 28495 9862
rect 28494 9798 28500 9830
rect 28293 9454 28359 9455
rect 28293 9422 28294 9454
rect 28288 9390 28294 9422
rect 28358 9422 28359 9454
rect 28358 9390 28364 9422
rect 28152 8638 28228 8644
rect 28152 8574 28158 8638
rect 28222 8574 28228 8638
rect 28152 8230 28228 8574
rect 28288 8638 28364 9390
rect 28424 9318 28500 9798
rect 28424 9254 28430 9318
rect 28494 9254 28500 9318
rect 28424 9248 28500 9254
rect 28288 8574 28294 8638
rect 28358 8574 28364 8638
rect 28288 8568 28364 8574
rect 28152 8198 28158 8230
rect 28157 8166 28158 8198
rect 28222 8198 28228 8230
rect 28222 8166 28223 8198
rect 28157 8165 28223 8166
rect 28293 2926 28359 2927
rect 28293 2894 28294 2926
rect 28288 2862 28294 2894
rect 28358 2894 28359 2926
rect 28358 2862 28364 2894
rect 28288 0 28364 2862
rect 28973 1702 29039 1703
rect 28973 1670 28974 1702
rect 28968 1638 28974 1670
rect 29038 1670 29039 1702
rect 29038 1638 29044 1670
rect 28968 1294 29044 1638
rect 28968 1230 28974 1294
rect 29038 1230 29044 1294
rect 28968 1224 29044 1230
rect 29240 0 29316 10614
rect 29784 10614 29790 10678
rect 29854 10614 29860 10678
rect 30333 10678 30399 10679
rect 30333 10646 30334 10678
rect 29784 10134 29860 10614
rect 29784 10102 29790 10134
rect 29789 10070 29790 10102
rect 29854 10102 29860 10134
rect 30328 10614 30334 10646
rect 30398 10646 30399 10678
rect 30872 10678 30948 10684
rect 30398 10614 30404 10646
rect 29854 10070 29855 10102
rect 29789 10069 29855 10070
rect 29789 9862 29855 9863
rect 29789 9830 29790 9862
rect 29784 9798 29790 9830
rect 29854 9830 29855 9862
rect 29854 9798 29860 9830
rect 29653 9454 29719 9455
rect 29653 9422 29654 9454
rect 29648 9390 29654 9422
rect 29718 9422 29719 9454
rect 29718 9390 29724 9422
rect 29648 8638 29724 9390
rect 29784 9318 29860 9798
rect 29784 9254 29790 9318
rect 29854 9254 29860 9318
rect 29784 9248 29860 9254
rect 29648 8574 29654 8638
rect 29718 8574 29724 8638
rect 29648 8568 29724 8574
rect 29653 2926 29719 2927
rect 29653 2894 29654 2926
rect 29648 2862 29654 2894
rect 29718 2894 29719 2926
rect 29718 2862 29724 2894
rect 29648 0 29724 2862
rect 30328 0 30404 10614
rect 30872 10614 30878 10678
rect 30942 10614 30948 10678
rect 31965 10678 32031 10679
rect 31965 10646 31966 10678
rect 30872 10134 30948 10614
rect 30872 10102 30878 10134
rect 30877 10070 30878 10102
rect 30942 10102 30948 10134
rect 31960 10614 31966 10646
rect 32030 10646 32031 10678
rect 32232 10678 32308 10684
rect 32030 10614 32036 10646
rect 30942 10070 30943 10102
rect 30877 10069 30943 10070
rect 30877 9862 30943 9863
rect 30877 9830 30878 9862
rect 30872 9798 30878 9830
rect 30942 9830 30943 9862
rect 30942 9798 30948 9830
rect 30741 9454 30807 9455
rect 30741 9422 30742 9454
rect 30736 9390 30742 9422
rect 30806 9422 30807 9454
rect 30806 9390 30812 9422
rect 30736 8638 30812 9390
rect 30872 9318 30948 9798
rect 30872 9254 30878 9318
rect 30942 9254 30948 9318
rect 30872 9248 30948 9254
rect 30736 8574 30742 8638
rect 30806 8574 30812 8638
rect 30736 8568 30812 8574
rect 30741 2926 30807 2927
rect 30741 2894 30742 2926
rect 30736 2862 30742 2894
rect 30806 2894 30807 2926
rect 31829 2926 31895 2927
rect 31829 2894 31830 2926
rect 30806 2862 30812 2894
rect 30605 1702 30671 1703
rect 30605 1670 30606 1702
rect 30600 1638 30606 1670
rect 30670 1670 30671 1702
rect 30670 1638 30676 1670
rect 30600 1294 30676 1638
rect 30600 1230 30606 1294
rect 30670 1230 30676 1294
rect 30600 1224 30676 1230
rect 30736 0 30812 2862
rect 31824 2862 31830 2894
rect 31894 2894 31895 2926
rect 31894 2862 31900 2894
rect 31824 0 31900 2862
rect 31960 0 32036 10614
rect 32232 10614 32238 10678
rect 32302 10614 32308 10678
rect 33189 10678 33255 10679
rect 33189 10646 33190 10678
rect 32232 10134 32308 10614
rect 32232 10102 32238 10134
rect 32237 10070 32238 10102
rect 32302 10102 32308 10134
rect 33184 10614 33190 10646
rect 33254 10646 33255 10678
rect 33456 10678 33532 10684
rect 33254 10614 33260 10646
rect 32302 10070 32303 10102
rect 32237 10069 32303 10070
rect 32373 9862 32439 9863
rect 32373 9830 32374 9862
rect 32368 9798 32374 9830
rect 32438 9830 32439 9862
rect 32438 9798 32444 9830
rect 32237 9454 32303 9455
rect 32237 9422 32238 9454
rect 32232 9390 32238 9422
rect 32302 9422 32303 9454
rect 32302 9390 32308 9422
rect 32232 8638 32308 9390
rect 32368 9318 32444 9798
rect 32368 9254 32374 9318
rect 32438 9254 32444 9318
rect 32368 9248 32444 9254
rect 32232 8574 32238 8638
rect 32302 8574 32308 8638
rect 32232 8568 32308 8574
rect 33053 2926 33119 2927
rect 33053 2894 33054 2926
rect 33048 2862 33054 2894
rect 33118 2894 33119 2926
rect 33118 2862 33124 2894
rect 32373 1702 32439 1703
rect 32373 1670 32374 1702
rect 32368 1638 32374 1670
rect 32438 1670 32439 1702
rect 32438 1638 32444 1670
rect 32368 1294 32444 1638
rect 32368 1230 32374 1294
rect 32438 1230 32444 1294
rect 32368 1224 32444 1230
rect 33048 0 33124 2862
rect 33184 0 33260 10614
rect 33456 10614 33462 10678
rect 33526 10614 33532 10678
rect 34413 10678 34479 10679
rect 34413 10646 34414 10678
rect 33456 10134 33532 10614
rect 33456 10102 33462 10134
rect 33461 10070 33462 10102
rect 33526 10102 33532 10134
rect 34408 10614 34414 10646
rect 34478 10646 34479 10678
rect 34816 10678 34892 10684
rect 34478 10614 34484 10646
rect 33526 10070 33527 10102
rect 33461 10069 33527 10070
rect 33597 9862 33663 9863
rect 33597 9830 33598 9862
rect 33592 9798 33598 9830
rect 33662 9830 33663 9862
rect 33662 9798 33668 9830
rect 33461 9454 33527 9455
rect 33461 9422 33462 9454
rect 33456 9390 33462 9422
rect 33526 9422 33527 9454
rect 33526 9390 33532 9422
rect 33456 8638 33532 9390
rect 33592 9318 33668 9798
rect 33592 9254 33598 9318
rect 33662 9254 33668 9318
rect 33592 9248 33668 9254
rect 33456 8574 33462 8638
rect 33526 8574 33532 8638
rect 33456 8568 33532 8574
rect 34141 2926 34207 2927
rect 34141 2894 34142 2926
rect 34136 2862 34142 2894
rect 34206 2894 34207 2926
rect 34206 2862 34212 2894
rect 34005 1702 34071 1703
rect 34005 1670 34006 1702
rect 34000 1638 34006 1670
rect 34070 1670 34071 1702
rect 34070 1638 34076 1670
rect 34000 1294 34076 1638
rect 34000 1230 34006 1294
rect 34070 1230 34076 1294
rect 34000 1224 34076 1230
rect 34136 0 34212 2862
rect 34408 0 34484 10614
rect 34816 10614 34822 10678
rect 34886 10614 34892 10678
rect 35637 10678 35703 10679
rect 35637 10646 35638 10678
rect 34816 10134 34892 10614
rect 34816 10102 34822 10134
rect 34821 10070 34822 10102
rect 34886 10102 34892 10134
rect 35632 10614 35638 10646
rect 35702 10646 35703 10678
rect 36040 10678 36116 10684
rect 35702 10614 35708 10646
rect 34886 10070 34887 10102
rect 34821 10069 34887 10070
rect 34821 9862 34887 9863
rect 34821 9830 34822 9862
rect 34816 9798 34822 9830
rect 34886 9830 34887 9862
rect 34886 9798 34892 9830
rect 34685 9454 34751 9455
rect 34685 9422 34686 9454
rect 34680 9390 34686 9422
rect 34750 9422 34751 9454
rect 34750 9390 34756 9422
rect 34680 8638 34756 9390
rect 34816 9318 34892 9798
rect 34816 9254 34822 9318
rect 34886 9254 34892 9318
rect 34816 9248 34892 9254
rect 34680 8574 34686 8638
rect 34750 8574 34756 8638
rect 34680 8568 34756 8574
rect 35501 2926 35567 2927
rect 35501 2894 35502 2926
rect 35496 2862 35502 2894
rect 35566 2894 35567 2926
rect 35566 2862 35572 2894
rect 35496 0 35572 2862
rect 35632 0 35708 10614
rect 36040 10614 36046 10678
rect 36110 10614 36116 10678
rect 36861 10678 36927 10679
rect 36861 10646 36862 10678
rect 36040 10134 36116 10614
rect 36040 10102 36046 10134
rect 36045 10070 36046 10102
rect 36110 10102 36116 10134
rect 36856 10614 36862 10646
rect 36926 10646 36927 10678
rect 37128 10678 37204 10684
rect 36926 10614 36932 10646
rect 36110 10070 36111 10102
rect 36045 10069 36111 10070
rect 36045 9862 36111 9863
rect 36045 9830 36046 9862
rect 36040 9798 36046 9830
rect 36110 9830 36111 9862
rect 36110 9798 36116 9830
rect 35909 9454 35975 9455
rect 35909 9422 35910 9454
rect 35904 9390 35910 9422
rect 35974 9422 35975 9454
rect 35974 9390 35980 9422
rect 35904 8638 35980 9390
rect 36040 9318 36116 9798
rect 36040 9254 36046 9318
rect 36110 9254 36116 9318
rect 36040 9248 36116 9254
rect 35904 8574 35910 8638
rect 35974 8574 35980 8638
rect 35904 8568 35980 8574
rect 36589 2926 36655 2927
rect 36589 2894 36590 2926
rect 36584 2862 36590 2894
rect 36654 2894 36655 2926
rect 36654 2862 36660 2894
rect 35773 1702 35839 1703
rect 35773 1670 35774 1702
rect 35768 1638 35774 1670
rect 35838 1670 35839 1702
rect 35838 1638 35844 1670
rect 35768 1294 35844 1638
rect 35768 1230 35774 1294
rect 35838 1230 35844 1294
rect 35768 1224 35844 1230
rect 36584 0 36660 2862
rect 36856 0 36932 10614
rect 37128 10614 37134 10678
rect 37198 10614 37204 10678
rect 37813 10678 37879 10679
rect 37813 10646 37814 10678
rect 37128 10134 37204 10614
rect 37128 10102 37134 10134
rect 37133 10070 37134 10102
rect 37198 10102 37204 10134
rect 37808 10614 37814 10646
rect 37878 10646 37879 10678
rect 37878 10614 37884 10646
rect 37198 10070 37199 10102
rect 37133 10069 37199 10070
rect 37269 9862 37335 9863
rect 37269 9830 37270 9862
rect 37264 9798 37270 9830
rect 37334 9830 37335 9862
rect 37334 9798 37340 9830
rect 37133 9454 37199 9455
rect 37133 9422 37134 9454
rect 37128 9390 37134 9422
rect 37198 9422 37199 9454
rect 37198 9390 37204 9422
rect 37128 8638 37204 9390
rect 37264 9318 37340 9798
rect 37264 9254 37270 9318
rect 37334 9254 37340 9318
rect 37264 9248 37340 9254
rect 37128 8574 37134 8638
rect 37198 8574 37204 8638
rect 37128 8568 37204 8574
rect 37677 2926 37743 2927
rect 37677 2894 37678 2926
rect 37672 2862 37678 2894
rect 37742 2894 37743 2926
rect 37742 2862 37748 2894
rect 37405 1702 37471 1703
rect 37405 1670 37406 1702
rect 37400 1638 37406 1670
rect 37470 1670 37471 1702
rect 37470 1638 37476 1670
rect 37400 1294 37476 1638
rect 37400 1230 37406 1294
rect 37470 1230 37476 1294
rect 37400 1224 37476 1230
rect 37672 0 37748 2862
rect 37808 0 37884 10614
rect 38221 9862 38287 9863
rect 38221 9830 38222 9862
rect 38216 9798 38222 9830
rect 38286 9830 38287 9862
rect 38286 9798 38292 9830
rect 38216 9318 38292 9798
rect 38488 9590 38564 11022
rect 64600 11016 64812 11092
rect 64736 10814 64812 11016
rect 64736 10782 64742 10814
rect 64741 10750 64742 10782
rect 64806 10782 64812 10814
rect 64806 10750 64807 10782
rect 64741 10749 64807 10750
rect 38624 10678 38700 10684
rect 38624 10614 38630 10678
rect 38694 10614 38700 10678
rect 39309 10678 39375 10679
rect 39309 10646 39310 10678
rect 38624 10134 38700 10614
rect 38624 10102 38630 10134
rect 38629 10070 38630 10102
rect 38694 10102 38700 10134
rect 39304 10614 39310 10646
rect 39374 10646 39375 10678
rect 39712 10678 39788 10684
rect 39374 10614 39380 10646
rect 38694 10070 38695 10102
rect 38629 10069 38695 10070
rect 38488 9558 38494 9590
rect 38493 9526 38494 9558
rect 38558 9558 38564 9590
rect 38558 9526 38559 9558
rect 38493 9525 38559 9526
rect 38357 9454 38423 9455
rect 38357 9422 38358 9454
rect 38216 9254 38222 9318
rect 38286 9254 38292 9318
rect 38216 9248 38292 9254
rect 38352 9390 38358 9422
rect 38422 9422 38423 9454
rect 38422 9390 38428 9422
rect 38352 8638 38428 9390
rect 38352 8574 38358 8638
rect 38422 8574 38428 8638
rect 38352 8568 38428 8574
rect 38901 2926 38967 2927
rect 38901 2894 38902 2926
rect 38896 2862 38902 2894
rect 38966 2894 38967 2926
rect 38966 2862 38972 2894
rect 38896 0 38972 2862
rect 39173 1702 39239 1703
rect 39173 1670 39174 1702
rect 39168 1638 39174 1670
rect 39238 1670 39239 1702
rect 39238 1638 39244 1670
rect 39168 1294 39244 1638
rect 39168 1230 39174 1294
rect 39238 1230 39244 1294
rect 39168 1224 39244 1230
rect 39304 0 39380 10614
rect 39712 10614 39718 10678
rect 39782 10614 39788 10678
rect 40669 10678 40735 10679
rect 40669 10646 40670 10678
rect 39712 10134 39788 10614
rect 39712 10102 39718 10134
rect 39717 10070 39718 10102
rect 39782 10102 39788 10134
rect 40664 10614 40670 10646
rect 40734 10646 40735 10678
rect 40936 10678 41012 10684
rect 40734 10614 40740 10646
rect 39782 10070 39783 10102
rect 39717 10069 39783 10070
rect 39717 9862 39783 9863
rect 39717 9830 39718 9862
rect 39712 9798 39718 9830
rect 39782 9830 39783 9862
rect 39782 9798 39788 9830
rect 39581 9454 39647 9455
rect 39581 9422 39582 9454
rect 39576 9390 39582 9422
rect 39646 9422 39647 9454
rect 39646 9390 39652 9422
rect 39576 8638 39652 9390
rect 39712 9318 39788 9798
rect 39712 9254 39718 9318
rect 39782 9254 39788 9318
rect 39712 9248 39788 9254
rect 39576 8574 39582 8638
rect 39646 8574 39652 8638
rect 39576 8568 39652 8574
rect 40261 2926 40327 2927
rect 40261 2894 40262 2926
rect 40256 2862 40262 2894
rect 40326 2894 40327 2926
rect 40326 2862 40332 2894
rect 40256 0 40332 2862
rect 40533 1702 40599 1703
rect 40533 1670 40534 1702
rect 40528 1638 40534 1670
rect 40598 1670 40599 1702
rect 40598 1638 40604 1670
rect 40528 1294 40604 1638
rect 40528 1230 40534 1294
rect 40598 1230 40604 1294
rect 40528 1224 40604 1230
rect 40664 0 40740 10614
rect 40936 10614 40942 10678
rect 41006 10614 41012 10678
rect 41757 10678 41823 10679
rect 41757 10646 41758 10678
rect 40936 10134 41012 10614
rect 40936 10102 40942 10134
rect 40941 10070 40942 10102
rect 41006 10102 41012 10134
rect 41752 10614 41758 10646
rect 41822 10646 41823 10678
rect 41893 10678 41959 10679
rect 41893 10646 41894 10678
rect 41822 10614 41828 10646
rect 41752 10134 41828 10614
rect 41006 10070 41007 10102
rect 40941 10069 41007 10070
rect 41752 10070 41758 10134
rect 41822 10070 41828 10134
rect 41752 10064 41828 10070
rect 41888 10614 41894 10646
rect 41958 10646 41959 10678
rect 42296 10678 42372 10684
rect 41958 10614 41964 10646
rect 41077 9862 41143 9863
rect 41077 9830 41078 9862
rect 41072 9798 41078 9830
rect 41142 9830 41143 9862
rect 41142 9798 41148 9830
rect 40941 9454 41007 9455
rect 40941 9422 40942 9454
rect 40936 9390 40942 9422
rect 41006 9422 41007 9454
rect 41006 9390 41012 9422
rect 40936 8638 41012 9390
rect 41072 9318 41148 9798
rect 41072 9254 41078 9318
rect 41142 9254 41148 9318
rect 41072 9248 41148 9254
rect 40936 8574 40942 8638
rect 41006 8574 41012 8638
rect 40936 8568 41012 8574
rect 41349 2926 41415 2927
rect 41349 2894 41350 2926
rect 41344 2862 41350 2894
rect 41414 2894 41415 2926
rect 41414 2862 41420 2894
rect 41344 0 41420 2862
rect 41888 0 41964 10614
rect 42296 10614 42302 10678
rect 42366 10614 42372 10678
rect 43117 10678 43183 10679
rect 43117 10646 43118 10678
rect 42296 10134 42372 10614
rect 42296 10102 42302 10134
rect 42301 10070 42302 10102
rect 42366 10102 42372 10134
rect 43112 10614 43118 10646
rect 43182 10646 43183 10678
rect 43520 10678 43596 10684
rect 43182 10614 43188 10646
rect 42366 10070 42367 10102
rect 42301 10069 42367 10070
rect 42301 9862 42367 9863
rect 42301 9830 42302 9862
rect 42296 9798 42302 9830
rect 42366 9830 42367 9862
rect 42366 9798 42372 9830
rect 42165 9454 42231 9455
rect 42165 9422 42166 9454
rect 42160 9390 42166 9422
rect 42230 9422 42231 9454
rect 42230 9390 42236 9422
rect 42160 8638 42236 9390
rect 42296 9318 42372 9798
rect 42296 9254 42302 9318
rect 42366 9254 42372 9318
rect 42296 9248 42372 9254
rect 42160 8574 42166 8638
rect 42230 8574 42236 8638
rect 42160 8568 42236 8574
rect 42437 2926 42503 2927
rect 42437 2894 42438 2926
rect 42432 2862 42438 2894
rect 42502 2894 42503 2926
rect 42502 2862 42508 2894
rect 42301 1702 42367 1703
rect 42301 1670 42302 1702
rect 42296 1638 42302 1670
rect 42366 1670 42367 1702
rect 42366 1638 42372 1670
rect 42296 1294 42372 1638
rect 42296 1230 42302 1294
rect 42366 1230 42372 1294
rect 42296 1224 42372 1230
rect 42432 0 42508 2862
rect 43112 0 43188 10614
rect 43520 10614 43526 10678
rect 43590 10614 43596 10678
rect 44341 10678 44407 10679
rect 44341 10646 44342 10678
rect 43520 10134 43596 10614
rect 43520 10102 43526 10134
rect 43525 10070 43526 10102
rect 43590 10102 43596 10134
rect 44336 10614 44342 10646
rect 44406 10646 44407 10678
rect 44744 10678 44820 10684
rect 44406 10614 44412 10646
rect 43590 10070 43591 10102
rect 43525 10069 43591 10070
rect 43520 9862 43596 9868
rect 43520 9798 43526 9862
rect 43590 9798 43596 9862
rect 43389 9454 43455 9455
rect 43389 9422 43390 9454
rect 43384 9390 43390 9422
rect 43454 9422 43455 9454
rect 43454 9390 43460 9422
rect 43384 8638 43460 9390
rect 43520 9046 43596 9798
rect 43520 9014 43526 9046
rect 43525 8982 43526 9014
rect 43590 9014 43596 9046
rect 43590 8982 43591 9014
rect 43525 8981 43591 8982
rect 43384 8574 43390 8638
rect 43454 8574 43460 8638
rect 43384 8568 43460 8574
rect 43525 2926 43591 2927
rect 43525 2894 43526 2926
rect 43520 2862 43526 2894
rect 43590 2894 43591 2926
rect 43590 2862 43596 2894
rect 43520 0 43596 2862
rect 44205 1702 44271 1703
rect 44205 1670 44206 1702
rect 44200 1638 44206 1670
rect 44270 1670 44271 1702
rect 44270 1638 44276 1670
rect 44200 1294 44276 1638
rect 44200 1230 44206 1294
rect 44270 1230 44276 1294
rect 44200 1224 44276 1230
rect 44336 0 44412 10614
rect 44744 10614 44750 10678
rect 44814 10614 44820 10678
rect 45293 10678 45359 10679
rect 45293 10646 45294 10678
rect 44744 10134 44820 10614
rect 44744 10102 44750 10134
rect 44749 10070 44750 10102
rect 44814 10102 44820 10134
rect 45288 10614 45294 10646
rect 45358 10646 45359 10678
rect 45565 10678 45631 10679
rect 45565 10646 45566 10678
rect 45358 10614 45364 10646
rect 45288 10134 45364 10614
rect 44814 10070 44815 10102
rect 44749 10069 44815 10070
rect 45288 10070 45294 10134
rect 45358 10070 45364 10134
rect 45288 10064 45364 10070
rect 45560 10614 45566 10646
rect 45630 10646 45631 10678
rect 45968 10678 46044 10684
rect 45630 10614 45636 10646
rect 44749 9862 44815 9863
rect 44749 9830 44750 9862
rect 44744 9798 44750 9830
rect 44814 9830 44815 9862
rect 44814 9798 44820 9830
rect 44613 9454 44679 9455
rect 44613 9422 44614 9454
rect 44608 9390 44614 9422
rect 44678 9422 44679 9454
rect 44678 9390 44684 9422
rect 44608 8638 44684 9390
rect 44744 9318 44820 9798
rect 44744 9254 44750 9318
rect 44814 9254 44820 9318
rect 44744 9248 44820 9254
rect 44608 8574 44614 8638
rect 44678 8574 44684 8638
rect 44608 8568 44684 8574
rect 44885 2926 44951 2927
rect 44885 2894 44886 2926
rect 44880 2862 44886 2894
rect 44950 2894 44951 2926
rect 44950 2862 44956 2894
rect 44880 0 44956 2862
rect 45560 0 45636 10614
rect 45968 10614 45974 10678
rect 46038 10614 46044 10678
rect 46653 10678 46719 10679
rect 46653 10646 46654 10678
rect 45968 10134 46044 10614
rect 45968 10102 45974 10134
rect 45973 10070 45974 10102
rect 46038 10102 46044 10134
rect 46648 10614 46654 10646
rect 46718 10646 46719 10678
rect 47192 10678 47268 10684
rect 46718 10614 46724 10646
rect 46038 10070 46039 10102
rect 45973 10069 46039 10070
rect 45973 9862 46039 9863
rect 45973 9830 45974 9862
rect 45968 9798 45974 9830
rect 46038 9830 46039 9862
rect 46038 9798 46044 9830
rect 45837 9454 45903 9455
rect 45837 9422 45838 9454
rect 45832 9390 45838 9422
rect 45902 9422 45903 9454
rect 45902 9390 45908 9422
rect 45832 8638 45908 9390
rect 45968 9318 46044 9798
rect 45968 9254 45974 9318
rect 46038 9254 46044 9318
rect 45968 9248 46044 9254
rect 45832 8574 45838 8638
rect 45902 8574 45908 8638
rect 45832 8568 45908 8574
rect 45973 2926 46039 2927
rect 45973 2894 45974 2926
rect 45968 2862 45974 2894
rect 46038 2894 46039 2926
rect 46038 2862 46044 2894
rect 45837 1702 45903 1703
rect 45837 1670 45838 1702
rect 45832 1638 45838 1670
rect 45902 1670 45903 1702
rect 45902 1638 45908 1670
rect 45832 1294 45908 1638
rect 45832 1230 45838 1294
rect 45902 1230 45908 1294
rect 45832 1224 45908 1230
rect 45968 0 46044 2862
rect 46648 0 46724 10614
rect 47192 10614 47198 10678
rect 47262 10614 47268 10678
rect 47741 10678 47807 10679
rect 47741 10646 47742 10678
rect 47192 10134 47268 10614
rect 47192 10102 47198 10134
rect 47197 10070 47198 10102
rect 47262 10102 47268 10134
rect 47736 10614 47742 10646
rect 47806 10646 47807 10678
rect 47877 10678 47943 10679
rect 47877 10646 47878 10678
rect 47806 10614 47812 10646
rect 47736 10134 47812 10614
rect 47262 10070 47263 10102
rect 47197 10069 47263 10070
rect 47736 10070 47742 10134
rect 47806 10070 47812 10134
rect 47736 10064 47812 10070
rect 47872 10614 47878 10646
rect 47942 10646 47943 10678
rect 48416 10678 48492 10684
rect 47942 10614 47948 10646
rect 47197 9862 47263 9863
rect 47197 9830 47198 9862
rect 47192 9798 47198 9830
rect 47262 9830 47263 9862
rect 47262 9798 47268 9830
rect 47061 9454 47127 9455
rect 47061 9422 47062 9454
rect 47056 9390 47062 9422
rect 47126 9422 47127 9454
rect 47126 9390 47132 9422
rect 47056 8638 47132 9390
rect 47192 9318 47268 9798
rect 47192 9254 47198 9318
rect 47262 9254 47268 9318
rect 47192 9248 47268 9254
rect 47056 8574 47062 8638
rect 47126 8574 47132 8638
rect 47056 8568 47132 8574
rect 47061 2926 47127 2927
rect 47061 2894 47062 2926
rect 47056 2862 47062 2894
rect 47126 2894 47127 2926
rect 47126 2862 47132 2894
rect 47056 0 47132 2862
rect 47469 1702 47535 1703
rect 47469 1670 47470 1702
rect 47464 1638 47470 1670
rect 47534 1670 47535 1702
rect 47534 1638 47540 1670
rect 47464 1294 47540 1638
rect 47464 1230 47470 1294
rect 47534 1230 47540 1294
rect 47464 1224 47540 1230
rect 47872 0 47948 10614
rect 48416 10614 48422 10678
rect 48486 10614 48492 10678
rect 48965 10678 49031 10679
rect 48965 10646 48966 10678
rect 48416 10134 48492 10614
rect 48960 10614 48966 10646
rect 49030 10646 49031 10678
rect 49101 10678 49167 10679
rect 49101 10646 49102 10678
rect 49030 10614 49036 10646
rect 48960 10406 49036 10614
rect 48960 10342 48966 10406
rect 49030 10342 49036 10406
rect 48960 10336 49036 10342
rect 49096 10614 49102 10646
rect 49166 10646 49167 10678
rect 49640 10678 49716 10684
rect 49166 10614 49172 10646
rect 48416 10102 48422 10134
rect 48421 10070 48422 10102
rect 48486 10102 48492 10134
rect 48486 10070 48487 10102
rect 48421 10069 48487 10070
rect 48421 9862 48487 9863
rect 48421 9830 48422 9862
rect 48416 9798 48422 9830
rect 48486 9830 48487 9862
rect 48486 9798 48492 9830
rect 48285 9454 48351 9455
rect 48285 9422 48286 9454
rect 48280 9390 48286 9422
rect 48350 9422 48351 9454
rect 48350 9390 48356 9422
rect 48280 8638 48356 9390
rect 48416 9318 48492 9798
rect 48416 9254 48422 9318
rect 48486 9254 48492 9318
rect 48416 9248 48492 9254
rect 48280 8574 48286 8638
rect 48350 8574 48356 8638
rect 48280 8568 48356 8574
rect 48285 2926 48351 2927
rect 48285 2894 48286 2926
rect 48280 2862 48286 2894
rect 48350 2894 48351 2926
rect 48350 2862 48356 2894
rect 48280 0 48356 2862
rect 48965 1702 49031 1703
rect 48965 1670 48966 1702
rect 48960 1638 48966 1670
rect 49030 1670 49031 1702
rect 49030 1638 49036 1670
rect 48960 1294 49036 1638
rect 48960 1230 48966 1294
rect 49030 1230 49036 1294
rect 48960 1224 49036 1230
rect 49096 0 49172 10614
rect 49640 10614 49646 10678
rect 49710 10614 49716 10678
rect 49640 10406 49716 10614
rect 49640 10374 49646 10406
rect 49645 10342 49646 10374
rect 49710 10374 49716 10406
rect 49776 10678 49852 10684
rect 49776 10614 49782 10678
rect 49846 10614 49852 10678
rect 50597 10678 50663 10679
rect 50597 10646 50598 10678
rect 49710 10342 49711 10374
rect 49645 10341 49711 10342
rect 49776 10134 49852 10614
rect 49776 10102 49782 10134
rect 49781 10070 49782 10102
rect 49846 10102 49852 10134
rect 50592 10614 50598 10646
rect 50662 10646 50663 10678
rect 51000 10678 51076 10684
rect 50662 10614 50668 10646
rect 49846 10070 49847 10102
rect 49781 10069 49847 10070
rect 49781 9862 49847 9863
rect 49781 9830 49782 9862
rect 49776 9798 49782 9830
rect 49846 9830 49847 9862
rect 49846 9798 49852 9830
rect 49645 9454 49711 9455
rect 49645 9422 49646 9454
rect 49640 9390 49646 9422
rect 49710 9422 49711 9454
rect 49710 9390 49716 9422
rect 49640 8638 49716 9390
rect 49776 9318 49852 9798
rect 49776 9254 49782 9318
rect 49846 9254 49852 9318
rect 49776 9248 49852 9254
rect 49640 8574 49646 8638
rect 49710 8574 49716 8638
rect 49640 8568 49716 8574
rect 49373 2926 49439 2927
rect 49373 2894 49374 2926
rect 49368 2862 49374 2894
rect 49438 2894 49439 2926
rect 49438 2862 49444 2894
rect 49368 0 49444 2862
rect 50592 0 50668 10614
rect 51000 10614 51006 10678
rect 51070 10614 51076 10678
rect 51413 10678 51479 10679
rect 51413 10646 51414 10678
rect 51000 10134 51076 10614
rect 51000 10102 51006 10134
rect 51005 10070 51006 10102
rect 51070 10102 51076 10134
rect 51408 10614 51414 10646
rect 51478 10646 51479 10678
rect 52224 10678 52300 10684
rect 51478 10614 51484 10646
rect 51070 10070 51071 10102
rect 51005 10069 51071 10070
rect 50869 9862 50935 9863
rect 50869 9830 50870 9862
rect 50864 9798 50870 9830
rect 50934 9830 50935 9862
rect 50934 9798 50940 9830
rect 50733 9454 50799 9455
rect 50733 9422 50734 9454
rect 50728 9390 50734 9422
rect 50798 9422 50799 9454
rect 50798 9390 50804 9422
rect 50728 8638 50804 9390
rect 50864 9318 50940 9798
rect 50864 9254 50870 9318
rect 50934 9254 50940 9318
rect 50864 9248 50940 9254
rect 50728 8574 50734 8638
rect 50798 8574 50804 8638
rect 50728 8568 50804 8574
rect 50733 2926 50799 2927
rect 50733 2894 50734 2926
rect 50728 2862 50734 2894
rect 50798 2894 50799 2926
rect 50798 2862 50804 2894
rect 50728 0 50804 2862
rect 51005 1702 51071 1703
rect 51005 1670 51006 1702
rect 51000 1638 51006 1670
rect 51070 1670 51071 1702
rect 51070 1638 51076 1670
rect 51000 1294 51076 1638
rect 51000 1230 51006 1294
rect 51070 1230 51076 1294
rect 51000 1224 51076 1230
rect 51408 0 51484 10614
rect 52224 10614 52230 10678
rect 52294 10614 52300 10678
rect 53181 10678 53247 10679
rect 53181 10646 53182 10678
rect 52224 10134 52300 10614
rect 52224 10102 52230 10134
rect 52229 10070 52230 10102
rect 52294 10102 52300 10134
rect 53176 10614 53182 10646
rect 53246 10646 53247 10678
rect 53448 10678 53524 10684
rect 53246 10614 53252 10646
rect 52294 10070 52295 10102
rect 52229 10069 52295 10070
rect 52088 9862 52164 9868
rect 52088 9798 52094 9862
rect 52158 9798 52164 9862
rect 51957 9454 52023 9455
rect 51957 9422 51958 9454
rect 51952 9390 51958 9422
rect 52022 9422 52023 9454
rect 52022 9390 52028 9422
rect 51952 8638 52028 9390
rect 52088 9046 52164 9798
rect 52088 9014 52094 9046
rect 52093 8982 52094 9014
rect 52158 9014 52164 9046
rect 52158 8982 52159 9014
rect 52093 8981 52159 8982
rect 51952 8574 51958 8638
rect 52022 8574 52028 8638
rect 51952 8568 52028 8574
rect 51821 2926 51887 2927
rect 51821 2894 51822 2926
rect 51816 2862 51822 2894
rect 51886 2894 51887 2926
rect 52909 2926 52975 2927
rect 52909 2894 52910 2926
rect 51886 2862 51892 2894
rect 51816 0 51892 2862
rect 52904 2862 52910 2894
rect 52974 2894 52975 2926
rect 52974 2862 52980 2894
rect 52637 1702 52703 1703
rect 52637 1670 52638 1702
rect 52632 1638 52638 1670
rect 52702 1670 52703 1702
rect 52702 1638 52708 1670
rect 52632 1294 52708 1638
rect 52632 1230 52638 1294
rect 52702 1230 52708 1294
rect 52632 1224 52708 1230
rect 52904 0 52980 2862
rect 53176 0 53252 10614
rect 53448 10614 53454 10678
rect 53518 10614 53524 10678
rect 54405 10678 54471 10679
rect 54405 10646 54406 10678
rect 53448 10134 53524 10614
rect 53448 10102 53454 10134
rect 53453 10070 53454 10102
rect 53518 10102 53524 10134
rect 54400 10614 54406 10646
rect 54470 10646 54471 10678
rect 54672 10678 54748 10684
rect 54470 10614 54476 10646
rect 53518 10070 53519 10102
rect 53453 10069 53519 10070
rect 53589 9862 53655 9863
rect 53589 9830 53590 9862
rect 53584 9798 53590 9830
rect 53654 9830 53655 9862
rect 53654 9798 53660 9830
rect 53453 9454 53519 9455
rect 53453 9422 53454 9454
rect 53448 9390 53454 9422
rect 53518 9422 53519 9454
rect 53518 9390 53524 9422
rect 53448 8638 53524 9390
rect 53584 9318 53660 9798
rect 53584 9254 53590 9318
rect 53654 9254 53660 9318
rect 53584 9248 53660 9254
rect 53448 8574 53454 8638
rect 53518 8574 53524 8638
rect 53448 8568 53524 8574
rect 53997 2926 54063 2927
rect 53997 2894 53998 2926
rect 53992 2862 53998 2894
rect 54062 2894 54063 2926
rect 54062 2862 54068 2894
rect 53992 0 54068 2862
rect 54269 1702 54335 1703
rect 54269 1670 54270 1702
rect 54264 1638 54270 1670
rect 54334 1670 54335 1702
rect 54334 1638 54340 1670
rect 54264 1294 54340 1638
rect 54264 1230 54270 1294
rect 54334 1230 54340 1294
rect 54264 1224 54340 1230
rect 54400 0 54476 10614
rect 54672 10614 54678 10678
rect 54742 10614 54748 10678
rect 55629 10678 55695 10679
rect 55629 10646 55630 10678
rect 54672 10134 54748 10614
rect 54672 10102 54678 10134
rect 54677 10070 54678 10102
rect 54742 10102 54748 10134
rect 55624 10614 55630 10646
rect 55694 10646 55695 10678
rect 55896 10678 55972 10684
rect 55694 10614 55700 10646
rect 54742 10070 54743 10102
rect 54677 10069 54743 10070
rect 54677 9862 54743 9863
rect 54677 9830 54678 9862
rect 54672 9798 54678 9830
rect 54742 9830 54743 9862
rect 54742 9798 54748 9830
rect 54541 9454 54607 9455
rect 54541 9422 54542 9454
rect 54536 9390 54542 9422
rect 54606 9422 54607 9454
rect 54606 9390 54612 9422
rect 54536 8638 54612 9390
rect 54672 9318 54748 9798
rect 54672 9254 54678 9318
rect 54742 9254 54748 9318
rect 54672 9248 54748 9254
rect 54536 8574 54542 8638
rect 54606 8574 54612 8638
rect 54536 8568 54612 8574
rect 55221 2926 55287 2927
rect 55221 2894 55222 2926
rect 55216 2862 55222 2894
rect 55286 2894 55287 2926
rect 55286 2862 55292 2894
rect 55216 0 55292 2862
rect 55624 0 55700 10614
rect 55896 10614 55902 10678
rect 55966 10614 55972 10678
rect 56853 10678 56919 10679
rect 56853 10646 56854 10678
rect 55896 10134 55972 10614
rect 55896 10102 55902 10134
rect 55901 10070 55902 10102
rect 55966 10102 55972 10134
rect 56848 10614 56854 10646
rect 56918 10646 56919 10678
rect 57256 10678 57332 10684
rect 56918 10614 56924 10646
rect 55966 10070 55967 10102
rect 55901 10069 55967 10070
rect 56037 9862 56103 9863
rect 56037 9830 56038 9862
rect 56032 9798 56038 9830
rect 56102 9830 56103 9862
rect 56712 9862 56788 9868
rect 56102 9798 56108 9830
rect 55901 9454 55967 9455
rect 55901 9422 55902 9454
rect 55896 9390 55902 9422
rect 55966 9422 55967 9454
rect 55966 9390 55972 9422
rect 55896 8638 55972 9390
rect 56032 9318 56108 9798
rect 56032 9254 56038 9318
rect 56102 9254 56108 9318
rect 56712 9798 56718 9862
rect 56782 9798 56788 9862
rect 56712 9318 56788 9798
rect 56712 9286 56718 9318
rect 56032 9248 56108 9254
rect 56717 9254 56718 9286
rect 56782 9286 56788 9318
rect 56782 9254 56783 9286
rect 56717 9253 56783 9254
rect 55896 8574 55902 8638
rect 55966 8574 55972 8638
rect 55896 8568 55972 8574
rect 56581 2926 56647 2927
rect 56581 2894 56582 2926
rect 56576 2862 56582 2894
rect 56646 2894 56647 2926
rect 56646 2862 56652 2894
rect 55901 1702 55967 1703
rect 55901 1670 55902 1702
rect 55896 1638 55902 1670
rect 55966 1670 55967 1702
rect 55966 1638 55972 1670
rect 55896 1294 55972 1638
rect 55896 1230 55902 1294
rect 55966 1230 55972 1294
rect 55896 1224 55972 1230
rect 56576 0 56652 2862
rect 56848 0 56924 10614
rect 57256 10614 57262 10678
rect 57326 10614 57332 10678
rect 57805 10678 57871 10679
rect 57805 10646 57806 10678
rect 57256 10134 57332 10614
rect 57256 10102 57262 10134
rect 57261 10070 57262 10102
rect 57326 10102 57332 10134
rect 57800 10614 57806 10646
rect 57870 10646 57871 10678
rect 58480 10678 58556 10684
rect 57870 10614 57876 10646
rect 57326 10070 57327 10102
rect 57261 10069 57327 10070
rect 57125 9862 57191 9863
rect 57125 9830 57126 9862
rect 57120 9798 57126 9830
rect 57190 9830 57191 9862
rect 57190 9798 57196 9830
rect 56989 9454 57055 9455
rect 56989 9422 56990 9454
rect 56984 9390 56990 9422
rect 57054 9422 57055 9454
rect 57054 9390 57060 9422
rect 56984 8638 57060 9390
rect 57120 9318 57196 9798
rect 57120 9254 57126 9318
rect 57190 9254 57196 9318
rect 57120 9248 57196 9254
rect 56984 8574 56990 8638
rect 57054 8574 57060 8638
rect 56984 8568 57060 8574
rect 57669 2926 57735 2927
rect 57669 2894 57670 2926
rect 57664 2862 57670 2894
rect 57734 2894 57735 2926
rect 57734 2862 57740 2894
rect 57533 1702 57599 1703
rect 57533 1670 57534 1702
rect 57528 1638 57534 1670
rect 57598 1670 57599 1702
rect 57598 1638 57604 1670
rect 57528 1294 57604 1638
rect 57528 1230 57534 1294
rect 57598 1230 57604 1294
rect 57528 1224 57604 1230
rect 57664 0 57740 2862
rect 57800 0 57876 10614
rect 58480 10614 58486 10678
rect 58550 10614 58556 10678
rect 59165 10678 59231 10679
rect 59165 10646 59166 10678
rect 58480 10134 58556 10614
rect 58480 10102 58486 10134
rect 58485 10070 58486 10102
rect 58550 10102 58556 10134
rect 59160 10614 59166 10646
rect 59230 10646 59231 10678
rect 59301 10678 59367 10679
rect 59301 10646 59302 10678
rect 59230 10614 59236 10646
rect 59160 10134 59236 10614
rect 58550 10070 58551 10102
rect 58485 10069 58551 10070
rect 59160 10070 59166 10134
rect 59230 10070 59236 10134
rect 59160 10064 59236 10070
rect 59296 10614 59302 10646
rect 59366 10646 59367 10678
rect 59704 10678 59780 10684
rect 59366 10614 59372 10646
rect 58485 9862 58551 9863
rect 58485 9830 58486 9862
rect 58480 9798 58486 9830
rect 58550 9830 58551 9862
rect 58550 9798 58556 9830
rect 58349 9454 58415 9455
rect 58349 9422 58350 9454
rect 58344 9390 58350 9422
rect 58414 9422 58415 9454
rect 58414 9390 58420 9422
rect 58344 8638 58420 9390
rect 58480 9318 58556 9798
rect 58480 9254 58486 9318
rect 58550 9254 58556 9318
rect 58480 9248 58556 9254
rect 58344 8574 58350 8638
rect 58414 8574 58420 8638
rect 58344 8568 58420 8574
rect 59165 1702 59231 1703
rect 59165 1670 59166 1702
rect 59160 1638 59166 1670
rect 59230 1670 59231 1702
rect 59230 1638 59236 1670
rect 59160 1294 59236 1638
rect 59160 1230 59166 1294
rect 59230 1230 59236 1294
rect 59160 1224 59236 1230
rect 59296 0 59372 10614
rect 59704 10614 59710 10678
rect 59774 10614 59780 10678
rect 60525 10678 60591 10679
rect 60525 10646 60526 10678
rect 59704 10134 59780 10614
rect 59704 10102 59710 10134
rect 59709 10070 59710 10102
rect 59774 10102 59780 10134
rect 60520 10614 60526 10646
rect 60590 10646 60591 10678
rect 60928 10678 61004 10684
rect 60590 10614 60596 10646
rect 59774 10070 59775 10102
rect 59709 10069 59775 10070
rect 59709 9862 59775 9863
rect 59709 9830 59710 9862
rect 59704 9798 59710 9830
rect 59774 9830 59775 9862
rect 59774 9798 59780 9830
rect 59573 9454 59639 9455
rect 59573 9422 59574 9454
rect 59568 9390 59574 9422
rect 59638 9422 59639 9454
rect 59638 9390 59644 9422
rect 59568 8638 59644 9390
rect 59704 9318 59780 9798
rect 59704 9254 59710 9318
rect 59774 9254 59780 9318
rect 59704 9248 59780 9254
rect 59568 8574 59574 8638
rect 59638 8574 59644 8638
rect 59568 8568 59644 8574
rect 60520 0 60596 10614
rect 60928 10614 60934 10678
rect 60998 10614 61004 10678
rect 61749 10678 61815 10679
rect 61749 10646 61750 10678
rect 60928 10134 61004 10614
rect 60928 10102 60934 10134
rect 60933 10070 60934 10102
rect 60998 10102 61004 10134
rect 61744 10614 61750 10646
rect 61814 10646 61815 10678
rect 61885 10678 61951 10679
rect 61885 10646 61886 10678
rect 61814 10614 61820 10646
rect 61744 10134 61820 10614
rect 60998 10070 60999 10102
rect 60933 10069 60999 10070
rect 61744 10070 61750 10134
rect 61814 10070 61820 10134
rect 61744 10064 61820 10070
rect 61880 10614 61886 10646
rect 61950 10646 61951 10678
rect 62152 10678 62228 10684
rect 61950 10614 61956 10646
rect 60933 9862 60999 9863
rect 60933 9830 60934 9862
rect 60928 9798 60934 9830
rect 60998 9830 60999 9862
rect 60998 9798 61004 9830
rect 60797 9454 60863 9455
rect 60797 9422 60798 9454
rect 60792 9390 60798 9422
rect 60862 9422 60863 9454
rect 60862 9390 60868 9422
rect 60792 8638 60868 9390
rect 60928 9318 61004 9798
rect 60928 9254 60934 9318
rect 60998 9254 61004 9318
rect 60928 9248 61004 9254
rect 60792 8574 60798 8638
rect 60862 8574 60868 8638
rect 60792 8568 60868 8574
rect 60933 1702 60999 1703
rect 60933 1670 60934 1702
rect 60928 1638 60934 1670
rect 60998 1670 60999 1702
rect 60998 1638 61004 1670
rect 60928 1294 61004 1638
rect 60928 1230 60934 1294
rect 60998 1230 61004 1294
rect 60928 1224 61004 1230
rect 61880 0 61956 10614
rect 62152 10614 62158 10678
rect 62222 10614 62228 10678
rect 62973 10678 63039 10679
rect 62973 10646 62974 10678
rect 62152 10134 62228 10614
rect 62152 10102 62158 10134
rect 62157 10070 62158 10102
rect 62222 10102 62228 10134
rect 62968 10614 62974 10646
rect 63038 10646 63039 10678
rect 63109 10678 63175 10679
rect 63109 10646 63110 10678
rect 63038 10614 63044 10646
rect 62968 10134 63044 10614
rect 62222 10070 62223 10102
rect 62157 10069 62223 10070
rect 62968 10070 62974 10134
rect 63038 10070 63044 10134
rect 62968 10064 63044 10070
rect 63104 10614 63110 10646
rect 63174 10646 63175 10678
rect 63512 10678 63588 10684
rect 63174 10614 63180 10646
rect 62293 9862 62359 9863
rect 62293 9830 62294 9862
rect 62288 9798 62294 9830
rect 62358 9830 62359 9862
rect 62358 9798 62364 9830
rect 62157 9454 62223 9455
rect 62157 9422 62158 9454
rect 62152 9390 62158 9422
rect 62222 9422 62223 9454
rect 62222 9390 62228 9422
rect 62152 8638 62228 9390
rect 62288 9318 62364 9798
rect 62288 9254 62294 9318
rect 62358 9254 62364 9318
rect 62288 9248 62364 9254
rect 62152 8574 62158 8638
rect 62222 8574 62228 8638
rect 62152 8568 62228 8574
rect 62701 1702 62767 1703
rect 62701 1670 62702 1702
rect 62696 1638 62702 1670
rect 62766 1670 62767 1702
rect 62766 1638 62772 1670
rect 62696 1294 62772 1638
rect 62696 1230 62702 1294
rect 62766 1230 62772 1294
rect 62696 1224 62772 1230
rect 63104 0 63180 10614
rect 63512 10614 63518 10678
rect 63582 10614 63588 10678
rect 64333 10678 64399 10679
rect 64333 10646 64334 10678
rect 63512 10134 63588 10614
rect 63512 10102 63518 10134
rect 63517 10070 63518 10102
rect 63582 10102 63588 10134
rect 64328 10614 64334 10646
rect 64398 10646 64399 10678
rect 64736 10678 64812 10684
rect 64398 10614 64404 10646
rect 63582 10070 63583 10102
rect 63517 10069 63583 10070
rect 63517 9862 63583 9863
rect 63517 9830 63518 9862
rect 63512 9798 63518 9830
rect 63582 9830 63583 9862
rect 63582 9798 63588 9830
rect 63381 9454 63447 9455
rect 63381 9422 63382 9454
rect 63376 9390 63382 9422
rect 63446 9422 63447 9454
rect 63446 9390 63452 9422
rect 63376 8638 63452 9390
rect 63512 9318 63588 9798
rect 63512 9254 63518 9318
rect 63582 9254 63588 9318
rect 63512 9248 63588 9254
rect 63376 8574 63382 8638
rect 63446 8574 63452 8638
rect 63376 8568 63452 8574
rect 64061 1702 64127 1703
rect 64061 1670 64062 1702
rect 64056 1638 64062 1670
rect 64126 1670 64127 1702
rect 64126 1638 64132 1670
rect 64056 1294 64132 1638
rect 64056 1230 64062 1294
rect 64126 1230 64132 1294
rect 64056 1224 64132 1230
rect 64328 0 64404 10614
rect 64736 10614 64742 10678
rect 64806 10614 64812 10678
rect 65421 10678 65487 10679
rect 65421 10646 65422 10678
rect 64736 10134 64812 10614
rect 64736 10102 64742 10134
rect 64741 10070 64742 10102
rect 64806 10102 64812 10134
rect 65416 10614 65422 10646
rect 65486 10646 65487 10678
rect 65557 10678 65623 10679
rect 65557 10646 65558 10678
rect 65486 10614 65492 10646
rect 65416 10134 65492 10614
rect 64806 10070 64807 10102
rect 64741 10069 64807 10070
rect 65416 10070 65422 10134
rect 65486 10070 65492 10134
rect 65416 10064 65492 10070
rect 65552 10614 65558 10646
rect 65622 10646 65623 10678
rect 65960 10678 66036 10684
rect 65622 10614 65628 10646
rect 64736 9862 64812 9868
rect 64736 9798 64742 9862
rect 64806 9798 64812 9862
rect 64605 9454 64671 9455
rect 64605 9422 64606 9454
rect 64600 9390 64606 9422
rect 64670 9422 64671 9454
rect 64670 9390 64676 9422
rect 64600 8638 64676 9390
rect 64736 9046 64812 9798
rect 64736 9014 64742 9046
rect 64741 8982 64742 9014
rect 64806 9014 64812 9046
rect 64806 8982 64807 9014
rect 64741 8981 64807 8982
rect 64600 8574 64606 8638
rect 64670 8574 64676 8638
rect 64600 8568 64676 8574
rect 65552 0 65628 10614
rect 65960 10614 65966 10678
rect 66030 10614 66036 10678
rect 66781 10678 66847 10679
rect 66781 10646 66782 10678
rect 65960 10134 66036 10614
rect 65960 10102 65966 10134
rect 65965 10070 65966 10102
rect 66030 10102 66036 10134
rect 66776 10614 66782 10646
rect 66846 10646 66847 10678
rect 67048 10678 67124 10684
rect 66846 10614 66852 10646
rect 66030 10070 66031 10102
rect 65965 10069 66031 10070
rect 65829 9862 65895 9863
rect 65829 9830 65830 9862
rect 65824 9798 65830 9830
rect 65894 9830 65895 9862
rect 65894 9798 65900 9830
rect 65693 9454 65759 9455
rect 65693 9422 65694 9454
rect 65688 9390 65694 9422
rect 65758 9422 65759 9454
rect 65758 9390 65764 9422
rect 65688 8638 65764 9390
rect 65824 9318 65900 9798
rect 65824 9254 65830 9318
rect 65894 9254 65900 9318
rect 65824 9248 65900 9254
rect 65688 8574 65694 8638
rect 65758 8574 65764 8638
rect 65688 8568 65764 8574
rect 65965 1702 66031 1703
rect 65965 1670 65966 1702
rect 65960 1638 65966 1670
rect 66030 1670 66031 1702
rect 66030 1638 66036 1670
rect 65960 1294 66036 1638
rect 65960 1230 65966 1294
rect 66030 1230 66036 1294
rect 65960 1224 66036 1230
rect 66776 0 66852 10614
rect 67048 10614 67054 10678
rect 67118 10614 67124 10678
rect 67048 10134 67124 10614
rect 67048 10102 67054 10134
rect 67053 10070 67054 10102
rect 67118 10102 67124 10134
rect 82416 10134 82492 12790
rect 94656 12310 95004 13878
rect 94656 12246 94662 12310
rect 94726 12246 95004 12310
rect 83101 12038 83167 12039
rect 83101 12006 83102 12038
rect 83096 11974 83102 12006
rect 83166 12006 83167 12038
rect 83166 11974 83172 12006
rect 67118 10070 67119 10102
rect 67053 10069 67119 10070
rect 82416 10070 82422 10134
rect 82486 10070 82492 10134
rect 82416 10064 82492 10070
rect 82552 11494 82628 11500
rect 82552 11430 82558 11494
rect 82622 11430 82628 11494
rect 82416 9998 82492 10004
rect 82416 9934 82422 9998
rect 82486 9934 82492 9998
rect 67189 9862 67255 9863
rect 67189 9830 67190 9862
rect 67184 9798 67190 9830
rect 67254 9830 67255 9862
rect 67254 9798 67260 9830
rect 67053 9454 67119 9455
rect 67053 9422 67054 9454
rect 67048 9390 67054 9422
rect 67118 9422 67119 9454
rect 67118 9390 67124 9422
rect 67048 8638 67124 9390
rect 67184 9318 67260 9798
rect 67184 9254 67190 9318
rect 67254 9254 67260 9318
rect 67184 9248 67260 9254
rect 68005 8910 68071 8911
rect 68005 8878 68006 8910
rect 68000 8846 68006 8878
rect 68070 8878 68071 8910
rect 68070 8846 68076 8878
rect 67048 8574 67054 8638
rect 67118 8574 67124 8638
rect 67869 8638 67935 8639
rect 67869 8606 67870 8638
rect 67048 8568 67124 8574
rect 67864 8574 67870 8606
rect 67934 8606 67935 8638
rect 67934 8574 67940 8606
rect 67864 8230 67940 8574
rect 67864 8166 67870 8230
rect 67934 8166 67940 8230
rect 67864 8160 67940 8166
rect 68000 7142 68076 8846
rect 82416 7414 82492 9934
rect 82552 8774 82628 11430
rect 82693 10950 82759 10951
rect 82693 10918 82694 10950
rect 82552 8742 82558 8774
rect 82557 8710 82558 8742
rect 82622 8742 82628 8774
rect 82688 10886 82694 10918
rect 82758 10918 82759 10950
rect 82758 10886 82764 10918
rect 82622 8710 82623 8742
rect 82557 8709 82623 8710
rect 82416 7382 82422 7414
rect 82421 7350 82422 7382
rect 82486 7382 82492 7414
rect 82486 7350 82487 7382
rect 82421 7349 82487 7350
rect 68000 7078 68006 7142
rect 68070 7078 68076 7142
rect 68000 7072 68076 7078
rect 67733 1702 67799 1703
rect 67733 1670 67734 1702
rect 67728 1638 67734 1670
rect 67798 1670 67799 1702
rect 69229 1702 69295 1703
rect 69229 1670 69230 1702
rect 67798 1638 67804 1670
rect 67728 1294 67804 1638
rect 67728 1230 67734 1294
rect 67798 1230 67804 1294
rect 67728 1224 67804 1230
rect 69224 1638 69230 1670
rect 69294 1670 69295 1702
rect 70997 1702 71063 1703
rect 70997 1670 70998 1702
rect 69294 1638 69300 1670
rect 69224 1294 69300 1638
rect 69224 1230 69230 1294
rect 69294 1230 69300 1294
rect 69224 1224 69300 1230
rect 70992 1638 70998 1670
rect 71062 1670 71063 1702
rect 72629 1702 72695 1703
rect 72629 1670 72630 1702
rect 71062 1638 71068 1670
rect 70992 1294 71068 1638
rect 70992 1230 70998 1294
rect 71062 1230 71068 1294
rect 70992 1224 71068 1230
rect 72624 1638 72630 1670
rect 72694 1670 72695 1702
rect 74261 1702 74327 1703
rect 74261 1670 74262 1702
rect 72694 1638 72700 1670
rect 72624 1294 72700 1638
rect 72624 1230 72630 1294
rect 72694 1230 72700 1294
rect 72624 1224 72700 1230
rect 74256 1638 74262 1670
rect 74326 1670 74327 1702
rect 76165 1702 76231 1703
rect 76165 1670 76166 1702
rect 74326 1638 74332 1670
rect 74256 1294 74332 1638
rect 74256 1230 74262 1294
rect 74326 1230 74332 1294
rect 74256 1224 74332 1230
rect 76160 1638 76166 1670
rect 76230 1670 76231 1702
rect 77661 1702 77727 1703
rect 77661 1670 77662 1702
rect 76230 1638 76236 1670
rect 76160 1294 76236 1638
rect 76160 1230 76166 1294
rect 76230 1230 76236 1294
rect 76160 1224 76236 1230
rect 77656 1638 77662 1670
rect 77726 1670 77727 1702
rect 79429 1702 79495 1703
rect 79429 1670 79430 1702
rect 77726 1638 77732 1670
rect 77656 1294 77732 1638
rect 77656 1230 77662 1294
rect 77726 1230 77732 1294
rect 77656 1224 77732 1230
rect 79424 1638 79430 1670
rect 79494 1670 79495 1702
rect 81197 1702 81263 1703
rect 81197 1670 81198 1702
rect 79494 1638 79500 1670
rect 79424 1294 79500 1638
rect 79424 1230 79430 1294
rect 79494 1230 79500 1294
rect 79424 1224 79500 1230
rect 81192 1638 81198 1670
rect 81262 1670 81263 1702
rect 82557 1702 82623 1703
rect 82557 1670 82558 1702
rect 81262 1638 81268 1670
rect 81192 1294 81268 1638
rect 81192 1230 81198 1294
rect 81262 1230 81268 1294
rect 81192 1224 81268 1230
rect 82552 1638 82558 1670
rect 82622 1670 82623 1702
rect 82622 1638 82628 1670
rect 82552 1294 82628 1638
rect 82552 1230 82558 1294
rect 82622 1230 82628 1294
rect 82552 1224 82628 1230
rect 82688 0 82764 10886
rect 82829 9182 82895 9183
rect 82829 9150 82830 9182
rect 82824 9118 82830 9150
rect 82894 9150 82895 9182
rect 82894 9118 82900 9150
rect 82824 0 82900 9118
rect 82965 8094 83031 8095
rect 82965 8062 82966 8094
rect 82960 8030 82966 8062
rect 83030 8062 83031 8094
rect 83030 8030 83036 8062
rect 82960 0 83036 8030
rect 83096 0 83172 11974
rect 94656 10542 95004 12246
rect 94656 10478 94662 10542
rect 94726 10478 95004 10542
rect 94656 8910 95004 10478
rect 94656 8846 94662 8910
rect 94726 8846 95004 8910
rect 94656 7006 95004 8846
rect 94656 6942 94662 7006
rect 94726 6942 95004 7006
rect 94656 5374 95004 6942
rect 94656 5310 94662 5374
rect 94726 5310 95004 5374
rect 94656 3742 95004 5310
rect 94656 3678 94662 3742
rect 94726 3678 95004 3742
rect 94656 1974 95004 3678
rect 94656 1910 94662 1974
rect 94726 1910 95004 1974
rect 84461 1702 84527 1703
rect 84461 1670 84462 1702
rect 84456 1638 84462 1670
rect 84526 1670 84527 1702
rect 86229 1702 86295 1703
rect 86229 1670 86230 1702
rect 84526 1638 84532 1670
rect 84456 1294 84532 1638
rect 84456 1230 84462 1294
rect 84526 1230 84532 1294
rect 84456 1224 84532 1230
rect 86224 1638 86230 1670
rect 86294 1670 86295 1702
rect 87725 1702 87791 1703
rect 87725 1670 87726 1702
rect 86294 1638 86300 1670
rect 86224 1294 86300 1638
rect 86224 1230 86230 1294
rect 86294 1230 86300 1294
rect 86224 1224 86300 1230
rect 87720 1638 87726 1670
rect 87790 1670 87791 1702
rect 89493 1702 89559 1703
rect 89493 1670 89494 1702
rect 87790 1638 87796 1670
rect 87720 1294 87796 1638
rect 87720 1230 87726 1294
rect 87790 1230 87796 1294
rect 87720 1224 87796 1230
rect 89488 1638 89494 1670
rect 89558 1670 89559 1702
rect 91125 1702 91191 1703
rect 91125 1670 91126 1702
rect 89558 1638 89564 1670
rect 89488 1294 89564 1638
rect 89488 1230 89494 1294
rect 89558 1230 89564 1294
rect 89488 1224 89564 1230
rect 91120 1638 91126 1670
rect 91190 1670 91191 1702
rect 92757 1702 92823 1703
rect 92757 1670 92758 1702
rect 91190 1638 91196 1670
rect 91120 1294 91196 1638
rect 91120 1230 91126 1294
rect 91190 1230 91196 1294
rect 91120 1224 91196 1230
rect 92752 1638 92758 1670
rect 92822 1670 92823 1702
rect 92822 1638 92828 1670
rect 92752 1294 92828 1638
rect 92752 1230 92758 1294
rect 92822 1230 92828 1294
rect 92752 1224 92828 1230
rect 94656 1294 95004 1910
rect 94656 1230 94662 1294
rect 94726 1230 94798 1294
rect 94862 1230 94934 1294
rect 94998 1230 95004 1294
rect 94656 1158 95004 1230
rect 94656 1094 94662 1158
rect 94726 1094 94798 1158
rect 94862 1094 94934 1158
rect 94998 1094 95004 1158
rect 94656 1022 95004 1094
rect 94656 958 94662 1022
rect 94726 958 94798 1022
rect 94862 958 94934 1022
rect 94998 958 95004 1022
rect 94656 952 95004 958
rect 95336 77182 95684 78886
rect 95336 77118 95342 77182
rect 95406 77118 95684 77182
rect 95336 67254 95684 77118
rect 95336 67190 95342 67254
rect 95406 67190 95684 67254
rect 95336 61678 95684 67190
rect 95336 61614 95342 61678
rect 95406 61614 95684 61678
rect 95336 614 95684 61614
rect 95336 550 95342 614
rect 95406 550 95478 614
rect 95542 550 95614 614
rect 95678 550 95684 614
rect 95336 478 95684 550
rect 95336 414 95342 478
rect 95406 414 95478 478
rect 95542 414 95614 478
rect 95678 414 95684 478
rect 95336 342 95684 414
rect 95336 278 95342 342
rect 95406 278 95478 342
rect 95542 278 95614 342
rect 95678 278 95684 342
rect 95336 272 95684 278
use sky130_sram_1kbyte_1rw1r_32x256_8_bank  sky130_sram_1kbyte_1rw1r_32x256_8_bank_0
timestamp 1704896540
transform 1 0 14454 0 1 6974
box 0 0 67334 67312
use sky130_sram_1kbyte_1rw1r_32x256_8_col_addr_dff  sky130_sram_1kbyte_1rw1r_32x256_8_col_addr_dff_0
timestamp 1704896540
transform 1 0 15454 0 1 2388
box -36 -49 1204 1467
use sky130_sram_1kbyte_1rw1r_32x256_8_col_addr_dff  sky130_sram_1kbyte_1rw1r_32x256_8_col_addr_dff_1
timestamp 1704896540
transform -1 0 79620 0 -1 76383
box -36 -49 1204 1467
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_0
timestamp 1704896540
transform 1 0 94171 0 1 3695
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_1
timestamp 1704896540
transform 1 0 91189 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_2
timestamp 1704896540
transform 1 0 94171 0 1 2015
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_3
timestamp 1704896540
transform 1 0 92869 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_4
timestamp 1704896540
transform 1 0 84469 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_5
timestamp 1704896540
transform 1 0 89509 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_6
timestamp 1704896540
transform 1 0 87829 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_7
timestamp 1704896540
transform 1 0 86149 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_8
timestamp 1704896540
transform 1 0 94171 0 1 7055
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_9
timestamp 1704896540
transform 1 0 94171 0 1 5375
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_10
timestamp 1704896540
transform 1 0 94171 0 1 8735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_11
timestamp 1704896540
transform 1 0 81109 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_12
timestamp 1704896540
transform 1 0 79429 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_13
timestamp 1704896540
transform 1 0 82789 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_14
timestamp 1704896540
transform 1 0 72709 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_15
timestamp 1704896540
transform 1 0 76069 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_16
timestamp 1704896540
transform 1 0 74389 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_17
timestamp 1704896540
transform 1 0 81976 0 1 7994
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_18
timestamp 1704896540
transform 1 0 81238 0 1 9264
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_19
timestamp 1704896540
transform 1 0 81158 0 1 7994
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_20
timestamp 1704896540
transform 1 0 82921 0 1 8065
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_21
timestamp 1704896540
transform 1 0 82921 0 1 9193
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_22
timestamp 1704896540
transform 1 0 81976 0 1 9264
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_23
timestamp 1704896540
transform 1 0 77749 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_24
timestamp 1704896540
transform 1 0 81976 0 1 14920
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_25
timestamp 1704896540
transform 1 0 81638 0 1 16478
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_26
timestamp 1704896540
transform 1 0 81976 0 1 16478
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_27
timestamp 1704896540
transform 1 0 82921 0 1 10893
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_28
timestamp 1704896540
transform 1 0 82921 0 1 12021
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_29
timestamp 1704896540
transform 1 0 82921 0 1 13721
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_30
timestamp 1704896540
transform 1 0 82921 0 1 14849
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_31
timestamp 1704896540
transform 1 0 82921 0 1 16549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_32
timestamp 1704896540
transform 1 0 81318 0 1 10822
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_33
timestamp 1704896540
transform 1 0 81976 0 1 10822
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_34
timestamp 1704896540
transform 1 0 81398 0 1 12092
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_35
timestamp 1704896540
transform 1 0 81976 0 1 12092
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_36
timestamp 1704896540
transform 1 0 81478 0 1 13650
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_37
timestamp 1704896540
transform 1 0 81976 0 1 13650
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_38
timestamp 1704896540
transform 1 0 81558 0 1 14920
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_39
timestamp 1704896540
transform 1 0 94171 0 1 18815
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_40
timestamp 1704896540
transform 1 0 94171 0 1 17135
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_41
timestamp 1704896540
transform 1 0 94171 0 1 15455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_42
timestamp 1704896540
transform 1 0 94171 0 1 13775
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_43
timestamp 1704896540
transform 1 0 94171 0 1 12095
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_44
timestamp 1704896540
transform 1 0 94171 0 1 10415
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_45
timestamp 1704896540
transform 1 0 69349 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_46
timestamp 1704896540
transform 1 0 65989 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_47
timestamp 1704896540
transform 1 0 71029 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_48
timestamp 1704896540
transform 1 0 67669 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_49
timestamp 1704896540
transform 1 0 64309 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_50
timestamp 1704896540
transform 1 0 62629 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_51
timestamp 1704896540
transform 1 0 60949 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_52
timestamp 1704896540
transform 1 0 57639 0 1 2915
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_53
timestamp 1704896540
transform 1 0 56471 0 1 2915
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_54
timestamp 1704896540
transform 1 0 55303 0 1 2915
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_55
timestamp 1704896540
transform 1 0 54135 0 1 2915
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_56
timestamp 1704896540
transform 1 0 59269 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_57
timestamp 1704896540
transform 1 0 57589 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_58
timestamp 1704896540
transform 1 0 54229 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_59
timestamp 1704896540
transform 1 0 55909 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_60
timestamp 1704896540
transform 1 0 52967 0 1 2915
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_61
timestamp 1704896540
transform 1 0 50869 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_62
timestamp 1704896540
transform 1 0 51799 0 1 2915
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_63
timestamp 1704896540
transform 1 0 50631 0 1 2915
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_64
timestamp 1704896540
transform 1 0 49463 0 1 2915
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_65
timestamp 1704896540
transform 1 0 48295 0 1 2915
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_66
timestamp 1704896540
transform 1 0 49189 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_67
timestamp 1704896540
transform 1 0 52549 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_68
timestamp 1704896540
transform 1 0 48173 0 1 10748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_69
timestamp 1704896540
transform 1 0 53165 0 1 10748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_70
timestamp 1704896540
transform 1 0 51917 0 1 10748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_71
timestamp 1704896540
transform 1 0 59405 0 1 10748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_72
timestamp 1704896540
transform 1 0 49421 0 1 10748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_73
timestamp 1704896540
transform 1 0 58157 0 1 10748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_74
timestamp 1704896540
transform 1 0 56909 0 1 10748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_75
timestamp 1704896540
transform 1 0 50669 0 1 10748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_76
timestamp 1704896540
transform 1 0 55661 0 1 10748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_77
timestamp 1704896540
transform 1 0 54413 0 1 10748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_78
timestamp 1704896540
transform 1 0 66893 0 1 10748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_79
timestamp 1704896540
transform 1 0 65645 0 1 10748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_80
timestamp 1704896540
transform 1 0 64397 0 1 10748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_81
timestamp 1704896540
transform 1 0 63149 0 1 10748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_82
timestamp 1704896540
transform 1 0 61901 0 1 10748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_83
timestamp 1704896540
transform 1 0 60653 0 1 10748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_84
timestamp 1704896540
transform 1 0 94171 0 1 22175
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_85
timestamp 1704896540
transform 1 0 94171 0 1 28895
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_86
timestamp 1704896540
transform 1 0 94171 0 1 20495
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_87
timestamp 1704896540
transform 1 0 94171 0 1 27215
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_88
timestamp 1704896540
transform 1 0 94171 0 1 25535
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_89
timestamp 1704896540
transform 1 0 94171 0 1 23855
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_90
timestamp 1704896540
transform 1 0 94171 0 1 38975
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_91
timestamp 1704896540
transform 1 0 94171 0 1 37295
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_92
timestamp 1704896540
transform 1 0 94171 0 1 35615
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_93
timestamp 1704896540
transform 1 0 94171 0 1 33935
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_94
timestamp 1704896540
transform 1 0 94171 0 1 32255
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_95
timestamp 1704896540
transform 1 0 94171 0 1 30575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_96
timestamp 1704896540
transform 1 0 45959 0 1 2915
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_97
timestamp 1704896540
transform 1 0 43623 0 1 2915
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_98
timestamp 1704896540
transform 1 0 44149 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_99
timestamp 1704896540
transform 1 0 42455 0 1 2915
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_100
timestamp 1704896540
transform 1 0 47509 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_101
timestamp 1704896540
transform 1 0 47127 0 1 2915
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_102
timestamp 1704896540
transform 1 0 44791 0 1 2915
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_103
timestamp 1704896540
transform 1 0 45829 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_104
timestamp 1704896540
transform 1 0 42469 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_105
timestamp 1704896540
transform 1 0 40789 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_106
timestamp 1704896540
transform 1 0 37429 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_107
timestamp 1704896540
transform 1 0 39109 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_108
timestamp 1704896540
transform 1 0 41287 0 1 2915
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_109
timestamp 1704896540
transform 1 0 36615 0 1 2915
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_110
timestamp 1704896540
transform 1 0 40119 0 1 2915
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_111
timestamp 1704896540
transform 1 0 38951 0 1 2915
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_112
timestamp 1704896540
transform 1 0 37783 0 1 2915
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_113
timestamp 1704896540
transform 1 0 35749 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_114
timestamp 1704896540
transform 1 0 33111 0 1 2915
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_115
timestamp 1704896540
transform 1 0 32389 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_116
timestamp 1704896540
transform 1 0 31943 0 1 2915
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_117
timestamp 1704896540
transform 1 0 34279 0 1 2915
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_118
timestamp 1704896540
transform 1 0 30775 0 1 2915
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_119
timestamp 1704896540
transform 1 0 35447 0 1 2915
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_120
timestamp 1704896540
transform 1 0 30709 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_121
timestamp 1704896540
transform 1 0 34069 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_122
timestamp 1704896540
transform 1 0 25669 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_123
timestamp 1704896540
transform 1 0 24935 0 1 2915
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_124
timestamp 1704896540
transform 1 0 28439 0 1 2915
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_125
timestamp 1704896540
transform 1 0 27271 0 1 2915
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_126
timestamp 1704896540
transform 1 0 26103 0 1 2915
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_127
timestamp 1704896540
transform 1 0 29029 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_128
timestamp 1704896540
transform 1 0 27349 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_129
timestamp 1704896540
transform 1 0 29607 0 1 2915
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_130
timestamp 1704896540
transform 1 0 26222 0 1 9836
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_131
timestamp 1704896540
transform 1 0 34445 0 1 10748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_132
timestamp 1704896540
transform 1 0 33197 0 1 10748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_133
timestamp 1704896540
transform 1 0 31949 0 1 10748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_134
timestamp 1704896540
transform 1 0 30701 0 1 10748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_135
timestamp 1704896540
transform 1 0 29453 0 1 10748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_136
timestamp 1704896540
transform 1 0 35693 0 1 10748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_137
timestamp 1704896540
transform 1 0 28205 0 1 10748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_138
timestamp 1704896540
transform 1 0 26098 0 1 12664
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_139
timestamp 1704896540
transform 1 0 26346 0 1 11250
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_140
timestamp 1704896540
transform 1 0 44429 0 1 10748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_141
timestamp 1704896540
transform 1 0 43181 0 1 10748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_142
timestamp 1704896540
transform 1 0 41933 0 1 10748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_143
timestamp 1704896540
transform 1 0 40685 0 1 10748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_144
timestamp 1704896540
transform 1 0 39437 0 1 10748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_145
timestamp 1704896540
transform 1 0 38189 0 1 10748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_146
timestamp 1704896540
transform 1 0 36941 0 1 10748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_147
timestamp 1704896540
transform 1 0 46925 0 1 10748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_148
timestamp 1704896540
transform 1 0 45677 0 1 10748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_149
timestamp 1704896540
transform 1 0 22309 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_150
timestamp 1704896540
transform 1 0 18949 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_151
timestamp 1704896540
transform 1 0 20629 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_152
timestamp 1704896540
transform 1 0 20263 0 1 2915
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_153
timestamp 1704896540
transform 1 0 19095 0 1 2915
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_154
timestamp 1704896540
transform 1 0 23767 0 1 2915
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_155
timestamp 1704896540
transform 1 0 23989 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_156
timestamp 1704896540
transform 1 0 22599 0 1 2915
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_157
timestamp 1704896540
transform 1 0 21431 0 1 2915
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_158
timestamp 1704896540
transform 1 0 12229 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_159
timestamp 1704896540
transform 1 0 17269 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_160
timestamp 1704896540
transform 1 0 17927 0 1 2915
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_161
timestamp 1704896540
transform 1 0 16759 0 1 2915
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_162
timestamp 1704896540
transform 1 0 13909 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_163
timestamp 1704896540
transform 1 0 15591 0 1 2915
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_164
timestamp 1704896540
transform 1 0 15589 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_165
timestamp 1704896540
transform 1 0 14253 0 1 9836
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_166
timestamp 1704896540
transform 1 0 7189 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_167
timestamp 1704896540
transform 1 0 10549 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_168
timestamp 1704896540
transform 1 0 8869 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_169
timestamp 1704896540
transform 1 0 2149 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_170
timestamp 1704896540
transform 1 0 5509 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_171
timestamp 1704896540
transform 1 0 1813 0 1 3695
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_172
timestamp 1704896540
transform 1 0 3829 0 1 1679
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_173
timestamp 1704896540
transform 1 0 1813 0 1 2015
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_174
timestamp 1704896540
transform 1 0 1813 0 1 7055
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_175
timestamp 1704896540
transform 1 0 1813 0 1 5375
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_176
timestamp 1704896540
transform 1 0 1813 0 1 8735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_177
timestamp 1704896540
transform 1 0 2773 0 1 5451
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_178
timestamp 1704896540
transform 1 0 5994 0 1 5556
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_179
timestamp 1704896540
transform 1 0 2773 0 1 7151
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_180
timestamp 1704896540
transform 1 0 1813 0 1 10415
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_181
timestamp 1704896540
transform 1 0 1813 0 1 12095
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_182
timestamp 1704896540
transform 1 0 1813 0 1 13775
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_183
timestamp 1704896540
transform 1 0 1813 0 1 17135
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_184
timestamp 1704896540
transform 1 0 1813 0 1 15455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_185
timestamp 1704896540
transform 1 0 1813 0 1 18815
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_186
timestamp 1704896540
transform 1 0 14253 0 1 12664
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_187
timestamp 1704896540
transform 1 0 22395 0 1 15492
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_188
timestamp 1704896540
transform 1 0 14253 0 1 15492
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_189
timestamp 1704896540
transform 1 0 14253 0 1 11250
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_190
timestamp 1704896540
transform 1 0 14534 0 1 27206
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_191
timestamp 1704896540
transform 1 0 14200 0 1 27206
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_192
timestamp 1704896540
transform 1 0 14454 0 1 25648
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_193
timestamp 1704896540
transform 1 0 14200 0 1 28476
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_194
timestamp 1704896540
transform 1 0 14614 0 1 28476
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_195
timestamp 1704896540
transform 1 0 14200 0 1 25648
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_196
timestamp 1704896540
transform 1 0 13255 0 1 28405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_197
timestamp 1704896540
transform 1 0 13255 0 1 27277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_198
timestamp 1704896540
transform 1 0 13255 0 1 25577
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_199
timestamp 1704896540
transform 1 0 2560 0 1 22600
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_200
timestamp 1704896540
transform 1 0 1813 0 1 20495
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_201
timestamp 1704896540
transform 1 0 1813 0 1 23855
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_202
timestamp 1704896540
transform 1 0 1813 0 1 22175
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_203
timestamp 1704896540
transform 1 0 1813 0 1 27215
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_204
timestamp 1704896540
transform 1 0 1813 0 1 25535
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_205
timestamp 1704896540
transform 1 0 1813 0 1 28895
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_206
timestamp 1704896540
transform 1 0 1813 0 1 35615
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_207
timestamp 1704896540
transform 1 0 1813 0 1 33935
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_208
timestamp 1704896540
transform 1 0 1813 0 1 32255
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_209
timestamp 1704896540
transform 1 0 1813 0 1 38975
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_210
timestamp 1704896540
transform 1 0 1813 0 1 37295
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_211
timestamp 1704896540
transform 1 0 1813 0 1 30575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_212
timestamp 1704896540
transform 1 0 14854 0 1 32862
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_213
timestamp 1704896540
transform 1 0 14200 0 1 32862
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_214
timestamp 1704896540
transform 1 0 14774 0 1 31304
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_215
timestamp 1704896540
transform 1 0 14200 0 1 31304
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_216
timestamp 1704896540
transform 1 0 14694 0 1 30034
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_217
timestamp 1704896540
transform 1 0 14200 0 1 30034
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_218
timestamp 1704896540
transform 1 0 14934 0 1 34132
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_219
timestamp 1704896540
transform 1 0 14200 0 1 34132
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_220
timestamp 1704896540
transform 1 0 13255 0 1 34061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_221
timestamp 1704896540
transform 1 0 13255 0 1 32933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_222
timestamp 1704896540
transform 1 0 13255 0 1 31233
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_223
timestamp 1704896540
transform 1 0 13255 0 1 30105
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_224
timestamp 1704896540
transform 1 0 1813 0 1 45695
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_225
timestamp 1704896540
transform 1 0 1813 0 1 44015
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_226
timestamp 1704896540
transform 1 0 1813 0 1 49055
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_227
timestamp 1704896540
transform 1 0 1813 0 1 40655
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_228
timestamp 1704896540
transform 1 0 1813 0 1 42335
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_229
timestamp 1704896540
transform 1 0 1813 0 1 47375
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_230
timestamp 1704896540
transform 1 0 1813 0 1 59135
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_231
timestamp 1704896540
transform 1 0 1813 0 1 57455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_232
timestamp 1704896540
transform 1 0 1813 0 1 55775
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_233
timestamp 1704896540
transform 1 0 1813 0 1 54095
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_234
timestamp 1704896540
transform 1 0 1813 0 1 50735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_235
timestamp 1704896540
transform 1 0 1813 0 1 52415
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_236
timestamp 1704896540
transform 1 0 1813 0 1 69215
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_237
timestamp 1704896540
transform 1 0 1813 0 1 67535
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_238
timestamp 1704896540
transform 1 0 1813 0 1 65855
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_239
timestamp 1704896540
transform 1 0 1813 0 1 64175
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_240
timestamp 1704896540
transform 1 0 1813 0 1 62495
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_241
timestamp 1704896540
transform 1 0 1813 0 1 60815
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_242
timestamp 1704896540
transform 1 0 1813 0 1 70895
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_243
timestamp 1704896540
transform 1 0 1813 0 1 72575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_244
timestamp 1704896540
transform 1 0 3829 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_245
timestamp 1704896540
transform 1 0 1813 0 1 75935
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_246
timestamp 1704896540
transform 1 0 2149 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_247
timestamp 1704896540
transform 1 0 5509 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_248
timestamp 1704896540
transform 1 0 10549 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_249
timestamp 1704896540
transform 1 0 8869 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_250
timestamp 1704896540
transform 1 0 7189 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_251
timestamp 1704896540
transform 1 0 1813 0 1 74255
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_252
timestamp 1704896540
transform 1 0 15589 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_253
timestamp 1704896540
transform 1 0 13909 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_254
timestamp 1704896540
transform 1 0 12229 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_255
timestamp 1704896540
transform 1 0 17269 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_256
timestamp 1704896540
transform 1 0 23989 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_257
timestamp 1704896540
transform 1 0 22309 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_258
timestamp 1704896540
transform 1 0 20629 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_259
timestamp 1704896540
transform 1 0 18949 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_260
timestamp 1704896540
transform 1 0 35693 0 1 74038
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_261
timestamp 1704896540
transform 1 0 34445 0 1 74038
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_262
timestamp 1704896540
transform 1 0 33197 0 1 74038
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_263
timestamp 1704896540
transform 1 0 31949 0 1 74038
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_264
timestamp 1704896540
transform 1 0 30701 0 1 74038
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_265
timestamp 1704896540
transform 1 0 29453 0 1 74038
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_266
timestamp 1704896540
transform 1 0 28205 0 1 74038
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_267
timestamp 1704896540
transform 1 0 25669 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_268
timestamp 1704896540
transform 1 0 29029 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_269
timestamp 1704896540
transform 1 0 27349 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_270
timestamp 1704896540
transform 1 0 35749 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_271
timestamp 1704896540
transform 1 0 34069 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_272
timestamp 1704896540
transform 1 0 32389 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_273
timestamp 1704896540
transform 1 0 30709 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_274
timestamp 1704896540
transform 1 0 46925 0 1 74038
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_275
timestamp 1704896540
transform 1 0 45677 0 1 74038
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_276
timestamp 1704896540
transform 1 0 44429 0 1 74038
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_277
timestamp 1704896540
transform 1 0 43181 0 1 74038
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_278
timestamp 1704896540
transform 1 0 41933 0 1 74038
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_279
timestamp 1704896540
transform 1 0 40685 0 1 74038
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_280
timestamp 1704896540
transform 1 0 39437 0 1 74038
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_281
timestamp 1704896540
transform 1 0 38189 0 1 74038
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_282
timestamp 1704896540
transform 1 0 36941 0 1 74038
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_283
timestamp 1704896540
transform 1 0 40789 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_284
timestamp 1704896540
transform 1 0 39109 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_285
timestamp 1704896540
transform 1 0 37429 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_286
timestamp 1704896540
transform 1 0 42469 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_287
timestamp 1704896540
transform 1 0 47509 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_288
timestamp 1704896540
transform 1 0 45829 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_289
timestamp 1704896540
transform 1 0 44149 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_290
timestamp 1704896540
transform 1 0 94171 0 1 45695
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_291
timestamp 1704896540
transform 1 0 94171 0 1 44015
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_292
timestamp 1704896540
transform 1 0 94171 0 1 42335
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_293
timestamp 1704896540
transform 1 0 94171 0 1 40655
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_294
timestamp 1704896540
transform 1 0 94171 0 1 49055
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_295
timestamp 1704896540
transform 1 0 94171 0 1 47375
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_296
timestamp 1704896540
transform 1 0 94171 0 1 50735
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_297
timestamp 1704896540
transform 1 0 94171 0 1 54095
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_298
timestamp 1704896540
transform 1 0 94171 0 1 52415
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_299
timestamp 1704896540
transform 1 0 94171 0 1 55775
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_300
timestamp 1704896540
transform 1 0 93424 0 1 59358
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_301
timestamp 1704896540
transform 1 0 94171 0 1 59135
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_302
timestamp 1704896540
transform 1 0 94171 0 1 57455
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_303
timestamp 1704896540
transform 1 0 55661 0 1 74038
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_304
timestamp 1704896540
transform 1 0 54413 0 1 74038
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_305
timestamp 1704896540
transform 1 0 59405 0 1 74038
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_306
timestamp 1704896540
transform 1 0 58157 0 1 74038
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_307
timestamp 1704896540
transform 1 0 56909 0 1 74038
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_308
timestamp 1704896540
transform 1 0 49421 0 1 74038
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_309
timestamp 1704896540
transform 1 0 48173 0 1 74038
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_310
timestamp 1704896540
transform 1 0 50669 0 1 74038
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_311
timestamp 1704896540
transform 1 0 53165 0 1 74038
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_312
timestamp 1704896540
transform 1 0 51917 0 1 74038
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_313
timestamp 1704896540
transform 1 0 52549 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_314
timestamp 1704896540
transform 1 0 50869 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_315
timestamp 1704896540
transform 1 0 49189 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_316
timestamp 1704896540
transform 1 0 59269 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_317
timestamp 1704896540
transform 1 0 57589 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_318
timestamp 1704896540
transform 1 0 55909 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_319
timestamp 1704896540
transform 1 0 54229 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_320
timestamp 1704896540
transform 1 0 69836 0 1 70708
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_321
timestamp 1704896540
transform 1 0 66893 0 1 74038
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_322
timestamp 1704896540
transform 1 0 69712 0 1 72122
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_323
timestamp 1704896540
transform 1 0 65645 0 1 74038
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_324
timestamp 1704896540
transform 1 0 64397 0 1 74038
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_325
timestamp 1704896540
transform 1 0 63149 0 1 74038
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_326
timestamp 1704896540
transform 1 0 61901 0 1 74038
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_327
timestamp 1704896540
transform 1 0 60653 0 1 74038
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_328
timestamp 1704896540
transform 1 0 60949 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_329
timestamp 1704896540
transform 1 0 64309 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_330
timestamp 1704896540
transform 1 0 62629 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_331
timestamp 1704896540
transform 1 0 71029 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_332
timestamp 1704896540
transform 1 0 69349 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_333
timestamp 1704896540
transform 1 0 67669 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_334
timestamp 1704896540
transform 1 0 65989 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_335
timestamp 1704896540
transform 1 0 94171 0 1 64175
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_336
timestamp 1704896540
transform 1 0 94171 0 1 62495
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_337
timestamp 1704896540
transform 1 0 94171 0 1 60815
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_338
timestamp 1704896540
transform 1 0 94171 0 1 69215
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_339
timestamp 1704896540
transform 1 0 94171 0 1 67535
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_340
timestamp 1704896540
transform 1 0 94171 0 1 65855
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_341
timestamp 1704896540
transform 1 0 81923 0 1 70708
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_342
timestamp 1704896540
transform 1 0 81923 0 1 72122
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_343
timestamp 1704896540
transform 1 0 72709 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_344
timestamp 1704896540
transform 1 0 74389 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_345
timestamp 1704896540
transform 1 0 76069 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_346
timestamp 1704896540
transform 1 0 79417 0 1 75782
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_347
timestamp 1704896540
transform 1 0 82789 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_348
timestamp 1704896540
transform 1 0 81109 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_349
timestamp 1704896540
transform 1 0 79429 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_350
timestamp 1704896540
transform 1 0 77749 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_351
timestamp 1704896540
transform 1 0 94171 0 1 70895
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_352
timestamp 1704896540
transform 1 0 94171 0 1 72575
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_353
timestamp 1704896540
transform 1 0 84469 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_354
timestamp 1704896540
transform 1 0 89509 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_355
timestamp 1704896540
transform 1 0 87829 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_356
timestamp 1704896540
transform 1 0 86149 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_357
timestamp 1704896540
transform 1 0 94171 0 1 75935
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_358
timestamp 1704896540
transform 1 0 90074 0 1 76402
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_359
timestamp 1704896540
transform 1 0 93211 0 1 76507
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_360
timestamp 1704896540
transform 1 0 92869 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_361
timestamp 1704896540
transform 1 0 91189 0 1 77743
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_362
timestamp 1704896540
transform 1 0 94171 0 1 74255
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_363
timestamp 1704896540
transform 1 0 73697 0 1 69294
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_7  sky130_sram_1kbyte_1rw1r_32x256_8_contact_7_364
timestamp 1704896540
transform 1 0 81923 0 1 69294
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_0
timestamp 1704896540
transform 1 0 93213 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_1
timestamp 1704896540
transform 1 0 94179 0 1 4699
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_2
timestamp 1704896540
transform 1 0 94179 0 1 4363
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_3
timestamp 1704896540
transform 1 0 92205 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_4
timestamp 1704896540
transform 1 0 91869 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_5
timestamp 1704896540
transform 1 0 91533 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_6
timestamp 1704896540
transform 1 0 94179 0 1 4027
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_7
timestamp 1704896540
transform 1 0 94179 0 1 3691
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_8
timestamp 1704896540
transform 1 0 94179 0 1 3355
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_9
timestamp 1704896540
transform 1 0 94179 0 1 3019
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_10
timestamp 1704896540
transform 1 0 94179 0 1 2683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_11
timestamp 1704896540
transform 1 0 94179 0 1 2347
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_12
timestamp 1704896540
transform 1 0 94179 0 1 2011
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_13
timestamp 1704896540
transform 1 0 91197 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_14
timestamp 1704896540
transform 1 0 94179 0 1 5035
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_15
timestamp 1704896540
transform 1 0 90861 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_16
timestamp 1704896540
transform 1 0 89853 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_17
timestamp 1704896540
transform 1 0 90525 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_18
timestamp 1704896540
transform 1 0 92877 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_19
timestamp 1704896540
transform 1 0 92541 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_20
timestamp 1704896540
transform 1 0 90189 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_21
timestamp 1704896540
transform 1 0 93549 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_22
timestamp 1704896540
transform 1 0 89517 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_23
timestamp 1704896540
transform 1 0 84477 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_24
timestamp 1704896540
transform 1 0 89181 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_25
timestamp 1704896540
transform 1 0 84141 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_26
timestamp 1704896540
transform 1 0 88845 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_27
timestamp 1704896540
transform 1 0 88509 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_28
timestamp 1704896540
transform 1 0 88173 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_29
timestamp 1704896540
transform 1 0 87837 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_30
timestamp 1704896540
transform 1 0 87501 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_31
timestamp 1704896540
transform 1 0 87165 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_32
timestamp 1704896540
transform 1 0 86829 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_33
timestamp 1704896540
transform 1 0 86493 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_34
timestamp 1704896540
transform 1 0 86157 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_35
timestamp 1704896540
transform 1 0 85821 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_36
timestamp 1704896540
transform 1 0 85485 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_37
timestamp 1704896540
transform 1 0 85149 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_38
timestamp 1704896540
transform 1 0 84813 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_39
timestamp 1704896540
transform 1 0 94179 0 1 7387
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_40
timestamp 1704896540
transform 1 0 94179 0 1 7051
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_41
timestamp 1704896540
transform 1 0 94179 0 1 6715
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_42
timestamp 1704896540
transform 1 0 94179 0 1 5707
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_43
timestamp 1704896540
transform 1 0 94179 0 1 5371
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_44
timestamp 1704896540
transform 1 0 94179 0 1 6379
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_45
timestamp 1704896540
transform 1 0 94179 0 1 6043
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_46
timestamp 1704896540
transform 1 0 94179 0 1 9739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_47
timestamp 1704896540
transform 1 0 94179 0 1 9403
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_48
timestamp 1704896540
transform 1 0 94179 0 1 9067
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_49
timestamp 1704896540
transform 1 0 94179 0 1 8731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_50
timestamp 1704896540
transform 1 0 94179 0 1 8395
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_51
timestamp 1704896540
transform 1 0 94179 0 1 8059
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_52
timestamp 1704896540
transform 1 0 94179 0 1 7723
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_53
timestamp 1704896540
transform 1 0 78093 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_54
timestamp 1704896540
transform 1 0 82125 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_55
timestamp 1704896540
transform 1 0 81453 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_56
timestamp 1704896540
transform 1 0 81789 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_57
timestamp 1704896540
transform 1 0 82797 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_58
timestamp 1704896540
transform 1 0 78429 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_59
timestamp 1704896540
transform 1 0 83469 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_60
timestamp 1704896540
transform 1 0 81117 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_61
timestamp 1704896540
transform 1 0 80781 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_62
timestamp 1704896540
transform 1 0 80445 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_63
timestamp 1704896540
transform 1 0 80109 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_64
timestamp 1704896540
transform 1 0 79773 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_65
timestamp 1704896540
transform 1 0 82461 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_66
timestamp 1704896540
transform 1 0 83133 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_67
timestamp 1704896540
transform 1 0 79437 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_68
timestamp 1704896540
transform 1 0 79101 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_69
timestamp 1704896540
transform 1 0 78765 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_70
timestamp 1704896540
transform 1 0 76077 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_71
timestamp 1704896540
transform 1 0 75741 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_72
timestamp 1704896540
transform 1 0 73053 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_73
timestamp 1704896540
transform 1 0 74397 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_74
timestamp 1704896540
transform 1 0 72045 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_75
timestamp 1704896540
transform 1 0 72717 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_76
timestamp 1704896540
transform 1 0 75405 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_77
timestamp 1704896540
transform 1 0 77421 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_78
timestamp 1704896540
transform 1 0 74061 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_79
timestamp 1704896540
transform 1 0 77085 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_80
timestamp 1704896540
transform 1 0 75069 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_81
timestamp 1704896540
transform 1 0 73725 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_82
timestamp 1704896540
transform 1 0 74733 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_83
timestamp 1704896540
transform 1 0 76749 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_84
timestamp 1704896540
transform 1 0 72381 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_85
timestamp 1704896540
transform 1 0 73389 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_86
timestamp 1704896540
transform 1 0 76413 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_87
timestamp 1704896540
transform 1 0 77757 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_88
timestamp 1704896540
transform 1 0 94179 0 1 19819
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_89
timestamp 1704896540
transform 1 0 94179 0 1 19483
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_90
timestamp 1704896540
transform 1 0 94179 0 1 19147
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_91
timestamp 1704896540
transform 1 0 94179 0 1 18811
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_92
timestamp 1704896540
transform 1 0 94179 0 1 18475
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_93
timestamp 1704896540
transform 1 0 94179 0 1 18139
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_94
timestamp 1704896540
transform 1 0 94179 0 1 17803
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_95
timestamp 1704896540
transform 1 0 94179 0 1 17467
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_96
timestamp 1704896540
transform 1 0 94179 0 1 17131
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_97
timestamp 1704896540
transform 1 0 94179 0 1 16795
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_98
timestamp 1704896540
transform 1 0 94179 0 1 16459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_99
timestamp 1704896540
transform 1 0 94179 0 1 16123
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_100
timestamp 1704896540
transform 1 0 94179 0 1 15787
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_101
timestamp 1704896540
transform 1 0 94179 0 1 15451
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_102
timestamp 1704896540
transform 1 0 94179 0 1 15115
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_103
timestamp 1704896540
transform 1 0 94179 0 1 14779
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_104
timestamp 1704896540
transform 1 0 94179 0 1 14443
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_105
timestamp 1704896540
transform 1 0 94179 0 1 14107
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_106
timestamp 1704896540
transform 1 0 94179 0 1 13771
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_107
timestamp 1704896540
transform 1 0 94179 0 1 13435
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_108
timestamp 1704896540
transform 1 0 94179 0 1 13099
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_109
timestamp 1704896540
transform 1 0 94179 0 1 12763
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_110
timestamp 1704896540
transform 1 0 94179 0 1 12427
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_111
timestamp 1704896540
transform 1 0 94179 0 1 12091
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_112
timestamp 1704896540
transform 1 0 94179 0 1 11755
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_113
timestamp 1704896540
transform 1 0 94179 0 1 11419
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_114
timestamp 1704896540
transform 1 0 94179 0 1 11083
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_115
timestamp 1704896540
transform 1 0 94179 0 1 10747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_116
timestamp 1704896540
transform 1 0 94179 0 1 10411
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_117
timestamp 1704896540
transform 1 0 83805 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_118
timestamp 1704896540
transform 1 0 94179 0 1 10075
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_119
timestamp 1704896540
transform 1 0 65997 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_120
timestamp 1704896540
transform 1 0 67677 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_121
timestamp 1704896540
transform 1 0 69693 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_122
timestamp 1704896540
transform 1 0 66669 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_123
timestamp 1704896540
transform 1 0 69357 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_124
timestamp 1704896540
transform 1 0 71037 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_125
timestamp 1704896540
transform 1 0 66333 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_126
timestamp 1704896540
transform 1 0 69021 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_127
timestamp 1704896540
transform 1 0 71709 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_128
timestamp 1704896540
transform 1 0 67341 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_129
timestamp 1704896540
transform 1 0 70701 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_130
timestamp 1704896540
transform 1 0 68685 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_131
timestamp 1704896540
transform 1 0 71373 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_132
timestamp 1704896540
transform 1 0 70365 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_133
timestamp 1704896540
transform 1 0 67005 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_134
timestamp 1704896540
transform 1 0 70029 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_135
timestamp 1704896540
transform 1 0 68013 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_136
timestamp 1704896540
transform 1 0 68349 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_137
timestamp 1704896540
transform 1 0 65661 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_138
timestamp 1704896540
transform 1 0 65325 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_139
timestamp 1704896540
transform 1 0 64989 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_140
timestamp 1704896540
transform 1 0 64653 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_141
timestamp 1704896540
transform 1 0 63981 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_142
timestamp 1704896540
transform 1 0 63645 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_143
timestamp 1704896540
transform 1 0 62637 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_144
timestamp 1704896540
transform 1 0 63309 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_145
timestamp 1704896540
transform 1 0 62973 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_146
timestamp 1704896540
transform 1 0 62301 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_147
timestamp 1704896540
transform 1 0 61965 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_148
timestamp 1704896540
transform 1 0 61629 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_149
timestamp 1704896540
transform 1 0 61293 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_150
timestamp 1704896540
transform 1 0 64317 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_151
timestamp 1704896540
transform 1 0 60957 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_152
timestamp 1704896540
transform 1 0 60621 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_153
timestamp 1704896540
transform 1 0 60285 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_154
timestamp 1704896540
transform 1 0 55245 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_155
timestamp 1704896540
transform 1 0 59613 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_156
timestamp 1704896540
transform 1 0 54237 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_157
timestamp 1704896540
transform 1 0 54909 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_158
timestamp 1704896540
transform 1 0 59277 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_159
timestamp 1704896540
transform 1 0 58941 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_160
timestamp 1704896540
transform 1 0 58605 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_161
timestamp 1704896540
transform 1 0 58269 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_162
timestamp 1704896540
transform 1 0 57933 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_163
timestamp 1704896540
transform 1 0 54573 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_164
timestamp 1704896540
transform 1 0 57597 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_165
timestamp 1704896540
transform 1 0 57261 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_166
timestamp 1704896540
transform 1 0 56925 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_167
timestamp 1704896540
transform 1 0 56589 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_168
timestamp 1704896540
transform 1 0 56253 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_169
timestamp 1704896540
transform 1 0 55917 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_170
timestamp 1704896540
transform 1 0 55581 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_171
timestamp 1704896540
transform 1 0 50877 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_172
timestamp 1704896540
transform 1 0 50541 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_173
timestamp 1704896540
transform 1 0 48189 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_174
timestamp 1704896540
transform 1 0 48525 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_175
timestamp 1704896540
transform 1 0 52221 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_176
timestamp 1704896540
transform 1 0 50205 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_177
timestamp 1704896540
transform 1 0 51213 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_178
timestamp 1704896540
transform 1 0 51885 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_179
timestamp 1704896540
transform 1 0 49869 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_180
timestamp 1704896540
transform 1 0 51549 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_181
timestamp 1704896540
transform 1 0 49197 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_182
timestamp 1704896540
transform 1 0 53565 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_183
timestamp 1704896540
transform 1 0 48861 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_184
timestamp 1704896540
transform 1 0 49533 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_185
timestamp 1704896540
transform 1 0 53229 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_186
timestamp 1704896540
transform 1 0 52893 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_187
timestamp 1704896540
transform 1 0 52557 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_188
timestamp 1704896540
transform 1 0 53901 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_189
timestamp 1704896540
transform 1 0 59949 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_190
timestamp 1704896540
transform 1 0 94179 0 1 23515
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_191
timestamp 1704896540
transform 1 0 94179 0 1 23179
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_192
timestamp 1704896540
transform 1 0 94179 0 1 22843
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_193
timestamp 1704896540
transform 1 0 94179 0 1 22507
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_194
timestamp 1704896540
transform 1 0 94179 0 1 22171
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_195
timestamp 1704896540
transform 1 0 94179 0 1 29563
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_196
timestamp 1704896540
transform 1 0 94179 0 1 21835
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_197
timestamp 1704896540
transform 1 0 94179 0 1 21499
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_198
timestamp 1704896540
transform 1 0 94179 0 1 29227
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_199
timestamp 1704896540
transform 1 0 94179 0 1 28891
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_200
timestamp 1704896540
transform 1 0 94179 0 1 21163
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_201
timestamp 1704896540
transform 1 0 94179 0 1 20827
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_202
timestamp 1704896540
transform 1 0 94179 0 1 28555
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_203
timestamp 1704896540
transform 1 0 94179 0 1 20491
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_204
timestamp 1704896540
transform 1 0 94179 0 1 20155
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_205
timestamp 1704896540
transform 1 0 94179 0 1 28219
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_206
timestamp 1704896540
transform 1 0 94179 0 1 27883
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_207
timestamp 1704896540
transform 1 0 94179 0 1 27547
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_208
timestamp 1704896540
transform 1 0 94179 0 1 27211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_209
timestamp 1704896540
transform 1 0 94179 0 1 26875
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_210
timestamp 1704896540
transform 1 0 94179 0 1 26539
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_211
timestamp 1704896540
transform 1 0 94179 0 1 26203
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_212
timestamp 1704896540
transform 1 0 94179 0 1 25867
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_213
timestamp 1704896540
transform 1 0 94179 0 1 25531
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_214
timestamp 1704896540
transform 1 0 94179 0 1 25195
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_215
timestamp 1704896540
transform 1 0 94179 0 1 24859
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_216
timestamp 1704896540
transform 1 0 94179 0 1 24523
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_217
timestamp 1704896540
transform 1 0 94179 0 1 24187
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_218
timestamp 1704896540
transform 1 0 94179 0 1 23851
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_219
timestamp 1704896540
transform 1 0 94179 0 1 39307
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_220
timestamp 1704896540
transform 1 0 94179 0 1 38971
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_221
timestamp 1704896540
transform 1 0 94179 0 1 38635
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_222
timestamp 1704896540
transform 1 0 94179 0 1 38299
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_223
timestamp 1704896540
transform 1 0 94179 0 1 37963
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_224
timestamp 1704896540
transform 1 0 94179 0 1 37627
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_225
timestamp 1704896540
transform 1 0 94179 0 1 37291
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_226
timestamp 1704896540
transform 1 0 94179 0 1 36955
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_227
timestamp 1704896540
transform 1 0 94179 0 1 36619
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_228
timestamp 1704896540
transform 1 0 94179 0 1 36283
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_229
timestamp 1704896540
transform 1 0 94179 0 1 35947
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_230
timestamp 1704896540
transform 1 0 94179 0 1 35611
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_231
timestamp 1704896540
transform 1 0 94179 0 1 35275
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_232
timestamp 1704896540
transform 1 0 94179 0 1 34939
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_233
timestamp 1704896540
transform 1 0 94179 0 1 34603
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_234
timestamp 1704896540
transform 1 0 94179 0 1 34267
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_235
timestamp 1704896540
transform 1 0 94179 0 1 33931
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_236
timestamp 1704896540
transform 1 0 94179 0 1 33595
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_237
timestamp 1704896540
transform 1 0 94179 0 1 33259
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_238
timestamp 1704896540
transform 1 0 94179 0 1 32923
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_239
timestamp 1704896540
transform 1 0 94179 0 1 32587
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_240
timestamp 1704896540
transform 1 0 94179 0 1 32251
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_241
timestamp 1704896540
transform 1 0 94179 0 1 31915
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_242
timestamp 1704896540
transform 1 0 94179 0 1 31579
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_243
timestamp 1704896540
transform 1 0 94179 0 1 31243
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_244
timestamp 1704896540
transform 1 0 94179 0 1 30907
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_245
timestamp 1704896540
transform 1 0 94179 0 1 30571
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_246
timestamp 1704896540
transform 1 0 94179 0 1 30235
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_247
timestamp 1704896540
transform 1 0 94179 0 1 29899
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_248
timestamp 1704896540
transform 1 0 45165 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_249
timestamp 1704896540
transform 1 0 44829 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_250
timestamp 1704896540
transform 1 0 44493 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_251
timestamp 1704896540
transform 1 0 42141 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_252
timestamp 1704896540
transform 1 0 44157 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_253
timestamp 1704896540
transform 1 0 43821 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_254
timestamp 1704896540
transform 1 0 47853 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_255
timestamp 1704896540
transform 1 0 47517 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_256
timestamp 1704896540
transform 1 0 47181 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_257
timestamp 1704896540
transform 1 0 46845 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_258
timestamp 1704896540
transform 1 0 46509 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_259
timestamp 1704896540
transform 1 0 46173 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_260
timestamp 1704896540
transform 1 0 43485 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_261
timestamp 1704896540
transform 1 0 45837 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_262
timestamp 1704896540
transform 1 0 45501 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_263
timestamp 1704896540
transform 1 0 43149 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_264
timestamp 1704896540
transform 1 0 42813 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_265
timestamp 1704896540
transform 1 0 42477 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_266
timestamp 1704896540
transform 1 0 41133 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_267
timestamp 1704896540
transform 1 0 38109 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_268
timestamp 1704896540
transform 1 0 37773 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_269
timestamp 1704896540
transform 1 0 37437 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_270
timestamp 1704896540
transform 1 0 40797 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_271
timestamp 1704896540
transform 1 0 40461 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_272
timestamp 1704896540
transform 1 0 40125 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_273
timestamp 1704896540
transform 1 0 39789 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_274
timestamp 1704896540
transform 1 0 39453 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_275
timestamp 1704896540
transform 1 0 39117 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_276
timestamp 1704896540
transform 1 0 37101 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_277
timestamp 1704896540
transform 1 0 36765 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_278
timestamp 1704896540
transform 1 0 36429 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_279
timestamp 1704896540
transform 1 0 41805 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_280
timestamp 1704896540
transform 1 0 38781 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_281
timestamp 1704896540
transform 1 0 38445 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_282
timestamp 1704896540
transform 1 0 41469 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_283
timestamp 1704896540
transform 1 0 32733 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_284
timestamp 1704896540
transform 1 0 30717 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_285
timestamp 1704896540
transform 1 0 35757 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_286
timestamp 1704896540
transform 1 0 32397 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_287
timestamp 1704896540
transform 1 0 32061 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_288
timestamp 1704896540
transform 1 0 31725 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_289
timestamp 1704896540
transform 1 0 35421 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_290
timestamp 1704896540
transform 1 0 35085 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_291
timestamp 1704896540
transform 1 0 31389 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_292
timestamp 1704896540
transform 1 0 30381 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_293
timestamp 1704896540
transform 1 0 34749 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_294
timestamp 1704896540
transform 1 0 34413 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_295
timestamp 1704896540
transform 1 0 31053 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_296
timestamp 1704896540
transform 1 0 34077 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_297
timestamp 1704896540
transform 1 0 33741 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_298
timestamp 1704896540
transform 1 0 33405 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_299
timestamp 1704896540
transform 1 0 33069 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_300
timestamp 1704896540
transform 1 0 28701 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_301
timestamp 1704896540
transform 1 0 28365 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_302
timestamp 1704896540
transform 1 0 28029 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_303
timestamp 1704896540
transform 1 0 25341 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_304
timestamp 1704896540
transform 1 0 26349 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_305
timestamp 1704896540
transform 1 0 25005 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_306
timestamp 1704896540
transform 1 0 26013 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_307
timestamp 1704896540
transform 1 0 25677 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_308
timestamp 1704896540
transform 1 0 24669 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_309
timestamp 1704896540
transform 1 0 27357 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_310
timestamp 1704896540
transform 1 0 27021 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_311
timestamp 1704896540
transform 1 0 29709 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_312
timestamp 1704896540
transform 1 0 29373 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_313
timestamp 1704896540
transform 1 0 24333 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_314
timestamp 1704896540
transform 1 0 27693 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_315
timestamp 1704896540
transform 1 0 26685 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_316
timestamp 1704896540
transform 1 0 29037 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_317
timestamp 1704896540
transform 1 0 30045 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_318
timestamp 1704896540
transform 1 0 36093 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_319
timestamp 1704896540
transform 1 0 22653 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_320
timestamp 1704896540
transform 1 0 21309 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_321
timestamp 1704896540
transform 1 0 21645 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_322
timestamp 1704896540
transform 1 0 22317 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_323
timestamp 1704896540
transform 1 0 20637 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_324
timestamp 1704896540
transform 1 0 18285 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_325
timestamp 1704896540
transform 1 0 18621 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_326
timestamp 1704896540
transform 1 0 20973 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_327
timestamp 1704896540
transform 1 0 18957 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_328
timestamp 1704896540
transform 1 0 20301 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_329
timestamp 1704896540
transform 1 0 19965 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_330
timestamp 1704896540
transform 1 0 23997 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_331
timestamp 1704896540
transform 1 0 23661 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_332
timestamp 1704896540
transform 1 0 19629 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_333
timestamp 1704896540
transform 1 0 23325 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_334
timestamp 1704896540
transform 1 0 19293 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_335
timestamp 1704896540
transform 1 0 22989 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_336
timestamp 1704896540
transform 1 0 21981 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_337
timestamp 1704896540
transform 1 0 13245 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_338
timestamp 1704896540
transform 1 0 12909 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_339
timestamp 1704896540
transform 1 0 12573 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_340
timestamp 1704896540
transform 1 0 17949 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_341
timestamp 1704896540
transform 1 0 14253 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_342
timestamp 1704896540
transform 1 0 13917 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_343
timestamp 1704896540
transform 1 0 17277 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_344
timestamp 1704896540
transform 1 0 16941 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_345
timestamp 1704896540
transform 1 0 16605 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_346
timestamp 1704896540
transform 1 0 17613 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_347
timestamp 1704896540
transform 1 0 16269 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_348
timestamp 1704896540
transform 1 0 13581 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_349
timestamp 1704896540
transform 1 0 15933 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_350
timestamp 1704896540
transform 1 0 15597 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_351
timestamp 1704896540
transform 1 0 15261 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_352
timestamp 1704896540
transform 1 0 14925 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_353
timestamp 1704896540
transform 1 0 14589 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_354
timestamp 1704896540
transform 1 0 7197 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_355
timestamp 1704896540
transform 1 0 6861 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_356
timestamp 1704896540
transform 1 0 6525 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_357
timestamp 1704896540
transform 1 0 11901 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_358
timestamp 1704896540
transform 1 0 11565 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_359
timestamp 1704896540
transform 1 0 11229 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_360
timestamp 1704896540
transform 1 0 10893 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_361
timestamp 1704896540
transform 1 0 10557 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_362
timestamp 1704896540
transform 1 0 10221 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_363
timestamp 1704896540
transform 1 0 9885 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_364
timestamp 1704896540
transform 1 0 9549 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_365
timestamp 1704896540
transform 1 0 9213 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_366
timestamp 1704896540
transform 1 0 8877 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_367
timestamp 1704896540
transform 1 0 8541 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_368
timestamp 1704896540
transform 1 0 8205 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_369
timestamp 1704896540
transform 1 0 7869 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_370
timestamp 1704896540
transform 1 0 7533 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_371
timestamp 1704896540
transform 1 0 1821 0 1 2011
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_372
timestamp 1704896540
transform 1 0 3501 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_373
timestamp 1704896540
transform 1 0 3165 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_374
timestamp 1704896540
transform 1 0 2829 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_375
timestamp 1704896540
transform 1 0 2493 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_376
timestamp 1704896540
transform 1 0 5853 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_377
timestamp 1704896540
transform 1 0 2157 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_378
timestamp 1704896540
transform 1 0 1821 0 1 5035
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_379
timestamp 1704896540
transform 1 0 1821 0 1 4699
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_380
timestamp 1704896540
transform 1 0 1821 0 1 4363
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_381
timestamp 1704896540
transform 1 0 5517 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_382
timestamp 1704896540
transform 1 0 1821 0 1 4027
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_383
timestamp 1704896540
transform 1 0 1821 0 1 3691
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_384
timestamp 1704896540
transform 1 0 5181 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_385
timestamp 1704896540
transform 1 0 4845 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_386
timestamp 1704896540
transform 1 0 1821 0 1 3355
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_387
timestamp 1704896540
transform 1 0 1821 0 1 3019
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_388
timestamp 1704896540
transform 1 0 1821 0 1 2683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_389
timestamp 1704896540
transform 1 0 4509 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_390
timestamp 1704896540
transform 1 0 4173 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_391
timestamp 1704896540
transform 1 0 1821 0 1 2347
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_392
timestamp 1704896540
transform 1 0 3837 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_393
timestamp 1704896540
transform 1 0 1821 0 1 7387
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_394
timestamp 1704896540
transform 1 0 1821 0 1 7051
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_395
timestamp 1704896540
transform 1 0 1821 0 1 6715
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_396
timestamp 1704896540
transform 1 0 1821 0 1 6379
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_397
timestamp 1704896540
transform 1 0 1821 0 1 6043
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_398
timestamp 1704896540
transform 1 0 1821 0 1 5707
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_399
timestamp 1704896540
transform 1 0 1821 0 1 5371
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_400
timestamp 1704896540
transform 1 0 1821 0 1 9403
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_401
timestamp 1704896540
transform 1 0 1821 0 1 9067
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_402
timestamp 1704896540
transform 1 0 1821 0 1 8731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_403
timestamp 1704896540
transform 1 0 1821 0 1 8395
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_404
timestamp 1704896540
transform 1 0 1821 0 1 7723
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_405
timestamp 1704896540
transform 1 0 1821 0 1 8059
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_406
timestamp 1704896540
transform 1 0 1821 0 1 9739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_407
timestamp 1704896540
transform 1 0 6189 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_408
timestamp 1704896540
transform 1 0 1821 0 1 10747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_409
timestamp 1704896540
transform 1 0 1821 0 1 13435
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_410
timestamp 1704896540
transform 1 0 1821 0 1 13099
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_411
timestamp 1704896540
transform 1 0 1821 0 1 12763
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_412
timestamp 1704896540
transform 1 0 1821 0 1 12427
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_413
timestamp 1704896540
transform 1 0 1821 0 1 12091
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_414
timestamp 1704896540
transform 1 0 1821 0 1 11755
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_415
timestamp 1704896540
transform 1 0 1821 0 1 11419
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_416
timestamp 1704896540
transform 1 0 1821 0 1 11083
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_417
timestamp 1704896540
transform 1 0 1821 0 1 14779
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_418
timestamp 1704896540
transform 1 0 1821 0 1 14443
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_419
timestamp 1704896540
transform 1 0 1821 0 1 10411
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_420
timestamp 1704896540
transform 1 0 1821 0 1 14107
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_421
timestamp 1704896540
transform 1 0 1821 0 1 13771
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_422
timestamp 1704896540
transform 1 0 1821 0 1 17803
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_423
timestamp 1704896540
transform 1 0 1821 0 1 17467
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_424
timestamp 1704896540
transform 1 0 1821 0 1 17131
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_425
timestamp 1704896540
transform 1 0 1821 0 1 16795
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_426
timestamp 1704896540
transform 1 0 1821 0 1 16459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_427
timestamp 1704896540
transform 1 0 1821 0 1 16123
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_428
timestamp 1704896540
transform 1 0 1821 0 1 15787
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_429
timestamp 1704896540
transform 1 0 1821 0 1 15451
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_430
timestamp 1704896540
transform 1 0 1821 0 1 19819
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_431
timestamp 1704896540
transform 1 0 1821 0 1 19483
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_432
timestamp 1704896540
transform 1 0 1821 0 1 19147
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_433
timestamp 1704896540
transform 1 0 1821 0 1 18811
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_434
timestamp 1704896540
transform 1 0 1821 0 1 18475
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_435
timestamp 1704896540
transform 1 0 1821 0 1 18139
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_436
timestamp 1704896540
transform 1 0 1821 0 1 15115
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_437
timestamp 1704896540
transform 1 0 12237 0 1 1675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_438
timestamp 1704896540
transform 1 0 1821 0 1 10075
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_439
timestamp 1704896540
transform 1 0 1821 0 1 22171
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_440
timestamp 1704896540
transform 1 0 1821 0 1 21835
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_441
timestamp 1704896540
transform 1 0 1821 0 1 20155
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_442
timestamp 1704896540
transform 1 0 1821 0 1 21499
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_443
timestamp 1704896540
transform 1 0 1821 0 1 21163
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_444
timestamp 1704896540
transform 1 0 1821 0 1 20827
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_445
timestamp 1704896540
transform 1 0 1821 0 1 20491
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_446
timestamp 1704896540
transform 1 0 1821 0 1 24523
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_447
timestamp 1704896540
transform 1 0 1821 0 1 24187
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_448
timestamp 1704896540
transform 1 0 1821 0 1 23851
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_449
timestamp 1704896540
transform 1 0 1821 0 1 23515
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_450
timestamp 1704896540
transform 1 0 1821 0 1 23179
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_451
timestamp 1704896540
transform 1 0 1821 0 1 22843
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_452
timestamp 1704896540
transform 1 0 1821 0 1 22507
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_453
timestamp 1704896540
transform 1 0 1821 0 1 27211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_454
timestamp 1704896540
transform 1 0 1821 0 1 26875
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_455
timestamp 1704896540
transform 1 0 1821 0 1 26539
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_456
timestamp 1704896540
transform 1 0 1821 0 1 26203
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_457
timestamp 1704896540
transform 1 0 1821 0 1 25867
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_458
timestamp 1704896540
transform 1 0 1821 0 1 25531
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_459
timestamp 1704896540
transform 1 0 1821 0 1 25195
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_460
timestamp 1704896540
transform 1 0 1821 0 1 27547
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_461
timestamp 1704896540
transform 1 0 1821 0 1 29563
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_462
timestamp 1704896540
transform 1 0 1821 0 1 29227
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_463
timestamp 1704896540
transform 1 0 1821 0 1 28891
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_464
timestamp 1704896540
transform 1 0 1821 0 1 28555
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_465
timestamp 1704896540
transform 1 0 1821 0 1 28219
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_466
timestamp 1704896540
transform 1 0 1821 0 1 27883
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_467
timestamp 1704896540
transform 1 0 1821 0 1 24859
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_468
timestamp 1704896540
transform 1 0 1821 0 1 30571
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_469
timestamp 1704896540
transform 1 0 1821 0 1 35947
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_470
timestamp 1704896540
transform 1 0 1821 0 1 30235
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_471
timestamp 1704896540
transform 1 0 1821 0 1 35611
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_472
timestamp 1704896540
transform 1 0 1821 0 1 35275
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_473
timestamp 1704896540
transform 1 0 1821 0 1 34939
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_474
timestamp 1704896540
transform 1 0 1821 0 1 34603
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_475
timestamp 1704896540
transform 1 0 1821 0 1 34267
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_476
timestamp 1704896540
transform 1 0 1821 0 1 33931
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_477
timestamp 1704896540
transform 1 0 1821 0 1 33595
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_478
timestamp 1704896540
transform 1 0 1821 0 1 33259
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_479
timestamp 1704896540
transform 1 0 1821 0 1 32923
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_480
timestamp 1704896540
transform 1 0 1821 0 1 32587
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_481
timestamp 1704896540
transform 1 0 1821 0 1 32251
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_482
timestamp 1704896540
transform 1 0 1821 0 1 31915
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_483
timestamp 1704896540
transform 1 0 1821 0 1 31579
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_484
timestamp 1704896540
transform 1 0 1821 0 1 39307
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_485
timestamp 1704896540
transform 1 0 1821 0 1 38971
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_486
timestamp 1704896540
transform 1 0 1821 0 1 38635
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_487
timestamp 1704896540
transform 1 0 1821 0 1 38299
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_488
timestamp 1704896540
transform 1 0 1821 0 1 37963
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_489
timestamp 1704896540
transform 1 0 1821 0 1 37627
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_490
timestamp 1704896540
transform 1 0 1821 0 1 31243
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_491
timestamp 1704896540
transform 1 0 1821 0 1 37291
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_492
timestamp 1704896540
transform 1 0 1821 0 1 30907
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_493
timestamp 1704896540
transform 1 0 1821 0 1 36955
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_494
timestamp 1704896540
transform 1 0 1821 0 1 36619
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_495
timestamp 1704896540
transform 1 0 1821 0 1 36283
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_496
timestamp 1704896540
transform 1 0 1821 0 1 29899
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_497
timestamp 1704896540
transform 1 0 1821 0 1 46699
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_498
timestamp 1704896540
transform 1 0 1821 0 1 46363
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_499
timestamp 1704896540
transform 1 0 1821 0 1 46027
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_500
timestamp 1704896540
transform 1 0 1821 0 1 45691
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_501
timestamp 1704896540
transform 1 0 1821 0 1 45355
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_502
timestamp 1704896540
transform 1 0 1821 0 1 45019
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_503
timestamp 1704896540
transform 1 0 1821 0 1 44683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_504
timestamp 1704896540
transform 1 0 1821 0 1 44347
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_505
timestamp 1704896540
transform 1 0 1821 0 1 44011
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_506
timestamp 1704896540
transform 1 0 1821 0 1 49387
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_507
timestamp 1704896540
transform 1 0 1821 0 1 40315
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_508
timestamp 1704896540
transform 1 0 1821 0 1 39979
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_509
timestamp 1704896540
transform 1 0 1821 0 1 43339
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_510
timestamp 1704896540
transform 1 0 1821 0 1 41659
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_511
timestamp 1704896540
transform 1 0 1821 0 1 41323
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_512
timestamp 1704896540
transform 1 0 1821 0 1 41995
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_513
timestamp 1704896540
transform 1 0 1821 0 1 43003
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_514
timestamp 1704896540
transform 1 0 1821 0 1 43675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_515
timestamp 1704896540
transform 1 0 1821 0 1 47371
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_516
timestamp 1704896540
transform 1 0 1821 0 1 48379
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_517
timestamp 1704896540
transform 1 0 1821 0 1 40987
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_518
timestamp 1704896540
transform 1 0 1821 0 1 42667
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_519
timestamp 1704896540
transform 1 0 1821 0 1 48043
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_520
timestamp 1704896540
transform 1 0 1821 0 1 47035
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_521
timestamp 1704896540
transform 1 0 1821 0 1 47707
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_522
timestamp 1704896540
transform 1 0 1821 0 1 40651
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_523
timestamp 1704896540
transform 1 0 1821 0 1 42331
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_524
timestamp 1704896540
transform 1 0 1821 0 1 49051
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_525
timestamp 1704896540
transform 1 0 1821 0 1 48715
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_526
timestamp 1704896540
transform 1 0 1821 0 1 59131
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_527
timestamp 1704896540
transform 1 0 1821 0 1 58795
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_528
timestamp 1704896540
transform 1 0 1821 0 1 58459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_529
timestamp 1704896540
transform 1 0 1821 0 1 58123
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_530
timestamp 1704896540
transform 1 0 1821 0 1 57787
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_531
timestamp 1704896540
transform 1 0 1821 0 1 57451
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_532
timestamp 1704896540
transform 1 0 1821 0 1 57115
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_533
timestamp 1704896540
transform 1 0 1821 0 1 56779
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_534
timestamp 1704896540
transform 1 0 1821 0 1 56443
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_535
timestamp 1704896540
transform 1 0 1821 0 1 56107
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_536
timestamp 1704896540
transform 1 0 1821 0 1 55771
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_537
timestamp 1704896540
transform 1 0 1821 0 1 55435
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_538
timestamp 1704896540
transform 1 0 1821 0 1 55099
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_539
timestamp 1704896540
transform 1 0 1821 0 1 54763
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_540
timestamp 1704896540
transform 1 0 1821 0 1 54427
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_541
timestamp 1704896540
transform 1 0 1821 0 1 54091
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_542
timestamp 1704896540
transform 1 0 1821 0 1 50395
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_543
timestamp 1704896540
transform 1 0 1821 0 1 49723
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_544
timestamp 1704896540
transform 1 0 1821 0 1 50731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_545
timestamp 1704896540
transform 1 0 1821 0 1 50059
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_546
timestamp 1704896540
transform 1 0 1821 0 1 53755
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_547
timestamp 1704896540
transform 1 0 1821 0 1 52075
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_548
timestamp 1704896540
transform 1 0 1821 0 1 53419
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_549
timestamp 1704896540
transform 1 0 1821 0 1 51739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_550
timestamp 1704896540
transform 1 0 1821 0 1 51403
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_551
timestamp 1704896540
transform 1 0 1821 0 1 51067
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_552
timestamp 1704896540
transform 1 0 1821 0 1 53083
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_553
timestamp 1704896540
transform 1 0 1821 0 1 52747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_554
timestamp 1704896540
transform 1 0 1821 0 1 52411
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_555
timestamp 1704896540
transform 1 0 1821 0 1 60139
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_556
timestamp 1704896540
transform 1 0 1821 0 1 59803
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_557
timestamp 1704896540
transform 1 0 1821 0 1 69211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_558
timestamp 1704896540
transform 1 0 1821 0 1 68875
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_559
timestamp 1704896540
transform 1 0 1821 0 1 68539
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_560
timestamp 1704896540
transform 1 0 1821 0 1 68203
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_561
timestamp 1704896540
transform 1 0 1821 0 1 67867
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_562
timestamp 1704896540
transform 1 0 1821 0 1 67531
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_563
timestamp 1704896540
transform 1 0 1821 0 1 67195
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_564
timestamp 1704896540
transform 1 0 1821 0 1 66859
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_565
timestamp 1704896540
transform 1 0 1821 0 1 66523
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_566
timestamp 1704896540
transform 1 0 1821 0 1 66187
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_567
timestamp 1704896540
transform 1 0 1821 0 1 65851
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_568
timestamp 1704896540
transform 1 0 1821 0 1 65515
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_569
timestamp 1704896540
transform 1 0 1821 0 1 65179
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_570
timestamp 1704896540
transform 1 0 1821 0 1 64843
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_571
timestamp 1704896540
transform 1 0 1821 0 1 64507
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_572
timestamp 1704896540
transform 1 0 1821 0 1 64171
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_573
timestamp 1704896540
transform 1 0 1821 0 1 63835
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_574
timestamp 1704896540
transform 1 0 1821 0 1 63499
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_575
timestamp 1704896540
transform 1 0 1821 0 1 63163
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_576
timestamp 1704896540
transform 1 0 1821 0 1 62827
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_577
timestamp 1704896540
transform 1 0 1821 0 1 62491
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_578
timestamp 1704896540
transform 1 0 1821 0 1 62155
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_579
timestamp 1704896540
transform 1 0 1821 0 1 61819
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_580
timestamp 1704896540
transform 1 0 1821 0 1 61483
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_581
timestamp 1704896540
transform 1 0 1821 0 1 61147
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_582
timestamp 1704896540
transform 1 0 1821 0 1 60811
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_583
timestamp 1704896540
transform 1 0 1821 0 1 60475
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_584
timestamp 1704896540
transform 1 0 1821 0 1 70219
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_585
timestamp 1704896540
transform 1 0 1821 0 1 69883
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_586
timestamp 1704896540
transform 1 0 1821 0 1 69547
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_587
timestamp 1704896540
transform 1 0 1821 0 1 70555
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_588
timestamp 1704896540
transform 1 0 1821 0 1 71899
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_589
timestamp 1704896540
transform 1 0 1821 0 1 71563
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_590
timestamp 1704896540
transform 1 0 1821 0 1 73915
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_591
timestamp 1704896540
transform 1 0 1821 0 1 73579
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_592
timestamp 1704896540
transform 1 0 1821 0 1 73243
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_593
timestamp 1704896540
transform 1 0 1821 0 1 72907
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_594
timestamp 1704896540
transform 1 0 1821 0 1 72571
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_595
timestamp 1704896540
transform 1 0 1821 0 1 72235
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_596
timestamp 1704896540
transform 1 0 1821 0 1 71227
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_597
timestamp 1704896540
transform 1 0 1821 0 1 70891
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_598
timestamp 1704896540
transform 1 0 4173 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_599
timestamp 1704896540
transform 1 0 3837 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_600
timestamp 1704896540
transform 1 0 1821 0 1 77275
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_601
timestamp 1704896540
transform 1 0 1821 0 1 76939
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_602
timestamp 1704896540
transform 1 0 1821 0 1 76603
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_603
timestamp 1704896540
transform 1 0 1821 0 1 76267
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_604
timestamp 1704896540
transform 1 0 1821 0 1 75931
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_605
timestamp 1704896540
transform 1 0 1821 0 1 75595
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_606
timestamp 1704896540
transform 1 0 1821 0 1 75259
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_607
timestamp 1704896540
transform 1 0 1821 0 1 74923
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_608
timestamp 1704896540
transform 1 0 1821 0 1 74587
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_609
timestamp 1704896540
transform 1 0 3501 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_610
timestamp 1704896540
transform 1 0 3165 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_611
timestamp 1704896540
transform 1 0 2829 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_612
timestamp 1704896540
transform 1 0 2493 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_613
timestamp 1704896540
transform 1 0 2157 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_614
timestamp 1704896540
transform 1 0 5853 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_615
timestamp 1704896540
transform 1 0 5517 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_616
timestamp 1704896540
transform 1 0 5181 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_617
timestamp 1704896540
transform 1 0 4845 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_618
timestamp 1704896540
transform 1 0 4509 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_619
timestamp 1704896540
transform 1 0 6861 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_620
timestamp 1704896540
transform 1 0 6525 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_621
timestamp 1704896540
transform 1 0 11901 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_622
timestamp 1704896540
transform 1 0 11565 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_623
timestamp 1704896540
transform 1 0 11229 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_624
timestamp 1704896540
transform 1 0 10893 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_625
timestamp 1704896540
transform 1 0 10557 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_626
timestamp 1704896540
transform 1 0 10221 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_627
timestamp 1704896540
transform 1 0 9885 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_628
timestamp 1704896540
transform 1 0 9549 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_629
timestamp 1704896540
transform 1 0 9213 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_630
timestamp 1704896540
transform 1 0 8877 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_631
timestamp 1704896540
transform 1 0 8541 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_632
timestamp 1704896540
transform 1 0 8205 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_633
timestamp 1704896540
transform 1 0 7869 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_634
timestamp 1704896540
transform 1 0 7533 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_635
timestamp 1704896540
transform 1 0 7197 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_636
timestamp 1704896540
transform 1 0 1821 0 1 74251
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_637
timestamp 1704896540
transform 1 0 6189 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_638
timestamp 1704896540
transform 1 0 17277 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_639
timestamp 1704896540
transform 1 0 16941 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_640
timestamp 1704896540
transform 1 0 16605 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_641
timestamp 1704896540
transform 1 0 16269 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_642
timestamp 1704896540
transform 1 0 15933 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_643
timestamp 1704896540
transform 1 0 15597 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_644
timestamp 1704896540
transform 1 0 15261 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_645
timestamp 1704896540
transform 1 0 14925 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_646
timestamp 1704896540
transform 1 0 14589 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_647
timestamp 1704896540
transform 1 0 14253 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_648
timestamp 1704896540
transform 1 0 13917 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_649
timestamp 1704896540
transform 1 0 13581 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_650
timestamp 1704896540
transform 1 0 13245 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_651
timestamp 1704896540
transform 1 0 12909 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_652
timestamp 1704896540
transform 1 0 12573 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_653
timestamp 1704896540
transform 1 0 17949 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_654
timestamp 1704896540
transform 1 0 17613 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_655
timestamp 1704896540
transform 1 0 23997 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_656
timestamp 1704896540
transform 1 0 23661 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_657
timestamp 1704896540
transform 1 0 23325 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_658
timestamp 1704896540
transform 1 0 22989 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_659
timestamp 1704896540
transform 1 0 22653 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_660
timestamp 1704896540
transform 1 0 22317 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_661
timestamp 1704896540
transform 1 0 21981 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_662
timestamp 1704896540
transform 1 0 21645 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_663
timestamp 1704896540
transform 1 0 21309 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_664
timestamp 1704896540
transform 1 0 20973 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_665
timestamp 1704896540
transform 1 0 20637 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_666
timestamp 1704896540
transform 1 0 20301 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_667
timestamp 1704896540
transform 1 0 19965 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_668
timestamp 1704896540
transform 1 0 19629 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_669
timestamp 1704896540
transform 1 0 19293 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_670
timestamp 1704896540
transform 1 0 18957 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_671
timestamp 1704896540
transform 1 0 18621 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_672
timestamp 1704896540
transform 1 0 18285 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_673
timestamp 1704896540
transform 1 0 12237 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_674
timestamp 1704896540
transform 1 0 25677 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_675
timestamp 1704896540
transform 1 0 25341 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_676
timestamp 1704896540
transform 1 0 25005 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_677
timestamp 1704896540
transform 1 0 24669 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_678
timestamp 1704896540
transform 1 0 24333 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_679
timestamp 1704896540
transform 1 0 29709 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_680
timestamp 1704896540
transform 1 0 29373 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_681
timestamp 1704896540
transform 1 0 29037 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_682
timestamp 1704896540
transform 1 0 28701 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_683
timestamp 1704896540
transform 1 0 28365 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_684
timestamp 1704896540
transform 1 0 28029 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_685
timestamp 1704896540
transform 1 0 27693 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_686
timestamp 1704896540
transform 1 0 27357 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_687
timestamp 1704896540
transform 1 0 27021 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_688
timestamp 1704896540
transform 1 0 26685 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_689
timestamp 1704896540
transform 1 0 26349 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_690
timestamp 1704896540
transform 1 0 26013 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_691
timestamp 1704896540
transform 1 0 35757 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_692
timestamp 1704896540
transform 1 0 35421 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_693
timestamp 1704896540
transform 1 0 35085 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_694
timestamp 1704896540
transform 1 0 34749 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_695
timestamp 1704896540
transform 1 0 34413 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_696
timestamp 1704896540
transform 1 0 34077 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_697
timestamp 1704896540
transform 1 0 33741 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_698
timestamp 1704896540
transform 1 0 33405 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_699
timestamp 1704896540
transform 1 0 33069 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_700
timestamp 1704896540
transform 1 0 32733 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_701
timestamp 1704896540
transform 1 0 32397 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_702
timestamp 1704896540
transform 1 0 32061 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_703
timestamp 1704896540
transform 1 0 31725 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_704
timestamp 1704896540
transform 1 0 31389 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_705
timestamp 1704896540
transform 1 0 31053 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_706
timestamp 1704896540
transform 1 0 30717 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_707
timestamp 1704896540
transform 1 0 30381 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_708
timestamp 1704896540
transform 1 0 30045 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_709
timestamp 1704896540
transform 1 0 36429 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_710
timestamp 1704896540
transform 1 0 41805 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_711
timestamp 1704896540
transform 1 0 41469 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_712
timestamp 1704896540
transform 1 0 41133 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_713
timestamp 1704896540
transform 1 0 40797 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_714
timestamp 1704896540
transform 1 0 40461 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_715
timestamp 1704896540
transform 1 0 40125 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_716
timestamp 1704896540
transform 1 0 39789 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_717
timestamp 1704896540
transform 1 0 39453 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_718
timestamp 1704896540
transform 1 0 39117 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_719
timestamp 1704896540
transform 1 0 38781 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_720
timestamp 1704896540
transform 1 0 38445 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_721
timestamp 1704896540
transform 1 0 38109 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_722
timestamp 1704896540
transform 1 0 37773 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_723
timestamp 1704896540
transform 1 0 37437 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_724
timestamp 1704896540
transform 1 0 37101 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_725
timestamp 1704896540
transform 1 0 36765 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_726
timestamp 1704896540
transform 1 0 43149 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_727
timestamp 1704896540
transform 1 0 42813 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_728
timestamp 1704896540
transform 1 0 42477 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_729
timestamp 1704896540
transform 1 0 42141 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_730
timestamp 1704896540
transform 1 0 47853 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_731
timestamp 1704896540
transform 1 0 47517 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_732
timestamp 1704896540
transform 1 0 47181 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_733
timestamp 1704896540
transform 1 0 46845 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_734
timestamp 1704896540
transform 1 0 46509 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_735
timestamp 1704896540
transform 1 0 46173 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_736
timestamp 1704896540
transform 1 0 45837 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_737
timestamp 1704896540
transform 1 0 45501 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_738
timestamp 1704896540
transform 1 0 45165 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_739
timestamp 1704896540
transform 1 0 44829 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_740
timestamp 1704896540
transform 1 0 44493 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_741
timestamp 1704896540
transform 1 0 44157 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_742
timestamp 1704896540
transform 1 0 43821 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_743
timestamp 1704896540
transform 1 0 43485 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_744
timestamp 1704896540
transform 1 0 36093 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_745
timestamp 1704896540
transform 1 0 1821 0 1 59467
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_746
timestamp 1704896540
transform 1 0 94179 0 1 46363
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_747
timestamp 1704896540
transform 1 0 94179 0 1 46027
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_748
timestamp 1704896540
transform 1 0 94179 0 1 45691
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_749
timestamp 1704896540
transform 1 0 94179 0 1 45355
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_750
timestamp 1704896540
transform 1 0 94179 0 1 45019
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_751
timestamp 1704896540
transform 1 0 94179 0 1 44683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_752
timestamp 1704896540
transform 1 0 94179 0 1 44347
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_753
timestamp 1704896540
transform 1 0 94179 0 1 44011
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_754
timestamp 1704896540
transform 1 0 94179 0 1 43675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_755
timestamp 1704896540
transform 1 0 94179 0 1 43339
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_756
timestamp 1704896540
transform 1 0 94179 0 1 43003
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_757
timestamp 1704896540
transform 1 0 94179 0 1 42667
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_758
timestamp 1704896540
transform 1 0 94179 0 1 42331
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_759
timestamp 1704896540
transform 1 0 94179 0 1 41995
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_760
timestamp 1704896540
transform 1 0 94179 0 1 41659
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_761
timestamp 1704896540
transform 1 0 94179 0 1 41323
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_762
timestamp 1704896540
transform 1 0 94179 0 1 39979
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_763
timestamp 1704896540
transform 1 0 94179 0 1 40987
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_764
timestamp 1704896540
transform 1 0 94179 0 1 49387
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_765
timestamp 1704896540
transform 1 0 94179 0 1 49051
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_766
timestamp 1704896540
transform 1 0 94179 0 1 48715
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_767
timestamp 1704896540
transform 1 0 94179 0 1 48379
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_768
timestamp 1704896540
transform 1 0 94179 0 1 48043
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_769
timestamp 1704896540
transform 1 0 94179 0 1 47707
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_770
timestamp 1704896540
transform 1 0 94179 0 1 47371
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_771
timestamp 1704896540
transform 1 0 94179 0 1 40651
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_772
timestamp 1704896540
transform 1 0 94179 0 1 40315
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_773
timestamp 1704896540
transform 1 0 94179 0 1 47035
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_774
timestamp 1704896540
transform 1 0 94179 0 1 46699
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_775
timestamp 1704896540
transform 1 0 94179 0 1 50731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_776
timestamp 1704896540
transform 1 0 94179 0 1 50395
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_777
timestamp 1704896540
transform 1 0 94179 0 1 50059
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_778
timestamp 1704896540
transform 1 0 94179 0 1 49723
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_779
timestamp 1704896540
transform 1 0 94179 0 1 54427
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_780
timestamp 1704896540
transform 1 0 94179 0 1 54091
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_781
timestamp 1704896540
transform 1 0 94179 0 1 53755
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_782
timestamp 1704896540
transform 1 0 94179 0 1 53419
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_783
timestamp 1704896540
transform 1 0 94179 0 1 53083
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_784
timestamp 1704896540
transform 1 0 94179 0 1 52747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_785
timestamp 1704896540
transform 1 0 94179 0 1 52411
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_786
timestamp 1704896540
transform 1 0 94179 0 1 52075
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_787
timestamp 1704896540
transform 1 0 94179 0 1 51739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_788
timestamp 1704896540
transform 1 0 94179 0 1 51403
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_789
timestamp 1704896540
transform 1 0 94179 0 1 51067
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_790
timestamp 1704896540
transform 1 0 94179 0 1 55771
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_791
timestamp 1704896540
transform 1 0 94179 0 1 55435
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_792
timestamp 1704896540
transform 1 0 94179 0 1 55099
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_793
timestamp 1704896540
transform 1 0 94179 0 1 54763
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_794
timestamp 1704896540
transform 1 0 94179 0 1 59131
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_795
timestamp 1704896540
transform 1 0 94179 0 1 58795
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_796
timestamp 1704896540
transform 1 0 94179 0 1 58459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_797
timestamp 1704896540
transform 1 0 94179 0 1 58123
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_798
timestamp 1704896540
transform 1 0 94179 0 1 57787
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_799
timestamp 1704896540
transform 1 0 94179 0 1 57451
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_800
timestamp 1704896540
transform 1 0 94179 0 1 57115
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_801
timestamp 1704896540
transform 1 0 94179 0 1 56779
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_802
timestamp 1704896540
transform 1 0 94179 0 1 56443
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_803
timestamp 1704896540
transform 1 0 94179 0 1 56107
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_804
timestamp 1704896540
transform 1 0 48861 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_805
timestamp 1704896540
transform 1 0 48525 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_806
timestamp 1704896540
transform 1 0 48189 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_807
timestamp 1704896540
transform 1 0 53565 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_808
timestamp 1704896540
transform 1 0 53229 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_809
timestamp 1704896540
transform 1 0 52893 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_810
timestamp 1704896540
transform 1 0 52557 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_811
timestamp 1704896540
transform 1 0 52221 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_812
timestamp 1704896540
transform 1 0 51885 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_813
timestamp 1704896540
transform 1 0 51549 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_814
timestamp 1704896540
transform 1 0 51213 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_815
timestamp 1704896540
transform 1 0 50877 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_816
timestamp 1704896540
transform 1 0 50541 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_817
timestamp 1704896540
transform 1 0 50205 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_818
timestamp 1704896540
transform 1 0 49869 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_819
timestamp 1704896540
transform 1 0 49533 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_820
timestamp 1704896540
transform 1 0 49197 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_821
timestamp 1704896540
transform 1 0 59613 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_822
timestamp 1704896540
transform 1 0 59277 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_823
timestamp 1704896540
transform 1 0 58941 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_824
timestamp 1704896540
transform 1 0 58605 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_825
timestamp 1704896540
transform 1 0 58269 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_826
timestamp 1704896540
transform 1 0 57933 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_827
timestamp 1704896540
transform 1 0 57597 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_828
timestamp 1704896540
transform 1 0 57261 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_829
timestamp 1704896540
transform 1 0 56925 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_830
timestamp 1704896540
transform 1 0 56589 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_831
timestamp 1704896540
transform 1 0 56253 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_832
timestamp 1704896540
transform 1 0 55917 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_833
timestamp 1704896540
transform 1 0 55581 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_834
timestamp 1704896540
transform 1 0 55245 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_835
timestamp 1704896540
transform 1 0 54909 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_836
timestamp 1704896540
transform 1 0 54573 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_837
timestamp 1704896540
transform 1 0 54237 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_838
timestamp 1704896540
transform 1 0 53901 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_839
timestamp 1704896540
transform 1 0 62301 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_840
timestamp 1704896540
transform 1 0 61965 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_841
timestamp 1704896540
transform 1 0 61629 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_842
timestamp 1704896540
transform 1 0 61293 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_843
timestamp 1704896540
transform 1 0 60957 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_844
timestamp 1704896540
transform 1 0 60621 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_845
timestamp 1704896540
transform 1 0 60285 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_846
timestamp 1704896540
transform 1 0 62637 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_847
timestamp 1704896540
transform 1 0 64317 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_848
timestamp 1704896540
transform 1 0 63981 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_849
timestamp 1704896540
transform 1 0 65661 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_850
timestamp 1704896540
transform 1 0 65325 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_851
timestamp 1704896540
transform 1 0 64989 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_852
timestamp 1704896540
transform 1 0 64653 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_853
timestamp 1704896540
transform 1 0 63645 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_854
timestamp 1704896540
transform 1 0 63309 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_855
timestamp 1704896540
transform 1 0 62973 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_856
timestamp 1704896540
transform 1 0 71709 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_857
timestamp 1704896540
transform 1 0 71373 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_858
timestamp 1704896540
transform 1 0 71037 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_859
timestamp 1704896540
transform 1 0 70701 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_860
timestamp 1704896540
transform 1 0 70365 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_861
timestamp 1704896540
transform 1 0 70029 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_862
timestamp 1704896540
transform 1 0 69693 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_863
timestamp 1704896540
transform 1 0 69357 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_864
timestamp 1704896540
transform 1 0 69021 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_865
timestamp 1704896540
transform 1 0 68685 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_866
timestamp 1704896540
transform 1 0 68349 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_867
timestamp 1704896540
transform 1 0 68013 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_868
timestamp 1704896540
transform 1 0 67677 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_869
timestamp 1704896540
transform 1 0 67341 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_870
timestamp 1704896540
transform 1 0 67005 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_871
timestamp 1704896540
transform 1 0 66669 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_872
timestamp 1704896540
transform 1 0 66333 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_873
timestamp 1704896540
transform 1 0 65997 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_874
timestamp 1704896540
transform 1 0 59949 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_875
timestamp 1704896540
transform 1 0 94179 0 1 60811
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_876
timestamp 1704896540
transform 1 0 94179 0 1 59803
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_877
timestamp 1704896540
transform 1 0 94179 0 1 64171
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_878
timestamp 1704896540
transform 1 0 94179 0 1 63835
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_879
timestamp 1704896540
transform 1 0 94179 0 1 63499
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_880
timestamp 1704896540
transform 1 0 94179 0 1 63163
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_881
timestamp 1704896540
transform 1 0 94179 0 1 62827
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_882
timestamp 1704896540
transform 1 0 94179 0 1 62491
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_883
timestamp 1704896540
transform 1 0 94179 0 1 62155
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_884
timestamp 1704896540
transform 1 0 94179 0 1 61819
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_885
timestamp 1704896540
transform 1 0 94179 0 1 61483
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_886
timestamp 1704896540
transform 1 0 94179 0 1 60475
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_887
timestamp 1704896540
transform 1 0 94179 0 1 61147
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_888
timestamp 1704896540
transform 1 0 94179 0 1 60139
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_889
timestamp 1704896540
transform 1 0 94179 0 1 69211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_890
timestamp 1704896540
transform 1 0 94179 0 1 68875
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_891
timestamp 1704896540
transform 1 0 94179 0 1 68539
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_892
timestamp 1704896540
transform 1 0 94179 0 1 68203
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_893
timestamp 1704896540
transform 1 0 94179 0 1 67867
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_894
timestamp 1704896540
transform 1 0 94179 0 1 67531
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_895
timestamp 1704896540
transform 1 0 94179 0 1 67195
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_896
timestamp 1704896540
transform 1 0 94179 0 1 66859
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_897
timestamp 1704896540
transform 1 0 94179 0 1 66523
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_898
timestamp 1704896540
transform 1 0 94179 0 1 66187
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_899
timestamp 1704896540
transform 1 0 94179 0 1 65851
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_900
timestamp 1704896540
transform 1 0 94179 0 1 65515
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_901
timestamp 1704896540
transform 1 0 94179 0 1 65179
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_902
timestamp 1704896540
transform 1 0 94179 0 1 64843
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_903
timestamp 1704896540
transform 1 0 94179 0 1 64507
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_904
timestamp 1704896540
transform 1 0 76749 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_905
timestamp 1704896540
transform 1 0 72381 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_906
timestamp 1704896540
transform 1 0 76077 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_907
timestamp 1704896540
transform 1 0 75741 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_908
timestamp 1704896540
transform 1 0 75405 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_909
timestamp 1704896540
transform 1 0 75069 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_910
timestamp 1704896540
transform 1 0 74733 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_911
timestamp 1704896540
transform 1 0 74397 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_912
timestamp 1704896540
transform 1 0 74061 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_913
timestamp 1704896540
transform 1 0 73725 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_914
timestamp 1704896540
transform 1 0 73389 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_915
timestamp 1704896540
transform 1 0 72717 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_916
timestamp 1704896540
transform 1 0 76413 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_917
timestamp 1704896540
transform 1 0 77421 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_918
timestamp 1704896540
transform 1 0 77085 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_919
timestamp 1704896540
transform 1 0 73053 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_920
timestamp 1704896540
transform 1 0 72045 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_921
timestamp 1704896540
transform 1 0 83469 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_922
timestamp 1704896540
transform 1 0 83133 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_923
timestamp 1704896540
transform 1 0 82797 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_924
timestamp 1704896540
transform 1 0 78093 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_925
timestamp 1704896540
transform 1 0 82461 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_926
timestamp 1704896540
transform 1 0 82125 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_927
timestamp 1704896540
transform 1 0 81789 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_928
timestamp 1704896540
transform 1 0 81453 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_929
timestamp 1704896540
transform 1 0 81117 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_930
timestamp 1704896540
transform 1 0 80781 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_931
timestamp 1704896540
transform 1 0 80445 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_932
timestamp 1704896540
transform 1 0 80109 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_933
timestamp 1704896540
transform 1 0 79773 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_934
timestamp 1704896540
transform 1 0 79437 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_935
timestamp 1704896540
transform 1 0 79101 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_936
timestamp 1704896540
transform 1 0 78765 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_937
timestamp 1704896540
transform 1 0 78429 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_938
timestamp 1704896540
transform 1 0 77757 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_939
timestamp 1704896540
transform 1 0 94179 0 1 71899
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_940
timestamp 1704896540
transform 1 0 94179 0 1 71563
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_941
timestamp 1704896540
transform 1 0 94179 0 1 71227
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_942
timestamp 1704896540
transform 1 0 94179 0 1 70891
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_943
timestamp 1704896540
transform 1 0 94179 0 1 70555
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_944
timestamp 1704896540
transform 1 0 94179 0 1 70219
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_945
timestamp 1704896540
transform 1 0 94179 0 1 69883
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_946
timestamp 1704896540
transform 1 0 94179 0 1 69547
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_947
timestamp 1704896540
transform 1 0 94179 0 1 73915
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_948
timestamp 1704896540
transform 1 0 94179 0 1 73579
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_949
timestamp 1704896540
transform 1 0 94179 0 1 73243
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_950
timestamp 1704896540
transform 1 0 94179 0 1 72907
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_951
timestamp 1704896540
transform 1 0 94179 0 1 72571
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_952
timestamp 1704896540
transform 1 0 94179 0 1 72235
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_953
timestamp 1704896540
transform 1 0 84141 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_954
timestamp 1704896540
transform 1 0 84813 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_955
timestamp 1704896540
transform 1 0 84477 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_956
timestamp 1704896540
transform 1 0 89517 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_957
timestamp 1704896540
transform 1 0 89181 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_958
timestamp 1704896540
transform 1 0 88845 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_959
timestamp 1704896540
transform 1 0 88509 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_960
timestamp 1704896540
transform 1 0 88173 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_961
timestamp 1704896540
transform 1 0 87837 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_962
timestamp 1704896540
transform 1 0 87501 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_963
timestamp 1704896540
transform 1 0 87165 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_964
timestamp 1704896540
transform 1 0 86829 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_965
timestamp 1704896540
transform 1 0 86493 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_966
timestamp 1704896540
transform 1 0 86157 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_967
timestamp 1704896540
transform 1 0 85821 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_968
timestamp 1704896540
transform 1 0 85485 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_969
timestamp 1704896540
transform 1 0 85149 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_970
timestamp 1704896540
transform 1 0 90525 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_971
timestamp 1704896540
transform 1 0 94179 0 1 77275
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_972
timestamp 1704896540
transform 1 0 94179 0 1 76939
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_973
timestamp 1704896540
transform 1 0 94179 0 1 76603
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_974
timestamp 1704896540
transform 1 0 94179 0 1 76267
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_975
timestamp 1704896540
transform 1 0 94179 0 1 75931
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_976
timestamp 1704896540
transform 1 0 94179 0 1 75595
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_977
timestamp 1704896540
transform 1 0 94179 0 1 75259
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_978
timestamp 1704896540
transform 1 0 94179 0 1 74923
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_979
timestamp 1704896540
transform 1 0 94179 0 1 74587
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_980
timestamp 1704896540
transform 1 0 90189 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_981
timestamp 1704896540
transform 1 0 89853 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_982
timestamp 1704896540
transform 1 0 93549 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_983
timestamp 1704896540
transform 1 0 93213 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_984
timestamp 1704896540
transform 1 0 92877 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_985
timestamp 1704896540
transform 1 0 92541 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_986
timestamp 1704896540
transform 1 0 92205 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_987
timestamp 1704896540
transform 1 0 91869 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_988
timestamp 1704896540
transform 1 0 91533 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_989
timestamp 1704896540
transform 1 0 91197 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_990
timestamp 1704896540
transform 1 0 90861 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_991
timestamp 1704896540
transform 1 0 94179 0 1 74251
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_992
timestamp 1704896540
transform 1 0 83805 0 1 77739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_993
timestamp 1704896540
transform 1 0 94179 0 1 59467
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_994
timestamp 1704896540
transform 1 0 94179 0 1 39643
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_13  sky130_sram_1kbyte_1rw1r_32x256_8_contact_13_995
timestamp 1704896540
transform 1 0 1821 0 1 39643
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_0
timestamp 1704896540
transform 1 0 92201 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_1
timestamp 1704896540
transform 1 0 94175 0 1 4707
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_2
timestamp 1704896540
transform 1 0 94175 0 1 4371
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_3
timestamp 1704896540
transform 1 0 90857 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_4
timestamp 1704896540
transform 1 0 91865 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_5
timestamp 1704896540
transform 1 0 91529 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_6
timestamp 1704896540
transform 1 0 94175 0 1 4035
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_7
timestamp 1704896540
transform 1 0 94175 0 1 3699
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_8
timestamp 1704896540
transform 1 0 94175 0 1 3363
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_9
timestamp 1704896540
transform 1 0 94175 0 1 3027
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_10
timestamp 1704896540
transform 1 0 94175 0 1 2691
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_11
timestamp 1704896540
transform 1 0 94175 0 1 2355
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_12
timestamp 1704896540
transform 1 0 92537 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_13
timestamp 1704896540
transform 1 0 91193 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_14
timestamp 1704896540
transform 1 0 94175 0 1 2019
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_15
timestamp 1704896540
transform 1 0 94175 0 1 5043
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_16
timestamp 1704896540
transform 1 0 90521 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_17
timestamp 1704896540
transform 1 0 90185 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_18
timestamp 1704896540
transform 1 0 92873 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_19
timestamp 1704896540
transform 1 0 89849 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_20
timestamp 1704896540
transform 1 0 93545 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_21
timestamp 1704896540
transform 1 0 93209 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_22
timestamp 1704896540
transform 1 0 84473 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_23
timestamp 1704896540
transform 1 0 84137 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_24
timestamp 1704896540
transform 1 0 89177 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_25
timestamp 1704896540
transform 1 0 88841 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_26
timestamp 1704896540
transform 1 0 88505 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_27
timestamp 1704896540
transform 1 0 88169 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_28
timestamp 1704896540
transform 1 0 87833 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_29
timestamp 1704896540
transform 1 0 87497 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_30
timestamp 1704896540
transform 1 0 87161 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_31
timestamp 1704896540
transform 1 0 86825 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_32
timestamp 1704896540
transform 1 0 86489 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_33
timestamp 1704896540
transform 1 0 86153 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_34
timestamp 1704896540
transform 1 0 83801 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_35
timestamp 1704896540
transform 1 0 85817 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_36
timestamp 1704896540
transform 1 0 85481 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_37
timestamp 1704896540
transform 1 0 89513 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_38
timestamp 1704896540
transform 1 0 85145 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_39
timestamp 1704896540
transform 1 0 84809 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_40
timestamp 1704896540
transform 1 0 94175 0 1 7395
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_41
timestamp 1704896540
transform 1 0 94175 0 1 7059
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_42
timestamp 1704896540
transform 1 0 94175 0 1 6723
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_43
timestamp 1704896540
transform 1 0 94175 0 1 5715
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_44
timestamp 1704896540
transform 1 0 94175 0 1 5379
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_45
timestamp 1704896540
transform 1 0 94175 0 1 6387
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_46
timestamp 1704896540
transform 1 0 94175 0 1 6051
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_47
timestamp 1704896540
transform 1 0 94175 0 1 9747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_48
timestamp 1704896540
transform 1 0 94175 0 1 9411
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_49
timestamp 1704896540
transform 1 0 94175 0 1 9075
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_50
timestamp 1704896540
transform 1 0 94175 0 1 8739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_51
timestamp 1704896540
transform 1 0 94175 0 1 8403
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_52
timestamp 1704896540
transform 1 0 94175 0 1 8067
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_53
timestamp 1704896540
transform 1 0 94175 0 1 7731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_54
timestamp 1704896540
transform 1 0 78425 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_55
timestamp 1704896540
transform 1 0 82121 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_56
timestamp 1704896540
transform 1 0 81785 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_57
timestamp 1704896540
transform 1 0 81449 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_58
timestamp 1704896540
transform 1 0 81113 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_59
timestamp 1704896540
transform 1 0 80777 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_60
timestamp 1704896540
transform 1 0 80441 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_61
timestamp 1704896540
transform 1 0 80105 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_62
timestamp 1704896540
transform 1 0 79769 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_63
timestamp 1704896540
transform 1 0 83129 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_64
timestamp 1704896540
transform 1 0 78089 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_65
timestamp 1704896540
transform 1 0 82457 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_66
timestamp 1704896540
transform 1 0 79433 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_67
timestamp 1704896540
transform 1 0 79097 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_68
timestamp 1704896540
transform 1 0 83465 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_69
timestamp 1704896540
transform 1 0 78761 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_70
timestamp 1704896540
transform 1 0 82793 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_71
timestamp 1704896540
transform 1 0 72041 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_72
timestamp 1704896540
transform 1 0 76073 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_73
timestamp 1704896540
transform 1 0 75737 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_74
timestamp 1704896540
transform 1 0 75401 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_75
timestamp 1704896540
transform 1 0 73049 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_76
timestamp 1704896540
transform 1 0 72713 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_77
timestamp 1704896540
transform 1 0 77081 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_78
timestamp 1704896540
transform 1 0 74057 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_79
timestamp 1704896540
transform 1 0 76745 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_80
timestamp 1704896540
transform 1 0 73721 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_81
timestamp 1704896540
transform 1 0 75065 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_82
timestamp 1704896540
transform 1 0 74729 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_83
timestamp 1704896540
transform 1 0 72377 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_84
timestamp 1704896540
transform 1 0 73385 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_85
timestamp 1704896540
transform 1 0 76409 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_86
timestamp 1704896540
transform 1 0 77417 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_87
timestamp 1704896540
transform 1 0 74393 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_88
timestamp 1704896540
transform 1 0 77753 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_89
timestamp 1704896540
transform 1 0 94175 0 1 19827
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_90
timestamp 1704896540
transform 1 0 94175 0 1 19491
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_91
timestamp 1704896540
transform 1 0 94175 0 1 19155
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_92
timestamp 1704896540
transform 1 0 94175 0 1 18819
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_93
timestamp 1704896540
transform 1 0 94175 0 1 18483
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_94
timestamp 1704896540
transform 1 0 94175 0 1 18147
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_95
timestamp 1704896540
transform 1 0 94175 0 1 17811
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_96
timestamp 1704896540
transform 1 0 94175 0 1 17475
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_97
timestamp 1704896540
transform 1 0 94175 0 1 17139
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_98
timestamp 1704896540
transform 1 0 94175 0 1 16803
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_99
timestamp 1704896540
transform 1 0 94175 0 1 16467
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_100
timestamp 1704896540
transform 1 0 94175 0 1 16131
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_101
timestamp 1704896540
transform 1 0 94175 0 1 15795
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_102
timestamp 1704896540
transform 1 0 94175 0 1 15459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_103
timestamp 1704896540
transform 1 0 94175 0 1 15123
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_104
timestamp 1704896540
transform 1 0 94175 0 1 14787
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_105
timestamp 1704896540
transform 1 0 94175 0 1 14451
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_106
timestamp 1704896540
transform 1 0 94175 0 1 14115
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_107
timestamp 1704896540
transform 1 0 94175 0 1 13779
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_108
timestamp 1704896540
transform 1 0 94175 0 1 13443
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_109
timestamp 1704896540
transform 1 0 94175 0 1 13107
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_110
timestamp 1704896540
transform 1 0 94175 0 1 12771
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_111
timestamp 1704896540
transform 1 0 94175 0 1 12435
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_112
timestamp 1704896540
transform 1 0 94175 0 1 12099
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_113
timestamp 1704896540
transform 1 0 94175 0 1 11763
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_114
timestamp 1704896540
transform 1 0 94175 0 1 11427
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_115
timestamp 1704896540
transform 1 0 94175 0 1 11091
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_116
timestamp 1704896540
transform 1 0 94175 0 1 10755
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_117
timestamp 1704896540
transform 1 0 94175 0 1 10419
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_118
timestamp 1704896540
transform 1 0 94175 0 1 10083
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_119
timestamp 1704896540
transform 1 0 65993 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_120
timestamp 1704896540
transform 1 0 68009 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_121
timestamp 1704896540
transform 1 0 68345 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_122
timestamp 1704896540
transform 1 0 69689 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_123
timestamp 1704896540
transform 1 0 67673 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_124
timestamp 1704896540
transform 1 0 67337 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_125
timestamp 1704896540
transform 1 0 66329 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_126
timestamp 1704896540
transform 1 0 71033 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_127
timestamp 1704896540
transform 1 0 69017 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_128
timestamp 1704896540
transform 1 0 70697 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_129
timestamp 1704896540
transform 1 0 71705 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_130
timestamp 1704896540
transform 1 0 68681 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_131
timestamp 1704896540
transform 1 0 67001 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_132
timestamp 1704896540
transform 1 0 69353 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_133
timestamp 1704896540
transform 1 0 71369 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_134
timestamp 1704896540
transform 1 0 70361 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_135
timestamp 1704896540
transform 1 0 70025 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_136
timestamp 1704896540
transform 1 0 66665 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_137
timestamp 1704896540
transform 1 0 65657 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_138
timestamp 1704896540
transform 1 0 65321 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_139
timestamp 1704896540
transform 1 0 64985 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_140
timestamp 1704896540
transform 1 0 64649 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_141
timestamp 1704896540
transform 1 0 59945 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_142
timestamp 1704896540
transform 1 0 62633 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_143
timestamp 1704896540
transform 1 0 63977 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_144
timestamp 1704896540
transform 1 0 63641 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_145
timestamp 1704896540
transform 1 0 63305 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_146
timestamp 1704896540
transform 1 0 62969 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_147
timestamp 1704896540
transform 1 0 64313 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_148
timestamp 1704896540
transform 1 0 62297 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_149
timestamp 1704896540
transform 1 0 61961 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_150
timestamp 1704896540
transform 1 0 61625 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_151
timestamp 1704896540
transform 1 0 61289 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_152
timestamp 1704896540
transform 1 0 60953 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_153
timestamp 1704896540
transform 1 0 60617 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_154
timestamp 1704896540
transform 1 0 60281 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_155
timestamp 1704896540
transform 1 0 55241 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_156
timestamp 1704896540
transform 1 0 54233 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_157
timestamp 1704896540
transform 1 0 59609 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_158
timestamp 1704896540
transform 1 0 54905 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_159
timestamp 1704896540
transform 1 0 59273 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_160
timestamp 1704896540
transform 1 0 58937 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_161
timestamp 1704896540
transform 1 0 58601 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_162
timestamp 1704896540
transform 1 0 58265 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_163
timestamp 1704896540
transform 1 0 57929 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_164
timestamp 1704896540
transform 1 0 54569 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_165
timestamp 1704896540
transform 1 0 57593 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_166
timestamp 1704896540
transform 1 0 57257 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_167
timestamp 1704896540
transform 1 0 56921 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_168
timestamp 1704896540
transform 1 0 56585 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_169
timestamp 1704896540
transform 1 0 56249 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_170
timestamp 1704896540
transform 1 0 55913 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_171
timestamp 1704896540
transform 1 0 55577 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_172
timestamp 1704896540
transform 1 0 48521 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_173
timestamp 1704896540
transform 1 0 50873 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_174
timestamp 1704896540
transform 1 0 50537 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_175
timestamp 1704896540
transform 1 0 50201 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_176
timestamp 1704896540
transform 1 0 52217 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_177
timestamp 1704896540
transform 1 0 51209 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_178
timestamp 1704896540
transform 1 0 49193 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_179
timestamp 1704896540
transform 1 0 49865 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_180
timestamp 1704896540
transform 1 0 51881 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_181
timestamp 1704896540
transform 1 0 51545 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_182
timestamp 1704896540
transform 1 0 53561 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_183
timestamp 1704896540
transform 1 0 49529 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_184
timestamp 1704896540
transform 1 0 48857 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_185
timestamp 1704896540
transform 1 0 53225 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_186
timestamp 1704896540
transform 1 0 52889 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_187
timestamp 1704896540
transform 1 0 48185 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_188
timestamp 1704896540
transform 1 0 52553 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_189
timestamp 1704896540
transform 1 0 53897 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_190
timestamp 1704896540
transform 1 0 94175 0 1 23187
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_191
timestamp 1704896540
transform 1 0 94175 0 1 22851
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_192
timestamp 1704896540
transform 1 0 94175 0 1 22515
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_193
timestamp 1704896540
transform 1 0 94175 0 1 22179
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_194
timestamp 1704896540
transform 1 0 94175 0 1 21843
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_195
timestamp 1704896540
transform 1 0 94175 0 1 29571
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_196
timestamp 1704896540
transform 1 0 94175 0 1 21507
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_197
timestamp 1704896540
transform 1 0 94175 0 1 29235
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_198
timestamp 1704896540
transform 1 0 94175 0 1 28899
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_199
timestamp 1704896540
transform 1 0 94175 0 1 21171
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_200
timestamp 1704896540
transform 1 0 94175 0 1 20835
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_201
timestamp 1704896540
transform 1 0 94175 0 1 28563
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_202
timestamp 1704896540
transform 1 0 94175 0 1 20499
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_203
timestamp 1704896540
transform 1 0 94175 0 1 20163
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_204
timestamp 1704896540
transform 1 0 94175 0 1 28227
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_205
timestamp 1704896540
transform 1 0 94175 0 1 27891
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_206
timestamp 1704896540
transform 1 0 94175 0 1 27555
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_207
timestamp 1704896540
transform 1 0 94175 0 1 27219
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_208
timestamp 1704896540
transform 1 0 94175 0 1 26883
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_209
timestamp 1704896540
transform 1 0 94175 0 1 26547
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_210
timestamp 1704896540
transform 1 0 94175 0 1 26211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_211
timestamp 1704896540
transform 1 0 94175 0 1 25875
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_212
timestamp 1704896540
transform 1 0 94175 0 1 25539
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_213
timestamp 1704896540
transform 1 0 94175 0 1 25203
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_214
timestamp 1704896540
transform 1 0 94175 0 1 24867
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_215
timestamp 1704896540
transform 1 0 94175 0 1 24531
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_216
timestamp 1704896540
transform 1 0 94175 0 1 24195
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_217
timestamp 1704896540
transform 1 0 94175 0 1 23859
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_218
timestamp 1704896540
transform 1 0 94175 0 1 23523
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_219
timestamp 1704896540
transform 1 0 94175 0 1 39651
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_220
timestamp 1704896540
transform 1 0 94175 0 1 39315
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_221
timestamp 1704896540
transform 1 0 94175 0 1 38979
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_222
timestamp 1704896540
transform 1 0 94175 0 1 38643
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_223
timestamp 1704896540
transform 1 0 94175 0 1 38307
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_224
timestamp 1704896540
transform 1 0 94175 0 1 37971
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_225
timestamp 1704896540
transform 1 0 94175 0 1 37635
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_226
timestamp 1704896540
transform 1 0 94175 0 1 37299
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_227
timestamp 1704896540
transform 1 0 94175 0 1 36963
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_228
timestamp 1704896540
transform 1 0 94175 0 1 36627
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_229
timestamp 1704896540
transform 1 0 94175 0 1 36291
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_230
timestamp 1704896540
transform 1 0 94175 0 1 35955
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_231
timestamp 1704896540
transform 1 0 94175 0 1 35619
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_232
timestamp 1704896540
transform 1 0 94175 0 1 35283
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_233
timestamp 1704896540
transform 1 0 94175 0 1 34947
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_234
timestamp 1704896540
transform 1 0 94175 0 1 34611
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_235
timestamp 1704896540
transform 1 0 94175 0 1 34275
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_236
timestamp 1704896540
transform 1 0 94175 0 1 33939
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_237
timestamp 1704896540
transform 1 0 94175 0 1 33603
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_238
timestamp 1704896540
transform 1 0 94175 0 1 33267
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_239
timestamp 1704896540
transform 1 0 94175 0 1 32931
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_240
timestamp 1704896540
transform 1 0 94175 0 1 32595
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_241
timestamp 1704896540
transform 1 0 94175 0 1 32259
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_242
timestamp 1704896540
transform 1 0 94175 0 1 31923
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_243
timestamp 1704896540
transform 1 0 94175 0 1 31587
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_244
timestamp 1704896540
transform 1 0 94175 0 1 31251
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_245
timestamp 1704896540
transform 1 0 94175 0 1 30915
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_246
timestamp 1704896540
transform 1 0 94175 0 1 30579
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_247
timestamp 1704896540
transform 1 0 94175 0 1 30243
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_248
timestamp 1704896540
transform 1 0 94175 0 1 29907
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_249
timestamp 1704896540
transform 1 0 45161 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_250
timestamp 1704896540
transform 1 0 44825 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_251
timestamp 1704896540
transform 1 0 44489 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_252
timestamp 1704896540
transform 1 0 42137 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_253
timestamp 1704896540
transform 1 0 44153 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_254
timestamp 1704896540
transform 1 0 43817 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_255
timestamp 1704896540
transform 1 0 47849 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_256
timestamp 1704896540
transform 1 0 47513 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_257
timestamp 1704896540
transform 1 0 47177 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_258
timestamp 1704896540
transform 1 0 46841 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_259
timestamp 1704896540
transform 1 0 46505 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_260
timestamp 1704896540
transform 1 0 46169 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_261
timestamp 1704896540
transform 1 0 43481 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_262
timestamp 1704896540
transform 1 0 43145 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_263
timestamp 1704896540
transform 1 0 45833 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_264
timestamp 1704896540
transform 1 0 45497 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_265
timestamp 1704896540
transform 1 0 42809 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_266
timestamp 1704896540
transform 1 0 42473 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_267
timestamp 1704896540
transform 1 0 36089 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_268
timestamp 1704896540
transform 1 0 38105 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_269
timestamp 1704896540
transform 1 0 37769 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_270
timestamp 1704896540
transform 1 0 37433 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_271
timestamp 1704896540
transform 1 0 40793 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_272
timestamp 1704896540
transform 1 0 40457 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_273
timestamp 1704896540
transform 1 0 40121 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_274
timestamp 1704896540
transform 1 0 39785 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_275
timestamp 1704896540
transform 1 0 39449 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_276
timestamp 1704896540
transform 1 0 39113 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_277
timestamp 1704896540
transform 1 0 37097 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_278
timestamp 1704896540
transform 1 0 36761 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_279
timestamp 1704896540
transform 1 0 36425 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_280
timestamp 1704896540
transform 1 0 41801 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_281
timestamp 1704896540
transform 1 0 38777 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_282
timestamp 1704896540
transform 1 0 38441 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_283
timestamp 1704896540
transform 1 0 41465 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_284
timestamp 1704896540
transform 1 0 41129 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_285
timestamp 1704896540
transform 1 0 30713 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_286
timestamp 1704896540
transform 1 0 32729 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_287
timestamp 1704896540
transform 1 0 32393 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_288
timestamp 1704896540
transform 1 0 35753 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_289
timestamp 1704896540
transform 1 0 32057 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_290
timestamp 1704896540
transform 1 0 31721 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_291
timestamp 1704896540
transform 1 0 35417 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_292
timestamp 1704896540
transform 1 0 35081 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_293
timestamp 1704896540
transform 1 0 31385 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_294
timestamp 1704896540
transform 1 0 34745 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_295
timestamp 1704896540
transform 1 0 34409 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_296
timestamp 1704896540
transform 1 0 30377 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_297
timestamp 1704896540
transform 1 0 31049 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_298
timestamp 1704896540
transform 1 0 34073 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_299
timestamp 1704896540
transform 1 0 33737 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_300
timestamp 1704896540
transform 1 0 33401 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_301
timestamp 1704896540
transform 1 0 33065 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_302
timestamp 1704896540
transform 1 0 28361 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_303
timestamp 1704896540
transform 1 0 28025 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_304
timestamp 1704896540
transform 1 0 25001 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_305
timestamp 1704896540
transform 1 0 27689 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_306
timestamp 1704896540
transform 1 0 26009 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_307
timestamp 1704896540
transform 1 0 24665 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_308
timestamp 1704896540
transform 1 0 27353 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_309
timestamp 1704896540
transform 1 0 25673 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_310
timestamp 1704896540
transform 1 0 25337 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_311
timestamp 1704896540
transform 1 0 28697 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_312
timestamp 1704896540
transform 1 0 29705 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_313
timestamp 1704896540
transform 1 0 24329 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_314
timestamp 1704896540
transform 1 0 27017 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_315
timestamp 1704896540
transform 1 0 29369 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_316
timestamp 1704896540
transform 1 0 29033 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_317
timestamp 1704896540
transform 1 0 26681 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_318
timestamp 1704896540
transform 1 0 26345 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_319
timestamp 1704896540
transform 1 0 30041 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_320
timestamp 1704896540
transform 1 0 21305 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_321
timestamp 1704896540
transform 1 0 21641 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_322
timestamp 1704896540
transform 1 0 18281 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_323
timestamp 1704896540
transform 1 0 20969 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_324
timestamp 1704896540
transform 1 0 22313 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_325
timestamp 1704896540
transform 1 0 19289 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_326
timestamp 1704896540
transform 1 0 21977 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_327
timestamp 1704896540
transform 1 0 18953 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_328
timestamp 1704896540
transform 1 0 23993 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_329
timestamp 1704896540
transform 1 0 19961 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_330
timestamp 1704896540
transform 1 0 23657 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_331
timestamp 1704896540
transform 1 0 23321 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_332
timestamp 1704896540
transform 1 0 19625 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_333
timestamp 1704896540
transform 1 0 20297 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_334
timestamp 1704896540
transform 1 0 22985 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_335
timestamp 1704896540
transform 1 0 20633 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_336
timestamp 1704896540
transform 1 0 18617 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_337
timestamp 1704896540
transform 1 0 22649 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_338
timestamp 1704896540
transform 1 0 13241 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_339
timestamp 1704896540
transform 1 0 12905 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_340
timestamp 1704896540
transform 1 0 12569 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_341
timestamp 1704896540
transform 1 0 12233 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_342
timestamp 1704896540
transform 1 0 14249 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_343
timestamp 1704896540
transform 1 0 17945 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_344
timestamp 1704896540
transform 1 0 17609 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_345
timestamp 1704896540
transform 1 0 17273 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_346
timestamp 1704896540
transform 1 0 13913 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_347
timestamp 1704896540
transform 1 0 13577 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_348
timestamp 1704896540
transform 1 0 16937 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_349
timestamp 1704896540
transform 1 0 16601 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_350
timestamp 1704896540
transform 1 0 16265 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_351
timestamp 1704896540
transform 1 0 15929 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_352
timestamp 1704896540
transform 1 0 15593 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_353
timestamp 1704896540
transform 1 0 15257 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_354
timestamp 1704896540
transform 1 0 14921 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_355
timestamp 1704896540
transform 1 0 14585 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_356
timestamp 1704896540
transform 1 0 7193 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_357
timestamp 1704896540
transform 1 0 6857 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_358
timestamp 1704896540
transform 1 0 6521 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_359
timestamp 1704896540
transform 1 0 11897 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_360
timestamp 1704896540
transform 1 0 11561 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_361
timestamp 1704896540
transform 1 0 11225 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_362
timestamp 1704896540
transform 1 0 10889 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_363
timestamp 1704896540
transform 1 0 10553 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_364
timestamp 1704896540
transform 1 0 10217 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_365
timestamp 1704896540
transform 1 0 9881 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_366
timestamp 1704896540
transform 1 0 9545 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_367
timestamp 1704896540
transform 1 0 9209 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_368
timestamp 1704896540
transform 1 0 8873 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_369
timestamp 1704896540
transform 1 0 8537 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_370
timestamp 1704896540
transform 1 0 8201 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_371
timestamp 1704896540
transform 1 0 7865 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_372
timestamp 1704896540
transform 1 0 7529 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_373
timestamp 1704896540
transform 1 0 1817 0 1 2019
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_374
timestamp 1704896540
transform 1 0 3497 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_375
timestamp 1704896540
transform 1 0 3161 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_376
timestamp 1704896540
transform 1 0 2825 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_377
timestamp 1704896540
transform 1 0 2489 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_378
timestamp 1704896540
transform 1 0 5849 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_379
timestamp 1704896540
transform 1 0 2153 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_380
timestamp 1704896540
transform 1 0 1817 0 1 5043
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_381
timestamp 1704896540
transform 1 0 5513 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_382
timestamp 1704896540
transform 1 0 1817 0 1 4707
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_383
timestamp 1704896540
transform 1 0 1817 0 1 4371
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_384
timestamp 1704896540
transform 1 0 1817 0 1 4035
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_385
timestamp 1704896540
transform 1 0 1817 0 1 3699
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_386
timestamp 1704896540
transform 1 0 1817 0 1 3363
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_387
timestamp 1704896540
transform 1 0 5177 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_388
timestamp 1704896540
transform 1 0 4841 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_389
timestamp 1704896540
transform 1 0 4505 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_390
timestamp 1704896540
transform 1 0 1817 0 1 3027
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_391
timestamp 1704896540
transform 1 0 1817 0 1 2691
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_392
timestamp 1704896540
transform 1 0 1817 0 1 2355
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_393
timestamp 1704896540
transform 1 0 4169 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_394
timestamp 1704896540
transform 1 0 3833 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_395
timestamp 1704896540
transform 1 0 1817 0 1 7059
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_396
timestamp 1704896540
transform 1 0 1817 0 1 6723
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_397
timestamp 1704896540
transform 1 0 1817 0 1 6387
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_398
timestamp 1704896540
transform 1 0 1817 0 1 6051
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_399
timestamp 1704896540
transform 1 0 1817 0 1 5715
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_400
timestamp 1704896540
transform 1 0 1817 0 1 9411
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_401
timestamp 1704896540
transform 1 0 1817 0 1 5379
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_402
timestamp 1704896540
transform 1 0 1817 0 1 9075
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_403
timestamp 1704896540
transform 1 0 1817 0 1 8739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_404
timestamp 1704896540
transform 1 0 1817 0 1 8403
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_405
timestamp 1704896540
transform 1 0 1817 0 1 7731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_406
timestamp 1704896540
transform 1 0 1817 0 1 7395
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_407
timestamp 1704896540
transform 1 0 1817 0 1 8067
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_408
timestamp 1704896540
transform 1 0 1817 0 1 9747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_409
timestamp 1704896540
transform 1 0 6185 0 1 1683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_410
timestamp 1704896540
transform 1 0 1817 0 1 13443
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_411
timestamp 1704896540
transform 1 0 1817 0 1 13107
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_412
timestamp 1704896540
transform 1 0 1817 0 1 12771
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_413
timestamp 1704896540
transform 1 0 1817 0 1 12435
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_414
timestamp 1704896540
transform 1 0 1817 0 1 12099
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_415
timestamp 1704896540
transform 1 0 1817 0 1 11763
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_416
timestamp 1704896540
transform 1 0 1817 0 1 11427
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_417
timestamp 1704896540
transform 1 0 1817 0 1 10755
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_418
timestamp 1704896540
transform 1 0 1817 0 1 11091
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_419
timestamp 1704896540
transform 1 0 1817 0 1 14787
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_420
timestamp 1704896540
transform 1 0 1817 0 1 14451
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_421
timestamp 1704896540
transform 1 0 1817 0 1 10419
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_422
timestamp 1704896540
transform 1 0 1817 0 1 14115
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_423
timestamp 1704896540
transform 1 0 1817 0 1 13779
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_424
timestamp 1704896540
transform 1 0 1817 0 1 17811
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_425
timestamp 1704896540
transform 1 0 1817 0 1 17475
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_426
timestamp 1704896540
transform 1 0 1817 0 1 17139
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_427
timestamp 1704896540
transform 1 0 1817 0 1 16803
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_428
timestamp 1704896540
transform 1 0 1817 0 1 16467
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_429
timestamp 1704896540
transform 1 0 1817 0 1 16131
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_430
timestamp 1704896540
transform 1 0 1817 0 1 15795
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_431
timestamp 1704896540
transform 1 0 1817 0 1 15459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_432
timestamp 1704896540
transform 1 0 1817 0 1 15123
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_433
timestamp 1704896540
transform 1 0 1817 0 1 19827
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_434
timestamp 1704896540
transform 1 0 1817 0 1 19491
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_435
timestamp 1704896540
transform 1 0 1817 0 1 19155
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_436
timestamp 1704896540
transform 1 0 1817 0 1 18819
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_437
timestamp 1704896540
transform 1 0 1817 0 1 18483
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_438
timestamp 1704896540
transform 1 0 1817 0 1 18147
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_439
timestamp 1704896540
transform 1 0 1817 0 1 10083
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_440
timestamp 1704896540
transform 1 0 1817 0 1 22179
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_441
timestamp 1704896540
transform 1 0 1817 0 1 20163
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_442
timestamp 1704896540
transform 1 0 1817 0 1 21843
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_443
timestamp 1704896540
transform 1 0 1817 0 1 21507
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_444
timestamp 1704896540
transform 1 0 1817 0 1 21171
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_445
timestamp 1704896540
transform 1 0 1817 0 1 20835
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_446
timestamp 1704896540
transform 1 0 1817 0 1 20499
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_447
timestamp 1704896540
transform 1 0 1817 0 1 24867
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_448
timestamp 1704896540
transform 1 0 1817 0 1 24531
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_449
timestamp 1704896540
transform 1 0 1817 0 1 24195
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_450
timestamp 1704896540
transform 1 0 1817 0 1 23859
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_451
timestamp 1704896540
transform 1 0 1817 0 1 23523
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_452
timestamp 1704896540
transform 1 0 1817 0 1 23187
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_453
timestamp 1704896540
transform 1 0 1817 0 1 22851
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_454
timestamp 1704896540
transform 1 0 1817 0 1 22515
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_455
timestamp 1704896540
transform 1 0 1817 0 1 27219
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_456
timestamp 1704896540
transform 1 0 1817 0 1 26883
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_457
timestamp 1704896540
transform 1 0 1817 0 1 26547
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_458
timestamp 1704896540
transform 1 0 1817 0 1 26211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_459
timestamp 1704896540
transform 1 0 1817 0 1 25875
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_460
timestamp 1704896540
transform 1 0 1817 0 1 25539
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_461
timestamp 1704896540
transform 1 0 1817 0 1 25203
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_462
timestamp 1704896540
transform 1 0 1817 0 1 29571
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_463
timestamp 1704896540
transform 1 0 1817 0 1 29235
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_464
timestamp 1704896540
transform 1 0 1817 0 1 28899
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_465
timestamp 1704896540
transform 1 0 1817 0 1 28563
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_466
timestamp 1704896540
transform 1 0 1817 0 1 28227
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_467
timestamp 1704896540
transform 1 0 1817 0 1 27891
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_468
timestamp 1704896540
transform 1 0 1817 0 1 27555
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_469
timestamp 1704896540
transform 1 0 1817 0 1 30243
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_470
timestamp 1704896540
transform 1 0 1817 0 1 35955
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_471
timestamp 1704896540
transform 1 0 1817 0 1 29907
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_472
timestamp 1704896540
transform 1 0 1817 0 1 35619
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_473
timestamp 1704896540
transform 1 0 1817 0 1 35283
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_474
timestamp 1704896540
transform 1 0 1817 0 1 34947
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_475
timestamp 1704896540
transform 1 0 1817 0 1 34611
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_476
timestamp 1704896540
transform 1 0 1817 0 1 34275
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_477
timestamp 1704896540
transform 1 0 1817 0 1 33939
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_478
timestamp 1704896540
transform 1 0 1817 0 1 33603
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_479
timestamp 1704896540
transform 1 0 1817 0 1 33267
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_480
timestamp 1704896540
transform 1 0 1817 0 1 32931
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_481
timestamp 1704896540
transform 1 0 1817 0 1 32595
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_482
timestamp 1704896540
transform 1 0 1817 0 1 32259
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_483
timestamp 1704896540
transform 1 0 1817 0 1 31923
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_484
timestamp 1704896540
transform 1 0 1817 0 1 39651
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_485
timestamp 1704896540
transform 1 0 1817 0 1 31587
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_486
timestamp 1704896540
transform 1 0 1817 0 1 39315
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_487
timestamp 1704896540
transform 1 0 1817 0 1 38979
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_488
timestamp 1704896540
transform 1 0 1817 0 1 31251
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_489
timestamp 1704896540
transform 1 0 1817 0 1 38643
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_490
timestamp 1704896540
transform 1 0 1817 0 1 38307
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_491
timestamp 1704896540
transform 1 0 1817 0 1 37971
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_492
timestamp 1704896540
transform 1 0 1817 0 1 37635
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_493
timestamp 1704896540
transform 1 0 1817 0 1 37299
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_494
timestamp 1704896540
transform 1 0 1817 0 1 30915
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_495
timestamp 1704896540
transform 1 0 1817 0 1 36963
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_496
timestamp 1704896540
transform 1 0 1817 0 1 36627
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_497
timestamp 1704896540
transform 1 0 1817 0 1 36291
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_498
timestamp 1704896540
transform 1 0 1817 0 1 30579
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_499
timestamp 1704896540
transform 1 0 1817 0 1 46371
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_500
timestamp 1704896540
transform 1 0 1817 0 1 46035
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_501
timestamp 1704896540
transform 1 0 1817 0 1 45699
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_502
timestamp 1704896540
transform 1 0 1817 0 1 45363
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_503
timestamp 1704896540
transform 1 0 1817 0 1 45027
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_504
timestamp 1704896540
transform 1 0 1817 0 1 44691
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_505
timestamp 1704896540
transform 1 0 1817 0 1 44355
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_506
timestamp 1704896540
transform 1 0 1817 0 1 44019
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_507
timestamp 1704896540
transform 1 0 1817 0 1 43683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_508
timestamp 1704896540
transform 1 0 1817 0 1 40323
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_509
timestamp 1704896540
transform 1 0 1817 0 1 39987
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_510
timestamp 1704896540
transform 1 0 1817 0 1 49059
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_511
timestamp 1704896540
transform 1 0 1817 0 1 43347
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_512
timestamp 1704896540
transform 1 0 1817 0 1 41331
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_513
timestamp 1704896540
transform 1 0 1817 0 1 43011
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_514
timestamp 1704896540
transform 1 0 1817 0 1 41667
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_515
timestamp 1704896540
transform 1 0 1817 0 1 48387
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_516
timestamp 1704896540
transform 1 0 1817 0 1 42675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_517
timestamp 1704896540
transform 1 0 1817 0 1 40995
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_518
timestamp 1704896540
transform 1 0 1817 0 1 48051
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_519
timestamp 1704896540
transform 1 0 1817 0 1 47715
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_520
timestamp 1704896540
transform 1 0 1817 0 1 47043
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_521
timestamp 1704896540
transform 1 0 1817 0 1 46707
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_522
timestamp 1704896540
transform 1 0 1817 0 1 47379
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_523
timestamp 1704896540
transform 1 0 1817 0 1 42339
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_524
timestamp 1704896540
transform 1 0 1817 0 1 40659
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_525
timestamp 1704896540
transform 1 0 1817 0 1 42003
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_526
timestamp 1704896540
transform 1 0 1817 0 1 48723
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_527
timestamp 1704896540
transform 1 0 1817 0 1 49395
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_528
timestamp 1704896540
transform 1 0 1817 0 1 59139
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_529
timestamp 1704896540
transform 1 0 1817 0 1 58803
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_530
timestamp 1704896540
transform 1 0 1817 0 1 58467
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_531
timestamp 1704896540
transform 1 0 1817 0 1 58131
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_532
timestamp 1704896540
transform 1 0 1817 0 1 57795
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_533
timestamp 1704896540
transform 1 0 1817 0 1 57459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_534
timestamp 1704896540
transform 1 0 1817 0 1 57123
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_535
timestamp 1704896540
transform 1 0 1817 0 1 56787
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_536
timestamp 1704896540
transform 1 0 1817 0 1 56451
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_537
timestamp 1704896540
transform 1 0 1817 0 1 56115
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_538
timestamp 1704896540
transform 1 0 1817 0 1 55779
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_539
timestamp 1704896540
transform 1 0 1817 0 1 55443
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_540
timestamp 1704896540
transform 1 0 1817 0 1 55107
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_541
timestamp 1704896540
transform 1 0 1817 0 1 54771
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_542
timestamp 1704896540
transform 1 0 1817 0 1 54435
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_543
timestamp 1704896540
transform 1 0 1817 0 1 54099
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_544
timestamp 1704896540
transform 1 0 1817 0 1 53763
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_545
timestamp 1704896540
transform 1 0 1817 0 1 50739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_546
timestamp 1704896540
transform 1 0 1817 0 1 50403
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_547
timestamp 1704896540
transform 1 0 1817 0 1 49731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_548
timestamp 1704896540
transform 1 0 1817 0 1 50067
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_549
timestamp 1704896540
transform 1 0 1817 0 1 52083
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_550
timestamp 1704896540
transform 1 0 1817 0 1 53427
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_551
timestamp 1704896540
transform 1 0 1817 0 1 53091
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_552
timestamp 1704896540
transform 1 0 1817 0 1 51747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_553
timestamp 1704896540
transform 1 0 1817 0 1 51411
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_554
timestamp 1704896540
transform 1 0 1817 0 1 51075
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_555
timestamp 1704896540
transform 1 0 1817 0 1 52755
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_556
timestamp 1704896540
transform 1 0 1817 0 1 52419
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_557
timestamp 1704896540
transform 1 0 1817 0 1 59811
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_558
timestamp 1704896540
transform 1 0 1817 0 1 69219
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_559
timestamp 1704896540
transform 1 0 1817 0 1 68883
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_560
timestamp 1704896540
transform 1 0 1817 0 1 68547
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_561
timestamp 1704896540
transform 1 0 1817 0 1 68211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_562
timestamp 1704896540
transform 1 0 1817 0 1 67875
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_563
timestamp 1704896540
transform 1 0 1817 0 1 67539
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_564
timestamp 1704896540
transform 1 0 1817 0 1 67203
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_565
timestamp 1704896540
transform 1 0 1817 0 1 66867
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_566
timestamp 1704896540
transform 1 0 1817 0 1 66531
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_567
timestamp 1704896540
transform 1 0 1817 0 1 66195
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_568
timestamp 1704896540
transform 1 0 1817 0 1 65859
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_569
timestamp 1704896540
transform 1 0 1817 0 1 65523
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_570
timestamp 1704896540
transform 1 0 1817 0 1 65187
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_571
timestamp 1704896540
transform 1 0 1817 0 1 64851
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_572
timestamp 1704896540
transform 1 0 1817 0 1 64515
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_573
timestamp 1704896540
transform 1 0 1817 0 1 64179
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_574
timestamp 1704896540
transform 1 0 1817 0 1 63843
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_575
timestamp 1704896540
transform 1 0 1817 0 1 63507
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_576
timestamp 1704896540
transform 1 0 1817 0 1 63171
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_577
timestamp 1704896540
transform 1 0 1817 0 1 62835
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_578
timestamp 1704896540
transform 1 0 1817 0 1 62499
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_579
timestamp 1704896540
transform 1 0 1817 0 1 62163
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_580
timestamp 1704896540
transform 1 0 1817 0 1 61827
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_581
timestamp 1704896540
transform 1 0 1817 0 1 61491
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_582
timestamp 1704896540
transform 1 0 1817 0 1 61155
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_583
timestamp 1704896540
transform 1 0 1817 0 1 60819
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_584
timestamp 1704896540
transform 1 0 1817 0 1 60483
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_585
timestamp 1704896540
transform 1 0 1817 0 1 60147
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_586
timestamp 1704896540
transform 1 0 1817 0 1 70227
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_587
timestamp 1704896540
transform 1 0 1817 0 1 70563
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_588
timestamp 1704896540
transform 1 0 1817 0 1 69891
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_589
timestamp 1704896540
transform 1 0 1817 0 1 69555
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_590
timestamp 1704896540
transform 1 0 1817 0 1 70899
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_591
timestamp 1704896540
transform 1 0 1817 0 1 71571
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_592
timestamp 1704896540
transform 1 0 1817 0 1 73923
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_593
timestamp 1704896540
transform 1 0 1817 0 1 73587
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_594
timestamp 1704896540
transform 1 0 1817 0 1 73251
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_595
timestamp 1704896540
transform 1 0 1817 0 1 72915
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_596
timestamp 1704896540
transform 1 0 1817 0 1 72579
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_597
timestamp 1704896540
transform 1 0 1817 0 1 72243
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_598
timestamp 1704896540
transform 1 0 1817 0 1 71235
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_599
timestamp 1704896540
transform 1 0 1817 0 1 71907
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_600
timestamp 1704896540
transform 1 0 4169 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_601
timestamp 1704896540
transform 1 0 3833 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_602
timestamp 1704896540
transform 1 0 1817 0 1 77283
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_603
timestamp 1704896540
transform 1 0 1817 0 1 76947
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_604
timestamp 1704896540
transform 1 0 1817 0 1 76611
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_605
timestamp 1704896540
transform 1 0 1817 0 1 76275
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_606
timestamp 1704896540
transform 1 0 1817 0 1 75939
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_607
timestamp 1704896540
transform 1 0 1817 0 1 75603
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_608
timestamp 1704896540
transform 1 0 1817 0 1 75267
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_609
timestamp 1704896540
transform 1 0 1817 0 1 74931
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_610
timestamp 1704896540
transform 1 0 1817 0 1 74595
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_611
timestamp 1704896540
transform 1 0 3497 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_612
timestamp 1704896540
transform 1 0 3161 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_613
timestamp 1704896540
transform 1 0 2825 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_614
timestamp 1704896540
transform 1 0 2489 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_615
timestamp 1704896540
transform 1 0 2153 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_616
timestamp 1704896540
transform 1 0 5849 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_617
timestamp 1704896540
transform 1 0 5513 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_618
timestamp 1704896540
transform 1 0 5177 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_619
timestamp 1704896540
transform 1 0 4841 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_620
timestamp 1704896540
transform 1 0 4505 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_621
timestamp 1704896540
transform 1 0 6857 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_622
timestamp 1704896540
transform 1 0 6521 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_623
timestamp 1704896540
transform 1 0 11897 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_624
timestamp 1704896540
transform 1 0 11561 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_625
timestamp 1704896540
transform 1 0 11225 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_626
timestamp 1704896540
transform 1 0 10889 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_627
timestamp 1704896540
transform 1 0 10553 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_628
timestamp 1704896540
transform 1 0 10217 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_629
timestamp 1704896540
transform 1 0 9881 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_630
timestamp 1704896540
transform 1 0 9545 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_631
timestamp 1704896540
transform 1 0 9209 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_632
timestamp 1704896540
transform 1 0 8873 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_633
timestamp 1704896540
transform 1 0 8537 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_634
timestamp 1704896540
transform 1 0 8201 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_635
timestamp 1704896540
transform 1 0 7865 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_636
timestamp 1704896540
transform 1 0 7529 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_637
timestamp 1704896540
transform 1 0 7193 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_638
timestamp 1704896540
transform 1 0 1817 0 1 74259
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_639
timestamp 1704896540
transform 1 0 6185 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_640
timestamp 1704896540
transform 1 0 16937 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_641
timestamp 1704896540
transform 1 0 16601 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_642
timestamp 1704896540
transform 1 0 16265 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_643
timestamp 1704896540
transform 1 0 15929 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_644
timestamp 1704896540
transform 1 0 15593 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_645
timestamp 1704896540
transform 1 0 15257 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_646
timestamp 1704896540
transform 1 0 14921 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_647
timestamp 1704896540
transform 1 0 14585 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_648
timestamp 1704896540
transform 1 0 14249 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_649
timestamp 1704896540
transform 1 0 13913 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_650
timestamp 1704896540
transform 1 0 13577 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_651
timestamp 1704896540
transform 1 0 13241 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_652
timestamp 1704896540
transform 1 0 12905 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_653
timestamp 1704896540
transform 1 0 12569 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_654
timestamp 1704896540
transform 1 0 12233 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_655
timestamp 1704896540
transform 1 0 17945 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_656
timestamp 1704896540
transform 1 0 17609 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_657
timestamp 1704896540
transform 1 0 17273 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_658
timestamp 1704896540
transform 1 0 23993 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_659
timestamp 1704896540
transform 1 0 23657 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_660
timestamp 1704896540
transform 1 0 23321 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_661
timestamp 1704896540
transform 1 0 22985 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_662
timestamp 1704896540
transform 1 0 22649 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_663
timestamp 1704896540
transform 1 0 22313 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_664
timestamp 1704896540
transform 1 0 21977 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_665
timestamp 1704896540
transform 1 0 21641 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_666
timestamp 1704896540
transform 1 0 21305 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_667
timestamp 1704896540
transform 1 0 20969 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_668
timestamp 1704896540
transform 1 0 20633 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_669
timestamp 1704896540
transform 1 0 20297 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_670
timestamp 1704896540
transform 1 0 19961 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_671
timestamp 1704896540
transform 1 0 19625 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_672
timestamp 1704896540
transform 1 0 19289 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_673
timestamp 1704896540
transform 1 0 18953 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_674
timestamp 1704896540
transform 1 0 18617 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_675
timestamp 1704896540
transform 1 0 18281 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_676
timestamp 1704896540
transform 1 0 25673 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_677
timestamp 1704896540
transform 1 0 25337 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_678
timestamp 1704896540
transform 1 0 25001 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_679
timestamp 1704896540
transform 1 0 24665 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_680
timestamp 1704896540
transform 1 0 24329 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_681
timestamp 1704896540
transform 1 0 29705 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_682
timestamp 1704896540
transform 1 0 29369 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_683
timestamp 1704896540
transform 1 0 29033 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_684
timestamp 1704896540
transform 1 0 28697 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_685
timestamp 1704896540
transform 1 0 28361 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_686
timestamp 1704896540
transform 1 0 28025 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_687
timestamp 1704896540
transform 1 0 27689 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_688
timestamp 1704896540
transform 1 0 27353 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_689
timestamp 1704896540
transform 1 0 27017 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_690
timestamp 1704896540
transform 1 0 26681 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_691
timestamp 1704896540
transform 1 0 26345 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_692
timestamp 1704896540
transform 1 0 26009 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_693
timestamp 1704896540
transform 1 0 35753 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_694
timestamp 1704896540
transform 1 0 35417 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_695
timestamp 1704896540
transform 1 0 35081 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_696
timestamp 1704896540
transform 1 0 34745 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_697
timestamp 1704896540
transform 1 0 34409 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_698
timestamp 1704896540
transform 1 0 34073 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_699
timestamp 1704896540
transform 1 0 33737 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_700
timestamp 1704896540
transform 1 0 33401 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_701
timestamp 1704896540
transform 1 0 33065 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_702
timestamp 1704896540
transform 1 0 32729 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_703
timestamp 1704896540
transform 1 0 32393 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_704
timestamp 1704896540
transform 1 0 32057 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_705
timestamp 1704896540
transform 1 0 31721 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_706
timestamp 1704896540
transform 1 0 31385 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_707
timestamp 1704896540
transform 1 0 31049 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_708
timestamp 1704896540
transform 1 0 30713 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_709
timestamp 1704896540
transform 1 0 30377 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_710
timestamp 1704896540
transform 1 0 30041 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_711
timestamp 1704896540
transform 1 0 36425 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_712
timestamp 1704896540
transform 1 0 36089 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_713
timestamp 1704896540
transform 1 0 41801 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_714
timestamp 1704896540
transform 1 0 41465 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_715
timestamp 1704896540
transform 1 0 41129 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_716
timestamp 1704896540
transform 1 0 40793 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_717
timestamp 1704896540
transform 1 0 40457 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_718
timestamp 1704896540
transform 1 0 40121 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_719
timestamp 1704896540
transform 1 0 39785 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_720
timestamp 1704896540
transform 1 0 39449 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_721
timestamp 1704896540
transform 1 0 39113 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_722
timestamp 1704896540
transform 1 0 38777 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_723
timestamp 1704896540
transform 1 0 38441 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_724
timestamp 1704896540
transform 1 0 38105 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_725
timestamp 1704896540
transform 1 0 37769 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_726
timestamp 1704896540
transform 1 0 37433 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_727
timestamp 1704896540
transform 1 0 37097 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_728
timestamp 1704896540
transform 1 0 36761 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_729
timestamp 1704896540
transform 1 0 42809 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_730
timestamp 1704896540
transform 1 0 42473 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_731
timestamp 1704896540
transform 1 0 42137 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_732
timestamp 1704896540
transform 1 0 47849 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_733
timestamp 1704896540
transform 1 0 47513 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_734
timestamp 1704896540
transform 1 0 47177 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_735
timestamp 1704896540
transform 1 0 46841 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_736
timestamp 1704896540
transform 1 0 46505 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_737
timestamp 1704896540
transform 1 0 46169 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_738
timestamp 1704896540
transform 1 0 45833 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_739
timestamp 1704896540
transform 1 0 45497 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_740
timestamp 1704896540
transform 1 0 45161 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_741
timestamp 1704896540
transform 1 0 44825 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_742
timestamp 1704896540
transform 1 0 44489 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_743
timestamp 1704896540
transform 1 0 44153 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_744
timestamp 1704896540
transform 1 0 43817 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_745
timestamp 1704896540
transform 1 0 43481 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_746
timestamp 1704896540
transform 1 0 43145 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_747
timestamp 1704896540
transform 1 0 1817 0 1 59475
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_748
timestamp 1704896540
transform 1 0 94175 0 1 40323
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_749
timestamp 1704896540
transform 1 0 94175 0 1 46035
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_750
timestamp 1704896540
transform 1 0 94175 0 1 45699
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_751
timestamp 1704896540
transform 1 0 94175 0 1 45363
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_752
timestamp 1704896540
transform 1 0 94175 0 1 45027
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_753
timestamp 1704896540
transform 1 0 94175 0 1 44691
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_754
timestamp 1704896540
transform 1 0 94175 0 1 44355
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_755
timestamp 1704896540
transform 1 0 94175 0 1 44019
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_756
timestamp 1704896540
transform 1 0 94175 0 1 43683
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_757
timestamp 1704896540
transform 1 0 94175 0 1 43347
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_758
timestamp 1704896540
transform 1 0 94175 0 1 43011
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_759
timestamp 1704896540
transform 1 0 94175 0 1 42675
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_760
timestamp 1704896540
transform 1 0 94175 0 1 42339
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_761
timestamp 1704896540
transform 1 0 94175 0 1 42003
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_762
timestamp 1704896540
transform 1 0 94175 0 1 39987
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_763
timestamp 1704896540
transform 1 0 94175 0 1 41667
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_764
timestamp 1704896540
transform 1 0 94175 0 1 41331
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_765
timestamp 1704896540
transform 1 0 94175 0 1 40995
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_766
timestamp 1704896540
transform 1 0 94175 0 1 49395
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_767
timestamp 1704896540
transform 1 0 94175 0 1 49059
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_768
timestamp 1704896540
transform 1 0 94175 0 1 48723
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_769
timestamp 1704896540
transform 1 0 94175 0 1 48387
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_770
timestamp 1704896540
transform 1 0 94175 0 1 48051
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_771
timestamp 1704896540
transform 1 0 94175 0 1 47715
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_772
timestamp 1704896540
transform 1 0 94175 0 1 47379
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_773
timestamp 1704896540
transform 1 0 94175 0 1 40659
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_774
timestamp 1704896540
transform 1 0 94175 0 1 47043
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_775
timestamp 1704896540
transform 1 0 94175 0 1 46707
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_776
timestamp 1704896540
transform 1 0 94175 0 1 46371
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_777
timestamp 1704896540
transform 1 0 94175 0 1 50739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_778
timestamp 1704896540
transform 1 0 94175 0 1 50403
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_779
timestamp 1704896540
transform 1 0 94175 0 1 50067
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_780
timestamp 1704896540
transform 1 0 94175 0 1 49731
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_781
timestamp 1704896540
transform 1 0 94175 0 1 54435
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_782
timestamp 1704896540
transform 1 0 94175 0 1 54099
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_783
timestamp 1704896540
transform 1 0 94175 0 1 53763
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_784
timestamp 1704896540
transform 1 0 94175 0 1 53427
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_785
timestamp 1704896540
transform 1 0 94175 0 1 53091
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_786
timestamp 1704896540
transform 1 0 94175 0 1 52755
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_787
timestamp 1704896540
transform 1 0 94175 0 1 52419
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_788
timestamp 1704896540
transform 1 0 94175 0 1 52083
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_789
timestamp 1704896540
transform 1 0 94175 0 1 51747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_790
timestamp 1704896540
transform 1 0 94175 0 1 51411
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_791
timestamp 1704896540
transform 1 0 94175 0 1 51075
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_792
timestamp 1704896540
transform 1 0 94175 0 1 55779
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_793
timestamp 1704896540
transform 1 0 94175 0 1 55443
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_794
timestamp 1704896540
transform 1 0 94175 0 1 55107
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_795
timestamp 1704896540
transform 1 0 94175 0 1 54771
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_796
timestamp 1704896540
transform 1 0 94175 0 1 59139
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_797
timestamp 1704896540
transform 1 0 94175 0 1 58803
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_798
timestamp 1704896540
transform 1 0 94175 0 1 58467
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_799
timestamp 1704896540
transform 1 0 94175 0 1 58131
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_800
timestamp 1704896540
transform 1 0 94175 0 1 57795
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_801
timestamp 1704896540
transform 1 0 94175 0 1 57459
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_802
timestamp 1704896540
transform 1 0 94175 0 1 57123
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_803
timestamp 1704896540
transform 1 0 94175 0 1 56787
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_804
timestamp 1704896540
transform 1 0 94175 0 1 56451
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_805
timestamp 1704896540
transform 1 0 94175 0 1 56115
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_806
timestamp 1704896540
transform 1 0 48521 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_807
timestamp 1704896540
transform 1 0 48185 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_808
timestamp 1704896540
transform 1 0 53561 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_809
timestamp 1704896540
transform 1 0 53225 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_810
timestamp 1704896540
transform 1 0 52889 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_811
timestamp 1704896540
transform 1 0 52553 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_812
timestamp 1704896540
transform 1 0 52217 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_813
timestamp 1704896540
transform 1 0 51881 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_814
timestamp 1704896540
transform 1 0 51545 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_815
timestamp 1704896540
transform 1 0 51209 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_816
timestamp 1704896540
transform 1 0 50873 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_817
timestamp 1704896540
transform 1 0 50537 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_818
timestamp 1704896540
transform 1 0 50201 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_819
timestamp 1704896540
transform 1 0 49865 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_820
timestamp 1704896540
transform 1 0 49529 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_821
timestamp 1704896540
transform 1 0 49193 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_822
timestamp 1704896540
transform 1 0 48857 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_823
timestamp 1704896540
transform 1 0 59609 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_824
timestamp 1704896540
transform 1 0 59273 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_825
timestamp 1704896540
transform 1 0 58937 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_826
timestamp 1704896540
transform 1 0 58601 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_827
timestamp 1704896540
transform 1 0 58265 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_828
timestamp 1704896540
transform 1 0 57929 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_829
timestamp 1704896540
transform 1 0 57593 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_830
timestamp 1704896540
transform 1 0 57257 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_831
timestamp 1704896540
transform 1 0 56921 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_832
timestamp 1704896540
transform 1 0 56585 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_833
timestamp 1704896540
transform 1 0 56249 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_834
timestamp 1704896540
transform 1 0 55913 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_835
timestamp 1704896540
transform 1 0 55577 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_836
timestamp 1704896540
transform 1 0 55241 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_837
timestamp 1704896540
transform 1 0 54905 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_838
timestamp 1704896540
transform 1 0 54569 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_839
timestamp 1704896540
transform 1 0 54233 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_840
timestamp 1704896540
transform 1 0 53897 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_841
timestamp 1704896540
transform 1 0 62297 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_842
timestamp 1704896540
transform 1 0 61961 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_843
timestamp 1704896540
transform 1 0 61625 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_844
timestamp 1704896540
transform 1 0 61289 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_845
timestamp 1704896540
transform 1 0 60953 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_846
timestamp 1704896540
transform 1 0 60617 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_847
timestamp 1704896540
transform 1 0 60281 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_848
timestamp 1704896540
transform 1 0 59945 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_849
timestamp 1704896540
transform 1 0 62633 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_850
timestamp 1704896540
transform 1 0 64313 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_851
timestamp 1704896540
transform 1 0 63977 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_852
timestamp 1704896540
transform 1 0 63641 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_853
timestamp 1704896540
transform 1 0 65657 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_854
timestamp 1704896540
transform 1 0 65321 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_855
timestamp 1704896540
transform 1 0 64985 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_856
timestamp 1704896540
transform 1 0 64649 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_857
timestamp 1704896540
transform 1 0 63305 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_858
timestamp 1704896540
transform 1 0 62969 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_859
timestamp 1704896540
transform 1 0 71705 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_860
timestamp 1704896540
transform 1 0 71369 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_861
timestamp 1704896540
transform 1 0 71033 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_862
timestamp 1704896540
transform 1 0 70697 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_863
timestamp 1704896540
transform 1 0 70361 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_864
timestamp 1704896540
transform 1 0 70025 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_865
timestamp 1704896540
transform 1 0 69689 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_866
timestamp 1704896540
transform 1 0 69353 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_867
timestamp 1704896540
transform 1 0 69017 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_868
timestamp 1704896540
transform 1 0 68681 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_869
timestamp 1704896540
transform 1 0 68345 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_870
timestamp 1704896540
transform 1 0 68009 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_871
timestamp 1704896540
transform 1 0 67673 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_872
timestamp 1704896540
transform 1 0 67337 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_873
timestamp 1704896540
transform 1 0 67001 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_874
timestamp 1704896540
transform 1 0 66665 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_875
timestamp 1704896540
transform 1 0 66329 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_876
timestamp 1704896540
transform 1 0 65993 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_877
timestamp 1704896540
transform 1 0 94175 0 1 60819
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_878
timestamp 1704896540
transform 1 0 94175 0 1 59811
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_879
timestamp 1704896540
transform 1 0 94175 0 1 64179
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_880
timestamp 1704896540
transform 1 0 94175 0 1 63843
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_881
timestamp 1704896540
transform 1 0 94175 0 1 63507
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_882
timestamp 1704896540
transform 1 0 94175 0 1 63171
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_883
timestamp 1704896540
transform 1 0 94175 0 1 62835
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_884
timestamp 1704896540
transform 1 0 94175 0 1 62499
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_885
timestamp 1704896540
transform 1 0 94175 0 1 62163
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_886
timestamp 1704896540
transform 1 0 94175 0 1 61827
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_887
timestamp 1704896540
transform 1 0 94175 0 1 60483
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_888
timestamp 1704896540
transform 1 0 94175 0 1 61491
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_889
timestamp 1704896540
transform 1 0 94175 0 1 61155
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_890
timestamp 1704896540
transform 1 0 94175 0 1 60147
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_891
timestamp 1704896540
transform 1 0 94175 0 1 69219
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_892
timestamp 1704896540
transform 1 0 94175 0 1 68883
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_893
timestamp 1704896540
transform 1 0 94175 0 1 68547
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_894
timestamp 1704896540
transform 1 0 94175 0 1 68211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_895
timestamp 1704896540
transform 1 0 94175 0 1 67875
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_896
timestamp 1704896540
transform 1 0 94175 0 1 67539
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_897
timestamp 1704896540
transform 1 0 94175 0 1 67203
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_898
timestamp 1704896540
transform 1 0 94175 0 1 66867
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_899
timestamp 1704896540
transform 1 0 94175 0 1 66531
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_900
timestamp 1704896540
transform 1 0 94175 0 1 66195
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_901
timestamp 1704896540
transform 1 0 94175 0 1 65859
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_902
timestamp 1704896540
transform 1 0 94175 0 1 65523
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_903
timestamp 1704896540
transform 1 0 94175 0 1 65187
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_904
timestamp 1704896540
transform 1 0 94175 0 1 64851
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_905
timestamp 1704896540
transform 1 0 94175 0 1 64515
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_906
timestamp 1704896540
transform 1 0 76073 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_907
timestamp 1704896540
transform 1 0 72041 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_908
timestamp 1704896540
transform 1 0 75737 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_909
timestamp 1704896540
transform 1 0 75401 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_910
timestamp 1704896540
transform 1 0 75065 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_911
timestamp 1704896540
transform 1 0 74729 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_912
timestamp 1704896540
transform 1 0 74393 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_913
timestamp 1704896540
transform 1 0 74057 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_914
timestamp 1704896540
transform 1 0 73721 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_915
timestamp 1704896540
transform 1 0 73385 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_916
timestamp 1704896540
transform 1 0 73049 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_917
timestamp 1704896540
transform 1 0 72713 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_918
timestamp 1704896540
transform 1 0 72377 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_919
timestamp 1704896540
transform 1 0 76409 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_920
timestamp 1704896540
transform 1 0 77417 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_921
timestamp 1704896540
transform 1 0 77081 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_922
timestamp 1704896540
transform 1 0 76745 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_923
timestamp 1704896540
transform 1 0 78089 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_924
timestamp 1704896540
transform 1 0 83465 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_925
timestamp 1704896540
transform 1 0 83129 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_926
timestamp 1704896540
transform 1 0 82793 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_927
timestamp 1704896540
transform 1 0 82457 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_928
timestamp 1704896540
transform 1 0 82121 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_929
timestamp 1704896540
transform 1 0 81785 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_930
timestamp 1704896540
transform 1 0 81449 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_931
timestamp 1704896540
transform 1 0 81113 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_932
timestamp 1704896540
transform 1 0 80777 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_933
timestamp 1704896540
transform 1 0 80441 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_934
timestamp 1704896540
transform 1 0 80105 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_935
timestamp 1704896540
transform 1 0 79769 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_936
timestamp 1704896540
transform 1 0 79433 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_937
timestamp 1704896540
transform 1 0 79097 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_938
timestamp 1704896540
transform 1 0 78761 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_939
timestamp 1704896540
transform 1 0 78425 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_940
timestamp 1704896540
transform 1 0 77753 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_941
timestamp 1704896540
transform 1 0 94175 0 1 71907
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_942
timestamp 1704896540
transform 1 0 94175 0 1 71571
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_943
timestamp 1704896540
transform 1 0 94175 0 1 71235
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_944
timestamp 1704896540
transform 1 0 94175 0 1 70899
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_945
timestamp 1704896540
transform 1 0 94175 0 1 70563
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_946
timestamp 1704896540
transform 1 0 94175 0 1 70227
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_947
timestamp 1704896540
transform 1 0 94175 0 1 69891
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_948
timestamp 1704896540
transform 1 0 94175 0 1 69555
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_949
timestamp 1704896540
transform 1 0 94175 0 1 73923
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_950
timestamp 1704896540
transform 1 0 94175 0 1 73587
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_951
timestamp 1704896540
transform 1 0 94175 0 1 73251
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_952
timestamp 1704896540
transform 1 0 94175 0 1 72915
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_953
timestamp 1704896540
transform 1 0 94175 0 1 72579
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_954
timestamp 1704896540
transform 1 0 94175 0 1 72243
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_955
timestamp 1704896540
transform 1 0 84809 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_956
timestamp 1704896540
transform 1 0 84473 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_957
timestamp 1704896540
transform 1 0 84137 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_958
timestamp 1704896540
transform 1 0 83801 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_959
timestamp 1704896540
transform 1 0 89513 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_960
timestamp 1704896540
transform 1 0 89177 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_961
timestamp 1704896540
transform 1 0 88841 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_962
timestamp 1704896540
transform 1 0 88505 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_963
timestamp 1704896540
transform 1 0 88169 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_964
timestamp 1704896540
transform 1 0 87833 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_965
timestamp 1704896540
transform 1 0 87497 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_966
timestamp 1704896540
transform 1 0 87161 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_967
timestamp 1704896540
transform 1 0 86825 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_968
timestamp 1704896540
transform 1 0 86489 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_969
timestamp 1704896540
transform 1 0 86153 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_970
timestamp 1704896540
transform 1 0 85817 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_971
timestamp 1704896540
transform 1 0 85481 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_972
timestamp 1704896540
transform 1 0 85145 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_973
timestamp 1704896540
transform 1 0 94175 0 1 77283
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_974
timestamp 1704896540
transform 1 0 94175 0 1 76947
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_975
timestamp 1704896540
transform 1 0 94175 0 1 76611
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_976
timestamp 1704896540
transform 1 0 94175 0 1 76275
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_977
timestamp 1704896540
transform 1 0 94175 0 1 75939
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_978
timestamp 1704896540
transform 1 0 94175 0 1 75603
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_979
timestamp 1704896540
transform 1 0 94175 0 1 75267
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_980
timestamp 1704896540
transform 1 0 94175 0 1 74931
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_981
timestamp 1704896540
transform 1 0 94175 0 1 74595
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_982
timestamp 1704896540
transform 1 0 90185 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_983
timestamp 1704896540
transform 1 0 89849 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_984
timestamp 1704896540
transform 1 0 93545 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_985
timestamp 1704896540
transform 1 0 93209 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_986
timestamp 1704896540
transform 1 0 92873 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_987
timestamp 1704896540
transform 1 0 92537 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_988
timestamp 1704896540
transform 1 0 92201 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_989
timestamp 1704896540
transform 1 0 91865 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_990
timestamp 1704896540
transform 1 0 91529 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_991
timestamp 1704896540
transform 1 0 91193 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_992
timestamp 1704896540
transform 1 0 90857 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_993
timestamp 1704896540
transform 1 0 90521 0 1 77747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_994
timestamp 1704896540
transform 1 0 94175 0 1 74259
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_995
timestamp 1704896540
transform 1 0 94175 0 1 59475
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_0
timestamp 1704896540
transform 1 0 94172 0 1 4708
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_1
timestamp 1704896540
transform 1 0 94172 0 1 4372
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_2
timestamp 1704896540
transform 1 0 94172 0 1 4036
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_3
timestamp 1704896540
transform 1 0 94172 0 1 3700
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_4
timestamp 1704896540
transform 1 0 94172 0 1 3364
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_5
timestamp 1704896540
transform 1 0 94172 0 1 3028
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_6
timestamp 1704896540
transform 1 0 94172 0 1 2692
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_7
timestamp 1704896540
transform 1 0 94172 0 1 2356
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_8
timestamp 1704896540
transform 1 0 91190 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_9
timestamp 1704896540
transform 1 0 94172 0 1 2020
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_10
timestamp 1704896540
transform 1 0 94172 0 1 5044
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_11
timestamp 1704896540
transform 1 0 92870 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_12
timestamp 1704896540
transform 1 0 84470 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_13
timestamp 1704896540
transform 1 0 87830 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_14
timestamp 1704896540
transform 1 0 86150 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_15
timestamp 1704896540
transform 1 0 89510 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_16
timestamp 1704896540
transform 1 0 94172 0 1 7060
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_17
timestamp 1704896540
transform 1 0 94172 0 1 6724
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_18
timestamp 1704896540
transform 1 0 94172 0 1 5380
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_19
timestamp 1704896540
transform 1 0 94172 0 1 6388
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_20
timestamp 1704896540
transform 1 0 94172 0 1 6052
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_21
timestamp 1704896540
transform 1 0 94172 0 1 5716
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_22
timestamp 1704896540
transform 1 0 94172 0 1 9748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_23
timestamp 1704896540
transform 1 0 94172 0 1 9412
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_24
timestamp 1704896540
transform 1 0 94172 0 1 9076
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_25
timestamp 1704896540
transform 1 0 94172 0 1 8740
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_26
timestamp 1704896540
transform 1 0 94172 0 1 8404
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_27
timestamp 1704896540
transform 1 0 94172 0 1 8068
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_28
timestamp 1704896540
transform 1 0 94172 0 1 7732
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_29
timestamp 1704896540
transform 1 0 94172 0 1 7396
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_30
timestamp 1704896540
transform 1 0 81110 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_31
timestamp 1704896540
transform 1 0 79430 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_32
timestamp 1704896540
transform 1 0 82790 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_33
timestamp 1704896540
transform 1 0 72710 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_34
timestamp 1704896540
transform 1 0 74390 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_35
timestamp 1704896540
transform 1 0 76070 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_36
timestamp 1704896540
transform 1 0 81239 0 1 9269
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_37
timestamp 1704896540
transform 1 0 81159 0 1 7999
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_38
timestamp 1704896540
transform 1 0 77750 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_39
timestamp 1704896540
transform 1 0 81639 0 1 16483
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_40
timestamp 1704896540
transform 1 0 81319 0 1 10827
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_41
timestamp 1704896540
transform 1 0 81399 0 1 12097
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_42
timestamp 1704896540
transform 1 0 81479 0 1 13655
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_43
timestamp 1704896540
transform 1 0 81559 0 1 14925
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_44
timestamp 1704896540
transform 1 0 94172 0 1 19828
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_45
timestamp 1704896540
transform 1 0 94172 0 1 19492
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_46
timestamp 1704896540
transform 1 0 94172 0 1 19156
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_47
timestamp 1704896540
transform 1 0 94172 0 1 18820
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_48
timestamp 1704896540
transform 1 0 94172 0 1 18484
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_49
timestamp 1704896540
transform 1 0 94172 0 1 18148
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_50
timestamp 1704896540
transform 1 0 94172 0 1 17812
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_51
timestamp 1704896540
transform 1 0 94172 0 1 17476
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_52
timestamp 1704896540
transform 1 0 94172 0 1 17140
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_53
timestamp 1704896540
transform 1 0 94172 0 1 16804
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_54
timestamp 1704896540
transform 1 0 94172 0 1 16468
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_55
timestamp 1704896540
transform 1 0 94172 0 1 16132
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_56
timestamp 1704896540
transform 1 0 94172 0 1 15796
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_57
timestamp 1704896540
transform 1 0 94172 0 1 15460
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_58
timestamp 1704896540
transform 1 0 94172 0 1 15124
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_59
timestamp 1704896540
transform 1 0 94172 0 1 14788
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_60
timestamp 1704896540
transform 1 0 94172 0 1 14452
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_61
timestamp 1704896540
transform 1 0 94172 0 1 14116
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_62
timestamp 1704896540
transform 1 0 94172 0 1 13780
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_63
timestamp 1704896540
transform 1 0 94172 0 1 13444
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_64
timestamp 1704896540
transform 1 0 94172 0 1 13108
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_65
timestamp 1704896540
transform 1 0 94172 0 1 12772
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_66
timestamp 1704896540
transform 1 0 94172 0 1 12436
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_67
timestamp 1704896540
transform 1 0 94172 0 1 12100
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_68
timestamp 1704896540
transform 1 0 94172 0 1 11764
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_69
timestamp 1704896540
transform 1 0 94172 0 1 11428
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_70
timestamp 1704896540
transform 1 0 94172 0 1 11092
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_71
timestamp 1704896540
transform 1 0 94172 0 1 10756
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_72
timestamp 1704896540
transform 1 0 94172 0 1 10420
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_73
timestamp 1704896540
transform 1 0 94172 0 1 10084
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_74
timestamp 1704896540
transform 1 0 65990 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_75
timestamp 1704896540
transform 1 0 71030 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_76
timestamp 1704896540
transform 1 0 69350 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_77
timestamp 1704896540
transform 1 0 67670 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_78
timestamp 1704896540
transform 1 0 62630 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_79
timestamp 1704896540
transform 1 0 64310 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_80
timestamp 1704896540
transform 1 0 60950 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_81
timestamp 1704896540
transform 1 0 59270 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_82
timestamp 1704896540
transform 1 0 57590 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_83
timestamp 1704896540
transform 1 0 54230 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_84
timestamp 1704896540
transform 1 0 55910 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_85
timestamp 1704896540
transform 1 0 50870 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_86
timestamp 1704896540
transform 1 0 49190 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_87
timestamp 1704896540
transform 1 0 52550 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_88
timestamp 1704896540
transform 1 0 54414 0 1 10753
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_89
timestamp 1704896540
transform 1 0 48174 0 1 10753
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_90
timestamp 1704896540
transform 1 0 53166 0 1 10753
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_91
timestamp 1704896540
transform 1 0 51918 0 1 10753
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_92
timestamp 1704896540
transform 1 0 59406 0 1 10753
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_93
timestamp 1704896540
transform 1 0 58158 0 1 10753
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_94
timestamp 1704896540
transform 1 0 49422 0 1 10753
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_95
timestamp 1704896540
transform 1 0 56910 0 1 10753
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_96
timestamp 1704896540
transform 1 0 55662 0 1 10753
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_97
timestamp 1704896540
transform 1 0 50670 0 1 10753
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_98
timestamp 1704896540
transform 1 0 66894 0 1 10753
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_99
timestamp 1704896540
transform 1 0 65646 0 1 10753
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_100
timestamp 1704896540
transform 1 0 64398 0 1 10753
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_101
timestamp 1704896540
transform 1 0 63150 0 1 10753
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_102
timestamp 1704896540
transform 1 0 61902 0 1 10753
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_103
timestamp 1704896540
transform 1 0 60654 0 1 10753
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_104
timestamp 1704896540
transform 1 0 94172 0 1 23188
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_105
timestamp 1704896540
transform 1 0 94172 0 1 22852
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_106
timestamp 1704896540
transform 1 0 94172 0 1 22516
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_107
timestamp 1704896540
transform 1 0 94172 0 1 22180
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_108
timestamp 1704896540
transform 1 0 94172 0 1 21844
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_109
timestamp 1704896540
transform 1 0 94172 0 1 29572
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_110
timestamp 1704896540
transform 1 0 94172 0 1 21508
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_111
timestamp 1704896540
transform 1 0 94172 0 1 29236
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_112
timestamp 1704896540
transform 1 0 94172 0 1 28900
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_113
timestamp 1704896540
transform 1 0 94172 0 1 21172
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_114
timestamp 1704896540
transform 1 0 94172 0 1 20836
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_115
timestamp 1704896540
transform 1 0 94172 0 1 20500
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_116
timestamp 1704896540
transform 1 0 94172 0 1 28564
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_117
timestamp 1704896540
transform 1 0 94172 0 1 20164
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_118
timestamp 1704896540
transform 1 0 94172 0 1 28228
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_119
timestamp 1704896540
transform 1 0 94172 0 1 27892
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_120
timestamp 1704896540
transform 1 0 94172 0 1 27556
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_121
timestamp 1704896540
transform 1 0 94172 0 1 27220
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_122
timestamp 1704896540
transform 1 0 94172 0 1 26884
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_123
timestamp 1704896540
transform 1 0 94172 0 1 26548
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_124
timestamp 1704896540
transform 1 0 94172 0 1 26212
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_125
timestamp 1704896540
transform 1 0 94172 0 1 25876
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_126
timestamp 1704896540
transform 1 0 94172 0 1 25540
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_127
timestamp 1704896540
transform 1 0 94172 0 1 25204
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_128
timestamp 1704896540
transform 1 0 94172 0 1 24868
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_129
timestamp 1704896540
transform 1 0 94172 0 1 24532
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_130
timestamp 1704896540
transform 1 0 94172 0 1 24196
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_131
timestamp 1704896540
transform 1 0 94172 0 1 23860
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_132
timestamp 1704896540
transform 1 0 94172 0 1 23524
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_133
timestamp 1704896540
transform 1 0 94172 0 1 39652
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_134
timestamp 1704896540
transform 1 0 94172 0 1 39316
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_135
timestamp 1704896540
transform 1 0 94172 0 1 38980
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_136
timestamp 1704896540
transform 1 0 94172 0 1 38644
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_137
timestamp 1704896540
transform 1 0 94172 0 1 38308
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_138
timestamp 1704896540
transform 1 0 94172 0 1 37972
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_139
timestamp 1704896540
transform 1 0 94172 0 1 37636
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_140
timestamp 1704896540
transform 1 0 94172 0 1 37300
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_141
timestamp 1704896540
transform 1 0 94172 0 1 36964
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_142
timestamp 1704896540
transform 1 0 94172 0 1 36628
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_143
timestamp 1704896540
transform 1 0 94172 0 1 36292
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_144
timestamp 1704896540
transform 1 0 94172 0 1 35956
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_145
timestamp 1704896540
transform 1 0 94172 0 1 35620
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_146
timestamp 1704896540
transform 1 0 94172 0 1 35284
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_147
timestamp 1704896540
transform 1 0 94172 0 1 34948
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_148
timestamp 1704896540
transform 1 0 94172 0 1 34612
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_149
timestamp 1704896540
transform 1 0 94172 0 1 34276
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_150
timestamp 1704896540
transform 1 0 94172 0 1 33940
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_151
timestamp 1704896540
transform 1 0 94172 0 1 33604
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_152
timestamp 1704896540
transform 1 0 94172 0 1 33268
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_153
timestamp 1704896540
transform 1 0 94172 0 1 32932
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_154
timestamp 1704896540
transform 1 0 94172 0 1 32596
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_155
timestamp 1704896540
transform 1 0 94172 0 1 32260
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_156
timestamp 1704896540
transform 1 0 94172 0 1 31924
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_157
timestamp 1704896540
transform 1 0 94172 0 1 31588
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_158
timestamp 1704896540
transform 1 0 94172 0 1 31252
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_159
timestamp 1704896540
transform 1 0 94172 0 1 30916
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_160
timestamp 1704896540
transform 1 0 94172 0 1 30580
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_161
timestamp 1704896540
transform 1 0 94172 0 1 30244
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_162
timestamp 1704896540
transform 1 0 94172 0 1 29908
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_163
timestamp 1704896540
transform 1 0 44150 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_164
timestamp 1704896540
transform 1 0 47510 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_165
timestamp 1704896540
transform 1 0 45830 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_166
timestamp 1704896540
transform 1 0 42470 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_167
timestamp 1704896540
transform 1 0 40790 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_168
timestamp 1704896540
transform 1 0 37430 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_169
timestamp 1704896540
transform 1 0 39110 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_170
timestamp 1704896540
transform 1 0 30710 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_171
timestamp 1704896540
transform 1 0 35750 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_172
timestamp 1704896540
transform 1 0 32390 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_173
timestamp 1704896540
transform 1 0 34070 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_174
timestamp 1704896540
transform 1 0 27350 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_175
timestamp 1704896540
transform 1 0 25670 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_176
timestamp 1704896540
transform 1 0 29030 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_177
timestamp 1704896540
transform 1 0 34446 0 1 10753
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_178
timestamp 1704896540
transform 1 0 33198 0 1 10753
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_179
timestamp 1704896540
transform 1 0 31950 0 1 10753
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_180
timestamp 1704896540
transform 1 0 30702 0 1 10753
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_181
timestamp 1704896540
transform 1 0 29454 0 1 10753
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_182
timestamp 1704896540
transform 1 0 35694 0 1 10753
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_183
timestamp 1704896540
transform 1 0 28206 0 1 10753
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_184
timestamp 1704896540
transform 1 0 45678 0 1 10753
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_185
timestamp 1704896540
transform 1 0 44430 0 1 10753
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_186
timestamp 1704896540
transform 1 0 43182 0 1 10753
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_187
timestamp 1704896540
transform 1 0 41934 0 1 10753
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_188
timestamp 1704896540
transform 1 0 40686 0 1 10753
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_189
timestamp 1704896540
transform 1 0 39438 0 1 10753
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_190
timestamp 1704896540
transform 1 0 38190 0 1 10753
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_191
timestamp 1704896540
transform 1 0 36942 0 1 10753
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_192
timestamp 1704896540
transform 1 0 46926 0 1 10753
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_193
timestamp 1704896540
transform 1 0 22310 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_194
timestamp 1704896540
transform 1 0 18950 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_195
timestamp 1704896540
transform 1 0 20630 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_196
timestamp 1704896540
transform 1 0 23990 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_197
timestamp 1704896540
transform 1 0 12230 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_198
timestamp 1704896540
transform 1 0 13910 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_199
timestamp 1704896540
transform 1 0 17270 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_200
timestamp 1704896540
transform 1 0 15590 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_201
timestamp 1704896540
transform 1 0 7190 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_202
timestamp 1704896540
transform 1 0 10550 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_203
timestamp 1704896540
transform 1 0 8870 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_204
timestamp 1704896540
transform 1 0 2150 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_205
timestamp 1704896540
transform 1 0 5510 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_206
timestamp 1704896540
transform 1 0 1814 0 1 5044
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_207
timestamp 1704896540
transform 1 0 1814 0 1 4708
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_208
timestamp 1704896540
transform 1 0 1814 0 1 4372
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_209
timestamp 1704896540
transform 1 0 1814 0 1 4036
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_210
timestamp 1704896540
transform 1 0 1814 0 1 3700
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_211
timestamp 1704896540
transform 1 0 1814 0 1 3364
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_212
timestamp 1704896540
transform 1 0 1814 0 1 3028
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_213
timestamp 1704896540
transform 1 0 1814 0 1 2692
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_214
timestamp 1704896540
transform 1 0 1814 0 1 2356
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_215
timestamp 1704896540
transform 1 0 3830 0 1 1684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_216
timestamp 1704896540
transform 1 0 1814 0 1 2020
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_217
timestamp 1704896540
transform 1 0 1814 0 1 7060
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_218
timestamp 1704896540
transform 1 0 1814 0 1 6724
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_219
timestamp 1704896540
transform 1 0 1814 0 1 6388
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_220
timestamp 1704896540
transform 1 0 1814 0 1 6052
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_221
timestamp 1704896540
transform 1 0 1814 0 1 5716
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_222
timestamp 1704896540
transform 1 0 1814 0 1 5380
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_223
timestamp 1704896540
transform 1 0 1814 0 1 9076
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_224
timestamp 1704896540
transform 1 0 1814 0 1 8740
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_225
timestamp 1704896540
transform 1 0 1814 0 1 8404
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_226
timestamp 1704896540
transform 1 0 1814 0 1 7396
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_227
timestamp 1704896540
transform 1 0 1814 0 1 8068
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_228
timestamp 1704896540
transform 1 0 1814 0 1 7732
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_229
timestamp 1704896540
transform 1 0 1814 0 1 9412
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_230
timestamp 1704896540
transform 1 0 1814 0 1 9748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_231
timestamp 1704896540
transform 1 0 1814 0 1 13108
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_232
timestamp 1704896540
transform 1 0 1814 0 1 12772
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_233
timestamp 1704896540
transform 1 0 1814 0 1 12436
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_234
timestamp 1704896540
transform 1 0 1814 0 1 12100
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_235
timestamp 1704896540
transform 1 0 1814 0 1 11764
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_236
timestamp 1704896540
transform 1 0 1814 0 1 10420
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_237
timestamp 1704896540
transform 1 0 1814 0 1 11428
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_238
timestamp 1704896540
transform 1 0 1814 0 1 11092
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_239
timestamp 1704896540
transform 1 0 1814 0 1 10756
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_240
timestamp 1704896540
transform 1 0 1814 0 1 14788
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_241
timestamp 1704896540
transform 1 0 1814 0 1 14452
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_242
timestamp 1704896540
transform 1 0 1814 0 1 14116
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_243
timestamp 1704896540
transform 1 0 1814 0 1 13780
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_244
timestamp 1704896540
transform 1 0 1814 0 1 13444
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_245
timestamp 1704896540
transform 1 0 1814 0 1 17476
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_246
timestamp 1704896540
transform 1 0 1814 0 1 17140
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_247
timestamp 1704896540
transform 1 0 1814 0 1 16804
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_248
timestamp 1704896540
transform 1 0 1814 0 1 16468
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_249
timestamp 1704896540
transform 1 0 1814 0 1 16132
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_250
timestamp 1704896540
transform 1 0 1814 0 1 15796
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_251
timestamp 1704896540
transform 1 0 1814 0 1 15460
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_252
timestamp 1704896540
transform 1 0 1814 0 1 15124
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_253
timestamp 1704896540
transform 1 0 1814 0 1 17812
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_254
timestamp 1704896540
transform 1 0 1814 0 1 19828
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_255
timestamp 1704896540
transform 1 0 1814 0 1 19492
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_256
timestamp 1704896540
transform 1 0 1814 0 1 19156
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_257
timestamp 1704896540
transform 1 0 1814 0 1 18820
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_258
timestamp 1704896540
transform 1 0 1814 0 1 18484
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_259
timestamp 1704896540
transform 1 0 1814 0 1 18148
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_260
timestamp 1704896540
transform 1 0 1814 0 1 10084
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_261
timestamp 1704896540
transform 1 0 14535 0 1 27211
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_262
timestamp 1704896540
transform 1 0 14615 0 1 28481
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_263
timestamp 1704896540
transform 1 0 14455 0 1 25653
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_264
timestamp 1704896540
transform 1 0 1814 0 1 22180
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_265
timestamp 1704896540
transform 1 0 1814 0 1 21844
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_266
timestamp 1704896540
transform 1 0 1814 0 1 21508
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_267
timestamp 1704896540
transform 1 0 1814 0 1 21172
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_268
timestamp 1704896540
transform 1 0 1814 0 1 20836
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_269
timestamp 1704896540
transform 1 0 1814 0 1 20500
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_270
timestamp 1704896540
transform 1 0 1814 0 1 24868
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_271
timestamp 1704896540
transform 1 0 1814 0 1 24532
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_272
timestamp 1704896540
transform 1 0 1814 0 1 24196
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_273
timestamp 1704896540
transform 1 0 1814 0 1 23860
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_274
timestamp 1704896540
transform 1 0 1814 0 1 23524
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_275
timestamp 1704896540
transform 1 0 1814 0 1 23188
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_276
timestamp 1704896540
transform 1 0 1814 0 1 22852
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_277
timestamp 1704896540
transform 1 0 1814 0 1 22516
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_278
timestamp 1704896540
transform 1 0 1814 0 1 20164
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_279
timestamp 1704896540
transform 1 0 1814 0 1 27220
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_280
timestamp 1704896540
transform 1 0 1814 0 1 26884
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_281
timestamp 1704896540
transform 1 0 1814 0 1 26548
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_282
timestamp 1704896540
transform 1 0 1814 0 1 26212
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_283
timestamp 1704896540
transform 1 0 1814 0 1 25876
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_284
timestamp 1704896540
transform 1 0 1814 0 1 25540
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_285
timestamp 1704896540
transform 1 0 1814 0 1 25204
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_286
timestamp 1704896540
transform 1 0 1814 0 1 29572
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_287
timestamp 1704896540
transform 1 0 1814 0 1 29236
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_288
timestamp 1704896540
transform 1 0 1814 0 1 28900
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_289
timestamp 1704896540
transform 1 0 1814 0 1 28564
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_290
timestamp 1704896540
transform 1 0 1814 0 1 28228
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_291
timestamp 1704896540
transform 1 0 1814 0 1 27892
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_292
timestamp 1704896540
transform 1 0 1814 0 1 27556
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_293
timestamp 1704896540
transform 1 0 1814 0 1 30244
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_294
timestamp 1704896540
transform 1 0 1814 0 1 35956
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_295
timestamp 1704896540
transform 1 0 1814 0 1 29908
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_296
timestamp 1704896540
transform 1 0 1814 0 1 35620
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_297
timestamp 1704896540
transform 1 0 1814 0 1 35284
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_298
timestamp 1704896540
transform 1 0 1814 0 1 34948
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_299
timestamp 1704896540
transform 1 0 1814 0 1 34612
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_300
timestamp 1704896540
transform 1 0 1814 0 1 34276
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_301
timestamp 1704896540
transform 1 0 1814 0 1 33940
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_302
timestamp 1704896540
transform 1 0 1814 0 1 33604
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_303
timestamp 1704896540
transform 1 0 1814 0 1 33268
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_304
timestamp 1704896540
transform 1 0 1814 0 1 32932
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_305
timestamp 1704896540
transform 1 0 1814 0 1 32596
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_306
timestamp 1704896540
transform 1 0 1814 0 1 32260
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_307
timestamp 1704896540
transform 1 0 1814 0 1 31924
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_308
timestamp 1704896540
transform 1 0 1814 0 1 39652
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_309
timestamp 1704896540
transform 1 0 1814 0 1 31588
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_310
timestamp 1704896540
transform 1 0 1814 0 1 39316
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_311
timestamp 1704896540
transform 1 0 1814 0 1 38980
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_312
timestamp 1704896540
transform 1 0 1814 0 1 31252
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_313
timestamp 1704896540
transform 1 0 1814 0 1 38644
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_314
timestamp 1704896540
transform 1 0 1814 0 1 38308
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_315
timestamp 1704896540
transform 1 0 1814 0 1 37972
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_316
timestamp 1704896540
transform 1 0 1814 0 1 37636
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_317
timestamp 1704896540
transform 1 0 1814 0 1 30916
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_318
timestamp 1704896540
transform 1 0 1814 0 1 37300
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_319
timestamp 1704896540
transform 1 0 1814 0 1 36964
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_320
timestamp 1704896540
transform 1 0 1814 0 1 30580
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_321
timestamp 1704896540
transform 1 0 1814 0 1 36628
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_322
timestamp 1704896540
transform 1 0 1814 0 1 36292
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_323
timestamp 1704896540
transform 1 0 14855 0 1 32867
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_324
timestamp 1704896540
transform 1 0 14775 0 1 31309
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_325
timestamp 1704896540
transform 1 0 14695 0 1 30039
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_326
timestamp 1704896540
transform 1 0 14935 0 1 34137
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_327
timestamp 1704896540
transform 1 0 1814 0 1 46372
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_328
timestamp 1704896540
transform 1 0 1814 0 1 46036
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_329
timestamp 1704896540
transform 1 0 1814 0 1 45700
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_330
timestamp 1704896540
transform 1 0 1814 0 1 45364
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_331
timestamp 1704896540
transform 1 0 1814 0 1 45028
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_332
timestamp 1704896540
transform 1 0 1814 0 1 44692
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_333
timestamp 1704896540
transform 1 0 1814 0 1 44356
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_334
timestamp 1704896540
transform 1 0 1814 0 1 44020
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_335
timestamp 1704896540
transform 1 0 1814 0 1 43684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_336
timestamp 1704896540
transform 1 0 1814 0 1 40324
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_337
timestamp 1704896540
transform 1 0 1814 0 1 49060
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_338
timestamp 1704896540
transform 1 0 1814 0 1 41332
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_339
timestamp 1704896540
transform 1 0 1814 0 1 43012
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_340
timestamp 1704896540
transform 1 0 1814 0 1 40996
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_341
timestamp 1704896540
transform 1 0 1814 0 1 41668
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_342
timestamp 1704896540
transform 1 0 1814 0 1 48388
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_343
timestamp 1704896540
transform 1 0 1814 0 1 42676
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_344
timestamp 1704896540
transform 1 0 1814 0 1 47044
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_345
timestamp 1704896540
transform 1 0 1814 0 1 48052
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_346
timestamp 1704896540
transform 1 0 1814 0 1 42340
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_347
timestamp 1704896540
transform 1 0 1814 0 1 40660
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_348
timestamp 1704896540
transform 1 0 1814 0 1 47716
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_349
timestamp 1704896540
transform 1 0 1814 0 1 39988
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_350
timestamp 1704896540
transform 1 0 1814 0 1 46708
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_351
timestamp 1704896540
transform 1 0 1814 0 1 47380
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_352
timestamp 1704896540
transform 1 0 1814 0 1 42004
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_353
timestamp 1704896540
transform 1 0 1814 0 1 48724
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_354
timestamp 1704896540
transform 1 0 1814 0 1 49396
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_355
timestamp 1704896540
transform 1 0 1814 0 1 43348
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_356
timestamp 1704896540
transform 1 0 1814 0 1 59140
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_357
timestamp 1704896540
transform 1 0 1814 0 1 58804
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_358
timestamp 1704896540
transform 1 0 1814 0 1 58468
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_359
timestamp 1704896540
transform 1 0 1814 0 1 58132
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_360
timestamp 1704896540
transform 1 0 1814 0 1 57796
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_361
timestamp 1704896540
transform 1 0 1814 0 1 57460
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_362
timestamp 1704896540
transform 1 0 1814 0 1 57124
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_363
timestamp 1704896540
transform 1 0 1814 0 1 56788
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_364
timestamp 1704896540
transform 1 0 1814 0 1 56452
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_365
timestamp 1704896540
transform 1 0 1814 0 1 56116
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_366
timestamp 1704896540
transform 1 0 1814 0 1 55780
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_367
timestamp 1704896540
transform 1 0 1814 0 1 55444
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_368
timestamp 1704896540
transform 1 0 1814 0 1 55108
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_369
timestamp 1704896540
transform 1 0 1814 0 1 54772
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_370
timestamp 1704896540
transform 1 0 1814 0 1 54436
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_371
timestamp 1704896540
transform 1 0 1814 0 1 54100
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_372
timestamp 1704896540
transform 1 0 1814 0 1 53764
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_373
timestamp 1704896540
transform 1 0 1814 0 1 50068
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_374
timestamp 1704896540
transform 1 0 1814 0 1 50404
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_375
timestamp 1704896540
transform 1 0 1814 0 1 53428
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_376
timestamp 1704896540
transform 1 0 1814 0 1 49732
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_377
timestamp 1704896540
transform 1 0 1814 0 1 52084
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_378
timestamp 1704896540
transform 1 0 1814 0 1 53092
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_379
timestamp 1704896540
transform 1 0 1814 0 1 51748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_380
timestamp 1704896540
transform 1 0 1814 0 1 51412
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_381
timestamp 1704896540
transform 1 0 1814 0 1 51076
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_382
timestamp 1704896540
transform 1 0 1814 0 1 52756
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_383
timestamp 1704896540
transform 1 0 1814 0 1 52420
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_384
timestamp 1704896540
transform 1 0 1814 0 1 50740
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_385
timestamp 1704896540
transform 1 0 1814 0 1 59812
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_386
timestamp 1704896540
transform 1 0 1814 0 1 69220
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_387
timestamp 1704896540
transform 1 0 1814 0 1 68884
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_388
timestamp 1704896540
transform 1 0 1814 0 1 68548
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_389
timestamp 1704896540
transform 1 0 1814 0 1 68212
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_390
timestamp 1704896540
transform 1 0 1814 0 1 67876
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_391
timestamp 1704896540
transform 1 0 1814 0 1 67540
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_392
timestamp 1704896540
transform 1 0 1814 0 1 67204
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_393
timestamp 1704896540
transform 1 0 1814 0 1 66868
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_394
timestamp 1704896540
transform 1 0 1814 0 1 66532
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_395
timestamp 1704896540
transform 1 0 1814 0 1 66196
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_396
timestamp 1704896540
transform 1 0 1814 0 1 65860
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_397
timestamp 1704896540
transform 1 0 1814 0 1 65524
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_398
timestamp 1704896540
transform 1 0 1814 0 1 65188
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_399
timestamp 1704896540
transform 1 0 1814 0 1 64852
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_400
timestamp 1704896540
transform 1 0 1814 0 1 64516
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_401
timestamp 1704896540
transform 1 0 1814 0 1 64180
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_402
timestamp 1704896540
transform 1 0 1814 0 1 63844
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_403
timestamp 1704896540
transform 1 0 1814 0 1 63508
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_404
timestamp 1704896540
transform 1 0 1814 0 1 63172
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_405
timestamp 1704896540
transform 1 0 1814 0 1 62836
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_406
timestamp 1704896540
transform 1 0 1814 0 1 62500
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_407
timestamp 1704896540
transform 1 0 1814 0 1 62164
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_408
timestamp 1704896540
transform 1 0 1814 0 1 61828
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_409
timestamp 1704896540
transform 1 0 1814 0 1 61492
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_410
timestamp 1704896540
transform 1 0 1814 0 1 61156
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_411
timestamp 1704896540
transform 1 0 1814 0 1 60820
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_412
timestamp 1704896540
transform 1 0 1814 0 1 60484
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_413
timestamp 1704896540
transform 1 0 1814 0 1 60148
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_414
timestamp 1704896540
transform 1 0 1814 0 1 70228
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_415
timestamp 1704896540
transform 1 0 1814 0 1 69892
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_416
timestamp 1704896540
transform 1 0 1814 0 1 69556
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_417
timestamp 1704896540
transform 1 0 1814 0 1 70900
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_418
timestamp 1704896540
transform 1 0 1814 0 1 71572
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_419
timestamp 1704896540
transform 1 0 1814 0 1 73924
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_420
timestamp 1704896540
transform 1 0 1814 0 1 73588
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_421
timestamp 1704896540
transform 1 0 1814 0 1 73252
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_422
timestamp 1704896540
transform 1 0 1814 0 1 72916
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_423
timestamp 1704896540
transform 1 0 1814 0 1 72580
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_424
timestamp 1704896540
transform 1 0 1814 0 1 72244
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_425
timestamp 1704896540
transform 1 0 1814 0 1 71236
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_426
timestamp 1704896540
transform 1 0 1814 0 1 71908
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_427
timestamp 1704896540
transform 1 0 1814 0 1 70564
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_428
timestamp 1704896540
transform 1 0 3830 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_429
timestamp 1704896540
transform 1 0 1814 0 1 77284
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_430
timestamp 1704896540
transform 1 0 1814 0 1 76948
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_431
timestamp 1704896540
transform 1 0 1814 0 1 76612
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_432
timestamp 1704896540
transform 1 0 1814 0 1 76276
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_433
timestamp 1704896540
transform 1 0 1814 0 1 75940
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_434
timestamp 1704896540
transform 1 0 1814 0 1 75604
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_435
timestamp 1704896540
transform 1 0 1814 0 1 75268
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_436
timestamp 1704896540
transform 1 0 1814 0 1 74932
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_437
timestamp 1704896540
transform 1 0 1814 0 1 74596
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_438
timestamp 1704896540
transform 1 0 2150 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_439
timestamp 1704896540
transform 1 0 5510 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_440
timestamp 1704896540
transform 1 0 10550 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_441
timestamp 1704896540
transform 1 0 8870 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_442
timestamp 1704896540
transform 1 0 7190 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_443
timestamp 1704896540
transform 1 0 1814 0 1 74260
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_444
timestamp 1704896540
transform 1 0 15590 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_445
timestamp 1704896540
transform 1 0 13910 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_446
timestamp 1704896540
transform 1 0 12230 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_447
timestamp 1704896540
transform 1 0 17270 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_448
timestamp 1704896540
transform 1 0 23990 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_449
timestamp 1704896540
transform 1 0 22310 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_450
timestamp 1704896540
transform 1 0 20630 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_451
timestamp 1704896540
transform 1 0 18950 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_452
timestamp 1704896540
transform 1 0 35694 0 1 74043
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_453
timestamp 1704896540
transform 1 0 34446 0 1 74043
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_454
timestamp 1704896540
transform 1 0 33198 0 1 74043
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_455
timestamp 1704896540
transform 1 0 31950 0 1 74043
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_456
timestamp 1704896540
transform 1 0 30702 0 1 74043
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_457
timestamp 1704896540
transform 1 0 28206 0 1 74043
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_458
timestamp 1704896540
transform 1 0 29454 0 1 74043
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_459
timestamp 1704896540
transform 1 0 25670 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_460
timestamp 1704896540
transform 1 0 29030 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_461
timestamp 1704896540
transform 1 0 27350 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_462
timestamp 1704896540
transform 1 0 35750 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_463
timestamp 1704896540
transform 1 0 34070 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_464
timestamp 1704896540
transform 1 0 32390 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_465
timestamp 1704896540
transform 1 0 30710 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_466
timestamp 1704896540
transform 1 0 46926 0 1 74043
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_467
timestamp 1704896540
transform 1 0 45678 0 1 74043
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_468
timestamp 1704896540
transform 1 0 44430 0 1 74043
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_469
timestamp 1704896540
transform 1 0 43182 0 1 74043
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_470
timestamp 1704896540
transform 1 0 41934 0 1 74043
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_471
timestamp 1704896540
transform 1 0 40686 0 1 74043
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_472
timestamp 1704896540
transform 1 0 39438 0 1 74043
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_473
timestamp 1704896540
transform 1 0 38190 0 1 74043
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_474
timestamp 1704896540
transform 1 0 36942 0 1 74043
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_475
timestamp 1704896540
transform 1 0 40790 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_476
timestamp 1704896540
transform 1 0 39110 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_477
timestamp 1704896540
transform 1 0 37430 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_478
timestamp 1704896540
transform 1 0 42470 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_479
timestamp 1704896540
transform 1 0 47510 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_480
timestamp 1704896540
transform 1 0 45830 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_481
timestamp 1704896540
transform 1 0 44150 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_482
timestamp 1704896540
transform 1 0 1814 0 1 59476
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_483
timestamp 1704896540
transform 1 0 94172 0 1 46036
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_484
timestamp 1704896540
transform 1 0 94172 0 1 45700
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_485
timestamp 1704896540
transform 1 0 94172 0 1 45364
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_486
timestamp 1704896540
transform 1 0 94172 0 1 45028
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_487
timestamp 1704896540
transform 1 0 94172 0 1 44692
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_488
timestamp 1704896540
transform 1 0 94172 0 1 44356
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_489
timestamp 1704896540
transform 1 0 94172 0 1 44020
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_490
timestamp 1704896540
transform 1 0 94172 0 1 43684
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_491
timestamp 1704896540
transform 1 0 94172 0 1 43348
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_492
timestamp 1704896540
transform 1 0 94172 0 1 43012
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_493
timestamp 1704896540
transform 1 0 94172 0 1 42676
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_494
timestamp 1704896540
transform 1 0 94172 0 1 42340
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_495
timestamp 1704896540
transform 1 0 94172 0 1 42004
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_496
timestamp 1704896540
transform 1 0 94172 0 1 41668
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_497
timestamp 1704896540
transform 1 0 94172 0 1 40660
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_498
timestamp 1704896540
transform 1 0 94172 0 1 41332
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_499
timestamp 1704896540
transform 1 0 94172 0 1 40996
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_500
timestamp 1704896540
transform 1 0 94172 0 1 49396
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_501
timestamp 1704896540
transform 1 0 94172 0 1 49060
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_502
timestamp 1704896540
transform 1 0 94172 0 1 48724
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_503
timestamp 1704896540
transform 1 0 94172 0 1 48388
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_504
timestamp 1704896540
transform 1 0 94172 0 1 48052
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_505
timestamp 1704896540
transform 1 0 94172 0 1 47716
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_506
timestamp 1704896540
transform 1 0 94172 0 1 47380
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_507
timestamp 1704896540
transform 1 0 94172 0 1 47044
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_508
timestamp 1704896540
transform 1 0 94172 0 1 39988
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_509
timestamp 1704896540
transform 1 0 94172 0 1 46708
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_510
timestamp 1704896540
transform 1 0 94172 0 1 46372
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_511
timestamp 1704896540
transform 1 0 94172 0 1 40324
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_512
timestamp 1704896540
transform 1 0 94172 0 1 50740
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_513
timestamp 1704896540
transform 1 0 94172 0 1 50404
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_514
timestamp 1704896540
transform 1 0 94172 0 1 50068
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_515
timestamp 1704896540
transform 1 0 94172 0 1 49732
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_516
timestamp 1704896540
transform 1 0 94172 0 1 54436
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_517
timestamp 1704896540
transform 1 0 94172 0 1 54100
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_518
timestamp 1704896540
transform 1 0 94172 0 1 53764
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_519
timestamp 1704896540
transform 1 0 94172 0 1 53428
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_520
timestamp 1704896540
transform 1 0 94172 0 1 53092
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_521
timestamp 1704896540
transform 1 0 94172 0 1 52756
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_522
timestamp 1704896540
transform 1 0 94172 0 1 52420
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_523
timestamp 1704896540
transform 1 0 94172 0 1 52084
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_524
timestamp 1704896540
transform 1 0 94172 0 1 51748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_525
timestamp 1704896540
transform 1 0 94172 0 1 51412
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_526
timestamp 1704896540
transform 1 0 94172 0 1 51076
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_527
timestamp 1704896540
transform 1 0 94172 0 1 55780
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_528
timestamp 1704896540
transform 1 0 94172 0 1 55444
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_529
timestamp 1704896540
transform 1 0 94172 0 1 55108
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_530
timestamp 1704896540
transform 1 0 94172 0 1 54772
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_531
timestamp 1704896540
transform 1 0 94172 0 1 59140
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_532
timestamp 1704896540
transform 1 0 94172 0 1 58804
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_533
timestamp 1704896540
transform 1 0 94172 0 1 58468
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_534
timestamp 1704896540
transform 1 0 94172 0 1 58132
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_535
timestamp 1704896540
transform 1 0 94172 0 1 57796
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_536
timestamp 1704896540
transform 1 0 94172 0 1 57460
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_537
timestamp 1704896540
transform 1 0 94172 0 1 57124
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_538
timestamp 1704896540
transform 1 0 94172 0 1 56788
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_539
timestamp 1704896540
transform 1 0 94172 0 1 56452
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_540
timestamp 1704896540
transform 1 0 94172 0 1 56116
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_541
timestamp 1704896540
transform 1 0 55662 0 1 74043
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_542
timestamp 1704896540
transform 1 0 54414 0 1 74043
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_543
timestamp 1704896540
transform 1 0 59406 0 1 74043
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_544
timestamp 1704896540
transform 1 0 58158 0 1 74043
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_545
timestamp 1704896540
transform 1 0 56910 0 1 74043
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_546
timestamp 1704896540
transform 1 0 50670 0 1 74043
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_547
timestamp 1704896540
transform 1 0 49422 0 1 74043
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_548
timestamp 1704896540
transform 1 0 48174 0 1 74043
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_549
timestamp 1704896540
transform 1 0 53166 0 1 74043
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_550
timestamp 1704896540
transform 1 0 51918 0 1 74043
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_551
timestamp 1704896540
transform 1 0 52550 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_552
timestamp 1704896540
transform 1 0 50870 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_553
timestamp 1704896540
transform 1 0 49190 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_554
timestamp 1704896540
transform 1 0 59270 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_555
timestamp 1704896540
transform 1 0 57590 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_556
timestamp 1704896540
transform 1 0 55910 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_557
timestamp 1704896540
transform 1 0 54230 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_558
timestamp 1704896540
transform 1 0 66894 0 1 74043
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_559
timestamp 1704896540
transform 1 0 65646 0 1 74043
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_560
timestamp 1704896540
transform 1 0 64398 0 1 74043
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_561
timestamp 1704896540
transform 1 0 63150 0 1 74043
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_562
timestamp 1704896540
transform 1 0 61902 0 1 74043
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_563
timestamp 1704896540
transform 1 0 60654 0 1 74043
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_564
timestamp 1704896540
transform 1 0 60950 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_565
timestamp 1704896540
transform 1 0 62630 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_566
timestamp 1704896540
transform 1 0 64310 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_567
timestamp 1704896540
transform 1 0 71030 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_568
timestamp 1704896540
transform 1 0 69350 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_569
timestamp 1704896540
transform 1 0 67670 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_570
timestamp 1704896540
transform 1 0 65990 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_571
timestamp 1704896540
transform 1 0 94172 0 1 59812
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_572
timestamp 1704896540
transform 1 0 94172 0 1 60484
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_573
timestamp 1704896540
transform 1 0 94172 0 1 64180
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_574
timestamp 1704896540
transform 1 0 94172 0 1 63844
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_575
timestamp 1704896540
transform 1 0 94172 0 1 63508
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_576
timestamp 1704896540
transform 1 0 94172 0 1 63172
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_577
timestamp 1704896540
transform 1 0 94172 0 1 62836
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_578
timestamp 1704896540
transform 1 0 94172 0 1 62500
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_579
timestamp 1704896540
transform 1 0 94172 0 1 62164
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_580
timestamp 1704896540
transform 1 0 94172 0 1 61828
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_581
timestamp 1704896540
transform 1 0 94172 0 1 61492
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_582
timestamp 1704896540
transform 1 0 94172 0 1 60148
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_583
timestamp 1704896540
transform 1 0 94172 0 1 61156
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_584
timestamp 1704896540
transform 1 0 94172 0 1 60820
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_585
timestamp 1704896540
transform 1 0 94172 0 1 69220
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_586
timestamp 1704896540
transform 1 0 94172 0 1 68884
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_587
timestamp 1704896540
transform 1 0 94172 0 1 68548
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_588
timestamp 1704896540
transform 1 0 94172 0 1 68212
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_589
timestamp 1704896540
transform 1 0 94172 0 1 67876
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_590
timestamp 1704896540
transform 1 0 94172 0 1 67540
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_591
timestamp 1704896540
transform 1 0 94172 0 1 67204
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_592
timestamp 1704896540
transform 1 0 94172 0 1 66868
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_593
timestamp 1704896540
transform 1 0 94172 0 1 66532
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_594
timestamp 1704896540
transform 1 0 94172 0 1 66196
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_595
timestamp 1704896540
transform 1 0 94172 0 1 65860
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_596
timestamp 1704896540
transform 1 0 94172 0 1 65524
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_597
timestamp 1704896540
transform 1 0 94172 0 1 65188
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_598
timestamp 1704896540
transform 1 0 94172 0 1 64852
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_599
timestamp 1704896540
transform 1 0 94172 0 1 64516
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_600
timestamp 1704896540
transform 1 0 76070 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_601
timestamp 1704896540
transform 1 0 72710 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_602
timestamp 1704896540
transform 1 0 74390 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_603
timestamp 1704896540
transform 1 0 82790 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_604
timestamp 1704896540
transform 1 0 81110 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_605
timestamp 1704896540
transform 1 0 79430 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_606
timestamp 1704896540
transform 1 0 77750 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_607
timestamp 1704896540
transform 1 0 94172 0 1 71908
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_608
timestamp 1704896540
transform 1 0 94172 0 1 71572
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_609
timestamp 1704896540
transform 1 0 94172 0 1 71236
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_610
timestamp 1704896540
transform 1 0 94172 0 1 70900
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_611
timestamp 1704896540
transform 1 0 94172 0 1 70564
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_612
timestamp 1704896540
transform 1 0 94172 0 1 70228
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_613
timestamp 1704896540
transform 1 0 94172 0 1 69892
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_614
timestamp 1704896540
transform 1 0 94172 0 1 69556
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_615
timestamp 1704896540
transform 1 0 94172 0 1 73924
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_616
timestamp 1704896540
transform 1 0 94172 0 1 73588
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_617
timestamp 1704896540
transform 1 0 94172 0 1 73252
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_618
timestamp 1704896540
transform 1 0 94172 0 1 72916
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_619
timestamp 1704896540
transform 1 0 94172 0 1 72580
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_620
timestamp 1704896540
transform 1 0 94172 0 1 72244
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_621
timestamp 1704896540
transform 1 0 84470 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_622
timestamp 1704896540
transform 1 0 89510 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_623
timestamp 1704896540
transform 1 0 87830 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_624
timestamp 1704896540
transform 1 0 86150 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_625
timestamp 1704896540
transform 1 0 94172 0 1 77284
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_626
timestamp 1704896540
transform 1 0 94172 0 1 76948
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_627
timestamp 1704896540
transform 1 0 94172 0 1 76612
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_628
timestamp 1704896540
transform 1 0 94172 0 1 76276
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_629
timestamp 1704896540
transform 1 0 94172 0 1 75940
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_630
timestamp 1704896540
transform 1 0 94172 0 1 75604
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_631
timestamp 1704896540
transform 1 0 94172 0 1 75268
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_632
timestamp 1704896540
transform 1 0 94172 0 1 74932
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_633
timestamp 1704896540
transform 1 0 94172 0 1 74596
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_634
timestamp 1704896540
transform 1 0 92870 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_635
timestamp 1704896540
transform 1 0 91190 0 1 77748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_636
timestamp 1704896540
transform 1 0 94172 0 1 74260
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_637
timestamp 1704896540
transform 1 0 94172 0 1 59476
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_33  sky130_sram_1kbyte_1rw1r_32x256_8_contact_33_0
timestamp 1704896540
transform 1 0 81839 0 1 16805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_33  sky130_sram_1kbyte_1rw1r_32x256_8_contact_33_1
timestamp 1704896540
transform 1 0 14337 0 1 2659
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_33  sky130_sram_1kbyte_1rw1r_32x256_8_contact_33_2
timestamp 1704896540
transform 1 0 14337 0 1 25321
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_33  sky130_sram_1kbyte_1rw1r_32x256_8_contact_33_3
timestamp 1704896540
transform 1 0 81839 0 1 76038
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_0
timestamp 1704896540
transform 1 0 94656 0 1 3677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1
timestamp 1704896540
transform 1 0 94656 0 1 1909
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2
timestamp 1704896540
transform 1 0 92752 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_3
timestamp 1704896540
transform 1 0 92752 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_4
timestamp 1704896540
transform 1 0 91120 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_5
timestamp 1704896540
transform 1 0 91120 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_6
timestamp 1704896540
transform 1 0 89488 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_7
timestamp 1704896540
transform 1 0 89488 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_8
timestamp 1704896540
transform 1 0 87720 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_9
timestamp 1704896540
transform 1 0 87720 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_10
timestamp 1704896540
transform 1 0 86224 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_11
timestamp 1704896540
transform 1 0 86224 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_12
timestamp 1704896540
transform 1 0 84456 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_13
timestamp 1704896540
transform 1 0 84456 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_14
timestamp 1704896540
transform 1 0 94656 0 1 5309
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_15
timestamp 1704896540
transform 1 0 94656 0 1 6941
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_16
timestamp 1704896540
transform 1 0 94656 0 1 8845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_17
timestamp 1704896540
transform 1 0 82552 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_18
timestamp 1704896540
transform 1 0 82552 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_19
timestamp 1704896540
transform 1 0 81192 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_20
timestamp 1704896540
transform 1 0 81192 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_21
timestamp 1704896540
transform 1 0 79424 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_22
timestamp 1704896540
transform 1 0 79424 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_23
timestamp 1704896540
transform 1 0 74256 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_24
timestamp 1704896540
transform 1 0 74256 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_25
timestamp 1704896540
transform 1 0 72624 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_26
timestamp 1704896540
transform 1 0 72624 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_27
timestamp 1704896540
transform 1 0 77656 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_28
timestamp 1704896540
transform 1 0 77656 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_29
timestamp 1704896540
transform 1 0 76160 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_30
timestamp 1704896540
transform 1 0 76160 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_31
timestamp 1704896540
transform 1 0 82824 0 1 9117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_32
timestamp 1704896540
transform 1 0 82960 0 1 8029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_33
timestamp 1704896540
transform 1 0 82552 0 1 8709
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_34
timestamp 1704896540
transform 1 0 82416 0 1 10069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_35
timestamp 1704896540
transform 1 0 82416 0 1 9933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_36
timestamp 1704896540
transform 1 0 82416 0 1 7349
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_37
timestamp 1704896540
transform 1 0 82416 0 1 17005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_38
timestamp 1704896540
transform 1 0 82416 0 1 14421
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_39
timestamp 1704896540
transform 1 0 82280 0 1 11565
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_40
timestamp 1704896540
transform 1 0 82280 0 1 14149
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_41
timestamp 1704896540
transform 1 0 82552 0 1 11429
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_42
timestamp 1704896540
transform 1 0 82416 0 1 17141
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_43
timestamp 1704896540
transform 1 0 82416 0 1 17413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_44
timestamp 1704896540
transform 1 0 78608 0 1 17549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_45
timestamp 1704896540
transform 1 0 78608 0 1 18229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_46
timestamp 1704896540
transform 1 0 78608 0 1 18365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_47
timestamp 1704896540
transform 1 0 78608 0 1 19861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_48
timestamp 1704896540
transform 1 0 78472 0 1 18365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_49
timestamp 1704896540
transform 1 0 78472 0 1 18637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_50
timestamp 1704896540
transform 1 0 77928 0 1 18637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_51
timestamp 1704896540
transform 1 0 77928 0 1 18365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_52
timestamp 1704896540
transform 1 0 74392 0 1 18229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_53
timestamp 1704896540
transform 1 0 73984 0 1 18229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_54
timestamp 1704896540
transform 1 0 73984 0 1 17957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_55
timestamp 1704896540
transform 1 0 75616 0 1 18637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_56
timestamp 1704896540
transform 1 0 75616 0 1 18365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_57
timestamp 1704896540
transform 1 0 82416 0 1 12789
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_58
timestamp 1704896540
transform 1 0 82552 0 1 12925
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_59
timestamp 1704896540
transform 1 0 82552 0 1 15645
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_60
timestamp 1704896540
transform 1 0 79696 0 1 15781
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_61
timestamp 1704896540
transform 1 0 79696 0 1 17413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_62
timestamp 1704896540
transform 1 0 74392 0 1 17957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_63
timestamp 1704896540
transform 1 0 75072 0 1 18365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_64
timestamp 1704896540
transform 1 0 75072 0 1 17957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_65
timestamp 1704896540
transform 1 0 75072 0 1 18229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_66
timestamp 1704896540
transform 1 0 75616 0 1 17821
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_67
timestamp 1704896540
transform 1 0 75616 0 1 17549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_68
timestamp 1704896540
transform 1 0 79424 0 1 17549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_69
timestamp 1704896540
transform 1 0 79424 0 1 18093
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_70
timestamp 1704896540
transform 1 0 78200 0 1 19861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_71
timestamp 1704896540
transform 1 0 78200 0 1 18365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_72
timestamp 1704896540
transform 1 0 75616 0 1 19589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_73
timestamp 1704896540
transform 1 0 75616 0 1 19861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_74
timestamp 1704896540
transform 1 0 74800 0 1 17821
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_75
timestamp 1704896540
transform 1 0 75480 0 1 18773
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_76
timestamp 1704896540
transform 1 0 75480 0 1 19045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_77
timestamp 1704896540
transform 1 0 75480 0 1 19453
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_78
timestamp 1704896540
transform 1 0 75480 0 1 19181
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_79
timestamp 1704896540
transform 1 0 74664 0 1 17957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_80
timestamp 1704896540
transform 1 0 73848 0 1 17821
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_81
timestamp 1704896540
transform 1 0 73848 0 1 17549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_82
timestamp 1704896540
transform 1 0 74664 0 1 18229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_83
timestamp 1704896540
transform 1 0 77384 0 1 18229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_84
timestamp 1704896540
transform 1 0 77384 0 1 17549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_85
timestamp 1704896540
transform 1 0 73848 0 1 19045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_86
timestamp 1704896540
transform 1 0 73848 0 1 18773
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_87
timestamp 1704896540
transform 1 0 73848 0 1 18365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_88
timestamp 1704896540
transform 1 0 73848 0 1 18637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_89
timestamp 1704896540
transform 1 0 74800 0 1 17549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_90
timestamp 1704896540
transform 1 0 74936 0 1 17821
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_91
timestamp 1704896540
transform 1 0 74800 0 1 19045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_92
timestamp 1704896540
transform 1 0 75208 0 1 19181
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_93
timestamp 1704896540
transform 1 0 75208 0 1 19453
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_94
timestamp 1704896540
transform 1 0 74800 0 1 18773
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_95
timestamp 1704896540
transform 1 0 74256 0 1 19045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_96
timestamp 1704896540
transform 1 0 74256 0 1 18773
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_97
timestamp 1704896540
transform 1 0 74256 0 1 19589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_98
timestamp 1704896540
transform 1 0 74256 0 1 19861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_99
timestamp 1704896540
transform 1 0 73848 0 1 19861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_100
timestamp 1704896540
transform 1 0 73848 0 1 19589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_101
timestamp 1704896540
transform 1 0 73848 0 1 19181
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_102
timestamp 1704896540
transform 1 0 73848 0 1 19453
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_103
timestamp 1704896540
transform 1 0 74256 0 1 17821
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_104
timestamp 1704896540
transform 1 0 74256 0 1 17549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_105
timestamp 1704896540
transform 1 0 74256 0 1 19453
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_106
timestamp 1704896540
transform 1 0 74256 0 1 19181
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_107
timestamp 1704896540
transform 1 0 82688 0 1 10885
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_108
timestamp 1704896540
transform 1 0 75072 0 1 18637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_109
timestamp 1704896540
transform 1 0 83096 0 1 11973
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_110
timestamp 1704896540
transform 1 0 74256 0 1 18365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_111
timestamp 1704896540
transform 1 0 74936 0 1 17549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_112
timestamp 1704896540
transform 1 0 74256 0 1 18637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_113
timestamp 1704896540
transform 1 0 94656 0 1 13877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_114
timestamp 1704896540
transform 1 0 94656 0 1 18773
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_115
timestamp 1704896540
transform 1 0 94656 0 1 15373
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_116
timestamp 1704896540
transform 1 0 94656 0 1 17005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_117
timestamp 1704896540
transform 1 0 94656 0 1 12245
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_118
timestamp 1704896540
transform 1 0 94656 0 1 10477
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_119
timestamp 1704896540
transform 1 0 69224 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_120
timestamp 1704896540
transform 1 0 65960 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_121
timestamp 1704896540
transform 1 0 65960 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_122
timestamp 1704896540
transform 1 0 69224 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_123
timestamp 1704896540
transform 1 0 67728 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_124
timestamp 1704896540
transform 1 0 67728 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_125
timestamp 1704896540
transform 1 0 70992 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_126
timestamp 1704896540
transform 1 0 70992 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_127
timestamp 1704896540
transform 1 0 64056 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_128
timestamp 1704896540
transform 1 0 60928 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_129
timestamp 1704896540
transform 1 0 60928 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_130
timestamp 1704896540
transform 1 0 64056 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_131
timestamp 1704896540
transform 1 0 62696 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_132
timestamp 1704896540
transform 1 0 62696 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_133
timestamp 1704896540
transform 1 0 64736 0 1 10069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_134
timestamp 1704896540
transform 1 0 64736 0 1 9797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_135
timestamp 1704896540
transform 1 0 64736 0 1 8981
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_136
timestamp 1704896540
transform 1 0 62152 0 1 9389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_137
timestamp 1704896540
transform 1 0 63512 0 1 10069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_138
timestamp 1704896540
transform 1 0 63512 0 1 9253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_139
timestamp 1704896540
transform 1 0 63512 0 1 9797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_140
timestamp 1704896540
transform 1 0 62968 0 1 10069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_141
timestamp 1704896540
transform 1 0 62152 0 1 10069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_142
timestamp 1704896540
transform 1 0 62288 0 1 9253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_143
timestamp 1704896540
transform 1 0 62288 0 1 9797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_144
timestamp 1704896540
transform 1 0 61744 0 1 10069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_145
timestamp 1704896540
transform 1 0 65416 0 1 10069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_146
timestamp 1704896540
transform 1 0 60928 0 1 10069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_147
timestamp 1704896540
transform 1 0 60928 0 1 9253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_148
timestamp 1704896540
transform 1 0 60928 0 1 9797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_149
timestamp 1704896540
transform 1 0 63376 0 1 8573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_150
timestamp 1704896540
transform 1 0 63376 0 1 9389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_151
timestamp 1704896540
transform 1 0 64600 0 1 9389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_152
timestamp 1704896540
transform 1 0 60792 0 1 8573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_153
timestamp 1704896540
transform 1 0 65688 0 1 8573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_154
timestamp 1704896540
transform 1 0 60792 0 1 9389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_155
timestamp 1704896540
transform 1 0 64600 0 1 8573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_156
timestamp 1704896540
transform 1 0 65688 0 1 9389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_157
timestamp 1704896540
transform 1 0 62152 0 1 8573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_158
timestamp 1704896540
transform 1 0 68000 0 1 8845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_159
timestamp 1704896540
transform 1 0 65960 0 1 10069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_160
timestamp 1704896540
transform 1 0 68000 0 1 7077
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_161
timestamp 1704896540
transform 1 0 67048 0 1 9389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_162
timestamp 1704896540
transform 1 0 67048 0 1 10069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_163
timestamp 1704896540
transform 1 0 67184 0 1 9253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_164
timestamp 1704896540
transform 1 0 67184 0 1 9797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_165
timestamp 1704896540
transform 1 0 67864 0 1 8165
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_166
timestamp 1704896540
transform 1 0 67864 0 1 8573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_167
timestamp 1704896540
transform 1 0 67048 0 1 8573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_168
timestamp 1704896540
transform 1 0 65824 0 1 9253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_169
timestamp 1704896540
transform 1 0 65824 0 1 9797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_170
timestamp 1704896540
transform 1 0 55896 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_171
timestamp 1704896540
transform 1 0 55896 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_172
timestamp 1704896540
transform 1 0 59160 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_173
timestamp 1704896540
transform 1 0 59160 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_174
timestamp 1704896540
transform 1 0 57528 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_175
timestamp 1704896540
transform 1 0 57528 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_176
timestamp 1704896540
transform 1 0 57664 0 1 2861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_177
timestamp 1704896540
transform 1 0 56576 0 1 2861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_178
timestamp 1704896540
transform 1 0 55216 0 1 2861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_179
timestamp 1704896540
transform 1 0 53992 0 1 2861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_180
timestamp 1704896540
transform 1 0 54264 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_181
timestamp 1704896540
transform 1 0 54264 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_182
timestamp 1704896540
transform 1 0 51000 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_183
timestamp 1704896540
transform 1 0 51000 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_184
timestamp 1704896540
transform 1 0 52632 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_185
timestamp 1704896540
transform 1 0 52632 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_186
timestamp 1704896540
transform 1 0 48960 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_187
timestamp 1704896540
transform 1 0 48960 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_188
timestamp 1704896540
transform 1 0 52904 0 1 2861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_189
timestamp 1704896540
transform 1 0 51816 0 1 2861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_190
timestamp 1704896540
transform 1 0 50728 0 1 2861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_191
timestamp 1704896540
transform 1 0 49368 0 1 2861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_192
timestamp 1704896540
transform 1 0 48280 0 1 2861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_193
timestamp 1704896540
transform 1 0 48280 0 1 9389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_194
timestamp 1704896540
transform 1 0 51000 0 1 10069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_195
timestamp 1704896540
transform 1 0 50864 0 1 9253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_196
timestamp 1704896540
transform 1 0 50864 0 1 9797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_197
timestamp 1704896540
transform 1 0 49776 0 1 10069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_198
timestamp 1704896540
transform 1 0 49776 0 1 9253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_199
timestamp 1704896540
transform 1 0 49776 0 1 9797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_200
timestamp 1704896540
transform 1 0 48416 0 1 10069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_201
timestamp 1704896540
transform 1 0 48416 0 1 9253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_202
timestamp 1704896540
transform 1 0 48416 0 1 9797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_203
timestamp 1704896540
transform 1 0 49640 0 1 8573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_204
timestamp 1704896540
transform 1 0 49640 0 1 9389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_205
timestamp 1704896540
transform 1 0 48280 0 1 8573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_206
timestamp 1704896540
transform 1 0 53448 0 1 8573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_207
timestamp 1704896540
transform 1 0 53448 0 1 9389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_208
timestamp 1704896540
transform 1 0 51952 0 1 8573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_209
timestamp 1704896540
transform 1 0 51952 0 1 9389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_210
timestamp 1704896540
transform 1 0 50728 0 1 8573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_211
timestamp 1704896540
transform 1 0 50728 0 1 9389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_212
timestamp 1704896540
transform 1 0 53448 0 1 10069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_213
timestamp 1704896540
transform 1 0 53584 0 1 9253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_214
timestamp 1704896540
transform 1 0 53584 0 1 9797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_215
timestamp 1704896540
transform 1 0 52224 0 1 10069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_216
timestamp 1704896540
transform 1 0 52088 0 1 9797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_217
timestamp 1704896540
transform 1 0 52088 0 1 8981
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_218
timestamp 1704896540
transform 1 0 59704 0 1 10069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_219
timestamp 1704896540
transform 1 0 59704 0 1 9253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_220
timestamp 1704896540
transform 1 0 59704 0 1 9797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_221
timestamp 1704896540
transform 1 0 59160 0 1 10069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_222
timestamp 1704896540
transform 1 0 58480 0 1 10069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_223
timestamp 1704896540
transform 1 0 58480 0 1 9253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_224
timestamp 1704896540
transform 1 0 58480 0 1 9797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_225
timestamp 1704896540
transform 1 0 57256 0 1 10069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_226
timestamp 1704896540
transform 1 0 57120 0 1 9253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_227
timestamp 1704896540
transform 1 0 57120 0 1 9797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_228
timestamp 1704896540
transform 1 0 56712 0 1 9797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_229
timestamp 1704896540
transform 1 0 56712 0 1 9253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_230
timestamp 1704896540
transform 1 0 55896 0 1 10069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_231
timestamp 1704896540
transform 1 0 56032 0 1 9253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_232
timestamp 1704896540
transform 1 0 56032 0 1 9797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_233
timestamp 1704896540
transform 1 0 54672 0 1 10069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_234
timestamp 1704896540
transform 1 0 54672 0 1 9253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_235
timestamp 1704896540
transform 1 0 54672 0 1 9797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_236
timestamp 1704896540
transform 1 0 59568 0 1 8573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_237
timestamp 1704896540
transform 1 0 59568 0 1 9389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_238
timestamp 1704896540
transform 1 0 58344 0 1 8573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_239
timestamp 1704896540
transform 1 0 58344 0 1 9389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_240
timestamp 1704896540
transform 1 0 56984 0 1 8573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_241
timestamp 1704896540
transform 1 0 56984 0 1 9389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_242
timestamp 1704896540
transform 1 0 55896 0 1 8573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_243
timestamp 1704896540
transform 1 0 55896 0 1 9389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_244
timestamp 1704896540
transform 1 0 54536 0 1 8573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_245
timestamp 1704896540
transform 1 0 54536 0 1 9389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_246
timestamp 1704896540
transform 1 0 59296 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_247
timestamp 1704896540
transform 1 0 57800 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_248
timestamp 1704896540
transform 1 0 56848 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_249
timestamp 1704896540
transform 1 0 55624 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_250
timestamp 1704896540
transform 1 0 54400 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_251
timestamp 1704896540
transform 1 0 59704 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_252
timestamp 1704896540
transform 1 0 59160 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_253
timestamp 1704896540
transform 1 0 58480 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_254
timestamp 1704896540
transform 1 0 57256 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_255
timestamp 1704896540
transform 1 0 55896 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_256
timestamp 1704896540
transform 1 0 54672 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_257
timestamp 1704896540
transform 1 0 53448 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_258
timestamp 1704896540
transform 1 0 52224 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_259
timestamp 1704896540
transform 1 0 51000 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_260
timestamp 1704896540
transform 1 0 49776 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_261
timestamp 1704896540
transform 1 0 49640 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_262
timestamp 1704896540
transform 1 0 49640 0 1 10341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_263
timestamp 1704896540
transform 1 0 48960 0 1 10341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_264
timestamp 1704896540
transform 1 0 48960 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_265
timestamp 1704896540
transform 1 0 48416 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_266
timestamp 1704896540
transform 1 0 53176 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_267
timestamp 1704896540
transform 1 0 51408 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_268
timestamp 1704896540
transform 1 0 50592 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_269
timestamp 1704896540
transform 1 0 49096 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_270
timestamp 1704896540
transform 1 0 59704 0 1 11157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_271
timestamp 1704896540
transform 1 0 59704 0 1 11837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_272
timestamp 1704896540
transform 1 0 59568 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_273
timestamp 1704896540
transform 1 0 59568 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_274
timestamp 1704896540
transform 1 0 59024 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_275
timestamp 1704896540
transform 1 0 59024 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_276
timestamp 1704896540
transform 1 0 58480 0 1 11157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_277
timestamp 1704896540
transform 1 0 58480 0 1 11837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_278
timestamp 1704896540
transform 1 0 57936 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_279
timestamp 1704896540
transform 1 0 57936 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_280
timestamp 1704896540
transform 1 0 57800 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_281
timestamp 1704896540
transform 1 0 57800 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_282
timestamp 1704896540
transform 1 0 58072 0 1 15917
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_283
timestamp 1704896540
transform 1 0 58072 0 1 11973
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_284
timestamp 1704896540
transform 1 0 57120 0 1 11157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_285
timestamp 1704896540
transform 1 0 57120 0 1 11837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_286
timestamp 1704896540
transform 1 0 56984 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_287
timestamp 1704896540
transform 1 0 56984 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_288
timestamp 1704896540
transform 1 0 56440 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_289
timestamp 1704896540
transform 1 0 56440 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_290
timestamp 1704896540
transform 1 0 56032 0 1 11157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_291
timestamp 1704896540
transform 1 0 56032 0 1 11837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_292
timestamp 1704896540
transform 1 0 55760 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_293
timestamp 1704896540
transform 1 0 55760 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_294
timestamp 1704896540
transform 1 0 55352 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_295
timestamp 1704896540
transform 1 0 55352 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_296
timestamp 1704896540
transform 1 0 54536 0 1 11157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_297
timestamp 1704896540
transform 1 0 54536 0 1 11837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_298
timestamp 1704896540
transform 1 0 54536 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_299
timestamp 1704896540
transform 1 0 54536 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_300
timestamp 1704896540
transform 1 0 53992 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_301
timestamp 1704896540
transform 1 0 53992 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_302
timestamp 1704896540
transform 1 0 53448 0 1 11157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_303
timestamp 1704896540
transform 1 0 53448 0 1 11837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_304
timestamp 1704896540
transform 1 0 53312 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_305
timestamp 1704896540
transform 1 0 53312 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_306
timestamp 1704896540
transform 1 0 52088 0 1 11157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_307
timestamp 1704896540
transform 1 0 52088 0 1 11837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_308
timestamp 1704896540
transform 1 0 51952 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_309
timestamp 1704896540
transform 1 0 51952 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_310
timestamp 1704896540
transform 1 0 51544 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_311
timestamp 1704896540
transform 1 0 51544 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_312
timestamp 1704896540
transform 1 0 51000 0 1 11157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_313
timestamp 1704896540
transform 1 0 51000 0 1 11837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_314
timestamp 1704896540
transform 1 0 50728 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_315
timestamp 1704896540
transform 1 0 50728 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_316
timestamp 1704896540
transform 1 0 50320 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_317
timestamp 1704896540
transform 1 0 50320 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_318
timestamp 1704896540
transform 1 0 49776 0 1 11157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_319
timestamp 1704896540
transform 1 0 49776 0 1 11837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_320
timestamp 1704896540
transform 1 0 49368 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_321
timestamp 1704896540
transform 1 0 49368 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_322
timestamp 1704896540
transform 1 0 48416 0 1 11157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_323
timestamp 1704896540
transform 1 0 48416 0 1 11837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_324
timestamp 1704896540
transform 1 0 48280 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_325
timestamp 1704896540
transform 1 0 48280 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_326
timestamp 1704896540
transform 1 0 64736 0 1 10749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_327
timestamp 1704896540
transform 1 0 64736 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_328
timestamp 1704896540
transform 1 0 63512 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_329
timestamp 1704896540
transform 1 0 62968 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_330
timestamp 1704896540
transform 1 0 62152 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_331
timestamp 1704896540
transform 1 0 61744 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_332
timestamp 1704896540
transform 1 0 60928 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_333
timestamp 1704896540
transform 1 0 63376 0 1 11157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_334
timestamp 1704896540
transform 1 0 63376 0 1 11837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_335
timestamp 1704896540
transform 1 0 63240 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_336
timestamp 1704896540
transform 1 0 63240 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_337
timestamp 1704896540
transform 1 0 62152 0 1 11157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_338
timestamp 1704896540
transform 1 0 62152 0 1 11837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_339
timestamp 1704896540
transform 1 0 62016 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_340
timestamp 1704896540
transform 1 0 62016 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_341
timestamp 1704896540
transform 1 0 60792 0 1 11157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_342
timestamp 1704896540
transform 1 0 60792 0 1 11837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_343
timestamp 1704896540
transform 1 0 60792 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_344
timestamp 1704896540
transform 1 0 60792 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_345
timestamp 1704896540
transform 1 0 60248 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_346
timestamp 1704896540
transform 1 0 60248 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_347
timestamp 1704896540
transform 1 0 66776 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_348
timestamp 1704896540
transform 1 0 65552 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_349
timestamp 1704896540
transform 1 0 64328 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_350
timestamp 1704896540
transform 1 0 63104 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_351
timestamp 1704896540
transform 1 0 61880 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_352
timestamp 1704896540
transform 1 0 60520 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_353
timestamp 1704896540
transform 1 0 64600 0 1 12653
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_354
timestamp 1704896540
transform 1 0 68272 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_355
timestamp 1704896540
transform 1 0 68272 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_356
timestamp 1704896540
transform 1 0 67728 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_357
timestamp 1704896540
transform 1 0 67728 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_358
timestamp 1704896540
transform 1 0 67184 0 1 11157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_359
timestamp 1704896540
transform 1 0 67184 0 1 11837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_360
timestamp 1704896540
transform 1 0 67048 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_361
timestamp 1704896540
transform 1 0 67048 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_362
timestamp 1704896540
transform 1 0 66504 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_363
timestamp 1704896540
transform 1 0 66504 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_364
timestamp 1704896540
transform 1 0 65824 0 1 11157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_365
timestamp 1704896540
transform 1 0 65824 0 1 11837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_366
timestamp 1704896540
transform 1 0 65688 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_367
timestamp 1704896540
transform 1 0 65688 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_368
timestamp 1704896540
transform 1 0 65280 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_369
timestamp 1704896540
transform 1 0 65280 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_370
timestamp 1704896540
transform 1 0 64736 0 1 11157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_371
timestamp 1704896540
transform 1 0 64736 0 1 11837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_372
timestamp 1704896540
transform 1 0 64192 0 1 16597
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_373
timestamp 1704896540
transform 1 0 69088 0 1 19589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_374
timestamp 1704896540
transform 1 0 64192 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_375
timestamp 1704896540
transform 1 0 67048 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_376
timestamp 1704896540
transform 1 0 65960 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_377
timestamp 1704896540
transform 1 0 65416 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_378
timestamp 1704896540
transform 1 0 68952 0 1 28701
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_379
timestamp 1704896540
transform 1 0 68952 0 1 28429
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_380
timestamp 1704896540
transform 1 0 68952 0 1 21493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_381
timestamp 1704896540
transform 1 0 68952 0 1 21085
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_382
timestamp 1704896540
transform 1 0 69088 0 1 28701
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_383
timestamp 1704896540
transform 1 0 69088 0 1 28293
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_384
timestamp 1704896540
transform 1 0 69088 0 1 20541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_385
timestamp 1704896540
transform 1 0 69088 0 1 20813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_386
timestamp 1704896540
transform 1 0 69088 0 1 36181
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_387
timestamp 1704896540
transform 1 0 69088 0 1 35909
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_388
timestamp 1704896540
transform 1 0 68952 0 1 37133
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_389
timestamp 1704896540
transform 1 0 68952 0 1 37405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_390
timestamp 1704896540
transform 1 0 68952 0 1 23261
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_391
timestamp 1704896540
transform 1 0 68952 0 1 23533
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_392
timestamp 1704896540
transform 1 0 68952 0 1 36997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_393
timestamp 1704896540
transform 1 0 69088 0 1 21357
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_394
timestamp 1704896540
transform 1 0 69088 0 1 21765
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_395
timestamp 1704896540
transform 1 0 68952 0 1 24485
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_396
timestamp 1704896540
transform 1 0 68952 0 1 24757
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_397
timestamp 1704896540
transform 1 0 69088 0 1 27477
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_398
timestamp 1704896540
transform 1 0 69088 0 1 27205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_399
timestamp 1704896540
transform 1 0 68952 0 1 24077
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_400
timestamp 1704896540
transform 1 0 68952 0 1 24349
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_401
timestamp 1704896540
transform 1 0 68952 0 1 32781
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_402
timestamp 1704896540
transform 1 0 68952 0 1 33053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_403
timestamp 1704896540
transform 1 0 68952 0 1 28837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_404
timestamp 1704896540
transform 1 0 68952 0 1 29109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_405
timestamp 1704896540
transform 1 0 68952 0 1 36725
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_406
timestamp 1704896540
transform 1 0 94656 0 1 23805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_407
timestamp 1704896540
transform 1 0 94656 0 1 28973
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_408
timestamp 1704896540
transform 1 0 94656 0 1 20405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_409
timestamp 1704896540
transform 1 0 94656 0 1 22309
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_410
timestamp 1704896540
transform 1 0 94656 0 1 27341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_411
timestamp 1704896540
transform 1 0 94656 0 1 25437
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_412
timestamp 1704896540
transform 1 0 78064 0 1 24621
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_413
timestamp 1704896540
transform 1 0 78200 0 1 20541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_414
timestamp 1704896540
transform 1 0 79424 0 1 20405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_415
timestamp 1704896540
transform 1 0 79016 0 1 24621
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_416
timestamp 1704896540
transform 1 0 79016 0 1 23941
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_417
timestamp 1704896540
transform 1 0 79016 0 1 23805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_418
timestamp 1704896540
transform 1 0 79016 0 1 23125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_419
timestamp 1704896540
transform 1 0 78880 0 1 22309
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_420
timestamp 1704896540
transform 1 0 78880 0 1 22989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_421
timestamp 1704896540
transform 1 0 78608 0 1 22989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_422
timestamp 1704896540
transform 1 0 78608 0 1 20541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_423
timestamp 1704896540
transform 1 0 78608 0 1 22309
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_424
timestamp 1704896540
transform 1 0 78472 0 1 20813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_425
timestamp 1704896540
transform 1 0 78472 0 1 22037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_426
timestamp 1704896540
transform 1 0 78336 0 1 23125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_427
timestamp 1704896540
transform 1 0 78336 0 1 23805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_428
timestamp 1704896540
transform 1 0 78064 0 1 23941
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_429
timestamp 1704896540
transform 1 0 73848 0 1 22989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_430
timestamp 1704896540
transform 1 0 73848 0 1 22717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_431
timestamp 1704896540
transform 1 0 74664 0 1 24621
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_432
timestamp 1704896540
transform 1 0 75480 0 1 22581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_433
timestamp 1704896540
transform 1 0 75480 0 1 22309
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_434
timestamp 1704896540
transform 1 0 74392 0 1 21357
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_435
timestamp 1704896540
transform 1 0 74664 0 1 22309
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_436
timestamp 1704896540
transform 1 0 75480 0 1 20269
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_437
timestamp 1704896540
transform 1 0 74392 0 1 21085
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_438
timestamp 1704896540
transform 1 0 74936 0 1 24077
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_439
timestamp 1704896540
transform 1 0 74392 0 1 24213
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_440
timestamp 1704896540
transform 1 0 77656 0 1 20541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_441
timestamp 1704896540
transform 1 0 74392 0 1 23941
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_442
timestamp 1704896540
transform 1 0 77656 0 1 23805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_443
timestamp 1704896540
transform 1 0 77656 0 1 23261
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_444
timestamp 1704896540
transform 1 0 75616 0 1 22717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_445
timestamp 1704896540
transform 1 0 75616 0 1 22989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_446
timestamp 1704896540
transform 1 0 74392 0 1 23533
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_447
timestamp 1704896540
transform 1 0 74392 0 1 23805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_448
timestamp 1704896540
transform 1 0 74392 0 1 22989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_449
timestamp 1704896540
transform 1 0 74392 0 1 22717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_450
timestamp 1704896540
transform 1 0 74664 0 1 20677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_451
timestamp 1704896540
transform 1 0 74256 0 1 22309
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_452
timestamp 1704896540
transform 1 0 74256 0 1 22581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_453
timestamp 1704896540
transform 1 0 75480 0 1 24621
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_454
timestamp 1704896540
transform 1 0 75480 0 1 24349
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_455
timestamp 1704896540
transform 1 0 74936 0 1 23805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_456
timestamp 1704896540
transform 1 0 75480 0 1 20677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_457
timestamp 1704896540
transform 1 0 75480 0 1 20405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_458
timestamp 1704896540
transform 1 0 73984 0 1 23125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_459
timestamp 1704896540
transform 1 0 73984 0 1 23397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_460
timestamp 1704896540
transform 1 0 73984 0 1 23805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_461
timestamp 1704896540
transform 1 0 75616 0 1 24213
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_462
timestamp 1704896540
transform 1 0 75616 0 1 23941
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_463
timestamp 1704896540
transform 1 0 75616 0 1 24757
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_464
timestamp 1704896540
transform 1 0 73984 0 1 23533
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_465
timestamp 1704896540
transform 1 0 73848 0 1 23941
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_466
timestamp 1704896540
transform 1 0 74664 0 1 22581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_467
timestamp 1704896540
transform 1 0 73848 0 1 21765
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_468
timestamp 1704896540
transform 1 0 74664 0 1 20405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_469
timestamp 1704896540
transform 1 0 74256 0 1 23125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_470
timestamp 1704896540
transform 1 0 74256 0 1 23397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_471
timestamp 1704896540
transform 1 0 75480 0 1 20813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_472
timestamp 1704896540
transform 1 0 75480 0 1 21085
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_473
timestamp 1704896540
transform 1 0 74936 0 1 22173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_474
timestamp 1704896540
transform 1 0 74936 0 1 21901
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_475
timestamp 1704896540
transform 1 0 75208 0 1 23533
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_476
timestamp 1704896540
transform 1 0 74800 0 1 22173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_477
timestamp 1704896540
transform 1 0 74800 0 1 21901
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_478
timestamp 1704896540
transform 1 0 74800 0 1 23397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_479
timestamp 1704896540
transform 1 0 73848 0 1 24213
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_480
timestamp 1704896540
transform 1 0 74800 0 1 23125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_481
timestamp 1704896540
transform 1 0 73984 0 1 21357
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_482
timestamp 1704896540
transform 1 0 77248 0 1 22989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_483
timestamp 1704896540
transform 1 0 77248 0 1 22309
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_484
timestamp 1704896540
transform 1 0 77384 0 1 22173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_485
timestamp 1704896540
transform 1 0 77384 0 1 20813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_486
timestamp 1704896540
transform 1 0 75208 0 1 23805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_487
timestamp 1704896540
transform 1 0 74256 0 1 22173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_488
timestamp 1704896540
transform 1 0 74256 0 1 21901
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_489
timestamp 1704896540
transform 1 0 73984 0 1 22581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_490
timestamp 1704896540
transform 1 0 73984 0 1 22309
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_491
timestamp 1704896540
transform 1 0 75072 0 1 22581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_492
timestamp 1704896540
transform 1 0 75072 0 1 22309
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_493
timestamp 1704896540
transform 1 0 75208 0 1 22173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_494
timestamp 1704896540
transform 1 0 74392 0 1 21493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_495
timestamp 1704896540
transform 1 0 74392 0 1 21765
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_496
timestamp 1704896540
transform 1 0 75208 0 1 21901
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_497
timestamp 1704896540
transform 1 0 75072 0 1 21357
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_498
timestamp 1704896540
transform 1 0 75480 0 1 23125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_499
timestamp 1704896540
transform 1 0 75480 0 1 23397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_500
timestamp 1704896540
transform 1 0 75480 0 1 23805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_501
timestamp 1704896540
transform 1 0 75480 0 1 23533
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_502
timestamp 1704896540
transform 1 0 77248 0 1 23941
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_503
timestamp 1704896540
transform 1 0 77248 0 1 24485
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_504
timestamp 1704896540
transform 1 0 73984 0 1 21085
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_505
timestamp 1704896540
transform 1 0 73848 0 1 22173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_506
timestamp 1704896540
transform 1 0 75072 0 1 21085
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_507
timestamp 1704896540
transform 1 0 75208 0 1 22717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_508
timestamp 1704896540
transform 1 0 73848 0 1 21901
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_509
timestamp 1704896540
transform 1 0 73848 0 1 21493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_510
timestamp 1704896540
transform 1 0 75208 0 1 22989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_511
timestamp 1704896540
transform 1 0 74664 0 1 24349
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_512
timestamp 1704896540
transform 1 0 73984 0 1 28157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_513
timestamp 1704896540
transform 1 0 75616 0 1 29517
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_514
timestamp 1704896540
transform 1 0 74936 0 1 25301
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_515
timestamp 1704896540
transform 1 0 74936 0 1 25029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_516
timestamp 1704896540
transform 1 0 74936 0 1 28293
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_517
timestamp 1704896540
transform 1 0 73848 0 1 26525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_518
timestamp 1704896540
transform 1 0 73848 0 1 26253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_519
timestamp 1704896540
transform 1 0 73984 0 1 27885
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_520
timestamp 1704896540
transform 1 0 73984 0 1 27477
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_521
timestamp 1704896540
transform 1 0 73984 0 1 27749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_522
timestamp 1704896540
transform 1 0 73848 0 1 25845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_523
timestamp 1704896540
transform 1 0 74936 0 1 28565
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_524
timestamp 1704896540
transform 1 0 74392 0 1 25301
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_525
timestamp 1704896540
transform 1 0 74392 0 1 25029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_526
timestamp 1704896540
transform 1 0 74256 0 1 28157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_527
timestamp 1704896540
transform 1 0 74256 0 1 27885
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_528
timestamp 1704896540
transform 1 0 74256 0 1 27069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_529
timestamp 1704896540
transform 1 0 74256 0 1 27341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_530
timestamp 1704896540
transform 1 0 74256 0 1 27749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_531
timestamp 1704896540
transform 1 0 74256 0 1 27477
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_532
timestamp 1704896540
transform 1 0 75616 0 1 25029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_533
timestamp 1704896540
transform 1 0 73848 0 1 26117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_534
timestamp 1704896540
transform 1 0 75480 0 1 27477
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_535
timestamp 1704896540
transform 1 0 75480 0 1 27749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_536
timestamp 1704896540
transform 1 0 74664 0 1 26661
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_537
timestamp 1704896540
transform 1 0 74664 0 1 26933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_538
timestamp 1704896540
transform 1 0 74256 0 1 26525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_539
timestamp 1704896540
transform 1 0 74256 0 1 26253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_540
timestamp 1704896540
transform 1 0 75616 0 1 26525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_541
timestamp 1704896540
transform 1 0 75616 0 1 26253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_542
timestamp 1704896540
transform 1 0 74256 0 1 25437
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_543
timestamp 1704896540
transform 1 0 74256 0 1 25709
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_544
timestamp 1704896540
transform 1 0 75616 0 1 27885
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_545
timestamp 1704896540
transform 1 0 75616 0 1 28157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_546
timestamp 1704896540
transform 1 0 74256 0 1 26117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_547
timestamp 1704896540
transform 1 0 73848 0 1 29653
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_548
timestamp 1704896540
transform 1 0 73848 0 1 29381
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_549
timestamp 1704896540
transform 1 0 74256 0 1 25845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_550
timestamp 1704896540
transform 1 0 73848 0 1 25029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_551
timestamp 1704896540
transform 1 0 73848 0 1 25301
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_552
timestamp 1704896540
transform 1 0 74256 0 1 29789
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_553
timestamp 1704896540
transform 1 0 73984 0 1 29789
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_554
timestamp 1704896540
transform 1 0 75616 0 1 27341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_555
timestamp 1704896540
transform 1 0 75616 0 1 27069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_556
timestamp 1704896540
transform 1 0 75480 0 1 26661
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_557
timestamp 1704896540
transform 1 0 75480 0 1 26933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_558
timestamp 1704896540
transform 1 0 74256 0 1 26661
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_559
timestamp 1704896540
transform 1 0 73984 0 1 26661
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_560
timestamp 1704896540
transform 1 0 73984 0 1 26933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_561
timestamp 1704896540
transform 1 0 74256 0 1 26933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_562
timestamp 1704896540
transform 1 0 75616 0 1 28293
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_563
timestamp 1704896540
transform 1 0 75616 0 1 28565
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_564
timestamp 1704896540
transform 1 0 75480 0 1 28701
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_565
timestamp 1704896540
transform 1 0 75480 0 1 28973
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_566
timestamp 1704896540
transform 1 0 74936 0 1 26525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_567
timestamp 1704896540
transform 1 0 74936 0 1 26253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_568
timestamp 1704896540
transform 1 0 73984 0 1 25437
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_569
timestamp 1704896540
transform 1 0 73984 0 1 25709
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_570
timestamp 1704896540
transform 1 0 74664 0 1 28973
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_571
timestamp 1704896540
transform 1 0 74800 0 1 25301
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_572
timestamp 1704896540
transform 1 0 74936 0 1 29789
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_573
timestamp 1704896540
transform 1 0 74392 0 1 29653
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_574
timestamp 1704896540
transform 1 0 74392 0 1 29381
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_575
timestamp 1704896540
transform 1 0 74664 0 1 27477
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_576
timestamp 1704896540
transform 1 0 74664 0 1 27749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_577
timestamp 1704896540
transform 1 0 74800 0 1 25029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_578
timestamp 1704896540
transform 1 0 74664 0 1 29245
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_579
timestamp 1704896540
transform 1 0 74664 0 1 29789
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_580
timestamp 1704896540
transform 1 0 74664 0 1 26253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_581
timestamp 1704896540
transform 1 0 74664 0 1 26525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_582
timestamp 1704896540
transform 1 0 75072 0 1 26117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_583
timestamp 1704896540
transform 1 0 75072 0 1 25845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_584
timestamp 1704896540
transform 1 0 75208 0 1 27069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_585
timestamp 1704896540
transform 1 0 75208 0 1 27341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_586
timestamp 1704896540
transform 1 0 75072 0 1 26933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_587
timestamp 1704896540
transform 1 0 75072 0 1 26661
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_588
timestamp 1704896540
transform 1 0 73848 0 1 27069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_589
timestamp 1704896540
transform 1 0 73848 0 1 27341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_590
timestamp 1704896540
transform 1 0 75616 0 1 29789
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_591
timestamp 1704896540
transform 1 0 77792 0 1 22309
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_592
timestamp 1704896540
transform 1 0 77792 0 1 22989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_593
timestamp 1704896540
transform 1 0 77792 0 1 24485
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_594
timestamp 1704896540
transform 1 0 77792 0 1 23941
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_595
timestamp 1704896540
transform 1 0 77792 0 1 23125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_596
timestamp 1704896540
transform 1 0 77792 0 1 23805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_597
timestamp 1704896540
transform 1 0 73848 0 1 31693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_598
timestamp 1704896540
transform 1 0 73848 0 1 31421
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_599
timestamp 1704896540
transform 1 0 74664 0 1 32237
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_600
timestamp 1704896540
transform 1 0 73984 0 1 31285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_601
timestamp 1704896540
transform 1 0 75480 0 1 33733
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_602
timestamp 1704896540
transform 1 0 75480 0 1 33461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_603
timestamp 1704896540
transform 1 0 73984 0 1 31013
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_604
timestamp 1704896540
transform 1 0 74392 0 1 32509
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_605
timestamp 1704896540
transform 1 0 75616 0 1 32917
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_606
timestamp 1704896540
transform 1 0 73984 0 1 34549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_607
timestamp 1704896540
transform 1 0 74664 0 1 34141
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_608
timestamp 1704896540
transform 1 0 75616 0 1 32645
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_609
timestamp 1704896540
transform 1 0 74800 0 1 31829
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_610
timestamp 1704896540
transform 1 0 74936 0 1 30061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_611
timestamp 1704896540
transform 1 0 74256 0 1 32101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_612
timestamp 1704896540
transform 1 0 73984 0 1 31829
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_613
timestamp 1704896540
transform 1 0 75480 0 1 31829
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_614
timestamp 1704896540
transform 1 0 74664 0 1 34413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_615
timestamp 1704896540
transform 1 0 75480 0 1 32101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_616
timestamp 1704896540
transform 1 0 75480 0 1 32509
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_617
timestamp 1704896540
transform 1 0 75480 0 1 32237
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_618
timestamp 1704896540
transform 1 0 74392 0 1 30605
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_619
timestamp 1704896540
transform 1 0 73984 0 1 32101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_620
timestamp 1704896540
transform 1 0 73984 0 1 32509
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_621
timestamp 1704896540
transform 1 0 73984 0 1 32237
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_622
timestamp 1704896540
transform 1 0 75208 0 1 34413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_623
timestamp 1704896540
transform 1 0 74392 0 1 30877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_624
timestamp 1704896540
transform 1 0 74392 0 1 31285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_625
timestamp 1704896540
transform 1 0 74392 0 1 31013
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_626
timestamp 1704896540
transform 1 0 75208 0 1 34141
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_627
timestamp 1704896540
transform 1 0 75072 0 1 31285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_628
timestamp 1704896540
transform 1 0 75072 0 1 31013
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_629
timestamp 1704896540
transform 1 0 74936 0 1 34005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_630
timestamp 1704896540
transform 1 0 74936 0 1 33733
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_631
timestamp 1704896540
transform 1 0 74800 0 1 34005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_632
timestamp 1704896540
transform 1 0 73984 0 1 30061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_633
timestamp 1704896540
transform 1 0 74800 0 1 33733
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_634
timestamp 1704896540
transform 1 0 73848 0 1 30197
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_635
timestamp 1704896540
transform 1 0 74256 0 1 34549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_636
timestamp 1704896540
transform 1 0 75616 0 1 30877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_637
timestamp 1704896540
transform 1 0 75616 0 1 30605
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_638
timestamp 1704896540
transform 1 0 73848 0 1 34005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_639
timestamp 1704896540
transform 1 0 73848 0 1 33733
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_640
timestamp 1704896540
transform 1 0 73848 0 1 33325
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_641
timestamp 1704896540
transform 1 0 73848 0 1 33597
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_642
timestamp 1704896540
transform 1 0 73848 0 1 30469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_643
timestamp 1704896540
transform 1 0 73848 0 1 30877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_644
timestamp 1704896540
transform 1 0 73848 0 1 30605
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_645
timestamp 1704896540
transform 1 0 74256 0 1 31829
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_646
timestamp 1704896540
transform 1 0 74800 0 1 31421
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_647
timestamp 1704896540
transform 1 0 74664 0 1 30605
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_648
timestamp 1704896540
transform 1 0 74664 0 1 30877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_649
timestamp 1704896540
transform 1 0 74800 0 1 31693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_650
timestamp 1704896540
transform 1 0 75480 0 1 31013
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_651
timestamp 1704896540
transform 1 0 75480 0 1 31285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_652
timestamp 1704896540
transform 1 0 75616 0 1 31693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_653
timestamp 1704896540
transform 1 0 75616 0 1 31421
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_654
timestamp 1704896540
transform 1 0 74256 0 1 30061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_655
timestamp 1704896540
transform 1 0 74256 0 1 30469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_656
timestamp 1704896540
transform 1 0 74256 0 1 30197
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_657
timestamp 1704896540
transform 1 0 74664 0 1 30061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_658
timestamp 1704896540
transform 1 0 74800 0 1 32101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_659
timestamp 1704896540
transform 1 0 74256 0 1 33597
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_660
timestamp 1704896540
transform 1 0 74256 0 1 33325
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_661
timestamp 1704896540
transform 1 0 73984 0 1 34413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_662
timestamp 1704896540
transform 1 0 73984 0 1 34141
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_663
timestamp 1704896540
transform 1 0 74256 0 1 33733
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_664
timestamp 1704896540
transform 1 0 74256 0 1 34005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_665
timestamp 1704896540
transform 1 0 74392 0 1 34413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_666
timestamp 1704896540
transform 1 0 74392 0 1 34141
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_667
timestamp 1704896540
transform 1 0 74936 0 1 33189
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_668
timestamp 1704896540
transform 1 0 75480 0 1 30469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_669
timestamp 1704896540
transform 1 0 75480 0 1 30197
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_670
timestamp 1704896540
transform 1 0 74936 0 1 32917
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_671
timestamp 1704896540
transform 1 0 74800 0 1 33189
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_672
timestamp 1704896540
transform 1 0 74800 0 1 32917
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_673
timestamp 1704896540
transform 1 0 74392 0 1 31693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_674
timestamp 1704896540
transform 1 0 75480 0 1 34141
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_675
timestamp 1704896540
transform 1 0 75480 0 1 34413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_676
timestamp 1704896540
transform 1 0 74800 0 1 30197
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_677
timestamp 1704896540
transform 1 0 74800 0 1 30469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_678
timestamp 1704896540
transform 1 0 75072 0 1 34549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_679
timestamp 1704896540
transform 1 0 74392 0 1 31421
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_680
timestamp 1704896540
transform 1 0 74392 0 1 32237
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_681
timestamp 1704896540
transform 1 0 75208 0 1 31421
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_682
timestamp 1704896540
transform 1 0 75208 0 1 31693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_683
timestamp 1704896540
transform 1 0 74664 0 1 32509
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_684
timestamp 1704896540
transform 1 0 74800 0 1 35229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_685
timestamp 1704896540
transform 1 0 74800 0 1 34957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_686
timestamp 1704896540
transform 1 0 75616 0 1 35229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_687
timestamp 1704896540
transform 1 0 75616 0 1 34957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_688
timestamp 1704896540
transform 1 0 73984 0 1 34821
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_689
timestamp 1704896540
transform 1 0 75480 0 1 35365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_690
timestamp 1704896540
transform 1 0 75480 0 1 35637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_691
timestamp 1704896540
transform 1 0 75616 0 1 38901
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_692
timestamp 1704896540
transform 1 0 75616 0 1 39173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_693
timestamp 1704896540
transform 1 0 75616 0 1 39581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_694
timestamp 1704896540
transform 1 0 75616 0 1 39309
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_695
timestamp 1704896540
transform 1 0 75616 0 1 36589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_696
timestamp 1704896540
transform 1 0 75616 0 1 36861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_697
timestamp 1704896540
transform 1 0 74664 0 1 35365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_698
timestamp 1704896540
transform 1 0 75616 0 1 35773
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_699
timestamp 1704896540
transform 1 0 75616 0 1 36045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_700
timestamp 1704896540
transform 1 0 75616 0 1 36453
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_701
timestamp 1704896540
transform 1 0 75616 0 1 36181
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_702
timestamp 1704896540
transform 1 0 74664 0 1 35637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_703
timestamp 1704896540
transform 1 0 74392 0 1 37677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_704
timestamp 1704896540
transform 1 0 74392 0 1 37949
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_705
timestamp 1704896540
transform 1 0 74256 0 1 34821
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_706
timestamp 1704896540
transform 1 0 75480 0 1 37677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_707
timestamp 1704896540
transform 1 0 75480 0 1 37405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_708
timestamp 1704896540
transform 1 0 75616 0 1 36997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_709
timestamp 1704896540
transform 1 0 75616 0 1 37269
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_710
timestamp 1704896540
transform 1 0 74392 0 1 38765
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_711
timestamp 1704896540
transform 1 0 74392 0 1 38493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_712
timestamp 1704896540
transform 1 0 74256 0 1 38085
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_713
timestamp 1704896540
transform 1 0 74256 0 1 38357
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_714
timestamp 1704896540
transform 1 0 74256 0 1 35365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_715
timestamp 1704896540
transform 1 0 74256 0 1 35637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_716
timestamp 1704896540
transform 1 0 74392 0 1 36045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_717
timestamp 1704896540
transform 1 0 74392 0 1 35773
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_718
timestamp 1704896540
transform 1 0 74936 0 1 35229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_719
timestamp 1704896540
transform 1 0 74936 0 1 34957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_720
timestamp 1704896540
transform 1 0 75072 0 1 34821
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_721
timestamp 1704896540
transform 1 0 75072 0 1 36045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_722
timestamp 1704896540
transform 1 0 75072 0 1 35773
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_723
timestamp 1704896540
transform 1 0 73984 0 1 39173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_724
timestamp 1704896540
transform 1 0 73984 0 1 38901
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_725
timestamp 1704896540
transform 1 0 75072 0 1 36181
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_726
timestamp 1704896540
transform 1 0 75072 0 1 36453
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_727
timestamp 1704896540
transform 1 0 75208 0 1 39581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_728
timestamp 1704896540
transform 1 0 75208 0 1 39309
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_729
timestamp 1704896540
transform 1 0 75072 0 1 39173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_730
timestamp 1704896540
transform 1 0 75072 0 1 38901
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_731
timestamp 1704896540
transform 1 0 75072 0 1 35637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_732
timestamp 1704896540
transform 1 0 75072 0 1 35365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_733
timestamp 1704896540
transform 1 0 75072 0 1 38765
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_734
timestamp 1704896540
transform 1 0 75072 0 1 38493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_735
timestamp 1704896540
transform 1 0 73984 0 1 38765
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_736
timestamp 1704896540
transform 1 0 73984 0 1 38493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_737
timestamp 1704896540
transform 1 0 74936 0 1 36453
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_738
timestamp 1704896540
transform 1 0 74936 0 1 36181
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_739
timestamp 1704896540
transform 1 0 74664 0 1 38493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_740
timestamp 1704896540
transform 1 0 74664 0 1 38765
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_741
timestamp 1704896540
transform 1 0 73848 0 1 38357
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_742
timestamp 1704896540
transform 1 0 74256 0 1 39581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_743
timestamp 1704896540
transform 1 0 74256 0 1 39309
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_744
timestamp 1704896540
transform 1 0 73848 0 1 38085
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_745
timestamp 1704896540
transform 1 0 73848 0 1 36453
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_746
timestamp 1704896540
transform 1 0 73848 0 1 36181
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_747
timestamp 1704896540
transform 1 0 74936 0 1 39581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_748
timestamp 1704896540
transform 1 0 74936 0 1 39309
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_749
timestamp 1704896540
transform 1 0 73984 0 1 39309
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_750
timestamp 1704896540
transform 1 0 73984 0 1 39581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_751
timestamp 1704896540
transform 1 0 74664 0 1 39309
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_752
timestamp 1704896540
transform 1 0 74664 0 1 39581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_753
timestamp 1704896540
transform 1 0 74936 0 1 37269
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_754
timestamp 1704896540
transform 1 0 74936 0 1 36997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_755
timestamp 1704896540
transform 1 0 73848 0 1 36045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_756
timestamp 1704896540
transform 1 0 73848 0 1 35773
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_757
timestamp 1704896540
transform 1 0 73984 0 1 37949
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_758
timestamp 1704896540
transform 1 0 73984 0 1 37677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_759
timestamp 1704896540
transform 1 0 74664 0 1 37269
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_760
timestamp 1704896540
transform 1 0 74664 0 1 36997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_761
timestamp 1704896540
transform 1 0 74256 0 1 35229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_762
timestamp 1704896540
transform 1 0 74256 0 1 34957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_763
timestamp 1704896540
transform 1 0 73984 0 1 34957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_764
timestamp 1704896540
transform 1 0 73984 0 1 35229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_765
timestamp 1704896540
transform 1 0 73984 0 1 35637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_766
timestamp 1704896540
transform 1 0 74256 0 1 39173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_767
timestamp 1704896540
transform 1 0 74256 0 1 38901
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_768
timestamp 1704896540
transform 1 0 73984 0 1 35365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_769
timestamp 1704896540
transform 1 0 74664 0 1 37949
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_770
timestamp 1704896540
transform 1 0 74664 0 1 37677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_771
timestamp 1704896540
transform 1 0 74256 0 1 36453
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_772
timestamp 1704896540
transform 1 0 74256 0 1 36181
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_773
timestamp 1704896540
transform 1 0 94656 0 1 30605
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_774
timestamp 1704896540
transform 1 0 94656 0 1 32237
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_775
timestamp 1704896540
transform 1 0 94656 0 1 37405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_776
timestamp 1704896540
transform 1 0 94656 0 1 38901
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_777
timestamp 1704896540
transform 1 0 94656 0 1 35501
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_778
timestamp 1704896540
transform 1 0 94656 0 1 33869
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_779
timestamp 1704896540
transform 1 0 78608 0 1 19997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_780
timestamp 1704896540
transform 1 0 77656 0 1 19997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_781
timestamp 1704896540
transform 1 0 75480 0 1 19997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_782
timestamp 1704896540
transform 1 0 69088 0 1 19997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_783
timestamp 1704896540
transform 1 0 79424 0 1 19997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_784
timestamp 1704896540
transform 1 0 78200 0 1 19997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_785
timestamp 1704896540
transform 1 0 47056 0 1 2861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_786
timestamp 1704896540
transform 1 0 45968 0 1 2861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_787
timestamp 1704896540
transform 1 0 47464 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_788
timestamp 1704896540
transform 1 0 42432 0 1 2861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_789
timestamp 1704896540
transform 1 0 44880 0 1 2861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_790
timestamp 1704896540
transform 1 0 43520 0 1 2861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_791
timestamp 1704896540
transform 1 0 45832 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_792
timestamp 1704896540
transform 1 0 42296 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_793
timestamp 1704896540
transform 1 0 42296 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_794
timestamp 1704896540
transform 1 0 45832 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_795
timestamp 1704896540
transform 1 0 44200 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_796
timestamp 1704896540
transform 1 0 47464 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_797
timestamp 1704896540
transform 1 0 44200 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_798
timestamp 1704896540
transform 1 0 40256 0 1 2861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_799
timestamp 1704896540
transform 1 0 38896 0 1 2861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_800
timestamp 1704896540
transform 1 0 37672 0 1 2861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_801
timestamp 1704896540
transform 1 0 36584 0 1 2861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_802
timestamp 1704896540
transform 1 0 41344 0 1 2861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_803
timestamp 1704896540
transform 1 0 37400 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_804
timestamp 1704896540
transform 1 0 37400 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_805
timestamp 1704896540
transform 1 0 40528 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_806
timestamp 1704896540
transform 1 0 40528 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_807
timestamp 1704896540
transform 1 0 39168 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_808
timestamp 1704896540
transform 1 0 39168 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_809
timestamp 1704896540
transform 1 0 37128 0 1 10069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_810
timestamp 1704896540
transform 1 0 37264 0 1 9253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_811
timestamp 1704896540
transform 1 0 37264 0 1 9797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_812
timestamp 1704896540
transform 1 0 39576 0 1 9389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_813
timestamp 1704896540
transform 1 0 38352 0 1 8573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_814
timestamp 1704896540
transform 1 0 40936 0 1 8573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_815
timestamp 1704896540
transform 1 0 41752 0 1 10069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_816
timestamp 1704896540
transform 1 0 40936 0 1 9389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_817
timestamp 1704896540
transform 1 0 40936 0 1 10069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_818
timestamp 1704896540
transform 1 0 41072 0 1 9253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_819
timestamp 1704896540
transform 1 0 41072 0 1 9797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_820
timestamp 1704896540
transform 1 0 38352 0 1 9389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_821
timestamp 1704896540
transform 1 0 37128 0 1 8573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_822
timestamp 1704896540
transform 1 0 37128 0 1 9389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_823
timestamp 1704896540
transform 1 0 39712 0 1 10069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_824
timestamp 1704896540
transform 1 0 39712 0 1 9253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_825
timestamp 1704896540
transform 1 0 39712 0 1 9797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_826
timestamp 1704896540
transform 1 0 38624 0 1 10069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_827
timestamp 1704896540
transform 1 0 38216 0 1 9253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_828
timestamp 1704896540
transform 1 0 38488 0 1 9525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_829
timestamp 1704896540
transform 1 0 39576 0 1 8573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_830
timestamp 1704896540
transform 1 0 38216 0 1 9797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_831
timestamp 1704896540
transform 1 0 43520 0 1 10069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_832
timestamp 1704896540
transform 1 0 43520 0 1 9797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_833
timestamp 1704896540
transform 1 0 43520 0 1 8981
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_834
timestamp 1704896540
transform 1 0 42296 0 1 10069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_835
timestamp 1704896540
transform 1 0 42296 0 1 9253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_836
timestamp 1704896540
transform 1 0 42296 0 1 9797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_837
timestamp 1704896540
transform 1 0 47056 0 1 8573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_838
timestamp 1704896540
transform 1 0 47056 0 1 9389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_839
timestamp 1704896540
transform 1 0 42160 0 1 8573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_840
timestamp 1704896540
transform 1 0 42160 0 1 9389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_841
timestamp 1704896540
transform 1 0 43384 0 1 8573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_842
timestamp 1704896540
transform 1 0 43384 0 1 9389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_843
timestamp 1704896540
transform 1 0 44608 0 1 8573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_844
timestamp 1704896540
transform 1 0 44608 0 1 9389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_845
timestamp 1704896540
transform 1 0 47736 0 1 10069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_846
timestamp 1704896540
transform 1 0 45832 0 1 8573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_847
timestamp 1704896540
transform 1 0 47192 0 1 10069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_848
timestamp 1704896540
transform 1 0 47192 0 1 9253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_849
timestamp 1704896540
transform 1 0 47192 0 1 9797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_850
timestamp 1704896540
transform 1 0 45832 0 1 9389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_851
timestamp 1704896540
transform 1 0 45968 0 1 10069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_852
timestamp 1704896540
transform 1 0 45968 0 1 9253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_853
timestamp 1704896540
transform 1 0 45968 0 1 9797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_854
timestamp 1704896540
transform 1 0 45288 0 1 10069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_855
timestamp 1704896540
transform 1 0 44744 0 1 10069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_856
timestamp 1704896540
transform 1 0 44744 0 1 9253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_857
timestamp 1704896540
transform 1 0 44744 0 1 9797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_858
timestamp 1704896540
transform 1 0 35768 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_859
timestamp 1704896540
transform 1 0 30600 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_860
timestamp 1704896540
transform 1 0 35768 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_861
timestamp 1704896540
transform 1 0 34000 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_862
timestamp 1704896540
transform 1 0 35496 0 1 2861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_863
timestamp 1704896540
transform 1 0 34136 0 1 2861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_864
timestamp 1704896540
transform 1 0 33048 0 1 2861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_865
timestamp 1704896540
transform 1 0 31824 0 1 2861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_866
timestamp 1704896540
transform 1 0 30736 0 1 2861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_867
timestamp 1704896540
transform 1 0 34000 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_868
timestamp 1704896540
transform 1 0 32368 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_869
timestamp 1704896540
transform 1 0 32368 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_870
timestamp 1704896540
transform 1 0 30600 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_871
timestamp 1704896540
transform 1 0 29648 0 1 2861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_872
timestamp 1704896540
transform 1 0 28288 0 1 2861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_873
timestamp 1704896540
transform 1 0 27200 0 1 2861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_874
timestamp 1704896540
transform 1 0 26112 0 1 2861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_875
timestamp 1704896540
transform 1 0 25024 0 1 2861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_876
timestamp 1704896540
transform 1 0 26656 0 1 549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_877
timestamp 1704896540
transform 1 0 26656 0 1 2317
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_878
timestamp 1704896540
transform 1 0 27472 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_879
timestamp 1704896540
transform 1 0 27472 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_880
timestamp 1704896540
transform 1 0 28968 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_881
timestamp 1704896540
transform 1 0 28968 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_882
timestamp 1704896540
transform 1 0 25704 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_883
timestamp 1704896540
transform 1 0 25704 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_884
timestamp 1704896540
transform 1 0 27744 0 1 8845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_885
timestamp 1704896540
transform 1 0 27744 0 1 7077
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_886
timestamp 1704896540
transform 1 0 29648 0 1 8573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_887
timestamp 1704896540
transform 1 0 29648 0 1 9389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_888
timestamp 1704896540
transform 1 0 28288 0 1 9389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_889
timestamp 1704896540
transform 1 0 28560 0 1 10069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_890
timestamp 1704896540
transform 1 0 28424 0 1 9253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_891
timestamp 1704896540
transform 1 0 28424 0 1 9797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_892
timestamp 1704896540
transform 1 0 28152 0 1 8573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_893
timestamp 1704896540
transform 1 0 28152 0 1 8165
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_894
timestamp 1704896540
transform 1 0 29784 0 1 10069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_895
timestamp 1704896540
transform 1 0 29784 0 1 9253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_896
timestamp 1704896540
transform 1 0 29784 0 1 9797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_897
timestamp 1704896540
transform 1 0 28288 0 1 8573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_898
timestamp 1704896540
transform 1 0 32232 0 1 8573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_899
timestamp 1704896540
transform 1 0 32232 0 1 9389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_900
timestamp 1704896540
transform 1 0 34816 0 1 10069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_901
timestamp 1704896540
transform 1 0 34816 0 1 9253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_902
timestamp 1704896540
transform 1 0 34816 0 1 9797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_903
timestamp 1704896540
transform 1 0 33456 0 1 10069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_904
timestamp 1704896540
transform 1 0 33592 0 1 9253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_905
timestamp 1704896540
transform 1 0 33592 0 1 9797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_906
timestamp 1704896540
transform 1 0 30736 0 1 8573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_907
timestamp 1704896540
transform 1 0 32232 0 1 10069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_908
timestamp 1704896540
transform 1 0 32368 0 1 9253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_909
timestamp 1704896540
transform 1 0 32368 0 1 9797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_910
timestamp 1704896540
transform 1 0 30736 0 1 9389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_911
timestamp 1704896540
transform 1 0 30872 0 1 10069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_912
timestamp 1704896540
transform 1 0 30872 0 1 9253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_913
timestamp 1704896540
transform 1 0 30872 0 1 9797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_914
timestamp 1704896540
transform 1 0 35904 0 1 8573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_915
timestamp 1704896540
transform 1 0 35904 0 1 9389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_916
timestamp 1704896540
transform 1 0 33456 0 1 8573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_917
timestamp 1704896540
transform 1 0 33456 0 1 9389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_918
timestamp 1704896540
transform 1 0 34680 0 1 8573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_919
timestamp 1704896540
transform 1 0 34680 0 1 9389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_920
timestamp 1704896540
transform 1 0 27064 0 1 19861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_921
timestamp 1704896540
transform 1 0 30464 0 1 16597
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_922
timestamp 1704896540
transform 1 0 30464 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_923
timestamp 1704896540
transform 1 0 34680 0 1 11157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_924
timestamp 1704896540
transform 1 0 34680 0 1 11837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_925
timestamp 1704896540
transform 1 0 34544 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_926
timestamp 1704896540
transform 1 0 34544 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_927
timestamp 1704896540
transform 1 0 28560 0 1 14557
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_928
timestamp 1704896540
transform 1 0 28560 0 1 17005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_929
timestamp 1704896540
transform 1 0 29784 0 1 11157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_930
timestamp 1704896540
transform 1 0 32776 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_931
timestamp 1704896540
transform 1 0 29784 0 1 11837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_932
timestamp 1704896540
transform 1 0 29240 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_933
timestamp 1704896540
transform 1 0 32776 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_934
timestamp 1704896540
transform 1 0 33184 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_935
timestamp 1704896540
transform 1 0 31960 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_936
timestamp 1704896540
transform 1 0 32096 0 1 11157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_937
timestamp 1704896540
transform 1 0 29240 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_938
timestamp 1704896540
transform 1 0 30328 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_939
timestamp 1704896540
transform 1 0 29240 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_940
timestamp 1704896540
transform 1 0 32096 0 1 11837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_941
timestamp 1704896540
transform 1 0 32096 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_942
timestamp 1704896540
transform 1 0 27880 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_943
timestamp 1704896540
transform 1 0 31552 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_944
timestamp 1704896540
transform 1 0 31552 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_945
timestamp 1704896540
transform 1 0 31008 0 1 11157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_946
timestamp 1704896540
transform 1 0 32096 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_947
timestamp 1704896540
transform 1 0 28424 0 1 11157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_948
timestamp 1704896540
transform 1 0 31008 0 1 11837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_949
timestamp 1704896540
transform 1 0 35632 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_950
timestamp 1704896540
transform 1 0 28424 0 1 11837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_951
timestamp 1704896540
transform 1 0 34408 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_952
timestamp 1704896540
transform 1 0 34816 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_953
timestamp 1704896540
transform 1 0 33456 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_954
timestamp 1704896540
transform 1 0 32232 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_955
timestamp 1704896540
transform 1 0 31144 0 1 14285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_956
timestamp 1704896540
transform 1 0 31144 0 1 12653
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_957
timestamp 1704896540
transform 1 0 28288 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_958
timestamp 1704896540
transform 1 0 28288 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_959
timestamp 1704896540
transform 1 0 30872 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_960
timestamp 1704896540
transform 1 0 29784 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_961
timestamp 1704896540
transform 1 0 28560 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_962
timestamp 1704896540
transform 1 0 34136 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_963
timestamp 1704896540
transform 1 0 34136 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_964
timestamp 1704896540
transform 1 0 33456 0 1 11157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_965
timestamp 1704896540
transform 1 0 33456 0 1 11837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_966
timestamp 1704896540
transform 1 0 33320 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_967
timestamp 1704896540
transform 1 0 33320 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_968
timestamp 1704896540
transform 1 0 35768 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_969
timestamp 1704896540
transform 1 0 35768 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_970
timestamp 1704896540
transform 1 0 26520 0 1 16597
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_971
timestamp 1704896540
transform 1 0 26520 0 1 16869
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_972
timestamp 1704896540
transform 1 0 42160 0 1 11157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_973
timestamp 1704896540
transform 1 0 42160 0 1 11837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_974
timestamp 1704896540
transform 1 0 42024 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_975
timestamp 1704896540
transform 1 0 42024 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_976
timestamp 1704896540
transform 1 0 40800 0 1 11157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_977
timestamp 1704896540
transform 1 0 40800 0 1 11837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_978
timestamp 1704896540
transform 1 0 40800 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_979
timestamp 1704896540
transform 1 0 40800 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_980
timestamp 1704896540
transform 1 0 40256 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_981
timestamp 1704896540
transform 1 0 40256 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_982
timestamp 1704896540
transform 1 0 39712 0 1 11157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_983
timestamp 1704896540
transform 1 0 39712 0 1 11837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_984
timestamp 1704896540
transform 1 0 39576 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_985
timestamp 1704896540
transform 1 0 39576 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_986
timestamp 1704896540
transform 1 0 39032 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_987
timestamp 1704896540
transform 1 0 39032 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_988
timestamp 1704896540
transform 1 0 38488 0 1 11157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_989
timestamp 1704896540
transform 1 0 38488 0 1 11837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_990
timestamp 1704896540
transform 1 0 38488 0 1 11021
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_991
timestamp 1704896540
transform 1 0 38352 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_992
timestamp 1704896540
transform 1 0 38352 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_993
timestamp 1704896540
transform 1 0 44744 0 1 11837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_994
timestamp 1704896540
transform 1 0 37128 0 1 11157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_995
timestamp 1704896540
transform 1 0 37128 0 1 11837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_996
timestamp 1704896540
transform 1 0 36584 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_997
timestamp 1704896540
transform 1 0 36584 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_998
timestamp 1704896540
transform 1 0 44608 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_999
timestamp 1704896540
transform 1 0 44608 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1000
timestamp 1704896540
transform 1 0 47736 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1001
timestamp 1704896540
transform 1 0 47192 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1002
timestamp 1704896540
transform 1 0 45968 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1003
timestamp 1704896540
transform 1 0 45288 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1004
timestamp 1704896540
transform 1 0 44744 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1005
timestamp 1704896540
transform 1 0 43520 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1006
timestamp 1704896540
transform 1 0 42296 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1007
timestamp 1704896540
transform 1 0 41752 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1008
timestamp 1704896540
transform 1 0 40936 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1009
timestamp 1704896540
transform 1 0 39712 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1010
timestamp 1704896540
transform 1 0 38624 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1011
timestamp 1704896540
transform 1 0 37128 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1012
timestamp 1704896540
transform 1 0 43384 0 1 11157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1013
timestamp 1704896540
transform 1 0 43384 0 1 11837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1014
timestamp 1704896540
transform 1 0 42840 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1015
timestamp 1704896540
transform 1 0 42840 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1016
timestamp 1704896540
transform 1 0 47736 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1017
timestamp 1704896540
transform 1 0 47736 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1018
timestamp 1704896540
transform 1 0 47192 0 1 11157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1019
timestamp 1704896540
transform 1 0 47192 0 1 11837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1020
timestamp 1704896540
transform 1 0 47056 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1021
timestamp 1704896540
transform 1 0 47056 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1022
timestamp 1704896540
transform 1 0 46512 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1023
timestamp 1704896540
transform 1 0 46512 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1024
timestamp 1704896540
transform 1 0 45832 0 1 11157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1025
timestamp 1704896540
transform 1 0 45832 0 1 11837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1026
timestamp 1704896540
transform 1 0 47872 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1027
timestamp 1704896540
transform 1 0 46648 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1028
timestamp 1704896540
transform 1 0 45560 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1029
timestamp 1704896540
transform 1 0 44336 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1030
timestamp 1704896540
transform 1 0 43112 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1031
timestamp 1704896540
transform 1 0 41888 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1032
timestamp 1704896540
transform 1 0 40664 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1033
timestamp 1704896540
transform 1 0 39304 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1034
timestamp 1704896540
transform 1 0 37808 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1035
timestamp 1704896540
transform 1 0 36856 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1036
timestamp 1704896540
transform 1 0 45832 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1037
timestamp 1704896540
transform 1 0 45832 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1038
timestamp 1704896540
transform 1 0 45288 0 1 16053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1039
timestamp 1704896540
transform 1 0 45288 0 1 16461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1040
timestamp 1704896540
transform 1 0 44744 0 1 11157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1041
timestamp 1704896540
transform 1 0 36040 0 1 11157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1042
timestamp 1704896540
transform 1 0 36040 0 1 11837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1043
timestamp 1704896540
transform 1 0 36040 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1044
timestamp 1704896540
transform 1 0 36040 0 1 10069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1045
timestamp 1704896540
transform 1 0 36040 0 1 9253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1046
timestamp 1704896540
transform 1 0 36040 0 1 9797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1047
timestamp 1704896540
transform 1 0 18904 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1048
timestamp 1704896540
transform 1 0 18904 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1049
timestamp 1704896540
transform 1 0 22440 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1050
timestamp 1704896540
transform 1 0 20128 0 1 2861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1051
timestamp 1704896540
transform 1 0 19176 0 1 2861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1052
timestamp 1704896540
transform 1 0 23664 0 1 2861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1053
timestamp 1704896540
transform 1 0 22576 0 1 2861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1054
timestamp 1704896540
transform 1 0 21352 0 1 2861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1055
timestamp 1704896540
transform 1 0 22440 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1056
timestamp 1704896540
transform 1 0 20672 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1057
timestamp 1704896540
transform 1 0 23936 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1058
timestamp 1704896540
transform 1 0 23936 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1059
timestamp 1704896540
transform 1 0 20672 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1060
timestamp 1704896540
transform 1 0 17816 0 1 2861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1061
timestamp 1704896540
transform 1 0 16728 0 1 2861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1062
timestamp 1704896540
transform 1 0 15504 0 1 2861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1063
timestamp 1704896540
transform 1 0 14008 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1064
timestamp 1704896540
transform 1 0 14008 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1065
timestamp 1704896540
transform 1 0 17408 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1066
timestamp 1704896540
transform 1 0 16048 0 1 2453
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1067
timestamp 1704896540
transform 1 0 16048 0 1 4765
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1068
timestamp 1704896540
transform 1 0 17408 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1069
timestamp 1704896540
transform 1 0 14280 0 1 5037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1070
timestamp 1704896540
transform 1 0 17272 0 1 1773
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1071
timestamp 1704896540
transform 1 0 17272 0 1 3677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1072
timestamp 1704896540
transform 1 0 15776 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1073
timestamp 1704896540
transform 1 0 15776 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1074
timestamp 1704896540
transform 1 0 15912 0 1 3813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1075
timestamp 1704896540
transform 1 0 12240 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1076
timestamp 1704896540
transform 1 0 12240 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1077
timestamp 1704896540
transform 1 0 14280 0 1 7621
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1078
timestamp 1704896540
transform 1 0 14008 0 1 7757
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1079
timestamp 1704896540
transform 1 0 14280 0 1 9253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1080
timestamp 1704896540
transform 1 0 15912 0 1 6261
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1081
timestamp 1704896540
transform 1 0 14144 0 1 9117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1082
timestamp 1704896540
transform 1 0 14144 0 1 6397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1083
timestamp 1704896540
transform 1 0 8976 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1084
timestamp 1704896540
transform 1 0 10472 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1085
timestamp 1704896540
transform 1 0 10472 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1086
timestamp 1704896540
transform 1 0 8976 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1087
timestamp 1704896540
transform 1 0 7208 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1088
timestamp 1704896540
transform 1 0 7208 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1089
timestamp 1704896540
transform 1 0 5440 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1090
timestamp 1704896540
transform 1 0 3944 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1091
timestamp 1704896540
transform 1 0 3944 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1092
timestamp 1704896540
transform 1 0 2176 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1093
timestamp 1704896540
transform 1 0 2176 0 1 1637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1094
timestamp 1704896540
transform 1 0 1224 0 1 3677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1095
timestamp 1704896540
transform 1 0 5440 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1096
timestamp 1704896540
transform 1 0 544 0 1 5037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1097
timestamp 1704896540
transform 1 0 1224 0 1 6941
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1098
timestamp 1704896540
transform 1 0 2584 0 1 6397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1099
timestamp 1704896540
transform 1 0 2584 0 1 6941
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1100
timestamp 1704896540
transform 1 0 1224 0 1 8845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1101
timestamp 1704896540
transform 1 0 1224 0 1 5309
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1102
timestamp 1704896540
transform 1 0 544 0 1 7621
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1103
timestamp 1704896540
transform 1 0 5848 0 1 5445
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1104
timestamp 1704896540
transform 1 0 1224 0 1 11973
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1105
timestamp 1704896540
transform 1 0 1224 0 1 13741
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1106
timestamp 1704896540
transform 1 0 1224 0 1 10477
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1107
timestamp 1704896540
transform 1 0 3128 0 1 13469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1108
timestamp 1704896540
transform 1 0 3128 0 1 13741
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1109
timestamp 1704896540
transform 1 0 544 0 1 11837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1110
timestamp 1704896540
transform 1 0 3944 0 1 14693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1111
timestamp 1704896540
transform 1 0 3808 0 1 11973
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1112
timestamp 1704896540
transform 1 0 3808 0 1 14693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1113
timestamp 1704896540
transform 1 0 3808 0 1 17685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1114
timestamp 1704896540
transform 1 0 3808 0 1 17549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1115
timestamp 1704896540
transform 1 0 1224 0 1 18909
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1116
timestamp 1704896540
transform 1 0 1224 0 1 17277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1117
timestamp 1704896540
transform 1 0 2555 0 1 15197
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1118
timestamp 1704896540
transform 1 0 1224 0 1 15373
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1119
timestamp 1704896540
transform 1 0 2312 0 1 16189
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1120
timestamp 1704896540
transform 1 0 2312 0 1 15509
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1121
timestamp 1704896540
transform 1 0 20672 0 1 14693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1122
timestamp 1704896540
transform 1 0 20672 0 1 17413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1123
timestamp 1704896540
transform 1 0 20536 0 1 17821
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1124
timestamp 1704896540
transform 1 0 20536 0 1 17549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1125
timestamp 1704896540
transform 1 0 18224 0 1 18229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1126
timestamp 1704896540
transform 1 0 18224 0 1 17549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1127
timestamp 1704896540
transform 1 0 18224 0 1 18365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1128
timestamp 1704896540
transform 1 0 18224 0 1 19861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1129
timestamp 1704896540
transform 1 0 17544 0 1 18229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1130
timestamp 1704896540
transform 1 0 17544 0 1 17549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1131
timestamp 1704896540
transform 1 0 22032 0 1 19589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1132
timestamp 1704896540
transform 1 0 22032 0 1 19861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1133
timestamp 1704896540
transform 1 0 16184 0 1 17413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1134
timestamp 1704896540
transform 1 0 16184 0 1 16325
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1135
timestamp 1704896540
transform 1 0 14280 0 1 16189
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1136
timestamp 1704896540
transform 1 0 14280 0 1 13469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1137
timestamp 1704896540
transform 1 0 21488 0 1 19861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1138
timestamp 1704896540
transform 1 0 21488 0 1 19589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1139
timestamp 1704896540
transform 1 0 21216 0 1 18365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1140
timestamp 1704896540
transform 1 0 21216 0 1 18637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1141
timestamp 1704896540
transform 1 0 14008 0 1 13333
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1142
timestamp 1704896540
transform 1 0 14008 0 1 10613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1143
timestamp 1704896540
transform 1 0 14008 0 1 10477
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1144
timestamp 1704896540
transform 1 0 21352 0 1 18773
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1145
timestamp 1704896540
transform 1 0 21352 0 1 19045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1146
timestamp 1704896540
transform 1 0 22032 0 1 16869
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1147
timestamp 1704896540
transform 1 0 22032 0 1 13197
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1148
timestamp 1704896540
transform 1 0 20808 0 1 18365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1149
timestamp 1704896540
transform 1 0 20808 0 1 18637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1150
timestamp 1704896540
transform 1 0 20808 0 1 19589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1151
timestamp 1704896540
transform 1 0 20808 0 1 19861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1152
timestamp 1704896540
transform 1 0 20944 0 1 19453
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1153
timestamp 1704896540
transform 1 0 20944 0 1 19181
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1154
timestamp 1704896540
transform 1 0 20944 0 1 18229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1155
timestamp 1704896540
transform 1 0 20944 0 1 17957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1156
timestamp 1704896540
transform 1 0 20400 0 1 19045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1157
timestamp 1704896540
transform 1 0 21624 0 1 17821
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1158
timestamp 1704896540
transform 1 0 21624 0 1 17549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1159
timestamp 1704896540
transform 1 0 18768 0 1 17549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1160
timestamp 1704896540
transform 1 0 18768 0 1 18229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1161
timestamp 1704896540
transform 1 0 21624 0 1 19861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1162
timestamp 1704896540
transform 1 0 21624 0 1 19589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1163
timestamp 1704896540
transform 1 0 21624 0 1 19181
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1164
timestamp 1704896540
transform 1 0 21624 0 1 19453
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1165
timestamp 1704896540
transform 1 0 18632 0 1 18365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1166
timestamp 1704896540
transform 1 0 18632 0 1 19861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1167
timestamp 1704896540
transform 1 0 20400 0 1 19453
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1168
timestamp 1704896540
transform 1 0 22032 0 1 18637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1169
timestamp 1704896540
transform 1 0 22032 0 1 19045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1170
timestamp 1704896540
transform 1 0 22032 0 1 18773
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1171
timestamp 1704896540
transform 1 0 22168 0 1 19181
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1172
timestamp 1704896540
transform 1 0 22168 0 1 19453
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1173
timestamp 1704896540
transform 1 0 16592 0 1 17413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1174
timestamp 1704896540
transform 1 0 16592 0 1 14829
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1175
timestamp 1704896540
transform 1 0 14144 0 1 14693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1176
timestamp 1704896540
transform 1 0 22168 0 1 17549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1177
timestamp 1704896540
transform 1 0 14144 0 1 11973
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1178
timestamp 1704896540
transform 1 0 21624 0 1 19045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1179
timestamp 1704896540
transform 1 0 21624 0 1 18773
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1180
timestamp 1704896540
transform 1 0 14280 0 1 11837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1181
timestamp 1704896540
transform 1 0 22848 0 1 17005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1182
timestamp 1704896540
transform 1 0 22848 0 1 17413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1183
timestamp 1704896540
transform 1 0 22032 0 1 17005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1184
timestamp 1704896540
transform 1 0 22032 0 1 17413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1185
timestamp 1704896540
transform 1 0 22168 0 1 17821
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1186
timestamp 1704896540
transform 1 0 22168 0 1 18229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1187
timestamp 1704896540
transform 1 0 22168 0 1 17957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1188
timestamp 1704896540
transform 1 0 22032 0 1 18365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1189
timestamp 1704896540
transform 1 0 21760 0 1 17957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1190
timestamp 1704896540
transform 1 0 21760 0 1 18229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1191
timestamp 1704896540
transform 1 0 21624 0 1 18637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1192
timestamp 1704896540
transform 1 0 21624 0 1 18365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1193
timestamp 1704896540
transform 1 0 21080 0 1 11837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1194
timestamp 1704896540
transform 1 0 21080 0 1 14557
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1195
timestamp 1704896540
transform 1 0 20400 0 1 19589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1196
timestamp 1704896540
transform 1 0 20400 0 1 19861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1197
timestamp 1704896540
transform 1 0 20400 0 1 18365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1198
timestamp 1704896540
transform 1 0 20400 0 1 18637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1199
timestamp 1704896540
transform 1 0 20400 0 1 19181
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1200
timestamp 1704896540
transform 1 0 20400 0 1 18773
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1201
timestamp 1704896540
transform 1 0 18360 0 1 23125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1202
timestamp 1704896540
transform 1 0 22032 0 1 23805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1203
timestamp 1704896540
transform 1 0 18768 0 1 20541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1204
timestamp 1704896540
transform 1 0 21760 0 1 21901
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1205
timestamp 1704896540
transform 1 0 22032 0 1 23397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1206
timestamp 1704896540
transform 1 0 22032 0 1 23125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1207
timestamp 1704896540
transform 1 0 22032 0 1 22717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1208
timestamp 1704896540
transform 1 0 22032 0 1 22989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1209
timestamp 1704896540
transform 1 0 18360 0 1 23805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1210
timestamp 1704896540
transform 1 0 22032 0 1 23533
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1211
timestamp 1704896540
transform 1 0 21760 0 1 22173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1212
timestamp 1704896540
transform 1 0 21760 0 1 22581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1213
timestamp 1704896540
transform 1 0 21760 0 1 22309
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1214
timestamp 1704896540
transform 1 0 18360 0 1 23941
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1215
timestamp 1704896540
transform 1 0 20400 0 1 23125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1216
timestamp 1704896540
transform 1 0 22032 0 1 22581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1217
timestamp 1704896540
transform 1 0 20400 0 1 20269
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1218
timestamp 1704896540
transform 1 0 20400 0 1 20677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1219
timestamp 1704896540
transform 1 0 20400 0 1 20405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1220
timestamp 1704896540
transform 1 0 20400 0 1 23397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1221
timestamp 1704896540
transform 1 0 20536 0 1 23533
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1222
timestamp 1704896540
transform 1 0 18360 0 1 24485
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1223
timestamp 1704896540
transform 1 0 18496 0 1 21629
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1224
timestamp 1704896540
transform 1 0 18496 0 1 22173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1225
timestamp 1704896540
transform 1 0 18360 0 1 22989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1226
timestamp 1704896540
transform 1 0 21760 0 1 21357
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1227
timestamp 1704896540
transform 1 0 21760 0 1 21085
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1228
timestamp 1704896540
transform 1 0 20536 0 1 23805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1229
timestamp 1704896540
transform 1 0 20808 0 1 24485
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1230
timestamp 1704896540
transform 1 0 21080 0 1 21085
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1231
timestamp 1704896540
transform 1 0 21080 0 1 21357
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1232
timestamp 1704896540
transform 1 0 18360 0 1 22309
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1233
timestamp 1704896540
transform 1 0 22032 0 1 21765
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1234
timestamp 1704896540
transform 1 0 22032 0 1 21493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1235
timestamp 1704896540
transform 1 0 22032 0 1 21085
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1236
timestamp 1704896540
transform 1 0 22032 0 1 21357
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1237
timestamp 1704896540
transform 1 0 18360 0 1 20541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1238
timestamp 1704896540
transform 1 0 20944 0 1 23125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1239
timestamp 1704896540
transform 1 0 20944 0 1 23397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1240
timestamp 1704896540
transform 1 0 18632 0 1 23941
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1241
timestamp 1704896540
transform 1 0 18632 0 1 24485
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1242
timestamp 1704896540
transform 1 0 20536 0 1 24621
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1243
timestamp 1704896540
transform 1 0 20536 0 1 24349
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1244
timestamp 1704896540
transform 1 0 20808 0 1 23533
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1245
timestamp 1704896540
transform 1 0 18224 0 1 23941
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1246
timestamp 1704896540
transform 1 0 18224 0 1 24213
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1247
timestamp 1704896540
transform 1 0 22168 0 1 21901
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1248
timestamp 1704896540
transform 1 0 20400 0 1 23941
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1249
timestamp 1704896540
transform 1 0 20808 0 1 23805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1250
timestamp 1704896540
transform 1 0 21760 0 1 21765
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1251
timestamp 1704896540
transform 1 0 20808 0 1 22989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1252
timestamp 1704896540
transform 1 0 20808 0 1 22717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1253
timestamp 1704896540
transform 1 0 21488 0 1 24349
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1254
timestamp 1704896540
transform 1 0 21488 0 1 24621
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1255
timestamp 1704896540
transform 1 0 22168 0 1 24213
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1256
timestamp 1704896540
transform 1 0 22168 0 1 23941
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1257
timestamp 1704896540
transform 1 0 21488 0 1 20405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1258
timestamp 1704896540
transform 1 0 21488 0 1 20677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1259
timestamp 1704896540
transform 1 0 21760 0 1 21493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1260
timestamp 1704896540
transform 1 0 20400 0 1 24213
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1261
timestamp 1704896540
transform 1 0 22168 0 1 22173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1262
timestamp 1704896540
transform 1 0 18768 0 1 22989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1263
timestamp 1704896540
transform 1 0 20808 0 1 22173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1264
timestamp 1704896540
transform 1 0 20536 0 1 20813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1265
timestamp 1704896540
transform 1 0 20536 0 1 21085
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1266
timestamp 1704896540
transform 1 0 20808 0 1 21901
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1267
timestamp 1704896540
transform 1 0 18768 0 1 22309
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1268
timestamp 1704896540
transform 1 0 21624 0 1 23941
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1269
timestamp 1704896540
transform 1 0 21624 0 1 24213
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1270
timestamp 1704896540
transform 1 0 21760 0 1 23125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1271
timestamp 1704896540
transform 1 0 21488 0 1 21901
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1272
timestamp 1704896540
transform 1 0 21488 0 1 22173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1273
timestamp 1704896540
transform 1 0 21488 0 1 23397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1274
timestamp 1704896540
transform 1 0 21488 0 1 23125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1275
timestamp 1704896540
transform 1 0 21624 0 1 22989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1276
timestamp 1704896540
transform 1 0 21624 0 1 22717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1277
timestamp 1704896540
transform 1 0 21760 0 1 23397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1278
timestamp 1704896540
transform 1 0 21760 0 1 23805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1279
timestamp 1704896540
transform 1 0 21760 0 1 23533
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1280
timestamp 1704896540
transform 1 0 18632 0 1 22173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1281
timestamp 1704896540
transform 1 0 18632 0 1 20813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1282
timestamp 1704896540
transform 1 0 20400 0 1 24757
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1283
timestamp 1704896540
transform 1 0 20536 0 1 22989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1284
timestamp 1704896540
transform 1 0 20536 0 1 22717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1285
timestamp 1704896540
transform 1 0 20400 0 1 22309
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1286
timestamp 1704896540
transform 1 0 20400 0 1 22581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1287
timestamp 1704896540
transform 1 0 22032 0 1 22309
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1288
timestamp 1704896540
transform 1 0 17000 0 1 22309
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1289
timestamp 1704896540
transform 1 0 16456 0 1 20541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1290
timestamp 1704896540
transform 1 0 17816 0 1 23669
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1291
timestamp 1704896540
transform 1 0 17272 0 1 22173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1292
timestamp 1704896540
transform 1 0 17272 0 1 24213
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1293
timestamp 1704896540
transform 1 0 17000 0 1 22989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1294
timestamp 1704896540
transform 1 0 17272 0 1 23941
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1295
timestamp 1704896540
transform 1 0 17136 0 1 24621
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1296
timestamp 1704896540
transform 1 0 17680 0 1 22989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1297
timestamp 1704896540
transform 1 0 17136 0 1 23941
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1298
timestamp 1704896540
transform 1 0 15504 0 1 22309
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1299
timestamp 1704896540
transform 1 0 17680 0 1 22309
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1300
timestamp 1704896540
transform 1 0 17136 0 1 23125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1301
timestamp 1704896540
transform 1 0 17136 0 1 23805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1302
timestamp 1704896540
transform 1 0 17816 0 1 20541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1303
timestamp 1704896540
transform 1 0 17816 0 1 23125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1304
timestamp 1704896540
transform 1 0 17272 0 1 20813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1305
timestamp 1704896540
transform 1 0 17408 0 1 24757
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1306
timestamp 1704896540
transform 1 0 17408 0 1 20541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1307
timestamp 1704896540
transform 1 0 17952 0 1 24621
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1308
timestamp 1704896540
transform 1 0 17952 0 1 23941
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1309
timestamp 1704896540
transform 1 0 13736 0 1 25029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1310
timestamp 1704896540
transform 1 0 13464 0 1 27885
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1311
timestamp 1704896540
transform 1 0 13736 0 1 29381
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1312
timestamp 1704896540
transform 1 0 13600 0 1 29245
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1313
timestamp 1704896540
transform 1 0 13600 0 1 26525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1314
timestamp 1704896540
transform 1 0 13736 0 1 27749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1315
timestamp 1704896540
transform 1 0 17408 0 1 26389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1316
timestamp 1704896540
transform 1 0 22032 0 1 25029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1317
timestamp 1704896540
transform 1 0 22032 0 1 25301
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1318
timestamp 1704896540
transform 1 0 22032 0 1 27069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1319
timestamp 1704896540
transform 1 0 22032 0 1 27341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1320
timestamp 1704896540
transform 1 0 21760 0 1 26117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1321
timestamp 1704896540
transform 1 0 21760 0 1 25845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1322
timestamp 1704896540
transform 1 0 21760 0 1 25437
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1323
timestamp 1704896540
transform 1 0 22032 0 1 26525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1324
timestamp 1704896540
transform 1 0 22032 0 1 26253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1325
timestamp 1704896540
transform 1 0 22168 0 1 25845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1326
timestamp 1704896540
transform 1 0 22168 0 1 26117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1327
timestamp 1704896540
transform 1 0 21760 0 1 25709
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1328
timestamp 1704896540
transform 1 0 21760 0 1 26253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1329
timestamp 1704896540
transform 1 0 21760 0 1 26525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1330
timestamp 1704896540
transform 1 0 21760 0 1 26933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1331
timestamp 1704896540
transform 1 0 21760 0 1 26661
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1332
timestamp 1704896540
transform 1 0 22032 0 1 26661
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1333
timestamp 1704896540
transform 1 0 22032 0 1 26933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1334
timestamp 1704896540
transform 1 0 22032 0 1 28157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1335
timestamp 1704896540
transform 1 0 22032 0 1 27885
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1336
timestamp 1704896540
transform 1 0 22032 0 1 27477
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1337
timestamp 1704896540
transform 1 0 22032 0 1 27749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1338
timestamp 1704896540
transform 1 0 21760 0 1 29789
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1339
timestamp 1704896540
transform 1 0 21488 0 1 27749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1340
timestamp 1704896540
transform 1 0 21488 0 1 27477
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1341
timestamp 1704896540
transform 1 0 21488 0 1 26253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1342
timestamp 1704896540
transform 1 0 21488 0 1 26525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1343
timestamp 1704896540
transform 1 0 21216 0 1 29789
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1344
timestamp 1704896540
transform 1 0 21352 0 1 25029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1345
timestamp 1704896540
transform 1 0 21352 0 1 25301
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1346
timestamp 1704896540
transform 1 0 21080 0 1 28701
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1347
timestamp 1704896540
transform 1 0 20944 0 1 28837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1348
timestamp 1704896540
transform 1 0 21080 0 1 29245
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1349
timestamp 1704896540
transform 1 0 21080 0 1 28973
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1350
timestamp 1704896540
transform 1 0 21080 0 1 27341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1351
timestamp 1704896540
transform 1 0 21080 0 1 27069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1352
timestamp 1704896540
transform 1 0 21080 0 1 26661
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1353
timestamp 1704896540
transform 1 0 21080 0 1 26933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1354
timestamp 1704896540
transform 1 0 20944 0 1 26933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1355
timestamp 1704896540
transform 1 0 20944 0 1 26661
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1356
timestamp 1704896540
transform 1 0 20400 0 1 28701
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1357
timestamp 1704896540
transform 1 0 20400 0 1 28973
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1358
timestamp 1704896540
transform 1 0 20536 0 1 29789
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1359
timestamp 1704896540
transform 1 0 20536 0 1 29517
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1360
timestamp 1704896540
transform 1 0 20808 0 1 27069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1361
timestamp 1704896540
transform 1 0 20808 0 1 27341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1362
timestamp 1704896540
transform 1 0 20808 0 1 26525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1363
timestamp 1704896540
transform 1 0 20808 0 1 26253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1364
timestamp 1704896540
transform 1 0 20536 0 1 28565
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1365
timestamp 1704896540
transform 1 0 20536 0 1 28293
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1366
timestamp 1704896540
transform 1 0 20536 0 1 27885
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1367
timestamp 1704896540
transform 1 0 20536 0 1 28157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1368
timestamp 1704896540
transform 1 0 20808 0 1 28293
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1369
timestamp 1704896540
transform 1 0 20808 0 1 28565
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1370
timestamp 1704896540
transform 1 0 22168 0 1 25709
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1371
timestamp 1704896540
transform 1 0 20400 0 1 25029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1372
timestamp 1704896540
transform 1 0 22168 0 1 29653
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1373
timestamp 1704896540
transform 1 0 20400 0 1 27749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1374
timestamp 1704896540
transform 1 0 20400 0 1 27477
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1375
timestamp 1704896540
transform 1 0 22168 0 1 25437
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1376
timestamp 1704896540
transform 1 0 22032 0 1 29789
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1377
timestamp 1704896540
transform 1 0 20400 0 1 26661
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1378
timestamp 1704896540
transform 1 0 21624 0 1 25029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1379
timestamp 1704896540
transform 1 0 21624 0 1 25301
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1380
timestamp 1704896540
transform 1 0 20400 0 1 26933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1381
timestamp 1704896540
transform 1 0 20536 0 1 27341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1382
timestamp 1704896540
transform 1 0 21624 0 1 29381
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1383
timestamp 1704896540
transform 1 0 21624 0 1 29653
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1384
timestamp 1704896540
transform 1 0 20536 0 1 27069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1385
timestamp 1704896540
transform 1 0 22168 0 1 29381
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1386
timestamp 1704896540
transform 1 0 21760 0 1 28157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1387
timestamp 1704896540
transform 1 0 21760 0 1 27885
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1388
timestamp 1704896540
transform 1 0 20808 0 1 25301
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1389
timestamp 1704896540
transform 1 0 21624 0 1 27749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1390
timestamp 1704896540
transform 1 0 21624 0 1 27477
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1391
timestamp 1704896540
transform 1 0 21624 0 1 27069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1392
timestamp 1704896540
transform 1 0 21624 0 1 27341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1393
timestamp 1704896540
transform 1 0 20536 0 1 26253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1394
timestamp 1704896540
transform 1 0 20536 0 1 26525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1395
timestamp 1704896540
transform 1 0 15504 0 1 24893
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1396
timestamp 1704896540
transform 1 0 2555 0 1 22604
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1397
timestamp 1704896540
transform 1 0 3808 0 1 20405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1398
timestamp 1704896540
transform 1 0 544 0 1 23397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1399
timestamp 1704896540
transform 1 0 1224 0 1 22173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1400
timestamp 1704896540
transform 1 0 1224 0 1 20405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1401
timestamp 1704896540
transform 1 0 1224 0 1 23805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1402
timestamp 1704896540
transform 1 0 1224 0 1 28973
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1403
timestamp 1704896540
transform 1 0 1224 0 1 25437
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1404
timestamp 1704896540
transform 1 0 1224 0 1 27341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1405
timestamp 1704896540
transform 1 0 1224 0 1 33869
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1406
timestamp 1704896540
transform 1 0 1224 0 1 30605
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1407
timestamp 1704896540
transform 1 0 1224 0 1 38901
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1408
timestamp 1704896540
transform 1 0 1224 0 1 32237
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1409
timestamp 1704896540
transform 1 0 1224 0 1 37405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1410
timestamp 1704896540
transform 1 0 1224 0 1 35501
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1411
timestamp 1704896540
transform 1 0 22168 0 1 32237
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1412
timestamp 1704896540
transform 1 0 22168 0 1 32509
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1413
timestamp 1704896540
transform 1 0 20944 0 1 34549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1414
timestamp 1704896540
transform 1 0 20536 0 1 32237
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1415
timestamp 1704896540
transform 1 0 22168 0 1 30877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1416
timestamp 1704896540
transform 1 0 22168 0 1 30605
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1417
timestamp 1704896540
transform 1 0 22032 0 1 30197
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1418
timestamp 1704896540
transform 1 0 22032 0 1 30469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1419
timestamp 1704896540
transform 1 0 22032 0 1 34141
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1420
timestamp 1704896540
transform 1 0 22032 0 1 34413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1421
timestamp 1704896540
transform 1 0 20536 0 1 32509
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1422
timestamp 1704896540
transform 1 0 22032 0 1 34549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1423
timestamp 1704896540
transform 1 0 20400 0 1 30469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1424
timestamp 1704896540
transform 1 0 20400 0 1 30197
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1425
timestamp 1704896540
transform 1 0 21624 0 1 32237
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1426
timestamp 1704896540
transform 1 0 21624 0 1 32509
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1427
timestamp 1704896540
transform 1 0 22168 0 1 34005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1428
timestamp 1704896540
transform 1 0 22168 0 1 33733
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1429
timestamp 1704896540
transform 1 0 22168 0 1 33325
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1430
timestamp 1704896540
transform 1 0 22168 0 1 33597
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1431
timestamp 1704896540
transform 1 0 21760 0 1 30605
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1432
timestamp 1704896540
transform 1 0 21760 0 1 30877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1433
timestamp 1704896540
transform 1 0 20400 0 1 33733
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1434
timestamp 1704896540
transform 1 0 20400 0 1 33461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1435
timestamp 1704896540
transform 1 0 22032 0 1 32101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1436
timestamp 1704896540
transform 1 0 22032 0 1 31829
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1437
timestamp 1704896540
transform 1 0 21624 0 1 32101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1438
timestamp 1704896540
transform 1 0 21624 0 1 31829
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1439
timestamp 1704896540
transform 1 0 21488 0 1 34413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1440
timestamp 1704896540
transform 1 0 21488 0 1 34141
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1441
timestamp 1704896540
transform 1 0 21352 0 1 33733
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1442
timestamp 1704896540
transform 1 0 21352 0 1 34005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1443
timestamp 1704896540
transform 1 0 20536 0 1 34413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1444
timestamp 1704896540
transform 1 0 21760 0 1 34549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1445
timestamp 1704896540
transform 1 0 21488 0 1 32101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1446
timestamp 1704896540
transform 1 0 21488 0 1 31829
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1447
timestamp 1704896540
transform 1 0 21216 0 1 31421
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1448
timestamp 1704896540
transform 1 0 21216 0 1 31693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1449
timestamp 1704896540
transform 1 0 21216 0 1 30061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1450
timestamp 1704896540
transform 1 0 21488 0 1 30605
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1451
timestamp 1704896540
transform 1 0 21488 0 1 30877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1452
timestamp 1704896540
transform 1 0 22032 0 1 30061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1453
timestamp 1704896540
transform 1 0 21624 0 1 33733
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1454
timestamp 1704896540
transform 1 0 21624 0 1 34005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1455
timestamp 1704896540
transform 1 0 21760 0 1 34413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1456
timestamp 1704896540
transform 1 0 21080 0 1 31013
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1457
timestamp 1704896540
transform 1 0 21080 0 1 31285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1458
timestamp 1704896540
transform 1 0 20944 0 1 31013
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1459
timestamp 1704896540
transform 1 0 20944 0 1 31285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1460
timestamp 1704896540
transform 1 0 21760 0 1 34141
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1461
timestamp 1704896540
transform 1 0 21760 0 1 31013
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1462
timestamp 1704896540
transform 1 0 21760 0 1 31285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1463
timestamp 1704896540
transform 1 0 21624 0 1 31693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1464
timestamp 1704896540
transform 1 0 20944 0 1 31829
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1465
timestamp 1704896540
transform 1 0 20944 0 1 32101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1466
timestamp 1704896540
transform 1 0 21624 0 1 31421
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1467
timestamp 1704896540
transform 1 0 21760 0 1 33597
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1468
timestamp 1704896540
transform 1 0 20808 0 1 32237
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1469
timestamp 1704896540
transform 1 0 20808 0 1 32509
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1470
timestamp 1704896540
transform 1 0 20808 0 1 30877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1471
timestamp 1704896540
transform 1 0 20808 0 1 30605
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1472
timestamp 1704896540
transform 1 0 21760 0 1 33325
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1473
timestamp 1704896540
transform 1 0 20536 0 1 34141
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1474
timestamp 1704896540
transform 1 0 20400 0 1 30877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1475
timestamp 1704896540
transform 1 0 20400 0 1 30605
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1476
timestamp 1704896540
transform 1 0 20400 0 1 31013
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1477
timestamp 1704896540
transform 1 0 20400 0 1 31285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1478
timestamp 1704896540
transform 1 0 20536 0 1 31693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1479
timestamp 1704896540
transform 1 0 21760 0 1 30469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1480
timestamp 1704896540
transform 1 0 21760 0 1 30197
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1481
timestamp 1704896540
transform 1 0 21760 0 1 30061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1482
timestamp 1704896540
transform 1 0 21080 0 1 34549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1483
timestamp 1704896540
transform 1 0 20536 0 1 31421
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1484
timestamp 1704896540
transform 1 0 20400 0 1 31829
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1485
timestamp 1704896540
transform 1 0 20400 0 1 32101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1486
timestamp 1704896540
transform 1 0 20536 0 1 32917
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1487
timestamp 1704896540
transform 1 0 20536 0 1 32645
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1488
timestamp 1704896540
transform 1 0 22168 0 1 31693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1489
timestamp 1704896540
transform 1 0 22168 0 1 31421
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1490
timestamp 1704896540
transform 1 0 22032 0 1 31013
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1491
timestamp 1704896540
transform 1 0 22032 0 1 31285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1492
timestamp 1704896540
transform 1 0 13736 0 1 31965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1493
timestamp 1704896540
transform 1 0 13736 0 1 32101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1494
timestamp 1704896540
transform 1 0 13464 0 1 30605
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1495
timestamp 1704896540
transform 1 0 13600 0 1 30741
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1496
timestamp 1704896540
transform 1 0 13600 0 1 33461
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1497
timestamp 1704896540
transform 1 0 13736 0 1 34821
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1498
timestamp 1704896540
transform 1 0 22168 0 1 38765
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1499
timestamp 1704896540
transform 1 0 22168 0 1 38493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1500
timestamp 1704896540
transform 1 0 22032 0 1 34821
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1501
timestamp 1704896540
transform 1 0 22168 0 1 37677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1502
timestamp 1704896540
transform 1 0 22168 0 1 37949
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1503
timestamp 1704896540
transform 1 0 22168 0 1 38357
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1504
timestamp 1704896540
transform 1 0 22168 0 1 38085
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1505
timestamp 1704896540
transform 1 0 22032 0 1 35365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1506
timestamp 1704896540
transform 1 0 22032 0 1 35637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1507
timestamp 1704896540
transform 1 0 22168 0 1 36045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1508
timestamp 1704896540
transform 1 0 22168 0 1 35773
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1509
timestamp 1704896540
transform 1 0 21216 0 1 35773
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1510
timestamp 1704896540
transform 1 0 21216 0 1 36045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1511
timestamp 1704896540
transform 1 0 21352 0 1 36181
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1512
timestamp 1704896540
transform 1 0 21352 0 1 36453
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1513
timestamp 1704896540
transform 1 0 21488 0 1 38765
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1514
timestamp 1704896540
transform 1 0 21488 0 1 38493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1515
timestamp 1704896540
transform 1 0 21080 0 1 39173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1516
timestamp 1704896540
transform 1 0 21080 0 1 38901
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1517
timestamp 1704896540
transform 1 0 21080 0 1 37949
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1518
timestamp 1704896540
transform 1 0 21080 0 1 37677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1519
timestamp 1704896540
transform 1 0 20944 0 1 35365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1520
timestamp 1704896540
transform 1 0 20944 0 1 35637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1521
timestamp 1704896540
transform 1 0 20808 0 1 35229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1522
timestamp 1704896540
transform 1 0 20808 0 1 34957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1523
timestamp 1704896540
transform 1 0 22032 0 1 36181
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1524
timestamp 1704896540
transform 1 0 22032 0 1 36453
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1525
timestamp 1704896540
transform 1 0 20808 0 1 38901
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1526
timestamp 1704896540
transform 1 0 20808 0 1 39173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1527
timestamp 1704896540
transform 1 0 20808 0 1 39581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1528
timestamp 1704896540
transform 1 0 20808 0 1 39309
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1529
timestamp 1704896540
transform 1 0 20808 0 1 35773
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1530
timestamp 1704896540
transform 1 0 20808 0 1 36045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1531
timestamp 1704896540
transform 1 0 21080 0 1 34821
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1532
timestamp 1704896540
transform 1 0 22032 0 1 39173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1533
timestamp 1704896540
transform 1 0 22032 0 1 38901
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1534
timestamp 1704896540
transform 1 0 22168 0 1 39309
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1535
timestamp 1704896540
transform 1 0 20944 0 1 34821
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1536
timestamp 1704896540
transform 1 0 20808 0 1 36997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1537
timestamp 1704896540
transform 1 0 20808 0 1 37269
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1538
timestamp 1704896540
transform 1 0 21760 0 1 38765
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1539
timestamp 1704896540
transform 1 0 21760 0 1 38493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1540
timestamp 1704896540
transform 1 0 21760 0 1 34957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1541
timestamp 1704896540
transform 1 0 21760 0 1 35229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1542
timestamp 1704896540
transform 1 0 21760 0 1 35637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1543
timestamp 1704896540
transform 1 0 21760 0 1 35365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1544
timestamp 1704896540
transform 1 0 21760 0 1 34821
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1545
timestamp 1704896540
transform 1 0 21624 0 1 38357
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1546
timestamp 1704896540
transform 1 0 21624 0 1 38085
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1547
timestamp 1704896540
transform 1 0 21624 0 1 37677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1548
timestamp 1704896540
transform 1 0 21624 0 1 37949
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1549
timestamp 1704896540
transform 1 0 21624 0 1 38901
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1550
timestamp 1704896540
transform 1 0 21624 0 1 39173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1551
timestamp 1704896540
transform 1 0 21760 0 1 39309
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1552
timestamp 1704896540
transform 1 0 21760 0 1 39581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1553
timestamp 1704896540
transform 1 0 21624 0 1 36453
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1554
timestamp 1704896540
transform 1 0 21624 0 1 36181
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1555
timestamp 1704896540
transform 1 0 21624 0 1 35773
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1556
timestamp 1704896540
transform 1 0 21624 0 1 36045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1557
timestamp 1704896540
transform 1 0 20536 0 1 36589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1558
timestamp 1704896540
transform 1 0 20536 0 1 36861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1559
timestamp 1704896540
transform 1 0 20536 0 1 35637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1560
timestamp 1704896540
transform 1 0 20536 0 1 35365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1561
timestamp 1704896540
transform 1 0 20400 0 1 35229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1562
timestamp 1704896540
transform 1 0 20400 0 1 34957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1563
timestamp 1704896540
transform 1 0 20400 0 1 35773
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1564
timestamp 1704896540
transform 1 0 20400 0 1 36045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1565
timestamp 1704896540
transform 1 0 20400 0 1 36453
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1566
timestamp 1704896540
transform 1 0 20400 0 1 36181
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1567
timestamp 1704896540
transform 1 0 20536 0 1 37677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1568
timestamp 1704896540
transform 1 0 20536 0 1 37405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1569
timestamp 1704896540
transform 1 0 20400 0 1 36997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1570
timestamp 1704896540
transform 1 0 20400 0 1 37269
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1571
timestamp 1704896540
transform 1 0 20400 0 1 39173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1572
timestamp 1704896540
transform 1 0 20400 0 1 38901
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1573
timestamp 1704896540
transform 1 0 20536 0 1 39309
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1574
timestamp 1704896540
transform 1 0 20536 0 1 39581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1575
timestamp 1704896540
transform 1 0 22168 0 1 39581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1576
timestamp 1704896540
transform 1 0 22032 0 1 35229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1577
timestamp 1704896540
transform 1 0 22032 0 1 34957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1578
timestamp 1704896540
transform 1 0 27064 0 1 37133
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1579
timestamp 1704896540
transform 1 0 27064 0 1 37405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1580
timestamp 1704896540
transform 1 0 27200 0 1 20405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1581
timestamp 1704896540
transform 1 0 27200 0 1 20813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1582
timestamp 1704896540
transform 1 0 27200 0 1 25981
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1583
timestamp 1704896540
transform 1 0 27200 0 1 25709
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1584
timestamp 1704896540
transform 1 0 27064 0 1 20133
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1585
timestamp 1704896540
transform 1 0 26928 0 1 37541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1586
timestamp 1704896540
transform 1 0 26928 0 1 37813
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1587
timestamp 1704896540
transform 1 0 26928 0 1 20133
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1588
timestamp 1704896540
transform 1 0 26928 0 1 20405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1589
timestamp 1704896540
transform 1 0 27200 0 1 32237
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1590
timestamp 1704896540
transform 1 0 27200 0 1 31965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1591
timestamp 1704896540
transform 1 0 27200 0 1 33053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1592
timestamp 1704896540
transform 1 0 27200 0 1 32781
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1593
timestamp 1704896540
transform 1 0 26928 0 1 24485
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1594
timestamp 1704896540
transform 1 0 26928 0 1 24757
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1595
timestamp 1704896540
transform 1 0 27200 0 1 29109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1596
timestamp 1704896540
transform 1 0 27200 0 1 28837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1597
timestamp 1704896540
transform 1 0 27064 0 1 28429
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1598
timestamp 1704896540
transform 1 0 27064 0 1 28701
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1599
timestamp 1704896540
transform 1 0 27064 0 1 23941
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1600
timestamp 1704896540
transform 1 0 27064 0 1 23533
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1601
timestamp 1704896540
transform 1 0 27064 0 1 27205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1602
timestamp 1704896540
transform 1 0 27064 0 1 27477
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1603
timestamp 1704896540
transform 1 0 26928 0 1 22037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1604
timestamp 1704896540
transform 1 0 26928 0 1 21765
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1605
timestamp 1704896540
transform 1 0 18768 0 1 19997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1606
timestamp 1704896540
transform 1 0 17816 0 1 19997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1607
timestamp 1704896540
transform 1 0 20400 0 1 19997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1608
timestamp 1704896540
transform 1 0 18360 0 1 19997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1609
timestamp 1704896540
transform 1 0 17408 0 1 19997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1610
timestamp 1704896540
transform 1 0 16456 0 1 19997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1611
timestamp 1704896540
transform 1 0 27200 0 1 58077
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1612
timestamp 1704896540
transform 1 0 27064 0 1 41349
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1613
timestamp 1704896540
transform 1 0 27064 0 1 41077
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1614
timestamp 1704896540
transform 1 0 27200 0 1 49645
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1615
timestamp 1704896540
transform 1 0 27200 0 1 49373
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1616
timestamp 1704896540
transform 1 0 26928 0 1 53589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1617
timestamp 1704896540
transform 1 0 26928 0 1 53317
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1618
timestamp 1704896540
transform 1 0 27064 0 1 53997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1619
timestamp 1704896540
transform 1 0 27064 0 1 53589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1620
timestamp 1704896540
transform 1 0 26928 0 1 58349
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1621
timestamp 1704896540
transform 1 0 26928 0 1 58077
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1622
timestamp 1704896540
transform 1 0 25432 0 1 42845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1623
timestamp 1704896540
transform 1 0 25432 0 1 42437
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1624
timestamp 1704896540
transform 1 0 27200 0 1 52773
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1625
timestamp 1704896540
transform 1 0 27200 0 1 52501
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1626
timestamp 1704896540
transform 1 0 27200 0 1 45293
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1627
timestamp 1704896540
transform 1 0 27200 0 1 45021
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1628
timestamp 1704896540
transform 1 0 27200 0 1 56717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1629
timestamp 1704896540
transform 1 0 27200 0 1 56445
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1630
timestamp 1704896540
transform 1 0 27200 0 1 40941
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1631
timestamp 1704896540
transform 1 0 27200 0 1 40669
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1632
timestamp 1704896540
transform 1 0 27200 0 1 53725
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1633
timestamp 1704896540
transform 1 0 27200 0 1 53997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1634
timestamp 1704896540
transform 1 0 27200 0 1 57669
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1635
timestamp 1704896540
transform 1 0 21760 0 1 43661
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1636
timestamp 1704896540
transform 1 0 21760 0 1 43933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1637
timestamp 1704896540
transform 1 0 22032 0 1 41893
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1638
timestamp 1704896540
transform 1 0 22032 0 1 41621
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1639
timestamp 1704896540
transform 1 0 22168 0 1 40397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1640
timestamp 1704896540
transform 1 0 22168 0 1 40125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1641
timestamp 1704896540
transform 1 0 21760 0 1 44341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1642
timestamp 1704896540
transform 1 0 22032 0 1 39989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1643
timestamp 1704896540
transform 1 0 21080 0 1 43661
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1644
timestamp 1704896540
transform 1 0 21080 0 1 43933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1645
timestamp 1704896540
transform 1 0 20400 0 1 40533
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1646
timestamp 1704896540
transform 1 0 22168 0 1 44477
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1647
timestamp 1704896540
transform 1 0 22032 0 1 44069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1648
timestamp 1704896540
transform 1 0 22032 0 1 44341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1649
timestamp 1704896540
transform 1 0 22168 0 1 40533
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1650
timestamp 1704896540
transform 1 0 22168 0 1 40805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1651
timestamp 1704896540
transform 1 0 21760 0 1 44069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1652
timestamp 1704896540
transform 1 0 21760 0 1 40533
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1653
timestamp 1704896540
transform 1 0 21760 0 1 40805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1654
timestamp 1704896540
transform 1 0 20536 0 1 43117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1655
timestamp 1704896540
transform 1 0 21488 0 1 41213
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1656
timestamp 1704896540
transform 1 0 21488 0 1 40941
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1657
timestamp 1704896540
transform 1 0 20536 0 1 42845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1658
timestamp 1704896540
transform 1 0 20536 0 1 41621
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1659
timestamp 1704896540
transform 1 0 20536 0 1 41349
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1660
timestamp 1704896540
transform 1 0 22032 0 1 42437
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1661
timestamp 1704896540
transform 1 0 22168 0 1 42029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1662
timestamp 1704896540
transform 1 0 22168 0 1 42301
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1663
timestamp 1704896540
transform 1 0 20400 0 1 43933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1664
timestamp 1704896540
transform 1 0 21352 0 1 42437
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1665
timestamp 1704896540
transform 1 0 21352 0 1 42709
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1666
timestamp 1704896540
transform 1 0 20400 0 1 43661
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1667
timestamp 1704896540
transform 1 0 22032 0 1 42709
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1668
timestamp 1704896540
transform 1 0 21760 0 1 42845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1669
timestamp 1704896540
transform 1 0 21760 0 1 43117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1670
timestamp 1704896540
transform 1 0 21760 0 1 43525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1671
timestamp 1704896540
transform 1 0 21760 0 1 43253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1672
timestamp 1704896540
transform 1 0 21760 0 1 42301
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1673
timestamp 1704896540
transform 1 0 21080 0 1 43525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1674
timestamp 1704896540
transform 1 0 21080 0 1 43253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1675
timestamp 1704896540
transform 1 0 20944 0 1 43525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1676
timestamp 1704896540
transform 1 0 21760 0 1 42029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1677
timestamp 1704896540
transform 1 0 21760 0 1 41621
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1678
timestamp 1704896540
transform 1 0 20944 0 1 43253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1679
timestamp 1704896540
transform 1 0 20400 0 1 43525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1680
timestamp 1704896540
transform 1 0 22168 0 1 43117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1681
timestamp 1704896540
transform 1 0 22168 0 1 42845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1682
timestamp 1704896540
transform 1 0 20400 0 1 43253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1683
timestamp 1704896540
transform 1 0 20944 0 1 39989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1684
timestamp 1704896540
transform 1 0 21216 0 1 42845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1685
timestamp 1704896540
transform 1 0 21216 0 1 43117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1686
timestamp 1704896540
transform 1 0 20808 0 1 42437
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1687
timestamp 1704896540
transform 1 0 21760 0 1 41893
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1688
timestamp 1704896540
transform 1 0 21624 0 1 44477
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1689
timestamp 1704896540
transform 1 0 22032 0 1 43933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1690
timestamp 1704896540
transform 1 0 21216 0 1 40397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1691
timestamp 1704896540
transform 1 0 21216 0 1 40125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1692
timestamp 1704896540
transform 1 0 20808 0 1 42709
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1693
timestamp 1704896540
transform 1 0 20536 0 1 44069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1694
timestamp 1704896540
transform 1 0 22032 0 1 43661
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1695
timestamp 1704896540
transform 1 0 22032 0 1 43253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1696
timestamp 1704896540
transform 1 0 22032 0 1 43525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1697
timestamp 1704896540
transform 1 0 20536 0 1 39989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1698
timestamp 1704896540
transform 1 0 20536 0 1 40397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1699
timestamp 1704896540
transform 1 0 21624 0 1 40397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1700
timestamp 1704896540
transform 1 0 20536 0 1 40941
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1701
timestamp 1704896540
transform 1 0 21080 0 1 41621
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1702
timestamp 1704896540
transform 1 0 21080 0 1 41893
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1703
timestamp 1704896540
transform 1 0 20400 0 1 40805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1704
timestamp 1704896540
transform 1 0 21624 0 1 40125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1705
timestamp 1704896540
transform 1 0 20536 0 1 41213
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1706
timestamp 1704896540
transform 1 0 21624 0 1 42709
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1707
timestamp 1704896540
transform 1 0 21624 0 1 42437
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1708
timestamp 1704896540
transform 1 0 20536 0 1 44341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1709
timestamp 1704896540
transform 1 0 21760 0 1 39989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1710
timestamp 1704896540
transform 1 0 20536 0 1 40125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1711
timestamp 1704896540
transform 1 0 20400 0 1 44477
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1712
timestamp 1704896540
transform 1 0 22168 0 1 44749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1713
timestamp 1704896540
transform 1 0 22032 0 1 46245
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1714
timestamp 1704896540
transform 1 0 22032 0 1 45973
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1715
timestamp 1704896540
transform 1 0 20400 0 1 47061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1716
timestamp 1704896540
transform 1 0 22032 0 1 48421
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1717
timestamp 1704896540
transform 1 0 22032 0 1 48693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1718
timestamp 1704896540
transform 1 0 22032 0 1 48285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1719
timestamp 1704896540
transform 1 0 22032 0 1 48013
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1720
timestamp 1704896540
transform 1 0 22032 0 1 47877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1721
timestamp 1704896540
transform 1 0 22032 0 1 47605
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1722
timestamp 1704896540
transform 1 0 20400 0 1 49237
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1723
timestamp 1704896540
transform 1 0 20400 0 1 49509
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1724
timestamp 1704896540
transform 1 0 21488 0 1 48013
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1725
timestamp 1704896540
transform 1 0 21488 0 1 48285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1726
timestamp 1704896540
transform 1 0 21488 0 1 47061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1727
timestamp 1704896540
transform 1 0 21488 0 1 46789
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1728
timestamp 1704896540
transform 1 0 20536 0 1 47469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1729
timestamp 1704896540
transform 1 0 20536 0 1 45293
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1730
timestamp 1704896540
transform 1 0 20536 0 1 45565
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1731
timestamp 1704896540
transform 1 0 20536 0 1 47197
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1732
timestamp 1704896540
transform 1 0 21216 0 1 48829
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1733
timestamp 1704896540
transform 1 0 21216 0 1 49101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1734
timestamp 1704896540
transform 1 0 20536 0 1 44885
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1735
timestamp 1704896540
transform 1 0 21352 0 1 47877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1736
timestamp 1704896540
transform 1 0 21352 0 1 47605
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1737
timestamp 1704896540
transform 1 0 20536 0 1 45157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1738
timestamp 1704896540
transform 1 0 21352 0 1 49509
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1739
timestamp 1704896540
transform 1 0 20400 0 1 47877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1740
timestamp 1704896540
transform 1 0 20400 0 1 47605
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1741
timestamp 1704896540
transform 1 0 21488 0 1 45837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1742
timestamp 1704896540
transform 1 0 21488 0 1 45565
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1743
timestamp 1704896540
transform 1 0 21352 0 1 44885
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1744
timestamp 1704896540
transform 1 0 21352 0 1 45157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1745
timestamp 1704896540
transform 1 0 20400 0 1 44749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1746
timestamp 1704896540
transform 1 0 20536 0 1 49101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1747
timestamp 1704896540
transform 1 0 20536 0 1 48829
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1748
timestamp 1704896540
transform 1 0 21760 0 1 48421
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1749
timestamp 1704896540
transform 1 0 21760 0 1 48693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1750
timestamp 1704896540
transform 1 0 21080 0 1 47877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1751
timestamp 1704896540
transform 1 0 21080 0 1 47605
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1752
timestamp 1704896540
transform 1 0 21080 0 1 47197
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1753
timestamp 1704896540
transform 1 0 21080 0 1 47469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1754
timestamp 1704896540
transform 1 0 20536 0 1 48013
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1755
timestamp 1704896540
transform 1 0 20536 0 1 48285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1756
timestamp 1704896540
transform 1 0 20536 0 1 48693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1757
timestamp 1704896540
transform 1 0 20536 0 1 48421
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1758
timestamp 1704896540
transform 1 0 21080 0 1 45429
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1759
timestamp 1704896540
transform 1 0 21080 0 1 45157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1760
timestamp 1704896540
transform 1 0 21760 0 1 48013
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1761
timestamp 1704896540
transform 1 0 21760 0 1 48285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1762
timestamp 1704896540
transform 1 0 20400 0 1 46789
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1763
timestamp 1704896540
transform 1 0 22032 0 1 46789
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1764
timestamp 1704896540
transform 1 0 22032 0 1 47061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1765
timestamp 1704896540
transform 1 0 22168 0 1 47469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1766
timestamp 1704896540
transform 1 0 22168 0 1 47197
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1767
timestamp 1704896540
transform 1 0 20808 0 1 46381
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1768
timestamp 1704896540
transform 1 0 20808 0 1 46653
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1769
timestamp 1704896540
transform 1 0 21760 0 1 47197
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1770
timestamp 1704896540
transform 1 0 21760 0 1 47469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1771
timestamp 1704896540
transform 1 0 21760 0 1 47877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1772
timestamp 1704896540
transform 1 0 21760 0 1 47605
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1773
timestamp 1704896540
transform 1 0 21624 0 1 47061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1774
timestamp 1704896540
transform 1 0 21624 0 1 46789
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1775
timestamp 1704896540
transform 1 0 20808 0 1 46789
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1776
timestamp 1704896540
transform 1 0 20808 0 1 47061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1777
timestamp 1704896540
transform 1 0 21760 0 1 45973
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1778
timestamp 1704896540
transform 1 0 21760 0 1 46245
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1779
timestamp 1704896540
transform 1 0 21760 0 1 46653
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1780
timestamp 1704896540
transform 1 0 21760 0 1 46381
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1781
timestamp 1704896540
transform 1 0 21624 0 1 44749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1782
timestamp 1704896540
transform 1 0 20808 0 1 48285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1783
timestamp 1704896540
transform 1 0 20808 0 1 48013
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1784
timestamp 1704896540
transform 1 0 22168 0 1 46381
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1785
timestamp 1704896540
transform 1 0 22168 0 1 46653
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1786
timestamp 1704896540
transform 1 0 1224 0 1 42301
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1787
timestamp 1704896540
transform 1 0 1224 0 1 49101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1788
timestamp 1704896540
transform 1 0 1224 0 1 43933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1789
timestamp 1704896540
transform 1 0 1224 0 1 47469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1790
timestamp 1704896540
transform 1 0 1224 0 1 40533
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1791
timestamp 1704896540
transform 1 0 1224 0 1 45837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1792
timestamp 1704896540
transform 1 0 1224 0 1 50733
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1793
timestamp 1704896540
transform 1 0 1224 0 1 53997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1794
timestamp 1704896540
transform 1 0 1224 0 1 52365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1795
timestamp 1704896540
transform 1 0 1224 0 1 59165
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1796
timestamp 1704896540
transform 1 0 1224 0 1 55901
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1797
timestamp 1704896540
transform 1 0 1224 0 1 57397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1798
timestamp 1704896540
transform 1 0 20536 0 1 53589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1799
timestamp 1704896540
transform 1 0 21080 0 1 53045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1800
timestamp 1704896540
transform 1 0 21216 0 1 50325
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1801
timestamp 1704896540
transform 1 0 21216 0 1 50597
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1802
timestamp 1704896540
transform 1 0 21216 0 1 51957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1803
timestamp 1704896540
transform 1 0 21216 0 1 52229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1804
timestamp 1704896540
transform 1 0 21080 0 1 52773
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1805
timestamp 1704896540
transform 1 0 20944 0 1 53045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1806
timestamp 1704896540
transform 1 0 21488 0 1 51821
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1807
timestamp 1704896540
transform 1 0 21488 0 1 51549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1808
timestamp 1704896540
transform 1 0 21352 0 1 51141
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1809
timestamp 1704896540
transform 1 0 21352 0 1 51413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1810
timestamp 1704896540
transform 1 0 21352 0 1 49781
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1811
timestamp 1704896540
transform 1 0 21488 0 1 54269
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1812
timestamp 1704896540
transform 1 0 20944 0 1 52773
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1813
timestamp 1704896540
transform 1 0 21488 0 1 53861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1814
timestamp 1704896540
transform 1 0 21488 0 1 53589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1815
timestamp 1704896540
transform 1 0 21080 0 1 52229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1816
timestamp 1704896540
transform 1 0 21080 0 1 51957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1817
timestamp 1704896540
transform 1 0 20944 0 1 52229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1818
timestamp 1704896540
transform 1 0 20944 0 1 51957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1819
timestamp 1704896540
transform 1 0 20536 0 1 53861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1820
timestamp 1704896540
transform 1 0 21624 0 1 51413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1821
timestamp 1704896540
transform 1 0 21624 0 1 51141
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1822
timestamp 1704896540
transform 1 0 21624 0 1 50733
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1823
timestamp 1704896540
transform 1 0 21624 0 1 51005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1824
timestamp 1704896540
transform 1 0 20400 0 1 54269
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1825
timestamp 1704896540
transform 1 0 20400 0 1 53997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1826
timestamp 1704896540
transform 1 0 20536 0 1 51957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1827
timestamp 1704896540
transform 1 0 20536 0 1 52229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1828
timestamp 1704896540
transform 1 0 20536 0 1 52637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1829
timestamp 1704896540
transform 1 0 21080 0 1 51005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1830
timestamp 1704896540
transform 1 0 21080 0 1 50733
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1831
timestamp 1704896540
transform 1 0 20808 0 1 50733
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1832
timestamp 1704896540
transform 1 0 20808 0 1 51005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1833
timestamp 1704896540
transform 1 0 21760 0 1 53045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1834
timestamp 1704896540
transform 1 0 21760 0 1 52773
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1835
timestamp 1704896540
transform 1 0 20808 0 1 51141
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1836
timestamp 1704896540
transform 1 0 20808 0 1 51413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1837
timestamp 1704896540
transform 1 0 20536 0 1 52365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1838
timestamp 1704896540
transform 1 0 20400 0 1 50053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1839
timestamp 1704896540
transform 1 0 20400 0 1 50325
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1840
timestamp 1704896540
transform 1 0 20536 0 1 53453
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1841
timestamp 1704896540
transform 1 0 20536 0 1 53181
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1842
timestamp 1704896540
transform 1 0 20400 0 1 52773
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1843
timestamp 1704896540
transform 1 0 22168 0 1 50189
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1844
timestamp 1704896540
transform 1 0 22168 0 1 49917
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1845
timestamp 1704896540
transform 1 0 21760 0 1 51549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1846
timestamp 1704896540
transform 1 0 21760 0 1 51821
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1847
timestamp 1704896540
transform 1 0 22032 0 1 54269
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1848
timestamp 1704896540
transform 1 0 20400 0 1 53045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1849
timestamp 1704896540
transform 1 0 20400 0 1 51005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1850
timestamp 1704896540
transform 1 0 21624 0 1 54269
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1851
timestamp 1704896540
transform 1 0 20400 0 1 50733
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1852
timestamp 1704896540
transform 1 0 20536 0 1 51821
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1853
timestamp 1704896540
transform 1 0 22032 0 1 51141
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1854
timestamp 1704896540
transform 1 0 22032 0 1 51413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1855
timestamp 1704896540
transform 1 0 22168 0 1 51821
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1856
timestamp 1704896540
transform 1 0 22168 0 1 51549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1857
timestamp 1704896540
transform 1 0 20536 0 1 51549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1858
timestamp 1704896540
transform 1 0 21624 0 1 50189
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1859
timestamp 1704896540
transform 1 0 21624 0 1 49917
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1860
timestamp 1704896540
transform 1 0 21624 0 1 52637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1861
timestamp 1704896540
transform 1 0 22032 0 1 52773
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1862
timestamp 1704896540
transform 1 0 22032 0 1 53045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1863
timestamp 1704896540
transform 1 0 21624 0 1 52365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1864
timestamp 1704896540
transform 1 0 21624 0 1 51957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1865
timestamp 1704896540
transform 1 0 21624 0 1 52229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1866
timestamp 1704896540
transform 1 0 21760 0 1 50325
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1867
timestamp 1704896540
transform 1 0 22032 0 1 51005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1868
timestamp 1704896540
transform 1 0 22032 0 1 50733
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1869
timestamp 1704896540
transform 1 0 22168 0 1 50325
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1870
timestamp 1704896540
transform 1 0 22168 0 1 50597
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1871
timestamp 1704896540
transform 1 0 22032 0 1 52637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1872
timestamp 1704896540
transform 1 0 22032 0 1 52365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1873
timestamp 1704896540
transform 1 0 22032 0 1 51957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1874
timestamp 1704896540
transform 1 0 22032 0 1 52229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1875
timestamp 1704896540
transform 1 0 21760 0 1 50597
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1876
timestamp 1704896540
transform 1 0 21488 0 1 56717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1877
timestamp 1704896540
transform 1 0 21488 0 1 56989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1878
timestamp 1704896540
transform 1 0 21488 0 1 55357
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1879
timestamp 1704896540
transform 1 0 21488 0 1 55085
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1880
timestamp 1704896540
transform 1 0 20400 0 1 56173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1881
timestamp 1704896540
transform 1 0 21080 0 1 59029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1882
timestamp 1704896540
transform 1 0 21080 0 1 59301
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1883
timestamp 1704896540
transform 1 0 20944 0 1 59029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1884
timestamp 1704896540
transform 1 0 20944 0 1 59301
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1885
timestamp 1704896540
transform 1 0 21080 0 1 55357
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1886
timestamp 1704896540
transform 1 0 21080 0 1 55085
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1887
timestamp 1704896540
transform 1 0 21080 0 1 54677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1888
timestamp 1704896540
transform 1 0 21080 0 1 54949
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1889
timestamp 1704896540
transform 1 0 20944 0 1 54677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1890
timestamp 1704896540
transform 1 0 20944 0 1 54949
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1891
timestamp 1704896540
transform 1 0 20808 0 1 57533
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1892
timestamp 1704896540
transform 1 0 20808 0 1 57805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1893
timestamp 1704896540
transform 1 0 20808 0 1 55765
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1894
timestamp 1704896540
transform 1 0 20808 0 1 55493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1895
timestamp 1704896540
transform 1 0 20808 0 1 55085
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1896
timestamp 1704896540
transform 1 0 20808 0 1 55357
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1897
timestamp 1704896540
transform 1 0 22168 0 1 58893
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1898
timestamp 1704896540
transform 1 0 22168 0 1 58621
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1899
timestamp 1704896540
transform 1 0 22032 0 1 54949
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1900
timestamp 1704896540
transform 1 0 22032 0 1 54677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1901
timestamp 1704896540
transform 1 0 20400 0 1 57941
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1902
timestamp 1704896540
transform 1 0 22168 0 1 58485
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1903
timestamp 1704896540
transform 1 0 22168 0 1 58213
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1904
timestamp 1704896540
transform 1 0 22168 0 1 55085
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1905
timestamp 1704896540
transform 1 0 22168 0 1 55357
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1906
timestamp 1704896540
transform 1 0 22168 0 1 56717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1907
timestamp 1704896540
transform 1 0 22168 0 1 56989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1908
timestamp 1704896540
transform 1 0 22032 0 1 59029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1909
timestamp 1704896540
transform 1 0 22032 0 1 59301
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1910
timestamp 1704896540
transform 1 0 22032 0 1 55493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1911
timestamp 1704896540
transform 1 0 22032 0 1 55765
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1912
timestamp 1704896540
transform 1 0 21080 0 1 58213
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1913
timestamp 1704896540
transform 1 0 21080 0 1 58485
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1914
timestamp 1704896540
transform 1 0 20808 0 1 58213
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1915
timestamp 1704896540
transform 1 0 20808 0 1 58485
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1916
timestamp 1704896540
transform 1 0 21080 0 1 55901
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1917
timestamp 1704896540
transform 1 0 21080 0 1 56173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1918
timestamp 1704896540
transform 1 0 22032 0 1 56581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1919
timestamp 1704896540
transform 1 0 22032 0 1 56309
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1920
timestamp 1704896540
transform 1 0 22032 0 1 55901
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1921
timestamp 1704896540
transform 1 0 22032 0 1 56173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1922
timestamp 1704896540
transform 1 0 20944 0 1 55901
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1923
timestamp 1704896540
transform 1 0 20944 0 1 56173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1924
timestamp 1704896540
transform 1 0 20944 0 1 56581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1925
timestamp 1704896540
transform 1 0 20944 0 1 56309
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1926
timestamp 1704896540
transform 1 0 21760 0 1 55901
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1927
timestamp 1704896540
transform 1 0 21760 0 1 56173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1928
timestamp 1704896540
transform 1 0 21624 0 1 56989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1929
timestamp 1704896540
transform 1 0 21624 0 1 56717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1930
timestamp 1704896540
transform 1 0 21624 0 1 56309
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1931
timestamp 1704896540
transform 1 0 21624 0 1 56581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1932
timestamp 1704896540
transform 1 0 21624 0 1 54949
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1933
timestamp 1704896540
transform 1 0 21624 0 1 54677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1934
timestamp 1704896540
transform 1 0 20400 0 1 58213
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1935
timestamp 1704896540
transform 1 0 21624 0 1 59301
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1936
timestamp 1704896540
transform 1 0 21624 0 1 59029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1937
timestamp 1704896540
transform 1 0 21624 0 1 58893
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1938
timestamp 1704896540
transform 1 0 21624 0 1 58621
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1939
timestamp 1704896540
transform 1 0 21760 0 1 58485
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1940
timestamp 1704896540
transform 1 0 21760 0 1 58213
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1941
timestamp 1704896540
transform 1 0 21624 0 1 55765
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1942
timestamp 1704896540
transform 1 0 21624 0 1 55493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1943
timestamp 1704896540
transform 1 0 21624 0 1 55085
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1944
timestamp 1704896540
transform 1 0 21624 0 1 55357
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1945
timestamp 1704896540
transform 1 0 20536 0 1 57805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1946
timestamp 1704896540
transform 1 0 20536 0 1 57533
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1947
timestamp 1704896540
transform 1 0 20536 0 1 56717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1948
timestamp 1704896540
transform 1 0 20536 0 1 56989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1949
timestamp 1704896540
transform 1 0 20536 0 1 57397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1950
timestamp 1704896540
transform 1 0 20536 0 1 57125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1951
timestamp 1704896540
transform 1 0 20400 0 1 55493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1952
timestamp 1704896540
transform 1 0 20400 0 1 55765
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1953
timestamp 1704896540
transform 1 0 20400 0 1 54949
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1954
timestamp 1704896540
transform 1 0 20400 0 1 54677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1955
timestamp 1704896540
transform 1 0 20400 0 1 56581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1956
timestamp 1704896540
transform 1 0 20400 0 1 56309
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1957
timestamp 1704896540
transform 1 0 20400 0 1 55901
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1958
timestamp 1704896540
transform 1 0 21488 0 1 54541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1959
timestamp 1704896540
transform 1 0 22032 0 1 54541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1960
timestamp 1704896540
transform 1 0 21624 0 1 54541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1961
timestamp 1704896540
transform 1 0 21488 0 1 62973
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1962
timestamp 1704896540
transform 1 0 21488 0 1 63245
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1963
timestamp 1704896540
transform 1 0 21624 0 1 60661
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1964
timestamp 1704896540
transform 1 0 21624 0 1 60933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1965
timestamp 1704896540
transform 1 0 21352 0 1 59845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1966
timestamp 1704896540
transform 1 0 21352 0 1 60117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1967
timestamp 1704896540
transform 1 0 21624 0 1 61341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1968
timestamp 1704896540
transform 1 0 21488 0 1 64197
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1969
timestamp 1704896540
transform 1 0 21216 0 1 63789
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1970
timestamp 1704896540
transform 1 0 21216 0 1 64061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1971
timestamp 1704896540
transform 1 0 21760 0 1 63381
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1972
timestamp 1704896540
transform 1 0 21760 0 1 63653
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1973
timestamp 1704896540
transform 1 0 21760 0 1 64061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1974
timestamp 1704896540
transform 1 0 21760 0 1 63789
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1975
timestamp 1704896540
transform 1 0 20536 0 1 60525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1976
timestamp 1704896540
transform 1 0 20536 0 1 60253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1977
timestamp 1704896540
transform 1 0 21624 0 1 61069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1978
timestamp 1704896540
transform 1 0 20536 0 1 64197
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1979
timestamp 1704896540
transform 1 0 20400 0 1 60661
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1980
timestamp 1704896540
transform 1 0 20400 0 1 60933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1981
timestamp 1704896540
transform 1 0 20536 0 1 60117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1982
timestamp 1704896540
transform 1 0 20536 0 1 59845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1983
timestamp 1704896540
transform 1 0 20536 0 1 61069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1984
timestamp 1704896540
transform 1 0 20536 0 1 61341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1985
timestamp 1704896540
transform 1 0 20536 0 1 59709
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1986
timestamp 1704896540
transform 1 0 20808 0 1 63245
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1987
timestamp 1704896540
transform 1 0 22032 0 1 60253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1988
timestamp 1704896540
transform 1 0 22032 0 1 60525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1989
timestamp 1704896540
transform 1 0 20400 0 1 61477
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1990
timestamp 1704896540
transform 1 0 20400 0 1 61749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1991
timestamp 1704896540
transform 1 0 20536 0 1 62157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1992
timestamp 1704896540
transform 1 0 20536 0 1 61885
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1993
timestamp 1704896540
transform 1 0 20536 0 1 64061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1994
timestamp 1704896540
transform 1 0 20536 0 1 63789
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1995
timestamp 1704896540
transform 1 0 20536 0 1 63381
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1996
timestamp 1704896540
transform 1 0 20536 0 1 63653
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1997
timestamp 1704896540
transform 1 0 22168 0 1 62837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1998
timestamp 1704896540
transform 1 0 22168 0 1 62565
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_1999
timestamp 1704896540
transform 1 0 21624 0 1 60117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2000
timestamp 1704896540
transform 1 0 21624 0 1 59845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2001
timestamp 1704896540
transform 1 0 20808 0 1 62973
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2002
timestamp 1704896540
transform 1 0 21624 0 1 59709
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2003
timestamp 1704896540
transform 1 0 22032 0 1 61341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2004
timestamp 1704896540
transform 1 0 21624 0 1 63245
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2005
timestamp 1704896540
transform 1 0 22168 0 1 60117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2006
timestamp 1704896540
transform 1 0 20808 0 1 59709
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2007
timestamp 1704896540
transform 1 0 22168 0 1 59845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2008
timestamp 1704896540
transform 1 0 22168 0 1 63245
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2009
timestamp 1704896540
transform 1 0 21624 0 1 62973
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2010
timestamp 1704896540
transform 1 0 21760 0 1 62565
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2011
timestamp 1704896540
transform 1 0 20808 0 1 63653
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2012
timestamp 1704896540
transform 1 0 20808 0 1 63381
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2013
timestamp 1704896540
transform 1 0 22168 0 1 62973
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2014
timestamp 1704896540
transform 1 0 22032 0 1 63381
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2015
timestamp 1704896540
transform 1 0 20808 0 1 62429
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2016
timestamp 1704896540
transform 1 0 21488 0 1 59709
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2017
timestamp 1704896540
transform 1 0 20808 0 1 62157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2018
timestamp 1704896540
transform 1 0 21352 0 1 60933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2019
timestamp 1704896540
transform 1 0 21352 0 1 60661
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2020
timestamp 1704896540
transform 1 0 22032 0 1 63653
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2021
timestamp 1704896540
transform 1 0 22032 0 1 64061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2022
timestamp 1704896540
transform 1 0 22032 0 1 63789
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2023
timestamp 1704896540
transform 1 0 22032 0 1 59709
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2024
timestamp 1704896540
transform 1 0 21080 0 1 59709
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2025
timestamp 1704896540
transform 1 0 20808 0 1 64197
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2026
timestamp 1704896540
transform 1 0 21080 0 1 60933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2027
timestamp 1704896540
transform 1 0 21080 0 1 60661
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2028
timestamp 1704896540
transform 1 0 21080 0 1 60253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2029
timestamp 1704896540
transform 1 0 21080 0 1 60525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2030
timestamp 1704896540
transform 1 0 20944 0 1 60253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2031
timestamp 1704896540
transform 1 0 20944 0 1 60525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2032
timestamp 1704896540
transform 1 0 21080 0 1 61477
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2033
timestamp 1704896540
transform 1 0 21080 0 1 61749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2034
timestamp 1704896540
transform 1 0 20944 0 1 61477
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2035
timestamp 1704896540
transform 1 0 20944 0 1 61749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2036
timestamp 1704896540
transform 1 0 21080 0 1 64061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2037
timestamp 1704896540
transform 1 0 21080 0 1 63789
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2038
timestamp 1704896540
transform 1 0 20944 0 1 64061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2039
timestamp 1704896540
transform 1 0 20944 0 1 63789
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2040
timestamp 1704896540
transform 1 0 21760 0 1 62837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2041
timestamp 1704896540
transform 1 0 21624 0 1 64197
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2042
timestamp 1704896540
transform 1 0 21760 0 1 60525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2043
timestamp 1704896540
transform 1 0 21760 0 1 60253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2044
timestamp 1704896540
transform 1 0 22032 0 1 64197
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2045
timestamp 1704896540
transform 1 0 22032 0 1 61069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2046
timestamp 1704896540
transform 1 0 22032 0 1 60933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2047
timestamp 1704896540
transform 1 0 22032 0 1 60661
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2048
timestamp 1704896540
transform 1 0 21352 0 1 66917
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2049
timestamp 1704896540
transform 1 0 21352 0 1 67189
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2050
timestamp 1704896540
transform 1 0 21488 0 1 64469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2051
timestamp 1704896540
transform 1 0 20536 0 1 64469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2052
timestamp 1704896540
transform 1 0 20536 0 1 66101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2053
timestamp 1704896540
transform 1 0 20536 0 1 65829
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2054
timestamp 1704896540
transform 1 0 20400 0 1 66917
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2055
timestamp 1704896540
transform 1 0 20400 0 1 66645
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2056
timestamp 1704896540
transform 1 0 20400 0 1 65693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2057
timestamp 1704896540
transform 1 0 20400 0 1 65421
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2058
timestamp 1704896540
transform 1 0 20400 0 1 64605
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2059
timestamp 1704896540
transform 1 0 20400 0 1 64877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2060
timestamp 1704896540
transform 1 0 20400 0 1 65285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2061
timestamp 1704896540
transform 1 0 20400 0 1 65013
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2062
timestamp 1704896540
transform 1 0 22032 0 1 66781
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2063
timestamp 1704896540
transform 1 0 22032 0 1 66509
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2064
timestamp 1704896540
transform 1 0 20808 0 1 65693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2065
timestamp 1704896540
transform 1 0 20808 0 1 65421
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2066
timestamp 1704896540
transform 1 0 21080 0 1 67189
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2067
timestamp 1704896540
transform 1 0 21080 0 1 66917
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2068
timestamp 1704896540
transform 1 0 20944 0 1 67189
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2069
timestamp 1704896540
transform 1 0 20944 0 1 66917
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2070
timestamp 1704896540
transform 1 0 21624 0 1 64469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2071
timestamp 1704896540
transform 1 0 21760 0 1 64605
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2072
timestamp 1704896540
transform 1 0 21760 0 1 64877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2073
timestamp 1704896540
transform 1 0 21760 0 1 65285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2074
timestamp 1704896540
transform 1 0 21760 0 1 65013
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2075
timestamp 1704896540
transform 1 0 21624 0 1 66781
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2076
timestamp 1704896540
transform 1 0 21624 0 1 66509
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2077
timestamp 1704896540
transform 1 0 21760 0 1 66917
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2078
timestamp 1704896540
transform 1 0 21760 0 1 67189
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2079
timestamp 1704896540
transform 1 0 20808 0 1 64469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2080
timestamp 1704896540
transform 1 0 22032 0 1 64469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2081
timestamp 1704896540
transform 1 0 22032 0 1 65285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2082
timestamp 1704896540
transform 1 0 22032 0 1 65013
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2083
timestamp 1704896540
transform 1 0 22032 0 1 64605
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2084
timestamp 1704896540
transform 1 0 22032 0 1 64877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2085
timestamp 1704896540
transform 1 0 22032 0 1 66917
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2086
timestamp 1704896540
transform 1 0 22032 0 1 67189
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2087
timestamp 1704896540
transform 1 0 21488 0 1 64877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2088
timestamp 1704896540
transform 1 0 21488 0 1 64605
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2089
timestamp 1704896540
transform 1 0 1224 0 1 64061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2090
timestamp 1704896540
transform 1 0 1224 0 1 60797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2091
timestamp 1704896540
transform 1 0 1224 0 1 69093
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2092
timestamp 1704896540
transform 1 0 1224 0 1 65965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2093
timestamp 1704896540
transform 1 0 1224 0 1 67597
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2094
timestamp 1704896540
transform 1 0 1224 0 1 62429
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2095
timestamp 1704896540
transform 1 0 1224 0 1 70861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2096
timestamp 1704896540
transform 1 0 1224 0 1 72493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2097
timestamp 1704896540
transform 1 0 5440 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2098
timestamp 1704896540
transform 1 0 5440 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2099
timestamp 1704896540
transform 1 0 3944 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2100
timestamp 1704896540
transform 1 0 3944 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2101
timestamp 1704896540
transform 1 0 2176 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2102
timestamp 1704896540
transform 1 0 2176 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2103
timestamp 1704896540
transform 1 0 1224 0 1 75893
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2104
timestamp 1704896540
transform 1 0 1224 0 1 74397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2105
timestamp 1704896540
transform 1 0 10472 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2106
timestamp 1704896540
transform 1 0 10472 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2107
timestamp 1704896540
transform 1 0 8976 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2108
timestamp 1704896540
transform 1 0 8976 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2109
timestamp 1704896540
transform 1 0 7208 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2110
timestamp 1704896540
transform 1 0 7208 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2111
timestamp 1704896540
transform 1 0 15640 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2112
timestamp 1704896540
transform 1 0 14008 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2113
timestamp 1704896540
transform 1 0 14008 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2114
timestamp 1704896540
transform 1 0 12240 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2115
timestamp 1704896540
transform 1 0 12240 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2116
timestamp 1704896540
transform 1 0 17408 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2117
timestamp 1704896540
transform 1 0 17408 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2118
timestamp 1704896540
transform 1 0 15640 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2119
timestamp 1704896540
transform 1 0 22168 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2120
timestamp 1704896540
transform 1 0 20672 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2121
timestamp 1704896540
transform 1 0 20672 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2122
timestamp 1704896540
transform 1 0 18904 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2123
timestamp 1704896540
transform 1 0 18904 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2124
timestamp 1704896540
transform 1 0 23936 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2125
timestamp 1704896540
transform 1 0 23936 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2126
timestamp 1704896540
transform 1 0 22168 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2127
timestamp 1704896540
transform 1 0 36584 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2128
timestamp 1704896540
transform 1 0 44064 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2129
timestamp 1704896540
transform 1 0 44064 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2130
timestamp 1704896540
transform 1 0 40256 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2131
timestamp 1704896540
transform 1 0 40256 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2132
timestamp 1704896540
transform 1 0 43384 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2133
timestamp 1704896540
transform 1 0 43384 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2134
timestamp 1704896540
transform 1 0 42840 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2135
timestamp 1704896540
transform 1 0 42840 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2136
timestamp 1704896540
transform 1 0 47736 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2137
timestamp 1704896540
transform 1 0 47736 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2138
timestamp 1704896540
transform 1 0 38352 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2139
timestamp 1704896540
transform 1 0 38352 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2140
timestamp 1704896540
transform 1 0 39304 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2141
timestamp 1704896540
transform 1 0 39304 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2142
timestamp 1704896540
transform 1 0 47056 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2143
timestamp 1704896540
transform 1 0 47056 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2144
timestamp 1704896540
transform 1 0 46512 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2145
timestamp 1704896540
transform 1 0 46512 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2146
timestamp 1704896540
transform 1 0 41888 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2147
timestamp 1704896540
transform 1 0 41888 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2148
timestamp 1704896540
transform 1 0 37808 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2149
timestamp 1704896540
transform 1 0 37808 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2150
timestamp 1704896540
transform 1 0 45832 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2151
timestamp 1704896540
transform 1 0 45832 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2152
timestamp 1704896540
transform 1 0 39032 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2153
timestamp 1704896540
transform 1 0 39032 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2154
timestamp 1704896540
transform 1 0 36584 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2155
timestamp 1704896540
transform 1 0 33320 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2156
timestamp 1704896540
transform 1 0 33320 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2157
timestamp 1704896540
transform 1 0 32776 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2158
timestamp 1704896540
transform 1 0 32776 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2159
timestamp 1704896540
transform 1 0 29240 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2160
timestamp 1704896540
transform 1 0 30600 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2161
timestamp 1704896540
transform 1 0 30600 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2162
timestamp 1704896540
transform 1 0 30328 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2163
timestamp 1704896540
transform 1 0 31688 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2164
timestamp 1704896540
transform 1 0 35768 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2165
timestamp 1704896540
transform 1 0 35768 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2166
timestamp 1704896540
transform 1 0 31688 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2167
timestamp 1704896540
transform 1 0 31552 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2168
timestamp 1704896540
transform 1 0 35224 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2169
timestamp 1704896540
transform 1 0 35224 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2170
timestamp 1704896540
transform 1 0 27064 0 1 62837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2171
timestamp 1704896540
transform 1 0 27064 0 1 62293
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2172
timestamp 1704896540
transform 1 0 26928 0 1 65557
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2173
timestamp 1704896540
transform 1 0 26928 0 1 65829
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2174
timestamp 1704896540
transform 1 0 27200 0 1 65421
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2175
timestamp 1704896540
transform 1 0 27200 0 1 65149
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2176
timestamp 1704896540
transform 1 0 27200 0 1 67053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2177
timestamp 1704896540
transform 1 0 27200 0 1 66781
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2178
timestamp 1704896540
transform 1 0 26928 0 1 61613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2179
timestamp 1704896540
transform 1 0 26928 0 1 61885
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2180
timestamp 1704896540
transform 1 0 26928 0 1 62293
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2181
timestamp 1704896540
transform 1 0 26928 0 1 62021
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2182
timestamp 1704896540
transform 1 0 27200 0 1 61477
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2183
timestamp 1704896540
transform 1 0 27200 0 1 61205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2184
timestamp 1704896540
transform 1 0 27200 0 1 62837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2185
timestamp 1704896540
transform 1 0 27200 0 1 63109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2186
timestamp 1704896540
transform 1 0 31552 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2187
timestamp 1704896540
transform 1 0 27608 0 1 68141
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2188
timestamp 1704896540
transform 1 0 26928 0 1 67733
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2189
timestamp 1704896540
transform 1 0 26928 0 1 68005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2190
timestamp 1704896540
transform 1 0 30328 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2191
timestamp 1704896540
transform 1 0 28288 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2192
timestamp 1704896540
transform 1 0 28288 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2193
timestamp 1704896540
transform 1 0 34136 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2194
timestamp 1704896540
transform 1 0 34136 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2195
timestamp 1704896540
transform 1 0 30872 0 1 68957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2196
timestamp 1704896540
transform 1 0 29240 0 1 68141
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2197
timestamp 1704896540
transform 1 0 33456 0 1 73037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2198
timestamp 1704896540
transform 1 0 32096 0 1 73717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2199
timestamp 1704896540
transform 1 0 32096 0 1 73037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2200
timestamp 1704896540
transform 1 0 31008 0 1 73717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2201
timestamp 1704896540
transform 1 0 31008 0 1 73037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2202
timestamp 1704896540
transform 1 0 30872 0 1 72765
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2203
timestamp 1704896540
transform 1 0 31144 0 1 73989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2204
timestamp 1704896540
transform 1 0 33456 0 1 73717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2205
timestamp 1704896540
transform 1 0 34680 0 1 73717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2206
timestamp 1704896540
transform 1 0 34680 0 1 73037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2207
timestamp 1704896540
transform 1 0 31144 0 1 72221
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2208
timestamp 1704896540
transform 1 0 34544 0 1 74125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2209
timestamp 1704896540
transform 1 0 35768 0 1 74125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2210
timestamp 1704896540
transform 1 0 33184 0 1 74125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2211
timestamp 1704896540
transform 1 0 31960 0 1 74125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2212
timestamp 1704896540
transform 1 0 30600 0 1 74125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2213
timestamp 1704896540
transform 1 0 29512 0 1 74125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2214
timestamp 1704896540
transform 1 0 28152 0 1 74125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2215
timestamp 1704896540
transform 1 0 28560 0 1 70453
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2216
timestamp 1704896540
transform 1 0 28560 0 1 72221
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2217
timestamp 1704896540
transform 1 0 27608 0 1 70317
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2218
timestamp 1704896540
transform 1 0 29784 0 1 73853
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2219
timestamp 1704896540
transform 1 0 28560 0 1 73717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2220
timestamp 1704896540
transform 1 0 28560 0 1 73037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2221
timestamp 1704896540
transform 1 0 29784 0 1 73717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2222
timestamp 1704896540
transform 1 0 29784 0 1 73037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2223
timestamp 1704896540
transform 1 0 28968 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2224
timestamp 1704896540
transform 1 0 28968 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2225
timestamp 1704896540
transform 1 0 29784 0 1 77661
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2226
timestamp 1704896540
transform 1 0 27472 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2227
timestamp 1704896540
transform 1 0 27472 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2228
timestamp 1704896540
transform 1 0 25704 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2229
timestamp 1704896540
transform 1 0 25704 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2230
timestamp 1704896540
transform 1 0 32504 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2231
timestamp 1704896540
transform 1 0 32504 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2232
timestamp 1704896540
transform 1 0 30872 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2233
timestamp 1704896540
transform 1 0 30872 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2234
timestamp 1704896540
transform 1 0 35496 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2235
timestamp 1704896540
transform 1 0 35496 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2236
timestamp 1704896540
transform 1 0 34136 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2237
timestamp 1704896540
transform 1 0 34136 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2238
timestamp 1704896540
transform 1 0 44744 0 1 73037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2239
timestamp 1704896540
transform 1 0 42024 0 1 73717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2240
timestamp 1704896540
transform 1 0 44336 0 1 74125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2241
timestamp 1704896540
transform 1 0 45560 0 1 74125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2242
timestamp 1704896540
transform 1 0 43384 0 1 73717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2243
timestamp 1704896540
transform 1 0 43384 0 1 73037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2244
timestamp 1704896540
transform 1 0 46920 0 1 74125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2245
timestamp 1704896540
transform 1 0 43248 0 1 74125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2246
timestamp 1704896540
transform 1 0 42296 0 1 73717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2247
timestamp 1704896540
transform 1 0 47192 0 1 73717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2248
timestamp 1704896540
transform 1 0 47192 0 1 73037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2249
timestamp 1704896540
transform 1 0 45968 0 1 73717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2250
timestamp 1704896540
transform 1 0 45968 0 1 73037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2251
timestamp 1704896540
transform 1 0 42296 0 1 73037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2252
timestamp 1704896540
transform 1 0 42024 0 1 73037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2253
timestamp 1704896540
transform 1 0 44744 0 1 73717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2254
timestamp 1704896540
transform 1 0 39712 0 1 73717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2255
timestamp 1704896540
transform 1 0 39712 0 1 73037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2256
timestamp 1704896540
transform 1 0 41888 0 1 74125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2257
timestamp 1704896540
transform 1 0 37264 0 1 73717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2258
timestamp 1704896540
transform 1 0 40664 0 1 74125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2259
timestamp 1704896540
transform 1 0 39304 0 1 74125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2260
timestamp 1704896540
transform 1 0 38488 0 1 73717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2261
timestamp 1704896540
transform 1 0 40800 0 1 73717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2262
timestamp 1704896540
transform 1 0 38216 0 1 74125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2263
timestamp 1704896540
transform 1 0 36856 0 1 74125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2264
timestamp 1704896540
transform 1 0 40800 0 1 73037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2265
timestamp 1704896540
transform 1 0 38488 0 1 73037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2266
timestamp 1704896540
transform 1 0 37264 0 1 73037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2267
timestamp 1704896540
transform 1 0 37400 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2268
timestamp 1704896540
transform 1 0 40528 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2269
timestamp 1704896540
transform 1 0 40528 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2270
timestamp 1704896540
transform 1 0 39168 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2271
timestamp 1704896540
transform 1 0 39168 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2272
timestamp 1704896540
transform 1 0 37400 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2273
timestamp 1704896540
transform 1 0 47464 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2274
timestamp 1704896540
transform 1 0 47464 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2275
timestamp 1704896540
transform 1 0 45832 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2276
timestamp 1704896540
transform 1 0 45832 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2277
timestamp 1704896540
transform 1 0 44200 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2278
timestamp 1704896540
transform 1 0 44200 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2279
timestamp 1704896540
transform 1 0 42432 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2280
timestamp 1704896540
transform 1 0 42432 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2281
timestamp 1704896540
transform 1 0 36040 0 1 73717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2282
timestamp 1704896540
transform 1 0 36040 0 1 73037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2283
timestamp 1704896540
transform 1 0 21624 0 1 59437
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2284
timestamp 1704896540
transform 1 0 20536 0 1 59437
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2285
timestamp 1704896540
transform 1 0 22032 0 1 59437
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2286
timestamp 1704896540
transform 1 0 21488 0 1 59437
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2287
timestamp 1704896540
transform 1 0 21080 0 1 59437
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2288
timestamp 1704896540
transform 1 0 20808 0 1 59437
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2289
timestamp 1704896540
transform 1 0 94656 0 1 47469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2290
timestamp 1704896540
transform 1 0 94656 0 1 42301
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2291
timestamp 1704896540
transform 1 0 94656 0 1 40669
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2292
timestamp 1704896540
transform 1 0 94656 0 1 49101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2293
timestamp 1704896540
transform 1 0 94656 0 1 43933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2294
timestamp 1704896540
transform 1 0 94656 0 1 45837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2295
timestamp 1704896540
transform 1 0 73848 0 1 40533
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2296
timestamp 1704896540
transform 1 0 74664 0 1 42845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2297
timestamp 1704896540
transform 1 0 74664 0 1 43117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2298
timestamp 1704896540
transform 1 0 73848 0 1 42301
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2299
timestamp 1704896540
transform 1 0 73848 0 1 40397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2300
timestamp 1704896540
transform 1 0 73848 0 1 41893
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2301
timestamp 1704896540
transform 1 0 73848 0 1 41621
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2302
timestamp 1704896540
transform 1 0 73848 0 1 40125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2303
timestamp 1704896540
transform 1 0 73848 0 1 44477
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2304
timestamp 1704896540
transform 1 0 74256 0 1 39989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2305
timestamp 1704896540
transform 1 0 74256 0 1 42437
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2306
timestamp 1704896540
transform 1 0 74256 0 1 42709
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2307
timestamp 1704896540
transform 1 0 74392 0 1 44341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2308
timestamp 1704896540
transform 1 0 74392 0 1 44069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2309
timestamp 1704896540
transform 1 0 74392 0 1 43661
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2310
timestamp 1704896540
transform 1 0 74392 0 1 43933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2311
timestamp 1704896540
transform 1 0 74256 0 1 40805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2312
timestamp 1704896540
transform 1 0 74256 0 1 40533
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2313
timestamp 1704896540
transform 1 0 74256 0 1 40125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2314
timestamp 1704896540
transform 1 0 74256 0 1 40397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2315
timestamp 1704896540
transform 1 0 74936 0 1 42437
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2316
timestamp 1704896540
transform 1 0 73984 0 1 44341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2317
timestamp 1704896540
transform 1 0 74256 0 1 44477
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2318
timestamp 1704896540
transform 1 0 75072 0 1 42301
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2319
timestamp 1704896540
transform 1 0 74800 0 1 42301
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2320
timestamp 1704896540
transform 1 0 73304 0 1 42709
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2321
timestamp 1704896540
transform 1 0 74256 0 1 42301
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2322
timestamp 1704896540
transform 1 0 74256 0 1 42029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2323
timestamp 1704896540
transform 1 0 73304 0 1 42437
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2324
timestamp 1704896540
transform 1 0 75208 0 1 40125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2325
timestamp 1704896540
transform 1 0 75480 0 1 39989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2326
timestamp 1704896540
transform 1 0 74936 0 1 42709
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2327
timestamp 1704896540
transform 1 0 74664 0 1 44069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2328
timestamp 1704896540
transform 1 0 74664 0 1 39989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2329
timestamp 1704896540
transform 1 0 75208 0 1 40397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2330
timestamp 1704896540
transform 1 0 73984 0 1 43117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2331
timestamp 1704896540
transform 1 0 75208 0 1 40941
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2332
timestamp 1704896540
transform 1 0 74664 0 1 44341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2333
timestamp 1704896540
transform 1 0 74256 0 1 43525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2334
timestamp 1704896540
transform 1 0 75616 0 1 41621
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2335
timestamp 1704896540
transform 1 0 75616 0 1 41349
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2336
timestamp 1704896540
transform 1 0 75616 0 1 40941
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2337
timestamp 1704896540
transform 1 0 75616 0 1 41213
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2338
timestamp 1704896540
transform 1 0 75480 0 1 44069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2339
timestamp 1704896540
transform 1 0 75480 0 1 44341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2340
timestamp 1704896540
transform 1 0 75208 0 1 41213
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2341
timestamp 1704896540
transform 1 0 75616 0 1 44477
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2342
timestamp 1704896540
transform 1 0 74256 0 1 43253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2343
timestamp 1704896540
transform 1 0 74256 0 1 42845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2344
timestamp 1704896540
transform 1 0 74256 0 1 43117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2345
timestamp 1704896540
transform 1 0 73848 0 1 40805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2346
timestamp 1704896540
transform 1 0 73984 0 1 39989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2347
timestamp 1704896540
transform 1 0 75072 0 1 43117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2348
timestamp 1704896540
transform 1 0 75616 0 1 43933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2349
timestamp 1704896540
transform 1 0 75616 0 1 43661
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2350
timestamp 1704896540
transform 1 0 75616 0 1 43253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2351
timestamp 1704896540
transform 1 0 75616 0 1 43525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2352
timestamp 1704896540
transform 1 0 75616 0 1 40805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2353
timestamp 1704896540
transform 1 0 75616 0 1 40533
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2354
timestamp 1704896540
transform 1 0 75616 0 1 40125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2355
timestamp 1704896540
transform 1 0 75616 0 1 40397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2356
timestamp 1704896540
transform 1 0 75072 0 1 42845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2357
timestamp 1704896540
transform 1 0 73984 0 1 43525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2358
timestamp 1704896540
transform 1 0 74936 0 1 44477
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2359
timestamp 1704896540
transform 1 0 74936 0 1 41893
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2360
timestamp 1704896540
transform 1 0 74800 0 1 43933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2361
timestamp 1704896540
transform 1 0 74800 0 1 43661
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2362
timestamp 1704896540
transform 1 0 74256 0 1 41893
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2363
timestamp 1704896540
transform 1 0 74256 0 1 41621
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2364
timestamp 1704896540
transform 1 0 73984 0 1 44069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2365
timestamp 1704896540
transform 1 0 73984 0 1 43661
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2366
timestamp 1704896540
transform 1 0 74936 0 1 41621
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2367
timestamp 1704896540
transform 1 0 75208 0 1 39989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2368
timestamp 1704896540
transform 1 0 73984 0 1 43253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2369
timestamp 1704896540
transform 1 0 73984 0 1 42845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2370
timestamp 1704896540
transform 1 0 75480 0 1 42845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2371
timestamp 1704896540
transform 1 0 75480 0 1 43117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2372
timestamp 1704896540
transform 1 0 73984 0 1 43933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2373
timestamp 1704896540
transform 1 0 73848 0 1 42709
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2374
timestamp 1704896540
transform 1 0 73848 0 1 42437
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2375
timestamp 1704896540
transform 1 0 73848 0 1 42029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2376
timestamp 1704896540
transform 1 0 74664 0 1 43525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2377
timestamp 1704896540
transform 1 0 74664 0 1 43253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2378
timestamp 1704896540
transform 1 0 74256 0 1 47061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2379
timestamp 1704896540
transform 1 0 74664 0 1 46653
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2380
timestamp 1704896540
transform 1 0 73984 0 1 48693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2381
timestamp 1704896540
transform 1 0 73984 0 1 48421
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2382
timestamp 1704896540
transform 1 0 74664 0 1 46381
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2383
timestamp 1704896540
transform 1 0 74800 0 1 48285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2384
timestamp 1704896540
transform 1 0 74800 0 1 48013
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2385
timestamp 1704896540
transform 1 0 74664 0 1 47197
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2386
timestamp 1704896540
transform 1 0 74664 0 1 47469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2387
timestamp 1704896540
transform 1 0 73848 0 1 48285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2388
timestamp 1704896540
transform 1 0 75616 0 1 49509
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2389
timestamp 1704896540
transform 1 0 75616 0 1 49237
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2390
timestamp 1704896540
transform 1 0 75616 0 1 49101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2391
timestamp 1704896540
transform 1 0 75616 0 1 48829
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2392
timestamp 1704896540
transform 1 0 75480 0 1 48693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2393
timestamp 1704896540
transform 1 0 75480 0 1 48421
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2394
timestamp 1704896540
transform 1 0 75616 0 1 47605
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2395
timestamp 1704896540
transform 1 0 75616 0 1 47877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2396
timestamp 1704896540
transform 1 0 75616 0 1 48285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2397
timestamp 1704896540
transform 1 0 75616 0 1 48013
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2398
timestamp 1704896540
transform 1 0 73848 0 1 48013
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2399
timestamp 1704896540
transform 1 0 73984 0 1 47197
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2400
timestamp 1704896540
transform 1 0 73984 0 1 47469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2401
timestamp 1704896540
transform 1 0 73984 0 1 47877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2402
timestamp 1704896540
transform 1 0 75480 0 1 47469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2403
timestamp 1704896540
transform 1 0 75480 0 1 47197
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2404
timestamp 1704896540
transform 1 0 75616 0 1 46789
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2405
timestamp 1704896540
transform 1 0 75616 0 1 47061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2406
timestamp 1704896540
transform 1 0 74936 0 1 44749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2407
timestamp 1704896540
transform 1 0 73984 0 1 47605
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2408
timestamp 1704896540
transform 1 0 73848 0 1 47061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2409
timestamp 1704896540
transform 1 0 73848 0 1 46789
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2410
timestamp 1704896540
transform 1 0 75208 0 1 48829
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2411
timestamp 1704896540
transform 1 0 75208 0 1 49101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2412
timestamp 1704896540
transform 1 0 75072 0 1 44885
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2413
timestamp 1704896540
transform 1 0 75072 0 1 45157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2414
timestamp 1704896540
transform 1 0 74392 0 1 47605
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2415
timestamp 1704896540
transform 1 0 74392 0 1 47877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2416
timestamp 1704896540
transform 1 0 75616 0 1 44749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2417
timestamp 1704896540
transform 1 0 74936 0 1 45565
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2418
timestamp 1704896540
transform 1 0 75480 0 1 44885
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2419
timestamp 1704896540
transform 1 0 75480 0 1 45157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2420
timestamp 1704896540
transform 1 0 75480 0 1 45565
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2421
timestamp 1704896540
transform 1 0 75480 0 1 45293
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2422
timestamp 1704896540
transform 1 0 75072 0 1 49509
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2423
timestamp 1704896540
transform 1 0 74256 0 1 46653
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2424
timestamp 1704896540
transform 1 0 74256 0 1 46381
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2425
timestamp 1704896540
transform 1 0 73984 0 1 45973
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2426
timestamp 1704896540
transform 1 0 74256 0 1 45973
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2427
timestamp 1704896540
transform 1 0 74256 0 1 46245
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2428
timestamp 1704896540
transform 1 0 74936 0 1 45837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2429
timestamp 1704896540
transform 1 0 74800 0 1 45565
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2430
timestamp 1704896540
transform 1 0 73984 0 1 46245
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2431
timestamp 1704896540
transform 1 0 73984 0 1 46653
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2432
timestamp 1704896540
transform 1 0 74800 0 1 45837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2433
timestamp 1704896540
transform 1 0 73848 0 1 44749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2434
timestamp 1704896540
transform 1 0 73984 0 1 46381
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2435
timestamp 1704896540
transform 1 0 74392 0 1 48693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2436
timestamp 1704896540
transform 1 0 74392 0 1 48421
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2437
timestamp 1704896540
transform 1 0 74392 0 1 48013
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2438
timestamp 1704896540
transform 1 0 74528 0 1 45021
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2439
timestamp 1704896540
transform 1 0 74528 0 1 45429
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2440
timestamp 1704896540
transform 1 0 74392 0 1 48285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2441
timestamp 1704896540
transform 1 0 74256 0 1 44749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2442
timestamp 1704896540
transform 1 0 75072 0 1 47877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2443
timestamp 1704896540
transform 1 0 75072 0 1 47605
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2444
timestamp 1704896540
transform 1 0 74936 0 1 47061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2445
timestamp 1704896540
transform 1 0 74936 0 1 46789
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2446
timestamp 1704896540
transform 1 0 74800 0 1 47061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2447
timestamp 1704896540
transform 1 0 74800 0 1 46789
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2448
timestamp 1704896540
transform 1 0 74392 0 1 47469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2449
timestamp 1704896540
transform 1 0 74392 0 1 47197
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2450
timestamp 1704896540
transform 1 0 74256 0 1 46789
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2451
timestamp 1704896540
transform 1 0 73848 0 1 51005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2452
timestamp 1704896540
transform 1 0 74800 0 1 51413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2453
timestamp 1704896540
transform 1 0 73848 0 1 52637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2454
timestamp 1704896540
transform 1 0 74800 0 1 51141
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2455
timestamp 1704896540
transform 1 0 73848 0 1 52365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2456
timestamp 1704896540
transform 1 0 74936 0 1 53181
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2457
timestamp 1704896540
transform 1 0 74936 0 1 53453
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2458
timestamp 1704896540
transform 1 0 74800 0 1 50597
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2459
timestamp 1704896540
transform 1 0 75208 0 1 50733
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2460
timestamp 1704896540
transform 1 0 73848 0 1 54269
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2461
timestamp 1704896540
transform 1 0 74392 0 1 51821
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2462
timestamp 1704896540
transform 1 0 74392 0 1 51549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2463
timestamp 1704896540
transform 1 0 74392 0 1 52365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2464
timestamp 1704896540
transform 1 0 74392 0 1 52637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2465
timestamp 1704896540
transform 1 0 75208 0 1 51005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2466
timestamp 1704896540
transform 1 0 75072 0 1 49781
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2467
timestamp 1704896540
transform 1 0 75480 0 1 52365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2468
timestamp 1704896540
transform 1 0 75480 0 1 52637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2469
timestamp 1704896540
transform 1 0 74800 0 1 50325
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2470
timestamp 1704896540
transform 1 0 74664 0 1 53861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2471
timestamp 1704896540
transform 1 0 75208 0 1 54269
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2472
timestamp 1704896540
transform 1 0 73848 0 1 50733
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2473
timestamp 1704896540
transform 1 0 74664 0 1 53589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2474
timestamp 1704896540
transform 1 0 73984 0 1 53045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2475
timestamp 1704896540
transform 1 0 73984 0 1 52773
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2476
timestamp 1704896540
transform 1 0 75480 0 1 52229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2477
timestamp 1704896540
transform 1 0 75480 0 1 51957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2478
timestamp 1704896540
transform 1 0 74800 0 1 52637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2479
timestamp 1704896540
transform 1 0 75616 0 1 50733
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2480
timestamp 1704896540
transform 1 0 75616 0 1 51005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2481
timestamp 1704896540
transform 1 0 74392 0 1 50733
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2482
timestamp 1704896540
transform 1 0 74392 0 1 51005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2483
timestamp 1704896540
transform 1 0 74392 0 1 51413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2484
timestamp 1704896540
transform 1 0 74392 0 1 51141
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2485
timestamp 1704896540
transform 1 0 75480 0 1 54269
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2486
timestamp 1704896540
transform 1 0 75480 0 1 53997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2487
timestamp 1704896540
transform 1 0 75480 0 1 53589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2488
timestamp 1704896540
transform 1 0 75480 0 1 53861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2489
timestamp 1704896540
transform 1 0 74800 0 1 52365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2490
timestamp 1704896540
transform 1 0 74664 0 1 52773
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2491
timestamp 1704896540
transform 1 0 75072 0 1 53589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2492
timestamp 1704896540
transform 1 0 75072 0 1 53861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2493
timestamp 1704896540
transform 1 0 73848 0 1 51141
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2494
timestamp 1704896540
transform 1 0 74256 0 1 52773
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2495
timestamp 1704896540
transform 1 0 74256 0 1 53045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2496
timestamp 1704896540
transform 1 0 74936 0 1 51549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2497
timestamp 1704896540
transform 1 0 75616 0 1 50053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2498
timestamp 1704896540
transform 1 0 75616 0 1 50325
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2499
timestamp 1704896540
transform 1 0 74936 0 1 51821
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2500
timestamp 1704896540
transform 1 0 75480 0 1 52773
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2501
timestamp 1704896540
transform 1 0 75480 0 1 53045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2502
timestamp 1704896540
transform 1 0 75616 0 1 53453
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2503
timestamp 1704896540
transform 1 0 75616 0 1 53181
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2504
timestamp 1704896540
transform 1 0 75480 0 1 51821
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2505
timestamp 1704896540
transform 1 0 75480 0 1 51549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2506
timestamp 1704896540
transform 1 0 73984 0 1 51549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2507
timestamp 1704896540
transform 1 0 73984 0 1 51821
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2508
timestamp 1704896540
transform 1 0 73984 0 1 52229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2509
timestamp 1704896540
transform 1 0 73984 0 1 51957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2510
timestamp 1704896540
transform 1 0 74256 0 1 54269
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2511
timestamp 1704896540
transform 1 0 74664 0 1 52229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2512
timestamp 1704896540
transform 1 0 74664 0 1 53045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2513
timestamp 1704896540
transform 1 0 74664 0 1 51957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2514
timestamp 1704896540
transform 1 0 74256 0 1 52229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2515
timestamp 1704896540
transform 1 0 74256 0 1 51957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2516
timestamp 1704896540
transform 1 0 73848 0 1 50597
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2517
timestamp 1704896540
transform 1 0 74256 0 1 49917
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2518
timestamp 1704896540
transform 1 0 74256 0 1 50189
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2519
timestamp 1704896540
transform 1 0 73848 0 1 50325
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2520
timestamp 1704896540
transform 1 0 73848 0 1 49917
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2521
timestamp 1704896540
transform 1 0 73848 0 1 50189
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2522
timestamp 1704896540
transform 1 0 75072 0 1 50325
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2523
timestamp 1704896540
transform 1 0 75072 0 1 50597
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2524
timestamp 1704896540
transform 1 0 73848 0 1 51413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2525
timestamp 1704896540
transform 1 0 74256 0 1 50325
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2526
timestamp 1704896540
transform 1 0 74256 0 1 50597
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2527
timestamp 1704896540
transform 1 0 73848 0 1 54949
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2528
timestamp 1704896540
transform 1 0 73848 0 1 54677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2529
timestamp 1704896540
transform 1 0 73984 0 1 55901
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2530
timestamp 1704896540
transform 1 0 73848 0 1 58621
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2531
timestamp 1704896540
transform 1 0 73848 0 1 58893
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2532
timestamp 1704896540
transform 1 0 73848 0 1 59301
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2533
timestamp 1704896540
transform 1 0 75616 0 1 56309
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2534
timestamp 1704896540
transform 1 0 75616 0 1 56581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2535
timestamp 1704896540
transform 1 0 73848 0 1 59029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2536
timestamp 1704896540
transform 1 0 75480 0 1 56173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2537
timestamp 1704896540
transform 1 0 75480 0 1 55901
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2538
timestamp 1704896540
transform 1 0 74664 0 1 55901
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2539
timestamp 1704896540
transform 1 0 74664 0 1 56173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2540
timestamp 1704896540
transform 1 0 75072 0 1 59029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2541
timestamp 1704896540
transform 1 0 75616 0 1 57533
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2542
timestamp 1704896540
transform 1 0 75616 0 1 57805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2543
timestamp 1704896540
transform 1 0 75616 0 1 58213
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2544
timestamp 1704896540
transform 1 0 75616 0 1 57941
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2545
timestamp 1704896540
transform 1 0 75616 0 1 55765
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2546
timestamp 1704896540
transform 1 0 75616 0 1 55493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2547
timestamp 1704896540
transform 1 0 73848 0 1 56309
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2548
timestamp 1704896540
transform 1 0 73848 0 1 56581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2549
timestamp 1704896540
transform 1 0 73848 0 1 56989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2550
timestamp 1704896540
transform 1 0 73848 0 1 56717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2551
timestamp 1704896540
transform 1 0 75616 0 1 54949
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2552
timestamp 1704896540
transform 1 0 75616 0 1 54677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2553
timestamp 1704896540
transform 1 0 75072 0 1 59301
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2554
timestamp 1704896540
transform 1 0 75480 0 1 56717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2555
timestamp 1704896540
transform 1 0 75480 0 1 56989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2556
timestamp 1704896540
transform 1 0 75480 0 1 57397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2557
timestamp 1704896540
transform 1 0 75480 0 1 57125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2558
timestamp 1704896540
transform 1 0 75208 0 1 57533
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2559
timestamp 1704896540
transform 1 0 75208 0 1 57805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2560
timestamp 1704896540
transform 1 0 75208 0 1 56309
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2561
timestamp 1704896540
transform 1 0 74392 0 1 58485
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2562
timestamp 1704896540
transform 1 0 74392 0 1 58213
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2563
timestamp 1704896540
transform 1 0 74256 0 1 58621
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2564
timestamp 1704896540
transform 1 0 74256 0 1 58893
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2565
timestamp 1704896540
transform 1 0 75208 0 1 56581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2566
timestamp 1704896540
transform 1 0 74392 0 1 55085
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2567
timestamp 1704896540
transform 1 0 74392 0 1 55357
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2568
timestamp 1704896540
transform 1 0 75072 0 1 56173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2569
timestamp 1704896540
transform 1 0 74256 0 1 54949
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2570
timestamp 1704896540
transform 1 0 74256 0 1 54677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2571
timestamp 1704896540
transform 1 0 73984 0 1 55357
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2572
timestamp 1704896540
transform 1 0 74392 0 1 56173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2573
timestamp 1704896540
transform 1 0 74392 0 1 55901
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2574
timestamp 1704896540
transform 1 0 74256 0 1 55493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2575
timestamp 1704896540
transform 1 0 74256 0 1 55765
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2576
timestamp 1704896540
transform 1 0 75072 0 1 55901
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2577
timestamp 1704896540
transform 1 0 73984 0 1 55085
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2578
timestamp 1704896540
transform 1 0 75208 0 1 55085
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2579
timestamp 1704896540
transform 1 0 75208 0 1 55357
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2580
timestamp 1704896540
transform 1 0 74392 0 1 56309
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2581
timestamp 1704896540
transform 1 0 74392 0 1 56581
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2582
timestamp 1704896540
transform 1 0 74256 0 1 56989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2583
timestamp 1704896540
transform 1 0 74256 0 1 56717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2584
timestamp 1704896540
transform 1 0 74664 0 1 58485
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2585
timestamp 1704896540
transform 1 0 74392 0 1 59029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2586
timestamp 1704896540
transform 1 0 74392 0 1 59301
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2587
timestamp 1704896540
transform 1 0 74664 0 1 58213
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2588
timestamp 1704896540
transform 1 0 74936 0 1 56989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2589
timestamp 1704896540
transform 1 0 74936 0 1 56717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2590
timestamp 1704896540
transform 1 0 74800 0 1 56989
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2591
timestamp 1704896540
transform 1 0 74800 0 1 56717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2592
timestamp 1704896540
transform 1 0 74936 0 1 58077
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2593
timestamp 1704896540
transform 1 0 74936 0 1 57805
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2594
timestamp 1704896540
transform 1 0 73984 0 1 58485
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2595
timestamp 1704896540
transform 1 0 73984 0 1 58213
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2596
timestamp 1704896540
transform 1 0 74664 0 1 54677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2597
timestamp 1704896540
transform 1 0 74664 0 1 54949
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2598
timestamp 1704896540
transform 1 0 73848 0 1 55493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2599
timestamp 1704896540
transform 1 0 73848 0 1 55765
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2600
timestamp 1704896540
transform 1 0 73984 0 1 56173
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2601
timestamp 1704896540
transform 1 0 73848 0 1 54541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2602
timestamp 1704896540
transform 1 0 74256 0 1 54541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2603
timestamp 1704896540
transform 1 0 75208 0 1 54541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2604
timestamp 1704896540
transform 1 0 94656 0 1 53997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2605
timestamp 1704896540
transform 1 0 94656 0 1 50597
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2606
timestamp 1704896540
transform 1 0 94656 0 1 52365
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2607
timestamp 1704896540
transform 1 0 91936 0 1 58757
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2608
timestamp 1704896540
transform 1 0 93419 0 1 59362
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2609
timestamp 1704896540
transform 1 0 94656 0 1 59029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2610
timestamp 1704896540
transform 1 0 94656 0 1 57397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2611
timestamp 1704896540
transform 1 0 94656 0 1 55901
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2612
timestamp 1704896540
transform 1 0 68952 0 1 40669
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2613
timestamp 1704896540
transform 1 0 68952 0 1 40941
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2614
timestamp 1704896540
transform 1 0 69088 0 1 42573
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2615
timestamp 1704896540
transform 1 0 69088 0 1 42301
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2616
timestamp 1704896540
transform 1 0 69088 0 1 44069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2617
timestamp 1704896540
transform 1 0 69088 0 1 43797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2618
timestamp 1704896540
transform 1 0 69088 0 1 52773
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2619
timestamp 1704896540
transform 1 0 69088 0 1 52501
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2620
timestamp 1704896540
transform 1 0 69088 0 1 44885
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2621
timestamp 1704896540
transform 1 0 69088 0 1 44613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2622
timestamp 1704896540
transform 1 0 69088 0 1 49917
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2623
timestamp 1704896540
transform 1 0 69088 0 1 49645
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2624
timestamp 1704896540
transform 1 0 69088 0 1 41077
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2625
timestamp 1704896540
transform 1 0 69088 0 1 41349
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2626
timestamp 1704896540
transform 1 0 68952 0 1 45973
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2627
timestamp 1704896540
transform 1 0 68952 0 1 45701
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2628
timestamp 1704896540
transform 1 0 68952 0 1 46245
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2629
timestamp 1704896540
transform 1 0 68952 0 1 46517
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2630
timestamp 1704896540
transform 1 0 69088 0 1 57941
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2631
timestamp 1704896540
transform 1 0 69088 0 1 57669
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2632
timestamp 1704896540
transform 1 0 69088 0 1 48557
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2633
timestamp 1704896540
transform 1 0 69088 0 1 48829
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2634
timestamp 1704896540
transform 1 0 69088 0 1 39853
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2635
timestamp 1704896540
transform 1 0 69088 0 1 40125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2636
timestamp 1704896540
transform 1 0 68952 0 1 45021
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2637
timestamp 1704896540
transform 1 0 68952 0 1 45293
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2638
timestamp 1704896540
transform 1 0 68952 0 1 53997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2639
timestamp 1704896540
transform 1 0 68952 0 1 53725
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2640
timestamp 1704896540
transform 1 0 68952 0 1 49373
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2641
timestamp 1704896540
transform 1 0 68952 0 1 49645
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2642
timestamp 1704896540
transform 1 0 68952 0 1 58077
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2643
timestamp 1704896540
transform 1 0 68952 0 1 58349
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2644
timestamp 1704896540
transform 1 0 69088 0 1 53589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2645
timestamp 1704896540
transform 1 0 69088 0 1 53317
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2646
timestamp 1704896540
transform 1 0 69088 0 1 45429
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2647
timestamp 1704896540
transform 1 0 69088 0 1 45701
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2648
timestamp 1704896540
transform 1 0 62696 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2649
timestamp 1704896540
transform 1 0 62696 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2650
timestamp 1704896540
transform 1 0 65280 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2651
timestamp 1704896540
transform 1 0 65280 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2652
timestamp 1704896540
transform 1 0 60792 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2653
timestamp 1704896540
transform 1 0 60792 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2654
timestamp 1704896540
transform 1 0 70312 0 1 68005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2655
timestamp 1704896540
transform 1 0 70312 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2656
timestamp 1704896540
transform 1 0 68272 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2657
timestamp 1704896540
transform 1 0 68272 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2658
timestamp 1704896540
transform 1 0 69360 0 1 68005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2659
timestamp 1704896540
transform 1 0 69360 0 1 67733
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2660
timestamp 1704896540
transform 1 0 68952 0 1 61885
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2661
timestamp 1704896540
transform 1 0 68952 0 1 61613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2662
timestamp 1704896540
transform 1 0 69088 0 1 67053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2663
timestamp 1704896540
transform 1 0 69088 0 1 66781
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2664
timestamp 1704896540
transform 1 0 68952 0 1 66237
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2665
timestamp 1704896540
transform 1 0 68952 0 1 65965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2666
timestamp 1704896540
transform 1 0 68952 0 1 65557
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2667
timestamp 1704896540
transform 1 0 68952 0 1 65829
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2668
timestamp 1704896540
transform 1 0 69088 0 1 66509
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2669
timestamp 1704896540
transform 1 0 69088 0 1 66237
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2670
timestamp 1704896540
transform 1 0 68952 0 1 67733
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2671
timestamp 1704896540
transform 1 0 67728 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2672
timestamp 1704896540
transform 1 0 67728 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2673
timestamp 1704896540
transform 1 0 60248 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2674
timestamp 1704896540
transform 1 0 60248 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2675
timestamp 1704896540
transform 1 0 64056 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2676
timestamp 1704896540
transform 1 0 64056 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2677
timestamp 1704896540
transform 1 0 67048 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2678
timestamp 1704896540
transform 1 0 67048 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2679
timestamp 1704896540
transform 1 0 66504 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2680
timestamp 1704896540
transform 1 0 66504 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2681
timestamp 1704896540
transform 1 0 61472 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2682
timestamp 1704896540
transform 1 0 61472 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2683
timestamp 1704896540
transform 1 0 50592 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2684
timestamp 1704896540
transform 1 0 50592 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2685
timestamp 1704896540
transform 1 0 55760 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2686
timestamp 1704896540
transform 1 0 55760 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2687
timestamp 1704896540
transform 1 0 55216 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2688
timestamp 1704896540
transform 1 0 55216 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2689
timestamp 1704896540
transform 1 0 48960 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2690
timestamp 1704896540
transform 1 0 48960 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2691
timestamp 1704896540
transform 1 0 59568 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2692
timestamp 1704896540
transform 1 0 59568 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2693
timestamp 1704896540
transform 1 0 52088 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2694
timestamp 1704896540
transform 1 0 52088 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2695
timestamp 1704896540
transform 1 0 59024 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2696
timestamp 1704896540
transform 1 0 59024 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2697
timestamp 1704896540
transform 1 0 53992 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2698
timestamp 1704896540
transform 1 0 53992 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2699
timestamp 1704896540
transform 1 0 57936 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2700
timestamp 1704896540
transform 1 0 57936 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2701
timestamp 1704896540
transform 1 0 57800 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2702
timestamp 1704896540
transform 1 0 57800 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2703
timestamp 1704896540
transform 1 0 51544 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2704
timestamp 1704896540
transform 1 0 51544 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2705
timestamp 1704896540
transform 1 0 53040 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2706
timestamp 1704896540
transform 1 0 53040 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2707
timestamp 1704896540
transform 1 0 56848 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2708
timestamp 1704896540
transform 1 0 56848 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2709
timestamp 1704896540
transform 1 0 52768 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2710
timestamp 1704896540
transform 1 0 52768 0 1 68277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2711
timestamp 1704896540
transform 1 0 59704 0 1 73037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2712
timestamp 1704896540
transform 1 0 58480 0 1 73717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2713
timestamp 1704896540
transform 1 0 58480 0 1 73037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2714
timestamp 1704896540
transform 1 0 57256 0 1 73717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2715
timestamp 1704896540
transform 1 0 57256 0 1 73037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2716
timestamp 1704896540
transform 1 0 59296 0 1 74125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2717
timestamp 1704896540
transform 1 0 58208 0 1 74125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2718
timestamp 1704896540
transform 1 0 56848 0 1 74125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2719
timestamp 1704896540
transform 1 0 55624 0 1 74125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2720
timestamp 1704896540
transform 1 0 54264 0 1 74125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2721
timestamp 1704896540
transform 1 0 56032 0 1 73717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2722
timestamp 1704896540
transform 1 0 56032 0 1 73037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2723
timestamp 1704896540
transform 1 0 54672 0 1 73717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2724
timestamp 1704896540
transform 1 0 54672 0 1 73037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2725
timestamp 1704896540
transform 1 0 59704 0 1 73717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2726
timestamp 1704896540
transform 1 0 51000 0 1 73717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2727
timestamp 1704896540
transform 1 0 51000 0 1 73037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2728
timestamp 1704896540
transform 1 0 52088 0 1 73717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2729
timestamp 1704896540
transform 1 0 49776 0 1 73717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2730
timestamp 1704896540
transform 1 0 53040 0 1 74125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2731
timestamp 1704896540
transform 1 0 51952 0 1 74125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2732
timestamp 1704896540
transform 1 0 50592 0 1 74125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2733
timestamp 1704896540
transform 1 0 49504 0 1 74125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2734
timestamp 1704896540
transform 1 0 48144 0 1 74125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2735
timestamp 1704896540
transform 1 0 49776 0 1 73037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2736
timestamp 1704896540
transform 1 0 48552 0 1 73717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2737
timestamp 1704896540
transform 1 0 48552 0 1 73037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2738
timestamp 1704896540
transform 1 0 52088 0 1 73037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2739
timestamp 1704896540
transform 1 0 53448 0 1 73717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2740
timestamp 1704896540
transform 1 0 53448 0 1 73037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2741
timestamp 1704896540
transform 1 0 50728 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2742
timestamp 1704896540
transform 1 0 50728 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2743
timestamp 1704896540
transform 1 0 49232 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2744
timestamp 1704896540
transform 1 0 49232 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2745
timestamp 1704896540
transform 1 0 52632 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2746
timestamp 1704896540
transform 1 0 52632 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2747
timestamp 1704896540
transform 1 0 59160 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2748
timestamp 1704896540
transform 1 0 59160 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2749
timestamp 1704896540
transform 1 0 57664 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2750
timestamp 1704896540
transform 1 0 57664 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2751
timestamp 1704896540
transform 1 0 54128 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2752
timestamp 1704896540
transform 1 0 54128 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2753
timestamp 1704896540
transform 1 0 55896 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2754
timestamp 1704896540
transform 1 0 55896 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2755
timestamp 1704896540
transform 1 0 65960 0 1 73717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2756
timestamp 1704896540
transform 1 0 67184 0 1 73717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2757
timestamp 1704896540
transform 1 0 67184 0 1 73037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2758
timestamp 1704896540
transform 1 0 66912 0 1 74125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2759
timestamp 1704896540
transform 1 0 65960 0 1 73037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2760
timestamp 1704896540
transform 1 0 68952 0 1 70317
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2761
timestamp 1704896540
transform 1 0 65552 0 1 74125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2762
timestamp 1704896540
transform 1 0 64328 0 1 74125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2763
timestamp 1704896540
transform 1 0 63240 0 1 74125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2764
timestamp 1704896540
transform 1 0 61880 0 1 74125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2765
timestamp 1704896540
transform 1 0 60656 0 1 74125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2766
timestamp 1704896540
transform 1 0 63512 0 1 73717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2767
timestamp 1704896540
transform 1 0 63512 0 1 73037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2768
timestamp 1704896540
transform 1 0 60792 0 1 73717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2769
timestamp 1704896540
transform 1 0 60792 0 1 73037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2770
timestamp 1704896540
transform 1 0 64736 0 1 73717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2771
timestamp 1704896540
transform 1 0 64736 0 1 73037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2772
timestamp 1704896540
transform 1 0 62152 0 1 73717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2773
timestamp 1704896540
transform 1 0 62152 0 1 73037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2774
timestamp 1704896540
transform 1 0 64056 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2775
timestamp 1704896540
transform 1 0 64056 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2776
timestamp 1704896540
transform 1 0 62696 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2777
timestamp 1704896540
transform 1 0 62696 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2778
timestamp 1704896540
transform 1 0 60928 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2779
timestamp 1704896540
transform 1 0 60928 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2780
timestamp 1704896540
transform 1 0 71128 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2781
timestamp 1704896540
transform 1 0 71128 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2782
timestamp 1704896540
transform 1 0 69224 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2783
timestamp 1704896540
transform 1 0 69224 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2784
timestamp 1704896540
transform 1 0 67728 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2785
timestamp 1704896540
transform 1 0 67728 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2786
timestamp 1704896540
transform 1 0 65960 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2787
timestamp 1704896540
transform 1 0 65960 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2788
timestamp 1704896540
transform 1 0 95336 0 1 61613
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2789
timestamp 1704896540
transform 1 0 91936 0 1 61477
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2790
timestamp 1704896540
transform 1 0 94656 0 1 60797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2791
timestamp 1704896540
transform 1 0 94656 0 1 64061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2792
timestamp 1704896540
transform 1 0 94656 0 1 62429
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2793
timestamp 1704896540
transform 1 0 94112 0 1 60797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2794
timestamp 1704896540
transform 1 0 94112 0 1 60253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2795
timestamp 1704896540
transform 1 0 94112 0 1 62565
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2796
timestamp 1704896540
transform 1 0 94112 0 1 62837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2797
timestamp 1704896540
transform 1 0 95336 0 1 67189
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2798
timestamp 1704896540
transform 1 0 92480 0 1 67189
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2799
timestamp 1704896540
transform 1 0 92616 0 1 67053
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2800
timestamp 1704896540
transform 1 0 92480 0 1 64469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2801
timestamp 1704896540
transform 1 0 94656 0 1 65965
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2802
timestamp 1704896540
transform 1 0 94656 0 1 67597
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2803
timestamp 1704896540
transform 1 0 94656 0 1 69229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2804
timestamp 1704896540
transform 1 0 94112 0 1 69093
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2805
timestamp 1704896540
transform 1 0 94112 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2806
timestamp 1704896540
transform 1 0 75072 0 1 60933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2807
timestamp 1704896540
transform 1 0 75072 0 1 60661
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2808
timestamp 1704896540
transform 1 0 74936 0 1 62429
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2809
timestamp 1704896540
transform 1 0 74936 0 1 62157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2810
timestamp 1704896540
transform 1 0 74664 0 1 61477
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2811
timestamp 1704896540
transform 1 0 74936 0 1 63653
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2812
timestamp 1704896540
transform 1 0 74936 0 1 63381
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2813
timestamp 1704896540
transform 1 0 74664 0 1 61749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2814
timestamp 1704896540
transform 1 0 74800 0 1 64197
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2815
timestamp 1704896540
transform 1 0 74936 0 1 60525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2816
timestamp 1704896540
transform 1 0 74936 0 1 60253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2817
timestamp 1704896540
transform 1 0 74800 0 1 59845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2818
timestamp 1704896540
transform 1 0 75480 0 1 61749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2819
timestamp 1704896540
transform 1 0 75480 0 1 61477
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2820
timestamp 1704896540
transform 1 0 74664 0 1 60253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2821
timestamp 1704896540
transform 1 0 74664 0 1 60525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2822
timestamp 1704896540
transform 1 0 75480 0 1 60525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2823
timestamp 1704896540
transform 1 0 75480 0 1 60253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2824
timestamp 1704896540
transform 1 0 75616 0 1 61341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2825
timestamp 1704896540
transform 1 0 75616 0 1 61069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2826
timestamp 1704896540
transform 1 0 75616 0 1 60661
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2827
timestamp 1704896540
transform 1 0 75616 0 1 60933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2828
timestamp 1704896540
transform 1 0 73984 0 1 61341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2829
timestamp 1704896540
transform 1 0 75208 0 1 62973
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2830
timestamp 1704896540
transform 1 0 74664 0 1 59709
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2831
timestamp 1704896540
transform 1 0 75072 0 1 61749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2832
timestamp 1704896540
transform 1 0 73984 0 1 60933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2833
timestamp 1704896540
transform 1 0 73984 0 1 60661
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2834
timestamp 1704896540
transform 1 0 74800 0 1 60117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2835
timestamp 1704896540
transform 1 0 75616 0 1 59709
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2836
timestamp 1704896540
transform 1 0 75616 0 1 60117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2837
timestamp 1704896540
transform 1 0 75616 0 1 59845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2838
timestamp 1704896540
transform 1 0 73984 0 1 62837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2839
timestamp 1704896540
transform 1 0 75616 0 1 64197
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2840
timestamp 1704896540
transform 1 0 75616 0 1 63789
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2841
timestamp 1704896540
transform 1 0 75616 0 1 64061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2842
timestamp 1704896540
transform 1 0 75616 0 1 61885
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2843
timestamp 1704896540
transform 1 0 75616 0 1 62157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2844
timestamp 1704896540
transform 1 0 75616 0 1 63653
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2845
timestamp 1704896540
transform 1 0 75616 0 1 63381
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2846
timestamp 1704896540
transform 1 0 73984 0 1 62565
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2847
timestamp 1704896540
transform 1 0 73984 0 1 60253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2848
timestamp 1704896540
transform 1 0 74800 0 1 63245
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2849
timestamp 1704896540
transform 1 0 74800 0 1 62973
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2850
timestamp 1704896540
transform 1 0 73984 0 1 60525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2851
timestamp 1704896540
transform 1 0 73848 0 1 62973
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2852
timestamp 1704896540
transform 1 0 73848 0 1 63245
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2853
timestamp 1704896540
transform 1 0 73984 0 1 63381
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2854
timestamp 1704896540
transform 1 0 74392 0 1 63245
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2855
timestamp 1704896540
transform 1 0 74392 0 1 62973
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2856
timestamp 1704896540
transform 1 0 74256 0 1 63381
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2857
timestamp 1704896540
transform 1 0 74256 0 1 63653
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2858
timestamp 1704896540
transform 1 0 74392 0 1 62837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2859
timestamp 1704896540
transform 1 0 74392 0 1 62565
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2860
timestamp 1704896540
transform 1 0 73984 0 1 63653
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2861
timestamp 1704896540
transform 1 0 73984 0 1 64061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2862
timestamp 1704896540
transform 1 0 73984 0 1 63789
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2863
timestamp 1704896540
transform 1 0 75072 0 1 61477
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2864
timestamp 1704896540
transform 1 0 74392 0 1 60525
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2865
timestamp 1704896540
transform 1 0 74392 0 1 60253
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2866
timestamp 1704896540
transform 1 0 74256 0 1 59845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2867
timestamp 1704896540
transform 1 0 74256 0 1 60117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2868
timestamp 1704896540
transform 1 0 74256 0 1 60661
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2869
timestamp 1704896540
transform 1 0 74256 0 1 60933
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2870
timestamp 1704896540
transform 1 0 74256 0 1 61341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2871
timestamp 1704896540
transform 1 0 74256 0 1 61069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2872
timestamp 1704896540
transform 1 0 74392 0 1 63789
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2873
timestamp 1704896540
transform 1 0 74392 0 1 64061
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2874
timestamp 1704896540
transform 1 0 73848 0 1 64197
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2875
timestamp 1704896540
transform 1 0 74392 0 1 64197
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2876
timestamp 1704896540
transform 1 0 73848 0 1 60117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2877
timestamp 1704896540
transform 1 0 73848 0 1 59845
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2878
timestamp 1704896540
transform 1 0 74392 0 1 59709
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2879
timestamp 1704896540
transform 1 0 75208 0 1 63245
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2880
timestamp 1704896540
transform 1 0 73848 0 1 59709
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2881
timestamp 1704896540
transform 1 0 73984 0 1 61069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2882
timestamp 1704896540
transform 1 0 75072 0 1 66101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2883
timestamp 1704896540
transform 1 0 74800 0 1 64469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2884
timestamp 1704896540
transform 1 0 75480 0 1 64605
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2885
timestamp 1704896540
transform 1 0 75480 0 1 64877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2886
timestamp 1704896540
transform 1 0 75616 0 1 65013
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2887
timestamp 1704896540
transform 1 0 75616 0 1 65285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2888
timestamp 1704896540
transform 1 0 75480 0 1 66101
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2889
timestamp 1704896540
transform 1 0 75480 0 1 65829
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2890
timestamp 1704896540
transform 1 0 75480 0 1 65421
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2891
timestamp 1704896540
transform 1 0 75480 0 1 65693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2892
timestamp 1704896540
transform 1 0 75616 0 1 64469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2893
timestamp 1704896540
transform 1 0 75616 0 1 66917
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2894
timestamp 1704896540
transform 1 0 75616 0 1 66645
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2895
timestamp 1704896540
transform 1 0 74936 0 1 65693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2896
timestamp 1704896540
transform 1 0 74528 0 1 67325
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2897
timestamp 1704896540
transform 1 0 74392 0 1 67189
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2898
timestamp 1704896540
transform 1 0 74392 0 1 66917
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2899
timestamp 1704896540
transform 1 0 74256 0 1 64605
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2900
timestamp 1704896540
transform 1 0 74256 0 1 64877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2901
timestamp 1704896540
transform 1 0 74256 0 1 65285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2902
timestamp 1704896540
transform 1 0 74256 0 1 65013
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2903
timestamp 1704896540
transform 1 0 74392 0 1 64469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2904
timestamp 1704896540
transform 1 0 74256 0 1 66781
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2905
timestamp 1704896540
transform 1 0 74256 0 1 66509
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2906
timestamp 1704896540
transform 1 0 74936 0 1 65421
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2907
timestamp 1704896540
transform 1 0 74664 0 1 65421
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2908
timestamp 1704896540
transform 1 0 74664 0 1 65693
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2909
timestamp 1704896540
transform 1 0 74664 0 1 66917
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2910
timestamp 1704896540
transform 1 0 74664 0 1 67189
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2911
timestamp 1704896540
transform 1 0 73984 0 1 64877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2912
timestamp 1704896540
transform 1 0 73984 0 1 64605
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2913
timestamp 1704896540
transform 1 0 73848 0 1 67733
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2914
timestamp 1704896540
transform 1 0 73984 0 1 66509
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2915
timestamp 1704896540
transform 1 0 73984 0 1 66781
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2916
timestamp 1704896540
transform 1 0 73984 0 1 66917
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2917
timestamp 1704896540
transform 1 0 73984 0 1 67189
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2918
timestamp 1704896540
transform 1 0 74664 0 1 68005
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2919
timestamp 1704896540
transform 1 0 73848 0 1 65013
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2920
timestamp 1704896540
transform 1 0 73848 0 1 65285
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2921
timestamp 1704896540
transform 1 0 73848 0 1 67325
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2922
timestamp 1704896540
transform 1 0 73848 0 1 64469
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2923
timestamp 1704896540
transform 1 0 75072 0 1 64605
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2924
timestamp 1704896540
transform 1 0 75072 0 1 64877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2925
timestamp 1704896540
transform 1 0 75072 0 1 66373
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2926
timestamp 1704896540
transform 1 0 82008 0 1 68685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2927
timestamp 1704896540
transform 1 0 82144 0 1 70045
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2928
timestamp 1704896540
transform 1 0 82144 0 1 72765
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2929
timestamp 1704896540
transform 1 0 82008 0 1 74125
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2930
timestamp 1704896540
transform 1 0 82008 0 1 71541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2931
timestamp 1704896540
transform 1 0 82008 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2932
timestamp 1704896540
transform 1 0 81872 0 1 72901
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2933
timestamp 1704896540
transform 1 0 74664 0 1 71541
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2934
timestamp 1704896540
transform 1 0 74800 0 1 70317
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2935
timestamp 1704896540
transform 1 0 74800 0 1 72901
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2936
timestamp 1704896540
transform 1 0 74528 0 1 70181
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2937
timestamp 1704896540
transform 1 0 74392 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2938
timestamp 1704896540
transform 1 0 72760 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2939
timestamp 1704896540
transform 1 0 72760 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2940
timestamp 1704896540
transform 1 0 77656 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2941
timestamp 1704896540
transform 1 0 77656 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2942
timestamp 1704896540
transform 1 0 76160 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2943
timestamp 1704896540
transform 1 0 76160 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2944
timestamp 1704896540
transform 1 0 74392 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2945
timestamp 1704896540
transform 1 0 82144 0 1 78885
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2946
timestamp 1704896540
transform 1 0 82144 0 1 77117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2947
timestamp 1704896540
transform 1 0 82008 0 1 76981
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2948
timestamp 1704896540
transform 1 0 78880 0 1 78885
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2949
timestamp 1704896540
transform 1 0 78880 0 1 76437
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2950
timestamp 1704896540
transform 1 0 82688 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2951
timestamp 1704896540
transform 1 0 82688 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2952
timestamp 1704896540
transform 1 0 81872 0 1 75621
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2953
timestamp 1704896540
transform 1 0 81192 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2954
timestamp 1704896540
transform 1 0 81192 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2955
timestamp 1704896540
transform 1 0 81872 0 1 75757
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2956
timestamp 1704896540
transform 1 0 81872 0 1 77661
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2957
timestamp 1704896540
transform 1 0 79288 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2958
timestamp 1704896540
transform 1 0 79288 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2959
timestamp 1704896540
transform 1 0 79288 0 1 77661
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2960
timestamp 1704896540
transform 1 0 79288 0 1 75077
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2961
timestamp 1704896540
transform 1 0 79424 0 1 75893
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2962
timestamp 1704896540
transform 1 0 82008 0 1 74261
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2963
timestamp 1704896540
transform 1 0 92480 0 1 69909
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2964
timestamp 1704896540
transform 1 0 93419 0 1 69597
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2965
timestamp 1704896540
transform 1 0 94656 0 1 70861
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2966
timestamp 1704896540
transform 1 0 94656 0 1 72493
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2967
timestamp 1704896540
transform 1 0 94112 0 1 70997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2968
timestamp 1704896540
transform 1 0 94112 0 1 71405
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2969
timestamp 1704896540
transform 1 0 89624 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2970
timestamp 1704896540
transform 1 0 89624 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2971
timestamp 1704896540
transform 1 0 87720 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2972
timestamp 1704896540
transform 1 0 87720 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2973
timestamp 1704896540
transform 1 0 86224 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2974
timestamp 1704896540
transform 1 0 86224 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2975
timestamp 1704896540
transform 1 0 84456 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2976
timestamp 1704896540
transform 1 0 84456 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2977
timestamp 1704896540
transform 1 0 95336 0 1 77117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2978
timestamp 1704896540
transform 1 0 94656 0 1 75893
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2979
timestamp 1704896540
transform 1 0 92888 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2980
timestamp 1704896540
transform 1 0 92888 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2981
timestamp 1704896540
transform 1 0 91256 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2982
timestamp 1704896540
transform 1 0 91256 0 1 77797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2983
timestamp 1704896540
transform 1 0 90032 0 1 76437
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2984
timestamp 1704896540
transform 1 0 94656 0 1 74261
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2985
timestamp 1704896540
transform 1 0 75616 0 1 59437
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2986
timestamp 1704896540
transform 1 0 74392 0 1 59437
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2987
timestamp 1704896540
transform 1 0 74664 0 1 59437
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2988
timestamp 1704896540
transform 1 0 73848 0 1 59437
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2989
timestamp 1704896540
transform 1 0 75480 0 1 39717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2990
timestamp 1704896540
transform 1 0 74256 0 1 39717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2991
timestamp 1704896540
transform 1 0 21760 0 1 39717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2992
timestamp 1704896540
transform 1 0 20536 0 1 39717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2993
timestamp 1704896540
transform 1 0 75208 0 1 39717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2994
timestamp 1704896540
transform 1 0 74664 0 1 39717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2995
timestamp 1704896540
transform 1 0 73984 0 1 39717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2996
timestamp 1704896540
transform 1 0 22032 0 1 39717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_34  sky130_sram_1kbyte_1rw1r_32x256_8_contact_34_2997
timestamp 1704896540
transform 1 0 20944 0 1 39717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_39  sky130_sram_1kbyte_1rw1r_32x256_8_contact_39_0
timestamp 1704896540
transform 1 0 94108 0 1 1620
box 0 0 192 192
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_39  sky130_sram_1kbyte_1rw1r_32x256_8_contact_39_1
timestamp 1704896540
transform 1 0 1750 0 1 1620
box 0 0 192 192
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_39  sky130_sram_1kbyte_1rw1r_32x256_8_contact_39_2
timestamp 1704896540
transform 1 0 1750 0 1 77684
box 0 0 192 192
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_39  sky130_sram_1kbyte_1rw1r_32x256_8_contact_39_3
timestamp 1704896540
transform 1 0 94108 0 1 77684
box 0 0 192 192
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_0
timestamp 1704896540
transform 1 0 94928 0 1 957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_1
timestamp 1704896540
transform 1 0 94656 0 1 1093
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_2
timestamp 1704896540
transform 1 0 94928 0 1 1093
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_3
timestamp 1704896540
transform 1 0 94656 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_4
timestamp 1704896540
transform 1 0 95608 0 1 549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_5
timestamp 1704896540
transform 1 0 94792 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_6
timestamp 1704896540
transform 1 0 95472 0 1 549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_7
timestamp 1704896540
transform 1 0 94792 0 1 957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_8
timestamp 1704896540
transform 1 0 95472 0 1 413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_9
timestamp 1704896540
transform 1 0 95472 0 1 277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_10
timestamp 1704896540
transform 1 0 95336 0 1 549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_11
timestamp 1704896540
transform 1 0 95608 0 1 277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_12
timestamp 1704896540
transform 1 0 94928 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_13
timestamp 1704896540
transform 1 0 94656 0 1 957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_14
timestamp 1704896540
transform 1 0 94792 0 1 1093
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_15
timestamp 1704896540
transform 1 0 95336 0 1 413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_16
timestamp 1704896540
transform 1 0 95336 0 1 277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_17
timestamp 1704896540
transform 1 0 95608 0 1 413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_18
timestamp 1704896540
transform 1 0 1088 0 1 1093
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_19
timestamp 1704896540
transform 1 0 952 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_20
timestamp 1704896540
transform 1 0 1088 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_21
timestamp 1704896540
transform 1 0 1224 0 1 1229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_22
timestamp 1704896540
transform 1 0 1224 0 1 957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_23
timestamp 1704896540
transform 1 0 1224 0 1 1093
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_24
timestamp 1704896540
transform 1 0 952 0 1 1093
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_25
timestamp 1704896540
transform 1 0 544 0 1 413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_26
timestamp 1704896540
transform 1 0 408 0 1 413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_27
timestamp 1704896540
transform 1 0 272 0 1 549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_28
timestamp 1704896540
transform 1 0 272 0 1 413
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_29
timestamp 1704896540
transform 1 0 408 0 1 277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_30
timestamp 1704896540
transform 1 0 544 0 1 277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_31
timestamp 1704896540
transform 1 0 952 0 1 957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_32
timestamp 1704896540
transform 1 0 544 0 1 549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_33
timestamp 1704896540
transform 1 0 1088 0 1 957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_34
timestamp 1704896540
transform 1 0 408 0 1 549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_35
timestamp 1704896540
transform 1 0 272 0 1 277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_36
timestamp 1704896540
transform 1 0 1224 0 1 78341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_37
timestamp 1704896540
transform 1 0 272 0 1 78885
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_38
timestamp 1704896540
transform 1 0 544 0 1 78885
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_39
timestamp 1704896540
transform 1 0 544 0 1 79021
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_40
timestamp 1704896540
transform 1 0 408 0 1 78885
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_41
timestamp 1704896540
transform 1 0 272 0 1 79157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_42
timestamp 1704896540
transform 1 0 408 0 1 79021
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_43
timestamp 1704896540
transform 1 0 544 0 1 79157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_44
timestamp 1704896540
transform 1 0 272 0 1 79021
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_45
timestamp 1704896540
transform 1 0 408 0 1 79157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_46
timestamp 1704896540
transform 1 0 1224 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_47
timestamp 1704896540
transform 1 0 1088 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_48
timestamp 1704896540
transform 1 0 952 0 1 78341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_49
timestamp 1704896540
transform 1 0 952 0 1 78477
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_50
timestamp 1704896540
transform 1 0 1224 0 1 78477
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_51
timestamp 1704896540
transform 1 0 952 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_52
timestamp 1704896540
transform 1 0 1088 0 1 78341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_53
timestamp 1704896540
transform 1 0 1088 0 1 78477
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_54
timestamp 1704896540
transform 1 0 95608 0 1 79021
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_55
timestamp 1704896540
transform 1 0 95336 0 1 79157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_56
timestamp 1704896540
transform 1 0 95472 0 1 79021
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_57
timestamp 1704896540
transform 1 0 95608 0 1 79157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_58
timestamp 1704896540
transform 1 0 95472 0 1 78885
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_59
timestamp 1704896540
transform 1 0 95336 0 1 79021
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_60
timestamp 1704896540
transform 1 0 95336 0 1 78885
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_61
timestamp 1704896540
transform 1 0 95608 0 1 78885
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_62
timestamp 1704896540
transform 1 0 95472 0 1 79157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_63
timestamp 1704896540
transform 1 0 94656 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_64
timestamp 1704896540
transform 1 0 94928 0 1 78477
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_65
timestamp 1704896540
transform 1 0 94928 0 1 78341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_66
timestamp 1704896540
transform 1 0 94792 0 1 78477
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_67
timestamp 1704896540
transform 1 0 94792 0 1 78341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_68
timestamp 1704896540
transform 1 0 94656 0 1 78341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_69
timestamp 1704896540
transform 1 0 94656 0 1 78477
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_70
timestamp 1704896540
transform 1 0 94928 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_40  sky130_sram_1kbyte_1rw1r_32x256_8_contact_40_71
timestamp 1704896540
transform 1 0 94792 0 1 78205
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_control_logic_r  sky130_sram_1kbyte_1rw1r_32x256_8_control_logic_r_0
timestamp 1704896540
transform -1 0 93414 0 -1 77108
box -75 -49 11458 18431
use sky130_sram_1kbyte_1rw1r_32x256_8_control_logic_rw  sky130_sram_1kbyte_1rw1r_32x256_8_control_logic_rw_0
timestamp 1704896540
transform 1 0 2636 0 1 4924
box -75 -49 11650 18431
use sky130_sram_1kbyte_1rw1r_32x256_8_cr_3  sky130_sram_1kbyte_1rw1r_32x256_8_cr_3_0
timestamp 1704896540
transform 1 0 14454 0 1 6974
box 2083 -3939 6102 5492
use sky130_sram_1kbyte_1rw1r_32x256_8_cr_4  sky130_sram_1kbyte_1rw1r_32x256_8_cr_4_0
timestamp 1704896540
transform 1 0 14454 0 1 6974
box 3208 -3962 52705 1462
use sky130_sram_1kbyte_1rw1r_32x256_8_cr_5  sky130_sram_1kbyte_1rw1r_32x256_8_cr_5_0
timestamp 1704896540
transform 1 0 14454 0 1 6974
box 61024 65420 64083 68762
use sky130_sram_1kbyte_1rw1r_32x256_8_data_dff  sky130_sram_1kbyte_1rw1r_32x256_8_data_dff_0
timestamp 1704896540
transform 1 0 21294 0 1 2388
box -36 -49 37412 1467
use sky130_sram_1kbyte_1rw1r_32x256_8_row_addr_dff  sky130_sram_1kbyte_1rw1r_32x256_8_row_addr_dff_0
timestamp 1704896540
transform -1 0 83124 0 -1 17150
box -36 -49 1204 9951
use sky130_sram_1kbyte_1rw1r_32x256_8_row_addr_dff  sky130_sram_1kbyte_1rw1r_32x256_8_row_addr_dff_1
timestamp 1704896540
transform 1 0 13118 0 1 25050
box -36 -49 1204 9951
use sky130_sram_1kbyte_1rw1r_32x256_8_wmask_dff  sky130_sram_1kbyte_1rw1r_32x256_8_wmask_dff_0
timestamp 1704896540
transform 1 0 16622 0 1 2388
box -36 -49 4708 1467
<< labels >>
rlabel metal3 s 0 5576 212 5652 4 csb0
port 49 nsew default input
rlabel metal3 s 0 7208 212 7284 4 web0
port 51 nsew default input
rlabel metal3 s 0 25704 212 25780 4 addr0[1]
port 39 nsew default input
rlabel metal3 s 0 27472 212 27548 4 addr0[2]
port 38 nsew default input
rlabel metal3 s 0 28424 212 28500 4 addr0[3]
port 37 nsew default input
rlabel metal3 s 0 30056 212 30132 4 addr0[4]
port 36 nsew default input
rlabel metal3 s 0 31144 212 31220 4 addr0[5]
port 35 nsew default input
rlabel metal3 s 0 32912 212 32988 4 addr0[6]
port 34 nsew default input
rlabel metal3 s 0 34136 212 34212 4 addr0[7]
port 33 nsew default input
rlabel metal3 s 95744 76432 95956 76508 4 csb1
port 50 nsew default input
rlabel metal3 s 95744 16592 95956 16668 4 addr1[1]
port 47 nsew default input
rlabel metal3 s 95744 14960 95956 15036 4 addr1[2]
port 46 nsew default input
rlabel metal3 s 95744 13600 95956 13676 4 addr1[3]
port 45 nsew default input
rlabel metal3 s 952 952 95004 1300 4 vccd1
port 122 nsew power bidirectional abutment
rlabel metal3 s 952 78200 95004 78548 4 vccd1
port 122 nsew power bidirectional abutment
rlabel metal3 s 272 78880 95684 79228 4 vssd1
port 123 nsew ground bidirectional abutment
rlabel metal3 s 272 272 95684 620 4 vssd1
port 123 nsew ground bidirectional abutment
rlabel metal4 s 90032 79288 90108 79500 4 clk1
port 53 nsew default input
rlabel metal4 s 48144 79288 48220 79500 4 dout1[16]
port 105 nsew default output
rlabel metal4 s 49504 79288 49580 79500 4 dout1[17]
port 104 nsew default output
rlabel metal4 s 50592 79288 50668 79500 4 dout1[18]
port 103 nsew default output
rlabel metal4 s 51952 79288 52028 79500 4 dout1[19]
port 102 nsew default output
rlabel metal4 s 53040 79288 53116 79500 4 dout1[20]
port 101 nsew default output
rlabel metal4 s 54264 79288 54340 79500 4 dout1[21]
port 100 nsew default output
rlabel metal4 s 55624 79288 55700 79500 4 dout1[22]
port 99 nsew default output
rlabel metal4 s 56848 79288 56924 79500 4 dout1[23]
port 98 nsew default output
rlabel metal4 s 58208 79288 58284 79500 4 dout1[24]
port 97 nsew default output
rlabel metal4 s 59296 79288 59372 79500 4 dout1[25]
port 96 nsew default output
rlabel metal4 s 60656 79288 60732 79500 4 dout1[26]
port 95 nsew default output
rlabel metal4 s 61880 79288 61956 79500 4 dout1[27]
port 94 nsew default output
rlabel metal4 s 63240 79288 63316 79500 4 dout1[28]
port 93 nsew default output
rlabel metal4 s 64328 79288 64404 79500 4 dout1[29]
port 92 nsew default output
rlabel metal4 s 65552 79288 65628 79500 4 dout1[30]
port 91 nsew default output
rlabel metal4 s 66912 79288 66988 79500 4 dout1[31]
port 90 nsew default output
rlabel metal4 s 79424 79288 79500 79500 4 addr1[0]
port 48 nsew default input
rlabel metal4 s 29512 79288 29588 79500 4 dout1[1]
port 120 nsew default output
rlabel metal4 s 30600 79288 30676 79500 4 dout1[2]
port 119 nsew default output
rlabel metal4 s 31960 79288 32036 79500 4 dout1[3]
port 118 nsew default output
rlabel metal4 s 33184 79288 33260 79500 4 dout1[4]
port 117 nsew default output
rlabel metal4 s 34544 79288 34620 79500 4 dout1[5]
port 116 nsew default output
rlabel metal4 s 35768 79288 35844 79500 4 dout1[6]
port 115 nsew default output
rlabel metal4 s 36856 79288 36932 79500 4 dout1[7]
port 114 nsew default output
rlabel metal4 s 38216 79288 38292 79500 4 dout1[8]
port 113 nsew default output
rlabel metal4 s 39304 79288 39380 79500 4 dout1[9]
port 112 nsew default output
rlabel metal4 s 40664 79288 40740 79500 4 dout1[10]
port 111 nsew default output
rlabel metal4 s 41888 79288 41964 79500 4 dout1[11]
port 110 nsew default output
rlabel metal4 s 43248 79288 43324 79500 4 dout1[12]
port 109 nsew default output
rlabel metal4 s 44336 79288 44412 79500 4 dout1[13]
port 108 nsew default output
rlabel metal4 s 45560 79288 45636 79500 4 dout1[14]
port 107 nsew default output
rlabel metal4 s 46920 79288 46996 79500 4 dout1[15]
port 106 nsew default output
rlabel metal4 s 28152 79288 28228 79500 4 dout1[0]
port 121 nsew default output
rlabel metal4 s 40664 0 40740 212 4 dout0[10]
port 79 nsew default output
rlabel metal4 s 41888 0 41964 212 4 dout0[11]
port 78 nsew default output
rlabel metal4 s 43112 0 43188 212 4 dout0[12]
port 77 nsew default output
rlabel metal4 s 44336 0 44412 212 4 dout0[13]
port 76 nsew default output
rlabel metal4 s 45560 0 45636 212 4 dout0[14]
port 75 nsew default output
rlabel metal4 s 46648 0 46724 212 4 dout0[15]
port 74 nsew default output
rlabel metal4 s 47872 0 47948 212 4 dout0[16]
port 73 nsew default output
rlabel metal4 s 15504 0 15580 212 4 addr0[0]
port 40 nsew default input
rlabel metal4 s 16728 0 16804 212 4 wmask0[0]
port 57 nsew default input
rlabel metal4 s 17816 0 17892 212 4 wmask0[1]
port 56 nsew default input
rlabel metal4 s 19176 0 19252 212 4 wmask0[2]
port 55 nsew default input
rlabel metal4 s 20128 0 20204 212 4 wmask0[3]
port 54 nsew default input
rlabel metal4 s 5848 0 5924 212 4 clk0
port 52 nsew default input
rlabel metal4 s 21352 0 21428 212 4 din0[0]
port 32 nsew default input
rlabel metal4 s 22576 0 22652 212 4 din0[1]
port 31 nsew default input
rlabel metal4 s 23664 0 23740 212 4 din0[2]
port 30 nsew default input
rlabel metal4 s 25024 0 25100 212 4 din0[3]
port 29 nsew default input
rlabel metal4 s 26112 0 26188 212 4 din0[4]
port 28 nsew default input
rlabel metal4 s 27200 0 27276 212 4 din0[5]
port 27 nsew default input
rlabel metal4 s 28288 0 28364 212 4 din0[6]
port 26 nsew default input
rlabel metal4 s 29648 0 29724 212 4 din0[7]
port 25 nsew default input
rlabel metal4 s 30736 0 30812 212 4 din0[8]
port 24 nsew default input
rlabel metal4 s 31824 0 31900 212 4 din0[9]
port 23 nsew default input
rlabel metal4 s 33048 0 33124 212 4 din0[10]
port 22 nsew default input
rlabel metal4 s 34136 0 34212 212 4 din0[11]
port 21 nsew default input
rlabel metal4 s 35496 0 35572 212 4 din0[12]
port 20 nsew default input
rlabel metal4 s 36584 0 36660 212 4 din0[13]
port 19 nsew default input
rlabel metal4 s 37672 0 37748 212 4 din0[14]
port 18 nsew default input
rlabel metal4 s 38896 0 38972 212 4 din0[15]
port 17 nsew default input
rlabel metal4 s 40256 0 40332 212 4 din0[16]
port 16 nsew default input
rlabel metal4 s 41344 0 41420 212 4 din0[17]
port 15 nsew default input
rlabel metal4 s 42432 0 42508 212 4 din0[18]
port 14 nsew default input
rlabel metal4 s 43520 0 43596 212 4 din0[19]
port 13 nsew default input
rlabel metal4 s 44880 0 44956 212 4 din0[20]
port 12 nsew default input
rlabel metal4 s 45968 0 46044 212 4 din0[21]
port 11 nsew default input
rlabel metal4 s 47056 0 47132 212 4 din0[22]
port 10 nsew default input
rlabel metal4 s 27880 0 27956 212 4 dout0[0]
port 89 nsew default output
rlabel metal4 s 29240 0 29316 212 4 dout0[1]
port 88 nsew default output
rlabel metal4 s 30328 0 30404 212 4 dout0[2]
port 87 nsew default output
rlabel metal4 s 31960 0 32036 212 4 dout0[3]
port 86 nsew default output
rlabel metal4 s 33184 0 33260 212 4 dout0[4]
port 85 nsew default output
rlabel metal4 s 34408 0 34484 212 4 dout0[5]
port 84 nsew default output
rlabel metal4 s 35632 0 35708 212 4 dout0[6]
port 83 nsew default output
rlabel metal4 s 36856 0 36932 212 4 dout0[7]
port 82 nsew default output
rlabel metal4 s 37808 0 37884 212 4 dout0[8]
port 81 nsew default output
rlabel metal4 s 39304 0 39380 212 4 dout0[9]
port 80 nsew default output
rlabel metal4 s 952 952 1300 78548 4 vccd1
port 122 nsew power bidirectional abutment
rlabel metal4 s 272 272 620 79228 4 vssd1
port 123 nsew ground bidirectional abutment
rlabel metal4 s 59296 0 59372 212 4 dout0[25]
port 64 nsew default output
rlabel metal4 s 60520 0 60596 212 4 dout0[26]
port 63 nsew default output
rlabel metal4 s 61880 0 61956 212 4 dout0[27]
port 62 nsew default output
rlabel metal4 s 63104 0 63180 212 4 dout0[28]
port 61 nsew default output
rlabel metal4 s 64328 0 64404 212 4 dout0[29]
port 60 nsew default output
rlabel metal4 s 65552 0 65628 212 4 dout0[30]
port 59 nsew default output
rlabel metal4 s 66776 0 66852 212 4 dout0[31]
port 58 nsew default output
rlabel metal4 s 57664 0 57740 212 4 din0[31]
port 1 nsew default input
rlabel metal4 s 48280 0 48356 212 4 din0[23]
port 9 nsew default input
rlabel metal4 s 49368 0 49444 212 4 din0[24]
port 8 nsew default input
rlabel metal4 s 50728 0 50804 212 4 din0[25]
port 7 nsew default input
rlabel metal4 s 51816 0 51892 212 4 din0[26]
port 6 nsew default input
rlabel metal4 s 52904 0 52980 212 4 din0[27]
port 5 nsew default input
rlabel metal4 s 53992 0 54068 212 4 din0[28]
port 4 nsew default input
rlabel metal4 s 55216 0 55292 212 4 din0[29]
port 3 nsew default input
rlabel metal4 s 56576 0 56652 212 4 din0[30]
port 2 nsew default input
rlabel metal4 s 49096 0 49172 212 4 dout0[17]
port 72 nsew default output
rlabel metal4 s 50592 0 50668 212 4 dout0[18]
port 71 nsew default output
rlabel metal4 s 51408 0 51484 212 4 dout0[19]
port 70 nsew default output
rlabel metal4 s 53176 0 53252 212 4 dout0[20]
port 69 nsew default output
rlabel metal4 s 54400 0 54476 212 4 dout0[21]
port 68 nsew default output
rlabel metal4 s 55624 0 55700 212 4 dout0[22]
port 67 nsew default output
rlabel metal4 s 83096 0 83172 212 4 addr1[4]
port 44 nsew default input
rlabel metal4 s 82688 0 82764 212 4 addr1[5]
port 43 nsew default input
rlabel metal4 s 82824 0 82900 212 4 addr1[6]
port 42 nsew default input
rlabel metal4 s 82960 0 83036 212 4 addr1[7]
port 41 nsew default input
rlabel metal4 s 94656 952 95004 78548 4 vccd1
port 122 nsew power bidirectional abutment
rlabel metal4 s 56848 0 56924 212 4 dout0[23]
port 66 nsew default output
rlabel metal4 s 57800 0 57876 212 4 dout0[24]
port 65 nsew default output
rlabel metal4 s 95336 272 95684 79228 4 vssd1
port 123 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 95956 79500
string GDS_END 9871762
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_32x256_8.gds
string GDS_START 8110160
string LEFclass BLOCK
string LEFsymmetry X Y R90
<< end >>
