magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< locali >>
rect 59870 65486 59904 65502
rect 59870 65436 59904 65452
<< viali >>
rect 59870 65452 59904 65486
<< metal1 >>
rect 59855 67389 59861 67441
rect 59913 67429 59919 67441
rect 63859 67429 63865 67441
rect 59913 67401 63865 67429
rect 59913 67389 59919 67401
rect 63859 67389 63865 67401
rect 63917 67389 63923 67441
rect 59855 65443 59861 65495
rect 59913 65443 59919 65495
<< via1 >>
rect 59861 67389 59913 67441
rect 63865 67389 63917 67441
rect 59861 65486 59913 65495
rect 59861 65452 59870 65486
rect 59870 65452 59904 65486
rect 59904 65452 59913 65486
rect 59861 65443 59913 65452
<< metal2 >>
rect 63877 67447 63905 69102
rect 59861 67441 59913 67447
rect 59861 67383 59913 67389
rect 63865 67441 63917 67447
rect 63865 67383 63917 67389
rect 59873 65501 59901 67383
rect 59861 65495 59913 65501
rect 59861 65437 59913 65443
use contact_7  contact_7_0
timestamp 1704896540
transform 1 0 59858 0 1 65436
box 0 0 1 1
use contact_8  contact_8_0
timestamp 1704896540
transform 1 0 63859 0 1 67383
box 0 0 1 1
use contact_8  contact_8_1
timestamp 1704896540
transform 1 0 59855 0 1 65437
box 0 0 1 1
use contact_8  contact_8_2
timestamp 1704896540
transform 1 0 59855 0 1 67383
box 0 0 1 1
<< properties >>
string FIXED_BBOX 59855 65436 63923 69102
string GDS_END 6490110
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 6489522
<< end >>
