magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -108 515 1517 1337
<< pwell >>
rect -67 367 67 455
rect 285 367 419 455
rect 637 367 771 455
rect 989 367 1123 455
rect 1341 367 1475 455
<< mvpsubdiff >>
rect -41 427 41 429
rect -41 393 -17 427
rect 17 393 41 427
rect 311 427 393 429
rect 311 393 335 427
rect 369 393 393 427
rect 663 427 745 429
rect 663 393 687 427
rect 721 393 745 427
rect 1015 427 1097 429
rect 1015 393 1039 427
rect 1073 393 1097 427
rect 1367 427 1449 429
rect 1367 393 1391 427
rect 1425 393 1449 427
<< mvnsubdiff >>
rect -41 583 -17 617
rect 17 583 41 617
rect -41 581 41 583
rect 311 583 335 617
rect 369 583 393 617
rect 311 581 393 583
rect 663 583 687 617
rect 721 583 745 617
rect 663 581 745 583
rect 1015 583 1039 617
rect 1073 583 1097 617
rect 1015 581 1097 583
rect 1367 583 1391 617
rect 1425 583 1449 617
rect 1367 581 1449 583
<< mvpsubdiffcont >>
rect -17 393 17 427
rect 335 393 369 427
rect 687 393 721 427
rect 1039 393 1073 427
rect 1391 393 1425 427
<< mvnsubdiffcont >>
rect -17 583 17 617
rect 335 583 369 617
rect 687 583 721 617
rect 1039 583 1073 617
rect 1391 583 1425 617
<< poly >>
rect 21 1353 1387 1369
rect 21 1319 37 1353
rect 71 1319 105 1353
rect 139 1319 213 1353
rect 247 1319 281 1353
rect 315 1319 389 1353
rect 423 1319 457 1353
rect 491 1319 565 1353
rect 599 1319 633 1353
rect 667 1319 741 1353
rect 775 1319 809 1353
rect 843 1319 916 1353
rect 950 1319 984 1353
rect 1018 1319 1093 1353
rect 1127 1319 1161 1353
rect 1195 1319 1269 1353
rect 1303 1319 1337 1353
rect 1371 1319 1387 1353
rect 21 1303 1387 1319
rect 28 1297 1387 1303
rect 52 345 147 645
rect 204 345 300 645
rect 404 345 500 645
rect 556 345 652 645
rect 756 345 852 645
rect 908 345 1004 645
rect 1108 345 1204 645
rect 1260 345 1356 645
rect 28 87 1387 93
rect 21 71 1387 87
rect 21 37 37 71
rect 71 37 105 71
rect 139 37 213 71
rect 247 37 281 71
rect 315 37 389 71
rect 423 37 457 71
rect 491 37 565 71
rect 599 37 633 71
rect 667 37 741 71
rect 775 37 809 71
rect 843 37 917 71
rect 951 37 985 71
rect 1019 37 1093 71
rect 1127 37 1161 71
rect 1195 37 1269 71
rect 1303 37 1337 71
rect 1371 37 1387 71
rect 21 21 1387 37
<< polycont >>
rect 37 1319 71 1353
rect 105 1319 139 1353
rect 213 1319 247 1353
rect 281 1319 315 1353
rect 389 1319 423 1353
rect 457 1319 491 1353
rect 565 1319 599 1353
rect 633 1319 667 1353
rect 741 1319 775 1353
rect 809 1319 843 1353
rect 916 1319 950 1353
rect 984 1319 1018 1353
rect 1093 1319 1127 1353
rect 1161 1319 1195 1353
rect 1269 1319 1303 1353
rect 1337 1319 1371 1353
rect 37 37 71 71
rect 105 37 139 71
rect 213 37 247 71
rect 281 37 315 71
rect 389 37 423 71
rect 457 37 491 71
rect 565 37 599 71
rect 633 37 667 71
rect 741 37 775 71
rect 809 37 843 71
rect 917 37 951 71
rect 985 37 1019 71
rect 1093 37 1127 71
rect 1161 37 1195 71
rect 1269 37 1303 71
rect 1337 37 1371 71
<< locali >>
rect 37 1353 139 1369
rect 71 1319 105 1353
rect 37 1303 139 1319
rect 213 1353 491 1369
rect 247 1319 281 1353
rect 315 1319 389 1353
rect 423 1319 457 1353
rect 213 1309 491 1319
rect 213 1303 315 1309
rect 389 1303 491 1309
rect 565 1353 843 1369
rect 599 1319 633 1353
rect 667 1319 741 1353
rect 775 1319 809 1353
rect 565 1309 843 1319
rect 565 1303 667 1309
rect 741 1303 843 1309
rect 916 1353 1195 1369
rect 950 1319 984 1353
rect 1018 1319 1093 1353
rect 1127 1319 1161 1353
rect 916 1309 1195 1319
rect 916 1303 1018 1309
rect 1093 1303 1195 1309
rect 1269 1353 1371 1369
rect 1303 1319 1337 1353
rect 1269 1303 1371 1319
rect -17 785 17 823
rect -17 713 17 751
rect -17 667 5 679
rect -17 567 17 583
rect -17 427 17 443
rect -17 259 17 297
rect -17 187 17 225
rect -17 121 17 153
rect 51 87 125 1303
rect 159 485 193 1269
rect 159 121 193 451
rect 227 87 301 1303
rect 335 785 369 823
rect 335 713 369 751
rect 335 567 369 583
rect 335 427 369 443
rect 335 259 369 297
rect 335 187 369 225
rect 403 87 477 1303
rect 511 485 545 1269
rect 511 121 545 451
rect 579 87 653 1303
rect 687 785 721 823
rect 687 713 721 751
rect 687 667 721 679
rect 687 567 721 583
rect 687 427 721 443
rect 687 259 721 297
rect 687 187 721 225
rect 755 87 829 1303
rect 863 485 897 1269
rect 863 121 897 451
rect 931 87 1005 1303
rect 1039 785 1073 823
rect 1039 713 1073 751
rect 1039 668 1073 679
rect 1039 567 1073 583
rect 1039 427 1073 443
rect 1039 259 1073 297
rect 1039 187 1073 225
rect 1039 121 1073 153
rect 1107 87 1181 1303
rect 1215 485 1249 1269
rect 1215 121 1249 451
rect 1283 87 1357 1303
rect 1391 857 1425 869
rect 1391 785 1425 823
rect 1391 713 1425 751
rect 1391 668 1425 679
rect 1391 567 1425 583
rect 1391 427 1425 443
rect 1391 259 1425 297
rect 1391 187 1425 225
rect 1391 121 1425 153
rect 37 71 139 87
rect 71 37 105 71
rect 37 21 139 37
rect 213 81 315 87
rect 389 81 491 87
rect 213 71 491 81
rect 247 37 281 71
rect 315 37 389 71
rect 423 37 457 71
rect 213 21 491 37
rect 565 81 667 87
rect 741 81 843 87
rect 565 71 843 81
rect 599 37 633 71
rect 667 37 741 71
rect 775 37 809 71
rect 565 21 843 37
rect 917 81 1019 87
rect 1093 81 1195 87
rect 917 71 1195 81
rect 951 37 985 71
rect 1019 37 1093 71
rect 1127 37 1161 71
rect 917 21 1195 37
rect 1269 71 1371 87
rect 1303 37 1337 71
rect 1269 21 1371 37
<< viali >>
rect -17 823 17 857
rect -17 751 17 785
rect -17 679 17 713
rect -17 617 17 633
rect -17 599 17 617
rect -17 393 17 411
rect -17 377 17 393
rect -17 297 17 331
rect -17 225 17 259
rect -17 153 17 187
rect 159 451 193 485
rect 335 823 369 857
rect 335 751 369 785
rect 335 679 369 713
rect 335 617 369 633
rect 335 599 369 617
rect 335 393 369 411
rect 335 377 369 393
rect 335 297 369 331
rect 335 225 369 259
rect 335 153 369 187
rect 511 451 545 485
rect 687 823 721 857
rect 687 751 721 785
rect 687 679 721 713
rect 687 617 721 633
rect 687 599 721 617
rect 687 393 721 411
rect 687 377 721 393
rect 687 297 721 331
rect 687 225 721 259
rect 687 153 721 187
rect 863 451 897 485
rect 1039 823 1073 857
rect 1039 751 1073 785
rect 1039 679 1073 713
rect 1039 617 1073 633
rect 1039 599 1073 617
rect 1039 393 1073 411
rect 1039 377 1073 393
rect 1039 297 1073 331
rect 1039 225 1073 259
rect 1039 153 1073 187
rect 1215 451 1249 485
rect 1391 823 1425 857
rect 1391 751 1425 785
rect 1391 679 1425 713
rect 1391 617 1425 633
rect 1391 599 1425 617
rect 1391 393 1425 411
rect 1391 377 1425 393
rect 1391 297 1425 331
rect 1391 225 1425 259
rect 1391 153 1425 187
<< metal1 >>
rect -29 857 1437 869
rect -29 823 -17 857
rect 17 823 335 857
rect 369 823 687 857
rect 721 823 1039 857
rect 1073 823 1391 857
rect 1425 823 1437 857
rect -29 785 1437 823
rect -29 751 -17 785
rect 17 751 335 785
rect 369 751 687 785
rect 721 751 1039 785
rect 1073 751 1391 785
rect 1425 751 1437 785
rect -29 713 1437 751
rect -29 679 -17 713
rect 17 679 335 713
rect 369 679 687 713
rect 721 679 1039 713
rect 1073 679 1391 713
rect 1425 679 1437 713
rect -29 667 1437 679
rect -29 633 1437 639
rect -29 599 -17 633
rect 17 599 335 633
rect 369 599 687 633
rect 721 599 1039 633
rect 1073 599 1391 633
rect 1425 599 1437 633
rect -29 593 1437 599
rect 147 485 1261 491
rect 147 451 159 485
rect 193 451 511 485
rect 545 451 863 485
rect 897 451 1215 485
rect 1249 451 1261 485
rect 147 445 1261 451
rect -29 411 1437 417
rect -29 377 -17 411
rect 17 377 335 411
rect 369 377 687 411
rect 721 377 1039 411
rect 1073 377 1391 411
rect 1425 377 1437 411
rect -29 371 1437 377
rect -29 331 1437 343
rect -29 297 -17 331
rect 17 297 335 331
rect 369 297 687 331
rect 721 297 1039 331
rect 1073 297 1391 331
rect 1425 297 1437 331
rect -29 259 1437 297
rect -29 225 -17 259
rect 17 225 335 259
rect 369 225 687 259
rect 721 225 1039 259
rect 1073 225 1391 259
rect 1425 225 1437 259
rect -29 187 1437 225
rect -29 153 -17 187
rect 17 153 335 187
rect 369 153 687 187
rect 721 153 1039 187
rect 1073 153 1391 187
rect 1425 153 1437 187
rect -29 141 1437 153
use hvnTran_CDNS_524688791851168  hvnTran_CDNS_524688791851168_0
timestamp 1704896540
transform 1 0 28 0 -1 319
box -79 -26 1431 226
use hvpTran_CDNS_524688791851169  hvpTran_CDNS_524688791851169_0
timestamp 1704896540
transform 1 0 28 0 1 671
box -119 -66 1471 666
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1704896540
transform 0 -1 17 -1 0 857
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_1
timestamp 1704896540
transform 0 -1 369 -1 0 857
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_2
timestamp 1704896540
transform 0 -1 721 -1 0 857
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_3
timestamp 1704896540
transform 0 -1 1073 -1 0 857
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_4
timestamp 1704896540
transform 0 -1 17 -1 0 331
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_5
timestamp 1704896540
transform 0 -1 369 -1 0 331
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_6
timestamp 1704896540
transform 0 -1 721 -1 0 331
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_7
timestamp 1704896540
transform 0 -1 1073 -1 0 331
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_8
timestamp 1704896540
transform 0 -1 1425 -1 0 331
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_9
timestamp 1704896540
transform 0 -1 1425 1 0 679
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_0
timestamp 1704896540
transform 1 0 687 0 1 377
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_1
timestamp 1704896540
transform 1 0 1391 0 1 377
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_2
timestamp 1704896540
transform 1 0 -17 0 1 599
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_3
timestamp 1704896540
transform 1 0 335 0 1 599
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_4
timestamp 1704896540
transform 1 0 687 0 1 599
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_5
timestamp 1704896540
transform 1 0 1039 0 1 599
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_6
timestamp 1704896540
transform 1 0 1391 0 1 599
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_7
timestamp 1704896540
transform 1 0 335 0 1 377
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_8
timestamp 1704896540
transform 1 0 1039 0 1 377
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_9
timestamp 1704896540
transform 1 0 863 0 1 451
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_10
timestamp 1704896540
transform 1 0 511 0 1 451
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_11
timestamp 1704896540
transform 1 0 1215 0 1 451
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_12
timestamp 1704896540
transform 1 0 159 0 1 451
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_13
timestamp 1704896540
transform 1 0 -17 0 1 377
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_0
timestamp 1704896540
transform 1 0 725 0 1 1303
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_1
timestamp 1704896540
transform 1 0 21 0 1 21
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_2
timestamp 1704896540
transform 1 0 197 0 1 21
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_3
timestamp 1704896540
transform 1 0 373 0 1 21
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_4
timestamp 1704896540
transform 1 0 549 0 1 21
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_5
timestamp 1704896540
transform 1 0 1077 0 1 21
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_6
timestamp 1704896540
transform 1 0 1253 0 1 21
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_7
timestamp 1704896540
transform 1 0 725 0 1 21
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_8
timestamp 1704896540
transform 1 0 901 0 1 21
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_9
timestamp 1704896540
transform 1 0 21 0 1 1303
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_10
timestamp 1704896540
transform 1 0 197 0 1 1303
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_11
timestamp 1704896540
transform 1 0 373 0 1 1303
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_12
timestamp 1704896540
transform 1 0 549 0 1 1303
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_13
timestamp 1704896540
transform 1 0 900 0 1 1303
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_14
timestamp 1704896540
transform 1 0 1077 0 1 1303
box 0 0 1 1
use PYL1_CDNS_5246887918526  PYL1_CDNS_5246887918526_15
timestamp 1704896540
transform 1 0 1253 0 1 1303
box 0 0 1 1
<< labels >>
flabel comment s 192 63 192 63 0 FreeSans 100 0 0 0 no_jumper_check
flabel comment s 369 63 369 63 0 FreeSans 100 0 0 0 no_jumper_check
flabel comment s 544 63 544 63 0 FreeSans 100 0 0 0 no_jumper_check
flabel comment s 723 63 723 63 0 FreeSans 100 0 0 0 no_jumper_check
flabel comment s 896 63 896 63 0 FreeSans 100 0 0 0 no_jumper_check
flabel comment s 1065 63 1065 63 0 FreeSans 100 0 0 0 no_jumper_check
flabel comment s 1244 63 1244 63 0 FreeSans 100 0 0 0 no_jumper_check
flabel metal1 s 1396 141 1408 343 3 FreeSans 200 180 0 0 vgnd
port 1 nsew
flabel metal1 s 1396 371 1408 417 3 FreeSans 200 180 0 0 vnb
port 2 nsew
flabel metal1 s 1396 593 1408 639 3 FreeSans 200 180 0 0 vpb
port 3 nsew
flabel metal1 s 1396 667 1408 869 3 FreeSans 200 180 0 0 vpwr
port 4 nsew
flabel metal1 s 0 141 12 343 3 FreeSans 200 0 0 0 vgnd
port 1 nsew
flabel metal1 s 0 371 12 417 3 FreeSans 200 0 0 0 vnb
port 2 nsew
flabel metal1 s 0 593 12 639 3 FreeSans 200 0 0 0 vpb
port 3 nsew
flabel metal1 s 0 667 12 869 3 FreeSans 200 0 0 0 vpwr
port 4 nsew
flabel locali s 950 1310 984 1360 0 FreeSans 200 0 0 0 in
port 6 nsew
flabel locali s 1303 1306 1337 1356 0 FreeSans 200 0 0 0 in
port 6 nsew
flabel locali s 423 1306 457 1356 0 FreeSans 200 0 0 0 in
port 6 nsew
flabel locali s 599 1306 633 1356 0 FreeSans 200 0 0 0 in
port 6 nsew
flabel locali s 247 1306 281 1356 0 FreeSans 200 0 0 0 in
port 6 nsew
flabel locali s 71 1306 105 1356 0 FreeSans 200 0 0 0 in
port 6 nsew
flabel locali s 1127 21 1161 71 0 FreeSans 200 0 0 0 in
port 6 nsew
flabel locali s 949 21 983 71 0 FreeSans 200 0 0 0 in
port 6 nsew
flabel locali s 775 21 809 71 0 FreeSans 200 0 0 0 in
port 6 nsew
flabel locali s 1303 21 1337 71 0 FreeSans 200 0 0 0 in
port 6 nsew
flabel locali s 423 21 457 71 0 FreeSans 200 0 0 0 in
port 6 nsew
flabel locali s 599 21 633 71 0 FreeSans 200 0 0 0 in
port 6 nsew
flabel locali s 247 21 281 71 0 FreeSans 200 0 0 0 in
port 6 nsew
flabel locali s 72 21 106 71 0 FreeSans 200 0 0 0 in
port 6 nsew
flabel locali s 511 121 545 171 0 FreeSans 200 0 0 0 out
port 7 nsew
flabel locali s 1215 1220 1249 1269 0 FreeSans 200 0 0 0 out
port 7 nsew
flabel locali s 863 1220 897 1269 0 FreeSans 200 0 0 0 out
port 7 nsew
flabel locali s 1215 121 1249 171 0 FreeSans 200 0 0 0 out
port 7 nsew
flabel locali s 159 121 193 171 0 FreeSans 200 0 0 0 out
port 7 nsew
flabel locali s 159 1220 193 1269 0 FreeSans 200 0 0 0 out
port 7 nsew
flabel locali s 863 121 897 171 0 FreeSans 200 0 0 0 out
port 7 nsew
flabel locali s 775 1306 809 1356 0 FreeSans 200 0 0 0 in
port 6 nsew
flabel locali s 511 1220 545 1269 0 FreeSans 200 0 0 0 out
port 7 nsew
flabel locali s 1127 1306 1161 1356 0 FreeSans 200 0 0 0 in
port 6 nsew
<< properties >>
string GDS_END 85328766
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85315956
<< end >>
