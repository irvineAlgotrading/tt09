magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< pwell >>
rect 0 89 883 1151
<< nmos >>
rect 194 115 224 1125
rect 348 115 378 1125
rect 502 115 532 1125
rect 656 115 686 1125
<< ndiff >>
rect 138 1113 194 1125
rect 138 1079 149 1113
rect 183 1079 194 1113
rect 138 1045 194 1079
rect 138 1011 149 1045
rect 183 1011 194 1045
rect 138 977 194 1011
rect 138 943 149 977
rect 183 943 194 977
rect 138 909 194 943
rect 138 875 149 909
rect 183 875 194 909
rect 138 841 194 875
rect 138 807 149 841
rect 183 807 194 841
rect 138 773 194 807
rect 138 739 149 773
rect 183 739 194 773
rect 138 705 194 739
rect 138 671 149 705
rect 183 671 194 705
rect 138 637 194 671
rect 138 603 149 637
rect 183 603 194 637
rect 138 569 194 603
rect 138 535 149 569
rect 183 535 194 569
rect 138 501 194 535
rect 138 467 149 501
rect 183 467 194 501
rect 138 433 194 467
rect 138 399 149 433
rect 183 399 194 433
rect 138 365 194 399
rect 138 331 149 365
rect 183 331 194 365
rect 138 297 194 331
rect 138 263 149 297
rect 183 263 194 297
rect 138 229 194 263
rect 138 195 149 229
rect 183 195 194 229
rect 138 161 194 195
rect 138 127 149 161
rect 183 127 194 161
rect 138 115 194 127
rect 224 1113 348 1125
rect 224 127 235 1113
rect 337 127 348 1113
rect 224 115 348 127
rect 378 1113 502 1125
rect 378 127 389 1113
rect 491 127 502 1113
rect 378 115 502 127
rect 532 1113 656 1125
rect 532 127 543 1113
rect 645 127 656 1113
rect 532 115 656 127
rect 686 1113 745 1125
rect 686 1079 697 1113
rect 731 1079 745 1113
rect 686 1045 745 1079
rect 686 1011 697 1045
rect 731 1011 745 1045
rect 686 977 745 1011
rect 686 943 697 977
rect 731 943 745 977
rect 686 909 745 943
rect 686 875 697 909
rect 731 875 745 909
rect 686 841 745 875
rect 686 807 697 841
rect 731 807 745 841
rect 686 773 745 807
rect 686 739 697 773
rect 731 739 745 773
rect 686 705 745 739
rect 686 671 697 705
rect 731 671 745 705
rect 686 637 745 671
rect 686 603 697 637
rect 731 603 745 637
rect 686 569 745 603
rect 686 535 697 569
rect 731 535 745 569
rect 686 501 745 535
rect 686 467 697 501
rect 731 467 745 501
rect 686 433 745 467
rect 686 399 697 433
rect 731 399 745 433
rect 686 365 745 399
rect 686 331 697 365
rect 731 331 745 365
rect 686 297 745 331
rect 686 263 697 297
rect 731 263 745 297
rect 686 229 745 263
rect 686 195 697 229
rect 731 195 745 229
rect 686 161 745 195
rect 686 127 697 161
rect 731 127 745 161
rect 686 115 745 127
<< ndiffc >>
rect 149 1079 183 1113
rect 149 1011 183 1045
rect 149 943 183 977
rect 149 875 183 909
rect 149 807 183 841
rect 149 739 183 773
rect 149 671 183 705
rect 149 603 183 637
rect 149 535 183 569
rect 149 467 183 501
rect 149 399 183 433
rect 149 331 183 365
rect 149 263 183 297
rect 149 195 183 229
rect 149 127 183 161
rect 235 127 337 1113
rect 389 127 491 1113
rect 543 127 645 1113
rect 697 1079 731 1113
rect 697 1011 731 1045
rect 697 943 731 977
rect 697 875 731 909
rect 697 807 731 841
rect 697 739 731 773
rect 697 671 731 705
rect 697 603 731 637
rect 697 535 731 569
rect 697 467 731 501
rect 697 399 731 433
rect 697 331 731 365
rect 697 263 731 297
rect 697 195 731 229
rect 697 127 731 161
<< psubdiff >>
rect 26 1079 84 1125
rect 26 1045 38 1079
rect 72 1045 84 1079
rect 26 1011 84 1045
rect 26 977 38 1011
rect 72 977 84 1011
rect 26 943 84 977
rect 26 909 38 943
rect 72 909 84 943
rect 26 875 84 909
rect 26 841 38 875
rect 72 841 84 875
rect 26 807 84 841
rect 26 773 38 807
rect 72 773 84 807
rect 26 739 84 773
rect 26 705 38 739
rect 72 705 84 739
rect 26 671 84 705
rect 26 637 38 671
rect 72 637 84 671
rect 26 603 84 637
rect 26 569 38 603
rect 72 569 84 603
rect 26 535 84 569
rect 26 501 38 535
rect 72 501 84 535
rect 26 467 84 501
rect 26 433 38 467
rect 72 433 84 467
rect 26 399 84 433
rect 26 365 38 399
rect 72 365 84 399
rect 26 331 84 365
rect 26 297 38 331
rect 72 297 84 331
rect 26 263 84 297
rect 26 229 38 263
rect 72 229 84 263
rect 26 195 84 229
rect 26 161 38 195
rect 72 161 84 195
rect 26 115 84 161
rect 799 1079 857 1125
rect 799 1045 811 1079
rect 845 1045 857 1079
rect 799 1011 857 1045
rect 799 977 811 1011
rect 845 977 857 1011
rect 799 943 857 977
rect 799 909 811 943
rect 845 909 857 943
rect 799 875 857 909
rect 799 841 811 875
rect 845 841 857 875
rect 799 807 857 841
rect 799 773 811 807
rect 845 773 857 807
rect 799 739 857 773
rect 799 705 811 739
rect 845 705 857 739
rect 799 671 857 705
rect 799 637 811 671
rect 845 637 857 671
rect 799 603 857 637
rect 799 569 811 603
rect 845 569 857 603
rect 799 535 857 569
rect 799 501 811 535
rect 845 501 857 535
rect 799 467 857 501
rect 799 433 811 467
rect 845 433 857 467
rect 799 399 857 433
rect 799 365 811 399
rect 845 365 857 399
rect 799 331 857 365
rect 799 297 811 331
rect 845 297 857 331
rect 799 263 857 297
rect 799 229 811 263
rect 845 229 857 263
rect 799 195 857 229
rect 799 161 811 195
rect 845 161 857 195
rect 799 115 857 161
<< psubdiffcont >>
rect 38 1045 72 1079
rect 38 977 72 1011
rect 38 909 72 943
rect 38 841 72 875
rect 38 773 72 807
rect 38 705 72 739
rect 38 637 72 671
rect 38 569 72 603
rect 38 501 72 535
rect 38 433 72 467
rect 38 365 72 399
rect 38 297 72 331
rect 38 229 72 263
rect 38 161 72 195
rect 811 1045 845 1079
rect 811 977 845 1011
rect 811 909 845 943
rect 811 841 845 875
rect 811 773 845 807
rect 811 705 845 739
rect 811 637 845 671
rect 811 569 845 603
rect 811 501 845 535
rect 811 433 845 467
rect 811 365 845 399
rect 811 297 845 331
rect 811 229 845 263
rect 811 161 845 195
<< poly >>
rect 194 1220 736 1236
rect 194 1186 210 1220
rect 244 1186 278 1220
rect 312 1186 346 1220
rect 380 1186 414 1220
rect 448 1186 482 1220
rect 516 1186 550 1220
rect 584 1186 618 1220
rect 652 1186 686 1220
rect 720 1186 736 1220
rect 194 1170 736 1186
rect 194 1125 224 1170
rect 348 1125 378 1170
rect 502 1125 532 1170
rect 656 1125 686 1170
rect 194 70 224 115
rect 348 70 378 115
rect 502 70 532 115
rect 656 70 686 115
rect 194 54 736 70
rect 194 20 210 54
rect 244 20 278 54
rect 312 20 346 54
rect 380 20 414 54
rect 448 20 482 54
rect 516 20 550 54
rect 584 20 618 54
rect 652 20 686 54
rect 720 20 736 54
rect 194 4 736 20
<< polycont >>
rect 210 1186 244 1220
rect 278 1186 312 1220
rect 346 1186 380 1220
rect 414 1186 448 1220
rect 482 1186 516 1220
rect 550 1186 584 1220
rect 618 1186 652 1220
rect 686 1186 720 1220
rect 210 20 244 54
rect 278 20 312 54
rect 346 20 380 54
rect 414 20 448 54
rect 482 20 516 54
rect 550 20 584 54
rect 618 20 652 54
rect 686 20 720 54
<< locali >>
rect 244 1186 266 1220
rect 312 1186 338 1220
rect 380 1186 410 1220
rect 448 1186 482 1220
rect 516 1186 550 1220
rect 588 1186 618 1220
rect 660 1186 686 1220
rect 732 1186 736 1220
rect 149 1113 183 1129
rect 38 1033 72 1045
rect 38 961 72 977
rect 38 889 72 909
rect 38 817 72 841
rect 38 745 72 773
rect 38 673 72 705
rect 38 603 72 637
rect 38 535 72 567
rect 38 467 72 495
rect 38 399 72 423
rect 38 331 72 351
rect 38 263 72 279
rect 38 195 72 207
rect 149 1045 183 1071
rect 149 977 183 999
rect 149 909 183 927
rect 149 841 183 855
rect 149 773 183 783
rect 149 705 183 711
rect 149 637 183 639
rect 149 601 183 603
rect 149 529 183 535
rect 149 457 183 467
rect 149 385 183 399
rect 149 313 183 331
rect 149 241 183 263
rect 149 169 183 195
rect 149 111 183 127
rect 233 1113 339 1129
rect 233 1105 235 1113
rect 337 1105 339 1113
rect 233 127 235 135
rect 337 127 339 135
rect 233 111 339 127
rect 387 1113 493 1129
rect 387 1105 389 1113
rect 491 1105 493 1113
rect 387 127 389 135
rect 491 127 493 135
rect 387 111 493 127
rect 541 1113 647 1129
rect 541 1105 543 1113
rect 645 1105 647 1113
rect 541 127 543 135
rect 645 127 647 135
rect 541 111 647 127
rect 697 1113 731 1129
rect 697 1045 731 1071
rect 697 977 731 999
rect 697 909 731 927
rect 697 841 731 855
rect 697 773 731 783
rect 697 705 731 711
rect 697 637 731 639
rect 697 601 731 603
rect 697 529 731 535
rect 697 457 731 467
rect 697 385 731 399
rect 697 313 731 331
rect 697 241 731 263
rect 697 169 731 195
rect 811 1033 845 1045
rect 811 961 845 977
rect 811 889 845 909
rect 811 817 845 841
rect 811 745 845 773
rect 811 673 845 705
rect 811 603 845 637
rect 811 535 845 567
rect 811 467 845 495
rect 811 399 845 423
rect 811 331 845 351
rect 811 263 845 279
rect 811 195 845 207
rect 697 111 731 127
rect 244 20 266 54
rect 312 20 338 54
rect 380 20 410 54
rect 448 20 482 54
rect 516 20 550 54
rect 588 20 618 54
rect 660 20 686 54
rect 732 20 736 54
<< viali >>
rect 194 1186 210 1220
rect 210 1186 228 1220
rect 266 1186 278 1220
rect 278 1186 300 1220
rect 338 1186 346 1220
rect 346 1186 372 1220
rect 410 1186 414 1220
rect 414 1186 444 1220
rect 482 1186 516 1220
rect 554 1186 584 1220
rect 584 1186 588 1220
rect 626 1186 652 1220
rect 652 1186 660 1220
rect 698 1186 720 1220
rect 720 1186 732 1220
rect 38 1079 72 1105
rect 38 1071 72 1079
rect 38 1011 72 1033
rect 38 999 72 1011
rect 38 943 72 961
rect 38 927 72 943
rect 38 875 72 889
rect 38 855 72 875
rect 38 807 72 817
rect 38 783 72 807
rect 38 739 72 745
rect 38 711 72 739
rect 38 671 72 673
rect 38 639 72 671
rect 38 569 72 601
rect 38 567 72 569
rect 38 501 72 529
rect 38 495 72 501
rect 38 433 72 457
rect 38 423 72 433
rect 38 365 72 385
rect 38 351 72 365
rect 38 297 72 313
rect 38 279 72 297
rect 38 229 72 241
rect 38 207 72 229
rect 38 161 72 169
rect 38 135 72 161
rect 149 1079 183 1105
rect 149 1071 183 1079
rect 149 1011 183 1033
rect 149 999 183 1011
rect 149 943 183 961
rect 149 927 183 943
rect 149 875 183 889
rect 149 855 183 875
rect 149 807 183 817
rect 149 783 183 807
rect 149 739 183 745
rect 149 711 183 739
rect 149 671 183 673
rect 149 639 183 671
rect 149 569 183 601
rect 149 567 183 569
rect 149 501 183 529
rect 149 495 183 501
rect 149 433 183 457
rect 149 423 183 433
rect 149 365 183 385
rect 149 351 183 365
rect 149 297 183 313
rect 149 279 183 297
rect 149 229 183 241
rect 149 207 183 229
rect 149 161 183 169
rect 149 135 183 161
rect 233 135 235 1105
rect 235 135 337 1105
rect 337 135 339 1105
rect 387 135 389 1105
rect 389 135 491 1105
rect 491 135 493 1105
rect 541 135 543 1105
rect 543 135 645 1105
rect 645 135 647 1105
rect 697 1079 731 1105
rect 697 1071 731 1079
rect 697 1011 731 1033
rect 697 999 731 1011
rect 697 943 731 961
rect 697 927 731 943
rect 697 875 731 889
rect 697 855 731 875
rect 697 807 731 817
rect 697 783 731 807
rect 697 739 731 745
rect 697 711 731 739
rect 697 671 731 673
rect 697 639 731 671
rect 697 569 731 601
rect 697 567 731 569
rect 697 501 731 529
rect 697 495 731 501
rect 697 433 731 457
rect 697 423 731 433
rect 697 365 731 385
rect 697 351 731 365
rect 697 297 731 313
rect 697 279 731 297
rect 697 229 731 241
rect 697 207 731 229
rect 697 161 731 169
rect 697 135 731 161
rect 811 1079 845 1105
rect 811 1071 845 1079
rect 811 1011 845 1033
rect 811 999 845 1011
rect 811 943 845 961
rect 811 927 845 943
rect 811 875 845 889
rect 811 855 845 875
rect 811 807 845 817
rect 811 783 845 807
rect 811 739 845 745
rect 811 711 845 739
rect 811 671 845 673
rect 811 639 845 671
rect 811 569 845 601
rect 811 567 845 569
rect 811 501 845 529
rect 811 495 845 501
rect 811 433 845 457
rect 811 423 845 433
rect 811 365 845 385
rect 811 351 845 365
rect 811 297 845 313
rect 811 279 845 297
rect 811 229 845 241
rect 811 207 845 229
rect 811 161 845 169
rect 811 135 845 161
rect 194 20 210 54
rect 210 20 228 54
rect 266 20 278 54
rect 278 20 300 54
rect 338 20 346 54
rect 346 20 372 54
rect 410 20 414 54
rect 414 20 444 54
rect 482 20 516 54
rect 554 20 584 54
rect 584 20 588 54
rect 626 20 652 54
rect 652 20 660 54
rect 698 20 720 54
rect 720 20 732 54
<< metal1 >>
rect 182 1220 744 1232
rect 182 1186 194 1220
rect 228 1186 266 1220
rect 300 1186 338 1220
rect 372 1186 410 1220
rect 444 1186 482 1220
rect 516 1186 554 1220
rect 588 1186 626 1220
rect 660 1186 698 1220
rect 732 1186 744 1220
rect 182 1174 744 1186
rect 140 1122 192 1128
rect 26 1105 84 1117
rect 26 1071 38 1105
rect 72 1071 84 1105
rect 26 1033 84 1071
rect 26 999 38 1033
rect 72 999 84 1033
rect 26 961 84 999
rect 26 927 38 961
rect 72 927 84 961
rect 26 889 84 927
rect 26 855 38 889
rect 72 855 84 889
rect 26 817 84 855
rect 26 783 38 817
rect 72 783 84 817
rect 26 745 84 783
rect 26 711 38 745
rect 72 711 84 745
rect 26 673 84 711
rect 26 639 38 673
rect 72 639 84 673
rect 26 601 84 639
rect 26 567 38 601
rect 72 567 84 601
rect 26 529 84 567
rect 26 495 38 529
rect 72 495 84 529
rect 26 457 84 495
rect 26 423 38 457
rect 72 423 84 457
rect 26 385 84 423
rect 26 351 38 385
rect 72 351 84 385
rect 26 313 84 351
rect 26 279 38 313
rect 72 279 84 313
rect 26 241 84 279
rect 26 207 38 241
rect 72 207 84 241
rect 26 169 84 207
rect 26 135 38 169
rect 72 135 84 169
rect 26 123 84 135
rect 382 1123 498 1129
rect 192 1070 195 1117
rect 140 1058 195 1070
rect 192 1006 195 1058
rect 140 999 149 1006
rect 183 999 195 1006
rect 140 994 195 999
rect 192 942 195 994
rect 140 930 149 942
rect 183 930 195 942
rect 192 878 195 930
rect 140 855 149 878
rect 183 855 195 878
rect 140 817 195 855
rect 140 783 149 817
rect 183 783 195 817
rect 140 745 195 783
rect 140 711 149 745
rect 183 711 195 745
rect 140 673 195 711
rect 140 639 149 673
rect 183 639 195 673
rect 140 601 195 639
rect 140 567 149 601
rect 183 567 195 601
rect 140 529 195 567
rect 140 495 149 529
rect 183 495 195 529
rect 140 457 195 495
rect 140 423 149 457
rect 183 423 195 457
rect 140 385 195 423
rect 140 362 149 385
rect 183 362 195 385
rect 192 310 195 362
rect 140 298 149 310
rect 183 298 195 310
rect 192 246 195 298
rect 140 241 195 246
rect 140 234 149 241
rect 183 234 195 241
rect 192 182 195 234
rect 140 170 195 182
rect 192 123 195 170
rect 223 1105 349 1117
rect 223 838 233 1105
rect 339 838 349 1105
rect 223 402 228 838
rect 344 402 349 838
rect 223 135 233 402
rect 339 135 349 402
rect 223 123 349 135
rect 377 879 382 1117
rect 688 1123 740 1129
rect 498 879 503 1117
rect 377 362 387 879
rect 493 362 503 879
rect 377 123 382 362
rect 140 112 192 118
rect 498 123 503 362
rect 531 1105 657 1117
rect 531 838 541 1105
rect 647 838 657 1105
rect 531 402 536 838
rect 652 402 657 838
rect 531 135 541 402
rect 647 135 657 402
rect 531 123 657 135
rect 685 1071 688 1117
rect 740 1071 743 1117
rect 685 1059 743 1071
rect 685 1007 688 1059
rect 740 1007 743 1059
rect 685 999 697 1007
rect 731 999 743 1007
rect 685 995 743 999
rect 685 943 688 995
rect 740 943 743 995
rect 685 931 697 943
rect 731 931 743 943
rect 685 879 688 931
rect 740 879 743 931
rect 685 855 697 879
rect 731 855 743 879
rect 685 817 743 855
rect 685 783 697 817
rect 731 783 743 817
rect 685 745 743 783
rect 685 711 697 745
rect 731 711 743 745
rect 685 673 743 711
rect 685 639 697 673
rect 731 639 743 673
rect 685 601 743 639
rect 685 567 697 601
rect 731 567 743 601
rect 685 529 743 567
rect 685 495 697 529
rect 731 495 743 529
rect 685 457 743 495
rect 685 423 697 457
rect 731 423 743 457
rect 685 385 743 423
rect 685 362 697 385
rect 731 362 743 385
rect 685 310 688 362
rect 740 310 743 362
rect 685 298 697 310
rect 731 298 743 310
rect 685 246 688 298
rect 740 246 743 298
rect 685 241 743 246
rect 685 234 697 241
rect 731 234 743 241
rect 685 182 688 234
rect 740 182 743 234
rect 685 170 743 182
rect 685 123 688 170
rect 382 112 498 118
rect 740 123 743 170
rect 799 1105 857 1117
rect 799 1071 811 1105
rect 845 1071 857 1105
rect 799 1033 857 1071
rect 799 999 811 1033
rect 845 999 857 1033
rect 799 961 857 999
rect 799 927 811 961
rect 845 927 857 961
rect 799 889 857 927
rect 799 855 811 889
rect 845 855 857 889
rect 799 817 857 855
rect 799 783 811 817
rect 845 783 857 817
rect 799 745 857 783
rect 799 711 811 745
rect 845 711 857 745
rect 799 673 857 711
rect 799 639 811 673
rect 845 639 857 673
rect 799 601 857 639
rect 799 567 811 601
rect 845 567 857 601
rect 799 529 857 567
rect 799 495 811 529
rect 845 495 857 529
rect 799 457 857 495
rect 799 423 811 457
rect 845 423 857 457
rect 799 385 857 423
rect 799 351 811 385
rect 845 351 857 385
rect 799 313 857 351
rect 799 279 811 313
rect 845 279 857 313
rect 799 241 857 279
rect 799 207 811 241
rect 845 207 857 241
rect 799 169 857 207
rect 799 135 811 169
rect 845 135 857 169
rect 799 123 857 135
rect 688 112 740 118
rect 182 54 744 66
rect 182 20 194 54
rect 228 20 266 54
rect 300 20 338 54
rect 372 20 410 54
rect 444 20 482 54
rect 516 20 554 54
rect 588 20 626 54
rect 660 20 698 54
rect 732 20 744 54
rect 182 8 744 20
<< via1 >>
rect 140 1105 192 1122
rect 140 1071 149 1105
rect 149 1071 183 1105
rect 183 1071 192 1105
rect 140 1070 192 1071
rect 140 1033 192 1058
rect 140 1006 149 1033
rect 149 1006 183 1033
rect 183 1006 192 1033
rect 140 961 192 994
rect 140 942 149 961
rect 149 942 183 961
rect 183 942 192 961
rect 140 927 149 930
rect 149 927 183 930
rect 183 927 192 930
rect 140 889 192 927
rect 140 878 149 889
rect 149 878 183 889
rect 183 878 192 889
rect 140 351 149 362
rect 149 351 183 362
rect 183 351 192 362
rect 140 313 192 351
rect 140 310 149 313
rect 149 310 183 313
rect 183 310 192 313
rect 140 279 149 298
rect 149 279 183 298
rect 183 279 192 298
rect 140 246 192 279
rect 140 207 149 234
rect 149 207 183 234
rect 183 207 192 234
rect 140 182 192 207
rect 140 169 192 170
rect 140 135 149 169
rect 149 135 183 169
rect 183 135 192 169
rect 140 118 192 135
rect 228 402 233 838
rect 233 402 339 838
rect 339 402 344 838
rect 382 1105 498 1123
rect 382 879 387 1105
rect 387 879 493 1105
rect 493 879 498 1105
rect 382 135 387 362
rect 387 135 493 362
rect 493 135 498 362
rect 382 118 498 135
rect 536 402 541 838
rect 541 402 647 838
rect 647 402 652 838
rect 688 1105 740 1123
rect 688 1071 697 1105
rect 697 1071 731 1105
rect 731 1071 740 1105
rect 688 1033 740 1059
rect 688 1007 697 1033
rect 697 1007 731 1033
rect 731 1007 740 1033
rect 688 961 740 995
rect 688 943 697 961
rect 697 943 731 961
rect 731 943 740 961
rect 688 927 697 931
rect 697 927 731 931
rect 731 927 740 931
rect 688 889 740 927
rect 688 879 697 889
rect 697 879 731 889
rect 731 879 740 889
rect 688 351 697 362
rect 697 351 731 362
rect 731 351 740 362
rect 688 313 740 351
rect 688 310 697 313
rect 697 310 731 313
rect 731 310 740 313
rect 688 279 697 298
rect 697 279 731 298
rect 731 279 740 298
rect 688 246 740 279
rect 688 207 697 234
rect 697 207 731 234
rect 731 207 740 234
rect 688 182 740 207
rect 688 169 740 170
rect 688 135 697 169
rect 697 135 731 169
rect 731 135 740 169
rect 688 118 740 135
<< metal2 >>
rect 0 1123 884 1129
rect 0 1122 382 1123
rect 0 1070 140 1122
rect 192 1070 382 1122
rect 0 1058 382 1070
rect 0 1006 140 1058
rect 192 1006 382 1058
rect 0 994 382 1006
rect 0 942 140 994
rect 192 942 382 994
rect 0 930 382 942
rect 0 878 140 930
rect 192 879 382 930
rect 498 1071 688 1123
rect 740 1071 884 1123
rect 498 1059 884 1071
rect 498 1007 688 1059
rect 740 1007 884 1059
rect 498 995 884 1007
rect 498 943 688 995
rect 740 943 884 995
rect 498 931 884 943
rect 498 879 688 931
rect 740 879 884 931
rect 192 878 884 879
rect 0 872 884 878
rect 0 838 884 844
rect 0 402 228 838
rect 344 402 536 838
rect 652 402 884 838
rect 0 396 884 402
rect 0 362 884 368
rect 0 310 140 362
rect 192 310 382 362
rect 0 298 382 310
rect 0 246 140 298
rect 192 246 382 298
rect 0 234 382 246
rect 0 182 140 234
rect 192 182 382 234
rect 0 170 382 182
rect 0 118 140 170
rect 192 118 382 170
rect 498 310 688 362
rect 740 310 884 362
rect 498 298 884 310
rect 498 246 688 298
rect 740 246 884 298
rect 498 234 884 246
rect 498 182 688 234
rect 740 182 884 234
rect 498 170 884 182
rect 498 118 688 170
rect 740 118 884 170
rect 0 112 884 118
<< labels >>
flabel comment s 737 655 737 655 0 FreeSans 300 0 0 0 S
flabel comment s 278 655 278 655 0 FreeSans 300 0 0 0 D
flabel comment s 586 655 586 655 0 FreeSans 300 0 0 0 D
flabel comment s 432 655 432 655 0 FreeSans 300 0 0 0 S
flabel comment s 158 655 158 655 0 FreeSans 300 180 0 0 S
flabel metal1 s 414 24 500 49 0 FreeSans 200 180 0 0 GATE
port 2 nsew
flabel metal2 s 0 1089 76 1114 0 FreeSans 200 0 0 0 SOURCE
port 5 nsew
flabel metal2 s 233 618 309 643 0 FreeSans 200 0 0 0 DRAIN
port 7 nsew
flabel metal1 s 39 594 74 674 0 FreeSans 400 90 0 0 SUBSTRATE
port 8 nsew
<< properties >>
string GDS_END 6758292
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 6728788
<< end >>
