magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< poly >>
rect -50 50 0 66
rect -50 16 -34 50
rect -50 0 0 16
rect 3127 50 3177 66
rect 3161 16 3177 50
rect 3127 0 3177 16
<< polycont >>
rect -34 16 0 50
rect 3127 16 3161 50
<< npolyres >>
rect 0 0 3127 66
<< locali >>
rect -34 50 0 66
rect -34 0 0 16
rect 3127 50 3161 66
rect 3127 0 3161 16
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_0
timestamp 1704896540
transform -1 0 16 0 1 0
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_1
timestamp 1704896540
transform 1 0 3111 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 6696272
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 6695838
<< end >>
