magic
tech sky130B
magscale 1 2
timestamp 1704896540
use sky130_fd_pr__dfm1sd__example_55959141808258  sky130_fd_pr__dfm1sd__example_55959141808258_0
timestamp 1704896540
transform 1 0 100 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 22091008
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 22090236
<< end >>
