magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< dnwell >>
rect -67 8739 1796 10364
<< nwell >>
rect 1516 9019 1876 10249
rect -147 8659 1876 9019
rect 1260 446 2609 616
rect 1260 170 1447 446
rect 2415 170 2609 446
rect 1260 0 2609 170
<< pwell >>
rect 1368 9167 1456 10398
rect -93 9079 1456 9167
<< nsubdiff >>
rect 1327 548 2573 549
rect 1327 515 1400 548
rect 1327 481 1328 515
rect 1362 514 1400 515
rect 1434 514 1468 548
rect 1502 514 1536 548
rect 1570 514 1604 548
rect 1638 514 1672 548
rect 1706 514 1740 548
rect 1774 514 1808 548
rect 1842 514 1876 548
rect 1910 514 1944 548
rect 1978 514 2012 548
rect 2046 514 2080 548
rect 2114 514 2148 548
rect 2182 514 2216 548
rect 2250 514 2284 548
rect 2318 514 2352 548
rect 2386 514 2420 548
rect 2454 514 2488 548
rect 2522 514 2573 548
rect 1362 513 2573 514
rect 1362 481 1363 513
rect 1327 447 1363 481
rect 1327 413 1328 447
rect 1362 413 1363 447
rect 1327 379 1363 413
rect 2537 478 2573 513
rect 2537 444 2538 478
rect 2572 444 2573 478
rect 2537 410 2573 444
rect 1327 345 1328 379
rect 1362 345 1363 379
rect 1327 311 1363 345
rect 1327 277 1328 311
rect 1362 277 1363 311
rect 1327 243 1363 277
rect 1327 209 1328 243
rect 1362 209 1363 243
rect 2537 376 2538 410
rect 2572 376 2573 410
rect 2537 342 2573 376
rect 2537 308 2538 342
rect 2572 308 2573 342
rect 2537 274 2573 308
rect 2537 240 2538 274
rect 2572 240 2573 274
rect 1327 103 1363 209
rect 2537 206 2573 240
rect 2537 172 2538 206
rect 2572 172 2573 206
rect 2537 138 2573 172
rect 2537 104 2538 138
rect 2572 104 2573 138
rect 2537 103 2573 104
rect 1327 102 2573 103
rect 1327 68 1361 102
rect 1395 68 1429 102
rect 1463 68 1497 102
rect 1531 68 1565 102
rect 1599 68 1633 102
rect 1667 68 1701 102
rect 1735 68 1769 102
rect 1803 68 1837 102
rect 1871 68 1905 102
rect 1939 68 1973 102
rect 2007 68 2041 102
rect 2075 68 2109 102
rect 2143 68 2177 102
rect 2211 68 2245 102
rect 2279 68 2313 102
rect 2347 68 2401 102
rect 2435 68 2469 102
rect 2503 68 2573 102
rect 1327 67 2573 68
<< mvpsubdiff >>
rect 1394 10329 1430 10372
rect 1394 10295 1395 10329
rect 1429 10295 1430 10329
rect 1394 10261 1430 10295
rect 1394 10227 1395 10261
rect 1429 10227 1430 10261
rect 1394 10193 1430 10227
rect 1394 10159 1395 10193
rect 1429 10159 1430 10193
rect 1394 10125 1430 10159
rect 1394 10091 1395 10125
rect 1429 10091 1430 10125
rect 1394 10057 1430 10091
rect 1394 10023 1395 10057
rect 1429 10023 1430 10057
rect 1394 9989 1430 10023
rect 1394 9955 1395 9989
rect 1429 9955 1430 9989
rect 1394 9921 1430 9955
rect 1394 9887 1395 9921
rect 1429 9887 1430 9921
rect 1394 9853 1430 9887
rect 1394 9819 1395 9853
rect 1429 9819 1430 9853
rect 1394 9785 1430 9819
rect 1394 9751 1395 9785
rect 1429 9751 1430 9785
rect 1394 9717 1430 9751
rect 1394 9683 1395 9717
rect 1429 9683 1430 9717
rect 1394 9649 1430 9683
rect 1394 9615 1395 9649
rect 1429 9615 1430 9649
rect 1394 9581 1430 9615
rect 1394 9547 1395 9581
rect 1429 9547 1430 9581
rect 1394 9513 1430 9547
rect 1394 9479 1395 9513
rect 1429 9479 1430 9513
rect 1394 9445 1430 9479
rect 1394 9411 1395 9445
rect 1429 9411 1430 9445
rect 1394 9377 1430 9411
rect 1394 9343 1395 9377
rect 1429 9343 1430 9377
rect 1394 9309 1430 9343
rect 1394 9275 1395 9309
rect 1429 9275 1430 9309
rect 1394 9241 1430 9275
rect 1394 9207 1395 9241
rect 1429 9207 1430 9241
rect 1394 9173 1430 9207
rect 1394 9141 1395 9173
rect -67 9140 1395 9141
rect -67 9106 -33 9140
rect 1 9106 35 9140
rect 69 9106 103 9140
rect 137 9106 171 9140
rect 205 9106 239 9140
rect 273 9106 307 9140
rect 341 9106 375 9140
rect 409 9106 443 9140
rect 477 9106 511 9140
rect 545 9106 579 9140
rect 613 9106 647 9140
rect 681 9106 715 9140
rect 749 9106 783 9140
rect 817 9106 851 9140
rect 885 9106 919 9140
rect 953 9106 987 9140
rect 1021 9106 1055 9140
rect 1089 9106 1123 9140
rect 1157 9106 1191 9140
rect 1225 9106 1259 9140
rect 1293 9106 1327 9140
rect 1361 9139 1395 9140
rect 1429 9139 1430 9173
rect 1361 9106 1430 9139
rect -67 9105 1430 9106
<< mvnsubdiff >>
rect 1583 10140 1619 10183
rect 1583 10106 1584 10140
rect 1618 10106 1619 10140
rect 1583 10072 1619 10106
rect 1583 10038 1584 10072
rect 1618 10038 1619 10072
rect 1583 10004 1619 10038
rect 1583 9970 1584 10004
rect 1618 9970 1619 10004
rect 1583 9936 1619 9970
rect 1583 9902 1584 9936
rect 1618 9902 1619 9936
rect 1583 9868 1619 9902
rect 1583 9834 1584 9868
rect 1618 9834 1619 9868
rect 1583 9800 1619 9834
rect 1583 9766 1584 9800
rect 1618 9766 1619 9800
rect 1583 9732 1619 9766
rect 1583 9698 1584 9732
rect 1618 9698 1619 9732
rect 1583 9664 1619 9698
rect 1583 9630 1584 9664
rect 1618 9630 1619 9664
rect 1583 9596 1619 9630
rect 1583 9562 1584 9596
rect 1618 9562 1619 9596
rect 1583 9528 1619 9562
rect 1583 9494 1584 9528
rect 1618 9494 1619 9528
rect 1583 9460 1619 9494
rect 1583 9426 1584 9460
rect 1618 9426 1619 9460
rect 1583 9392 1619 9426
rect 1583 9358 1584 9392
rect 1618 9358 1619 9392
rect 1583 9324 1619 9358
rect 1583 9290 1584 9324
rect 1618 9290 1619 9324
rect 1583 9256 1619 9290
rect 1583 9222 1584 9256
rect 1618 9222 1619 9256
rect 1583 9188 1619 9222
rect 1583 9154 1584 9188
rect 1618 9154 1619 9188
rect 1583 9120 1619 9154
rect 1583 9086 1584 9120
rect 1618 9086 1619 9120
rect 1583 9052 1619 9086
rect 1583 9018 1584 9052
rect 1618 9018 1619 9052
rect 1583 8984 1619 9018
rect 1583 8952 1584 8984
rect -67 8951 1584 8952
rect -67 8917 -33 8951
rect 1 8917 35 8951
rect 69 8917 103 8951
rect 137 8917 171 8951
rect 205 8917 239 8951
rect 273 8917 307 8951
rect 341 8917 375 8951
rect 409 8917 443 8951
rect 477 8917 511 8951
rect 545 8917 579 8951
rect 613 8917 647 8951
rect 681 8917 715 8951
rect 749 8917 783 8951
rect 817 8917 851 8951
rect 885 8917 919 8951
rect 953 8917 987 8951
rect 1021 8917 1055 8951
rect 1089 8917 1123 8951
rect 1157 8917 1191 8951
rect 1225 8917 1259 8951
rect 1293 8917 1327 8951
rect 1361 8917 1395 8951
rect 1429 8917 1508 8951
rect 1542 8950 1584 8951
rect 1618 8950 1619 8984
rect 1542 8917 1619 8950
rect -67 8916 1619 8917
<< nsubdiffcont >>
rect 1328 481 1362 515
rect 1400 514 1434 548
rect 1468 514 1502 548
rect 1536 514 1570 548
rect 1604 514 1638 548
rect 1672 514 1706 548
rect 1740 514 1774 548
rect 1808 514 1842 548
rect 1876 514 1910 548
rect 1944 514 1978 548
rect 2012 514 2046 548
rect 2080 514 2114 548
rect 2148 514 2182 548
rect 2216 514 2250 548
rect 2284 514 2318 548
rect 2352 514 2386 548
rect 2420 514 2454 548
rect 2488 514 2522 548
rect 1328 413 1362 447
rect 2538 444 2572 478
rect 1328 345 1362 379
rect 1328 277 1362 311
rect 1328 209 1362 243
rect 2538 376 2572 410
rect 2538 308 2572 342
rect 2538 240 2572 274
rect 2538 172 2572 206
rect 2538 104 2572 138
rect 1361 68 1395 102
rect 1429 68 1463 102
rect 1497 68 1531 102
rect 1565 68 1599 102
rect 1633 68 1667 102
rect 1701 68 1735 102
rect 1769 68 1803 102
rect 1837 68 1871 102
rect 1905 68 1939 102
rect 1973 68 2007 102
rect 2041 68 2075 102
rect 2109 68 2143 102
rect 2177 68 2211 102
rect 2245 68 2279 102
rect 2313 68 2347 102
rect 2401 68 2435 102
rect 2469 68 2503 102
<< mvpsubdiffcont >>
rect 1395 10295 1429 10329
rect 1395 10227 1429 10261
rect 1395 10159 1429 10193
rect 1395 10091 1429 10125
rect 1395 10023 1429 10057
rect 1395 9955 1429 9989
rect 1395 9887 1429 9921
rect 1395 9819 1429 9853
rect 1395 9751 1429 9785
rect 1395 9683 1429 9717
rect 1395 9615 1429 9649
rect 1395 9547 1429 9581
rect 1395 9479 1429 9513
rect 1395 9411 1429 9445
rect 1395 9343 1429 9377
rect 1395 9275 1429 9309
rect 1395 9207 1429 9241
rect -33 9106 1 9140
rect 35 9106 69 9140
rect 103 9106 137 9140
rect 171 9106 205 9140
rect 239 9106 273 9140
rect 307 9106 341 9140
rect 375 9106 409 9140
rect 443 9106 477 9140
rect 511 9106 545 9140
rect 579 9106 613 9140
rect 647 9106 681 9140
rect 715 9106 749 9140
rect 783 9106 817 9140
rect 851 9106 885 9140
rect 919 9106 953 9140
rect 987 9106 1021 9140
rect 1055 9106 1089 9140
rect 1123 9106 1157 9140
rect 1191 9106 1225 9140
rect 1259 9106 1293 9140
rect 1327 9106 1361 9140
rect 1395 9139 1429 9173
<< mvnsubdiffcont >>
rect 1584 10106 1618 10140
rect 1584 10038 1618 10072
rect 1584 9970 1618 10004
rect 1584 9902 1618 9936
rect 1584 9834 1618 9868
rect 1584 9766 1618 9800
rect 1584 9698 1618 9732
rect 1584 9630 1618 9664
rect 1584 9562 1618 9596
rect 1584 9494 1618 9528
rect 1584 9426 1618 9460
rect 1584 9358 1618 9392
rect 1584 9290 1618 9324
rect 1584 9222 1618 9256
rect 1584 9154 1618 9188
rect 1584 9086 1618 9120
rect 1584 9018 1618 9052
rect -33 8917 1 8951
rect 35 8917 69 8951
rect 103 8917 137 8951
rect 171 8917 205 8951
rect 239 8917 273 8951
rect 307 8917 341 8951
rect 375 8917 409 8951
rect 443 8917 477 8951
rect 511 8917 545 8951
rect 579 8917 613 8951
rect 647 8917 681 8951
rect 715 8917 749 8951
rect 783 8917 817 8951
rect 851 8917 885 8951
rect 919 8917 953 8951
rect 987 8917 1021 8951
rect 1055 8917 1089 8951
rect 1123 8917 1157 8951
rect 1191 8917 1225 8951
rect 1259 8917 1293 8951
rect 1327 8917 1361 8951
rect 1395 8917 1429 8951
rect 1508 8917 1542 8951
rect 1584 8950 1618 8984
<< poly >>
rect 1964 12487 4298 12553
rect -399 10322 -199 10338
rect -399 10288 -350 10322
rect -316 10288 -282 10322
rect -248 10288 -199 10322
rect -399 10272 -199 10288
rect -143 10322 57 10338
rect -143 10288 -94 10322
rect -60 10288 -26 10322
rect 8 10288 57 10322
rect -143 10272 57 10288
rect 113 10322 313 10338
rect 113 10288 162 10322
rect 196 10288 230 10322
rect 264 10288 313 10322
rect 113 10272 313 10288
rect 369 10322 569 10338
rect 369 10288 418 10322
rect 452 10288 486 10322
rect 520 10288 569 10322
rect 369 10272 569 10288
rect 625 10322 825 10338
rect 625 10288 674 10322
rect 708 10288 742 10322
rect 776 10288 825 10322
rect 625 10272 825 10288
rect 881 10322 1081 10338
rect 881 10288 930 10322
rect 964 10288 998 10322
rect 1032 10288 1081 10322
rect 881 10272 1081 10288
rect 1137 10322 1271 10338
rect 1137 10288 1153 10322
rect 1187 10288 1221 10322
rect 1255 10288 1271 10322
rect 1137 10272 1271 10288
rect 1964 8715 2030 12487
rect 2126 12375 2192 12391
rect 2126 12341 2142 12375
rect 2176 12341 2192 12375
rect 2126 12323 2192 12341
rect 2288 12375 2354 12391
rect 2288 12341 2304 12375
rect 2338 12341 2354 12375
rect 2288 12323 2354 12341
rect 2450 12375 2516 12391
rect 2450 12341 2466 12375
rect 2500 12341 2516 12375
rect 2450 12323 2516 12341
rect 2612 12375 2678 12391
rect 2612 12341 2628 12375
rect 2662 12341 2678 12375
rect 2612 12323 2678 12341
rect 2774 12375 2840 12391
rect 2774 12341 2790 12375
rect 2824 12341 2840 12375
rect 2774 12323 2840 12341
rect 2936 12375 3002 12391
rect 2936 12341 2952 12375
rect 2986 12341 3002 12375
rect 2936 12323 3002 12341
rect 3098 12375 3164 12391
rect 3098 12341 3114 12375
rect 3148 12341 3164 12375
rect 3098 12323 3164 12341
rect 3260 12375 3326 12391
rect 3260 12341 3276 12375
rect 3310 12341 3326 12375
rect 3260 12323 3326 12341
rect 3422 12375 3488 12391
rect 3422 12341 3438 12375
rect 3472 12341 3488 12375
rect 3422 12323 3488 12341
rect 3584 12375 3650 12391
rect 3584 12341 3600 12375
rect 3634 12341 3650 12375
rect 3584 12323 3650 12341
rect 3746 12375 3812 12391
rect 3746 12341 3762 12375
rect 3796 12341 3812 12375
rect 3746 12323 3812 12341
rect 3908 12375 3974 12391
rect 3908 12341 3924 12375
rect 3958 12341 3974 12375
rect 3908 12323 3974 12341
rect 4070 12375 4136 12391
rect 4070 12341 4086 12375
rect 4120 12341 4136 12375
rect 4070 12323 4136 12341
rect 182 8649 2030 8715
rect 182 647 248 8649
rect 344 8537 410 8553
rect 344 8503 360 8537
rect 394 8503 410 8537
rect 344 8469 410 8503
rect 344 8435 360 8469
rect 394 8435 410 8469
rect 344 8419 410 8435
rect 506 8537 572 8553
rect 506 8503 522 8537
rect 556 8503 572 8537
rect 506 8469 572 8503
rect 506 8435 522 8469
rect 556 8435 572 8469
rect 506 8419 572 8435
rect 668 8537 734 8553
rect 668 8503 684 8537
rect 718 8503 734 8537
rect 668 8469 734 8503
rect 668 8435 684 8469
rect 718 8435 734 8469
rect 668 8419 734 8435
rect 830 8537 896 8553
rect 830 8503 846 8537
rect 880 8503 896 8537
rect 830 8469 896 8503
rect 830 8435 846 8469
rect 880 8435 896 8469
rect 830 8419 896 8435
rect 992 8537 1058 8553
rect 992 8503 1008 8537
rect 1042 8503 1058 8537
rect 992 8469 1058 8503
rect 992 8435 1008 8469
rect 1042 8435 1058 8469
rect 992 8419 1058 8435
rect 1154 8537 1220 8553
rect 1154 8503 1170 8537
rect 1204 8503 1220 8537
rect 1154 8469 1220 8503
rect 1154 8435 1170 8469
rect 1204 8435 1220 8469
rect 1154 8419 1220 8435
rect 1316 8537 1382 8553
rect 1316 8503 1332 8537
rect 1366 8503 1382 8537
rect 1316 8469 1382 8503
rect 1316 8435 1332 8469
rect 1366 8435 1382 8469
rect 1316 8419 1382 8435
rect 1478 8537 1544 8553
rect 1478 8503 1494 8537
rect 1528 8503 1544 8537
rect 1478 8469 1544 8503
rect 1478 8435 1494 8469
rect 1528 8435 1544 8469
rect 1478 8419 1544 8435
rect 1640 8537 1706 8553
rect 1640 8503 1656 8537
rect 1690 8503 1706 8537
rect 1640 8469 1706 8503
rect 1640 8435 1656 8469
rect 1690 8435 1706 8469
rect 1640 8419 1706 8435
rect 1802 8537 1868 8553
rect 1802 8503 1818 8537
rect 1852 8503 1868 8537
rect 1802 8469 1868 8503
rect 1802 8435 1818 8469
rect 1852 8435 1868 8469
rect 1802 8419 1868 8435
rect 1964 8537 2030 8553
rect 1964 8503 1980 8537
rect 2014 8503 2030 8537
rect 1964 8469 2030 8503
rect 1964 8435 1980 8469
rect 2014 8435 2030 8469
rect 1964 8419 2030 8435
rect 2126 8537 2192 8553
rect 2126 8503 2142 8537
rect 2176 8503 2192 8537
rect 2126 8469 2192 8503
rect 2126 8435 2142 8469
rect 2176 8435 2192 8469
rect 2126 8419 2192 8435
rect 2288 8537 2354 8553
rect 2288 8503 2304 8537
rect 2338 8503 2354 8537
rect 2288 8469 2354 8503
rect 2288 8435 2304 8469
rect 2338 8435 2354 8469
rect 2288 8419 2354 8435
rect 2450 8537 2516 8553
rect 2450 8503 2466 8537
rect 2500 8503 2516 8537
rect 2450 8469 2516 8503
rect 2450 8435 2466 8469
rect 2500 8435 2516 8469
rect 2450 8419 2516 8435
rect 2612 8537 2678 8553
rect 2612 8503 2628 8537
rect 2662 8503 2678 8537
rect 2612 8469 2678 8503
rect 2612 8435 2628 8469
rect 2662 8435 2678 8469
rect 2612 8419 2678 8435
rect 2774 8537 2840 8553
rect 2774 8503 2790 8537
rect 2824 8503 2840 8537
rect 2774 8469 2840 8503
rect 2774 8435 2790 8469
rect 2824 8435 2840 8469
rect 2774 8419 2840 8435
rect 2936 8537 3002 8553
rect 2936 8503 2952 8537
rect 2986 8503 3002 8537
rect 2936 8469 3002 8503
rect 2936 8435 2952 8469
rect 2986 8435 3002 8469
rect 2936 8419 3002 8435
rect 3098 8537 3164 8553
rect 3098 8503 3114 8537
rect 3148 8503 3164 8537
rect 3098 8469 3164 8503
rect 3098 8435 3114 8469
rect 3148 8435 3164 8469
rect 3098 8419 3164 8435
rect 3260 8537 3326 8553
rect 3260 8503 3276 8537
rect 3310 8503 3326 8537
rect 3260 8469 3326 8503
rect 3422 8485 3488 8487
rect 3584 8485 3650 8487
rect 3746 8485 3812 8487
rect 3908 8485 3974 8487
rect 4070 8485 4136 8487
rect 3260 8435 3276 8469
rect 3310 8435 3326 8469
rect 3260 8419 3326 8435
rect 344 4647 410 4649
rect 506 4647 572 4649
rect 668 4647 734 4649
rect 830 4647 896 4649
rect 992 4647 1058 4649
rect 1154 4647 1220 4649
rect 1316 4647 1382 4649
rect 1478 4647 1544 4649
rect 1640 4647 1706 4649
rect 1802 4647 1868 4649
rect 1964 4647 2030 4649
rect 2126 4647 2192 4649
rect 2288 4647 2354 4649
rect 2450 4647 2516 4649
rect 2612 4647 2678 4649
rect 2774 4647 2840 4649
rect 2936 4647 3002 4649
rect 3098 4647 3164 4649
rect 3260 4647 3326 4649
rect 3422 4647 3488 4649
rect 3584 4647 3650 4649
rect 3746 4647 3812 4649
rect 3908 4647 3974 4649
rect 4070 4647 4136 4649
rect 344 793 410 811
rect 344 759 360 793
rect 394 759 410 793
rect 344 743 410 759
rect 506 793 572 811
rect 506 759 522 793
rect 556 759 572 793
rect 506 743 572 759
rect 668 793 734 811
rect 668 759 684 793
rect 718 759 734 793
rect 668 743 734 759
rect 830 793 896 811
rect 830 759 846 793
rect 880 759 896 793
rect 830 743 896 759
rect 992 793 1058 811
rect 992 759 1008 793
rect 1042 759 1058 793
rect 992 743 1058 759
rect 1154 793 1220 811
rect 1154 759 1170 793
rect 1204 759 1220 793
rect 1154 743 1220 759
rect 1316 793 1382 811
rect 1316 759 1332 793
rect 1366 759 1382 793
rect 1316 743 1382 759
rect 1478 793 1544 811
rect 1478 759 1494 793
rect 1528 759 1544 793
rect 1478 743 1544 759
rect 1640 793 1706 811
rect 1640 759 1656 793
rect 1690 759 1706 793
rect 1640 743 1706 759
rect 1802 793 1868 811
rect 1802 759 1818 793
rect 1852 759 1868 793
rect 1802 743 1868 759
rect 1964 793 2030 811
rect 1964 759 1980 793
rect 2014 759 2030 793
rect 1964 743 2030 759
rect 2126 793 2192 811
rect 2126 759 2142 793
rect 2176 759 2192 793
rect 2126 743 2192 759
rect 2288 793 2354 811
rect 2288 759 2304 793
rect 2338 759 2354 793
rect 2288 743 2354 759
rect 2450 793 2516 811
rect 2450 759 2466 793
rect 2500 759 2516 793
rect 2450 743 2516 759
rect 2612 793 2678 811
rect 2612 759 2628 793
rect 2662 759 2678 793
rect 2612 743 2678 759
rect 2774 793 2840 811
rect 2774 759 2790 793
rect 2824 759 2840 793
rect 2774 743 2840 759
rect 2936 793 3002 811
rect 2936 759 2952 793
rect 2986 759 3002 793
rect 2936 743 3002 759
rect 3098 793 3164 811
rect 3098 759 3114 793
rect 3148 759 3164 793
rect 3098 743 3164 759
rect 3260 793 3326 811
rect 3260 759 3276 793
rect 3310 759 3326 793
rect 3260 743 3326 759
rect 3422 793 3488 811
rect 3422 759 3438 793
rect 3472 759 3488 793
rect 3422 743 3488 759
rect 3584 793 3650 811
rect 3584 759 3600 793
rect 3634 759 3650 793
rect 3584 743 3650 759
rect 3746 793 3812 811
rect 3746 759 3762 793
rect 3796 759 3812 793
rect 3746 743 3812 759
rect 3908 793 3974 811
rect 3908 759 3924 793
rect 3958 759 3974 793
rect 3908 743 3974 759
rect 4070 793 4136 811
rect 4070 759 4086 793
rect 4120 759 4136 793
rect 4070 743 4136 759
rect 4232 647 4298 12487
rect 182 581 4298 647
rect 1385 359 1457 386
rect 1385 325 1401 359
rect 1435 336 1457 359
rect 1435 325 1451 336
rect 1385 291 1451 325
rect 1385 257 1401 291
rect 1435 280 1451 291
rect 1435 257 1457 280
rect 1385 230 1457 257
<< polycont >>
rect -350 10288 -316 10322
rect -282 10288 -248 10322
rect -94 10288 -60 10322
rect -26 10288 8 10322
rect 162 10288 196 10322
rect 230 10288 264 10322
rect 418 10288 452 10322
rect 486 10288 520 10322
rect 674 10288 708 10322
rect 742 10288 776 10322
rect 930 10288 964 10322
rect 998 10288 1032 10322
rect 1153 10288 1187 10322
rect 1221 10288 1255 10322
rect 2142 12341 2176 12375
rect 2304 12341 2338 12375
rect 2466 12341 2500 12375
rect 2628 12341 2662 12375
rect 2790 12341 2824 12375
rect 2952 12341 2986 12375
rect 3114 12341 3148 12375
rect 3276 12341 3310 12375
rect 3438 12341 3472 12375
rect 3600 12341 3634 12375
rect 3762 12341 3796 12375
rect 3924 12341 3958 12375
rect 4086 12341 4120 12375
rect 360 8503 394 8537
rect 360 8435 394 8469
rect 522 8503 556 8537
rect 522 8435 556 8469
rect 684 8503 718 8537
rect 684 8435 718 8469
rect 846 8503 880 8537
rect 846 8435 880 8469
rect 1008 8503 1042 8537
rect 1008 8435 1042 8469
rect 1170 8503 1204 8537
rect 1170 8435 1204 8469
rect 1332 8503 1366 8537
rect 1332 8435 1366 8469
rect 1494 8503 1528 8537
rect 1494 8435 1528 8469
rect 1656 8503 1690 8537
rect 1656 8435 1690 8469
rect 1818 8503 1852 8537
rect 1818 8435 1852 8469
rect 1980 8503 2014 8537
rect 1980 8435 2014 8469
rect 2142 8503 2176 8537
rect 2142 8435 2176 8469
rect 2304 8503 2338 8537
rect 2304 8435 2338 8469
rect 2466 8503 2500 8537
rect 2466 8435 2500 8469
rect 2628 8503 2662 8537
rect 2628 8435 2662 8469
rect 2790 8503 2824 8537
rect 2790 8435 2824 8469
rect 2952 8503 2986 8537
rect 2952 8435 2986 8469
rect 3114 8503 3148 8537
rect 3114 8435 3148 8469
rect 3276 8503 3310 8537
rect 3276 8435 3310 8469
rect 360 759 394 793
rect 522 759 556 793
rect 684 759 718 793
rect 846 759 880 793
rect 1008 759 1042 793
rect 1170 759 1204 793
rect 1332 759 1366 793
rect 1494 759 1528 793
rect 1656 759 1690 793
rect 1818 759 1852 793
rect 1980 759 2014 793
rect 2142 759 2176 793
rect 2304 759 2338 793
rect 2466 759 2500 793
rect 2628 759 2662 793
rect 2790 759 2824 793
rect 2952 759 2986 793
rect 3114 759 3148 793
rect 3276 759 3310 793
rect 3438 759 3472 793
rect 3600 759 3634 793
rect 3762 759 3796 793
rect 3924 759 3958 793
rect 4086 759 4120 793
rect 1401 325 1435 359
rect 1401 257 1435 291
<< locali >>
rect 1980 12502 2044 12537
rect 4218 12502 4282 12537
rect 1980 12470 2014 12502
rect 4248 12482 4282 12502
rect 2126 12377 2192 12389
rect 2126 12341 2142 12377
rect 2176 12341 2192 12377
rect 2126 12305 2192 12341
rect 2126 12271 2142 12305
rect 2176 12271 2192 12305
rect 2126 12259 2192 12271
rect 2288 12377 2354 12389
rect 2288 12341 2304 12377
rect 2338 12341 2354 12377
rect 2288 12305 2354 12341
rect 2288 12271 2304 12305
rect 2338 12271 2354 12305
rect 2288 12259 2354 12271
rect 2450 12377 2516 12389
rect 2450 12341 2466 12377
rect 2500 12341 2516 12377
rect 2450 12305 2516 12341
rect 2450 12271 2466 12305
rect 2500 12271 2516 12305
rect 2450 12259 2516 12271
rect 2612 12377 2678 12389
rect 2612 12341 2628 12377
rect 2662 12341 2678 12377
rect 2612 12305 2678 12341
rect 2612 12271 2628 12305
rect 2662 12271 2678 12305
rect 2612 12259 2678 12271
rect 2774 12377 2840 12389
rect 2774 12341 2790 12377
rect 2824 12341 2840 12377
rect 2774 12305 2840 12341
rect 2774 12271 2790 12305
rect 2824 12271 2840 12305
rect 2774 12259 2840 12271
rect 2936 12377 3002 12389
rect 2936 12341 2952 12377
rect 2986 12341 3002 12377
rect 2936 12305 3002 12341
rect 2936 12271 2952 12305
rect 2986 12271 3002 12305
rect 2936 12259 3002 12271
rect 3098 12377 3164 12389
rect 3098 12341 3114 12377
rect 3148 12341 3164 12377
rect 3098 12305 3164 12341
rect 3098 12271 3114 12305
rect 3148 12271 3164 12305
rect 3098 12259 3164 12271
rect 3260 12377 3326 12389
rect 3260 12341 3276 12377
rect 3310 12341 3326 12377
rect 3260 12305 3326 12341
rect 3260 12271 3276 12305
rect 3310 12271 3326 12305
rect 3260 12259 3326 12271
rect 3422 12377 3488 12389
rect 3422 12341 3438 12377
rect 3472 12341 3488 12377
rect 3422 12305 3488 12341
rect 3422 12271 3438 12305
rect 3472 12271 3488 12305
rect 3422 12259 3488 12271
rect 3584 12377 3650 12389
rect 3584 12341 3600 12377
rect 3634 12341 3650 12377
rect 3584 12305 3650 12341
rect 3584 12271 3600 12305
rect 3634 12271 3650 12305
rect 3584 12259 3650 12271
rect 3746 12377 3812 12389
rect 3746 12341 3762 12377
rect 3796 12341 3812 12377
rect 3746 12305 3812 12341
rect 3746 12271 3762 12305
rect 3796 12271 3812 12305
rect 3746 12259 3812 12271
rect 3908 12377 3974 12389
rect 3908 12341 3924 12377
rect 3958 12341 3974 12377
rect 3908 12305 3974 12341
rect 3908 12271 3924 12305
rect 3958 12271 3974 12305
rect 3908 12259 3974 12271
rect 4070 12377 4136 12389
rect 4070 12341 4086 12377
rect 4120 12341 4136 12377
rect 4070 12305 4136 12341
rect 4070 12271 4086 12305
rect 4120 12271 4136 12305
rect 4070 12259 4136 12271
rect 1394 10329 1430 10372
rect -366 10288 -350 10322
rect -316 10288 -282 10322
rect -248 10288 -232 10322
rect -110 10288 -94 10322
rect -60 10288 -26 10322
rect 8 10288 24 10322
rect 146 10288 162 10322
rect 196 10288 230 10322
rect 264 10288 280 10322
rect 402 10288 418 10322
rect 452 10288 486 10322
rect 520 10288 536 10322
rect 658 10288 674 10322
rect 708 10288 742 10322
rect 776 10288 792 10322
rect 914 10288 930 10322
rect 964 10288 998 10322
rect 1032 10288 1048 10322
rect 1137 10288 1153 10322
rect 1187 10288 1221 10322
rect 1255 10288 1356 10322
rect 1322 10242 1356 10288
rect 1322 10170 1356 10208
rect 1394 10295 1395 10329
rect 1429 10295 1430 10329
rect 1394 10261 1430 10295
rect 1394 10227 1395 10261
rect 1429 10227 1430 10261
rect 1394 10193 1430 10227
rect 1394 10159 1395 10193
rect 1429 10159 1430 10193
rect 1394 10125 1430 10159
rect 1394 10091 1395 10125
rect 1429 10091 1430 10125
rect 1394 10057 1430 10091
rect 1394 10023 1395 10057
rect 1429 10023 1430 10057
rect 1394 9989 1430 10023
rect 1394 9955 1395 9989
rect 1429 9955 1430 9989
rect 1394 9921 1430 9955
rect 1394 9887 1395 9921
rect 1429 9887 1430 9921
rect 1394 9853 1430 9887
rect 1394 9819 1395 9853
rect 1429 9819 1430 9853
rect 1394 9785 1430 9819
rect 1394 9751 1395 9785
rect 1429 9751 1430 9785
rect 1394 9717 1430 9751
rect 1394 9683 1395 9717
rect 1429 9683 1430 9717
rect 1394 9649 1430 9683
rect 1394 9615 1395 9649
rect 1429 9615 1430 9649
rect 1394 9581 1430 9615
rect 1394 9547 1395 9581
rect 1429 9547 1430 9581
rect 1394 9513 1430 9547
rect 1394 9479 1395 9513
rect 1429 9479 1430 9513
rect 1394 9445 1430 9479
rect 1394 9411 1395 9445
rect 1429 9411 1430 9445
rect 1394 9377 1430 9411
rect 1394 9343 1395 9377
rect 1429 9343 1430 9377
rect 1394 9309 1430 9343
rect 1394 9275 1395 9309
rect 1429 9275 1430 9309
rect 1394 9241 1430 9275
rect 1394 9207 1395 9241
rect 1429 9207 1430 9241
rect 1394 9173 1430 9207
rect 1394 9141 1395 9173
rect -67 9140 1395 9141
rect -67 9106 -33 9140
rect 1 9106 35 9140
rect 69 9106 103 9140
rect 137 9106 171 9140
rect 205 9106 239 9140
rect 273 9106 307 9140
rect 341 9106 375 9140
rect 409 9106 443 9140
rect 477 9106 511 9140
rect 545 9106 579 9140
rect 613 9106 647 9140
rect 681 9106 715 9140
rect 749 9106 783 9140
rect 817 9106 851 9140
rect 885 9106 919 9140
rect 953 9106 987 9140
rect 1021 9106 1055 9140
rect 1089 9106 1123 9140
rect 1157 9106 1191 9140
rect 1225 9106 1259 9140
rect 1293 9106 1327 9140
rect 1361 9139 1395 9140
rect 1429 9139 1430 9173
rect 1361 9106 1430 9139
rect -67 9105 1430 9106
rect 1583 10140 1631 10183
rect 1583 10106 1584 10140
rect 1618 10106 1631 10140
rect 1583 10072 1631 10106
rect 1583 10038 1584 10072
rect 1618 10038 1631 10072
rect 1583 10004 1631 10038
rect 1583 9970 1584 10004
rect 1618 9970 1631 10004
rect 1583 9936 1631 9970
rect 1583 9902 1584 9936
rect 1618 9902 1631 9936
rect 1583 9868 1631 9902
rect 1583 9834 1584 9868
rect 1618 9834 1631 9868
rect 1583 9800 1631 9834
rect 1583 9766 1584 9800
rect 1618 9766 1631 9800
rect 1583 9732 1631 9766
rect 1583 9698 1584 9732
rect 1618 9698 1631 9732
rect 1583 9664 1631 9698
rect 1583 9630 1584 9664
rect 1618 9630 1631 9664
rect 1583 9596 1631 9630
rect 1583 9562 1584 9596
rect 1618 9562 1631 9596
rect 1583 9528 1631 9562
rect 1583 9494 1584 9528
rect 1618 9494 1631 9528
rect 1583 9460 1631 9494
rect 1583 9426 1584 9460
rect 1618 9426 1631 9460
rect 1583 9392 1631 9426
rect 1583 9358 1584 9392
rect 1618 9358 1631 9392
rect 1583 9324 1631 9358
rect 1583 9290 1584 9324
rect 1618 9290 1631 9324
rect 1583 9256 1631 9290
rect 1583 9222 1584 9256
rect 1618 9222 1631 9256
rect 1583 9188 1631 9222
rect 1583 9154 1584 9188
rect 1618 9154 1631 9188
rect 1583 9120 1631 9154
rect 1583 9086 1584 9120
rect 1618 9086 1631 9120
rect 1583 9052 1631 9086
rect 1583 9018 1584 9052
rect 1618 9018 1631 9052
rect 1583 8984 1631 9018
rect 1583 8952 1584 8984
rect -67 8951 1584 8952
rect -67 8917 -42 8951
rect 1 8917 30 8951
rect 69 8917 102 8951
rect 137 8917 171 8951
rect 208 8917 239 8951
rect 280 8917 307 8951
rect 341 8917 375 8951
rect 409 8917 443 8951
rect 477 8917 511 8951
rect 545 8917 579 8951
rect 613 8917 647 8951
rect 681 8917 715 8951
rect 749 8917 783 8951
rect 817 8917 851 8951
rect 885 8917 919 8951
rect 953 8917 987 8951
rect 1021 8917 1055 8951
rect 1089 8917 1123 8951
rect 1157 8917 1191 8951
rect 1225 8917 1259 8951
rect 1293 8917 1327 8951
rect 1361 8917 1395 8951
rect 1429 8917 1508 8951
rect 1542 8950 1584 8951
rect 1618 8950 1631 8984
rect 1542 8917 1631 8950
rect -67 8916 1631 8917
rect 1980 8699 2014 8732
rect 198 8665 257 8699
rect 1955 8665 2014 8699
rect 344 8539 410 8551
rect 344 8503 360 8539
rect 394 8503 410 8539
rect 344 8469 410 8503
rect 344 8433 360 8469
rect 394 8433 410 8469
rect 344 8421 410 8433
rect 506 8539 572 8551
rect 506 8503 522 8539
rect 556 8503 572 8539
rect 506 8469 572 8503
rect 506 8433 522 8469
rect 556 8433 572 8469
rect 506 8421 572 8433
rect 668 8539 734 8551
rect 668 8503 684 8539
rect 718 8503 734 8539
rect 668 8469 734 8503
rect 668 8433 684 8469
rect 718 8433 734 8469
rect 668 8421 734 8433
rect 830 8539 896 8551
rect 830 8503 846 8539
rect 880 8503 896 8539
rect 830 8469 896 8503
rect 830 8433 846 8469
rect 880 8433 896 8469
rect 830 8421 896 8433
rect 992 8539 1058 8551
rect 992 8503 1008 8539
rect 1042 8503 1058 8539
rect 992 8469 1058 8503
rect 992 8433 1008 8469
rect 1042 8433 1058 8469
rect 992 8421 1058 8433
rect 1154 8539 1220 8551
rect 1154 8503 1170 8539
rect 1204 8503 1220 8539
rect 1154 8469 1220 8503
rect 1154 8433 1170 8469
rect 1204 8433 1220 8469
rect 1154 8421 1220 8433
rect 1316 8539 1382 8551
rect 1316 8503 1332 8539
rect 1366 8503 1382 8539
rect 1316 8469 1382 8503
rect 1316 8433 1332 8469
rect 1366 8433 1382 8469
rect 1316 8421 1382 8433
rect 1478 8539 1544 8551
rect 1478 8503 1494 8539
rect 1528 8503 1544 8539
rect 1478 8469 1544 8503
rect 1478 8433 1494 8469
rect 1528 8433 1544 8469
rect 1478 8421 1544 8433
rect 1640 8539 1706 8551
rect 1640 8503 1656 8539
rect 1690 8503 1706 8539
rect 1640 8469 1706 8503
rect 1640 8433 1656 8469
rect 1690 8433 1706 8469
rect 1640 8421 1706 8433
rect 1802 8539 1868 8551
rect 1802 8503 1818 8539
rect 1852 8503 1868 8539
rect 1802 8469 1868 8503
rect 1802 8433 1818 8469
rect 1852 8433 1868 8469
rect 1802 8421 1868 8433
rect 1964 8539 2030 8551
rect 1964 8503 1980 8539
rect 2014 8503 2030 8539
rect 1964 8469 2030 8503
rect 1964 8433 1980 8469
rect 2014 8433 2030 8469
rect 1964 8421 2030 8433
rect 2126 8539 2192 8551
rect 2126 8503 2142 8539
rect 2176 8503 2192 8539
rect 2126 8469 2192 8503
rect 2126 8433 2142 8469
rect 2176 8433 2192 8469
rect 2126 8421 2192 8433
rect 2288 8539 2354 8551
rect 2288 8503 2304 8539
rect 2338 8503 2354 8539
rect 2288 8469 2354 8503
rect 2288 8433 2304 8469
rect 2338 8433 2354 8469
rect 2288 8421 2354 8433
rect 2450 8539 2516 8551
rect 2450 8503 2466 8539
rect 2500 8503 2516 8539
rect 2450 8469 2516 8503
rect 2450 8433 2466 8469
rect 2500 8433 2516 8469
rect 2450 8421 2516 8433
rect 2612 8539 2678 8551
rect 2612 8503 2628 8539
rect 2662 8503 2678 8539
rect 2612 8469 2678 8503
rect 2612 8433 2628 8469
rect 2662 8433 2678 8469
rect 2612 8421 2678 8433
rect 2774 8539 2840 8551
rect 2774 8503 2790 8539
rect 2824 8503 2840 8539
rect 2774 8469 2840 8503
rect 2774 8433 2790 8469
rect 2824 8433 2840 8469
rect 2774 8421 2840 8433
rect 2936 8539 3002 8551
rect 2936 8503 2952 8539
rect 2986 8503 3002 8539
rect 2936 8469 3002 8503
rect 2936 8433 2952 8469
rect 2986 8433 3002 8469
rect 2936 8421 3002 8433
rect 3098 8539 3164 8551
rect 3098 8503 3114 8539
rect 3148 8503 3164 8539
rect 3098 8469 3164 8503
rect 3098 8433 3114 8469
rect 3148 8433 3164 8469
rect 3098 8421 3164 8433
rect 3260 8539 3326 8551
rect 3260 8503 3276 8539
rect 3310 8503 3326 8539
rect 3260 8469 3326 8503
rect 3260 8433 3276 8469
rect 3310 8433 3326 8469
rect 3260 8421 3326 8433
rect 3422 8539 3488 8551
rect 3422 8505 3438 8539
rect 3472 8505 3488 8539
rect 3422 8467 3488 8505
rect 3422 8433 3438 8467
rect 3472 8433 3488 8467
rect 3422 8421 3488 8433
rect 3584 8539 3650 8551
rect 3584 8505 3600 8539
rect 3634 8505 3650 8539
rect 3584 8467 3650 8505
rect 3584 8433 3600 8467
rect 3634 8433 3650 8467
rect 3584 8421 3650 8433
rect 3746 8539 3812 8551
rect 3746 8505 3762 8539
rect 3796 8505 3812 8539
rect 3746 8467 3812 8505
rect 3746 8433 3762 8467
rect 3796 8433 3812 8467
rect 3746 8421 3812 8433
rect 3908 8539 3974 8551
rect 3908 8505 3924 8539
rect 3958 8505 3974 8539
rect 3908 8467 3974 8505
rect 3908 8433 3924 8467
rect 3958 8433 3974 8467
rect 3908 8421 3974 8433
rect 4070 8539 4136 8551
rect 4070 8505 4086 8539
rect 4120 8505 4136 8539
rect 4070 8467 4136 8505
rect 4070 8433 4086 8467
rect 4120 8433 4136 8467
rect 4070 8421 4136 8433
rect 344 4701 410 4713
rect 344 4667 360 4701
rect 394 4667 410 4701
rect 344 4629 410 4667
rect 344 4595 360 4629
rect 394 4595 410 4629
rect 344 4583 410 4595
rect 506 4701 572 4713
rect 506 4667 522 4701
rect 556 4667 572 4701
rect 506 4629 572 4667
rect 506 4595 522 4629
rect 556 4595 572 4629
rect 506 4583 572 4595
rect 668 4701 734 4713
rect 668 4667 684 4701
rect 718 4667 734 4701
rect 668 4629 734 4667
rect 668 4595 684 4629
rect 718 4595 734 4629
rect 668 4583 734 4595
rect 830 4701 896 4713
rect 830 4667 846 4701
rect 880 4667 896 4701
rect 830 4629 896 4667
rect 830 4595 846 4629
rect 880 4595 896 4629
rect 830 4583 896 4595
rect 992 4701 1058 4713
rect 992 4667 1008 4701
rect 1042 4667 1058 4701
rect 992 4629 1058 4667
rect 992 4595 1008 4629
rect 1042 4595 1058 4629
rect 992 4583 1058 4595
rect 1154 4701 1220 4713
rect 1154 4667 1170 4701
rect 1204 4667 1220 4701
rect 1154 4629 1220 4667
rect 1154 4595 1170 4629
rect 1204 4595 1220 4629
rect 1154 4583 1220 4595
rect 1316 4701 1382 4713
rect 1316 4667 1332 4701
rect 1366 4667 1382 4701
rect 1316 4629 1382 4667
rect 1316 4595 1332 4629
rect 1366 4595 1382 4629
rect 1316 4583 1382 4595
rect 1478 4701 1544 4713
rect 1478 4667 1494 4701
rect 1528 4667 1544 4701
rect 1478 4629 1544 4667
rect 1478 4595 1494 4629
rect 1528 4595 1544 4629
rect 1478 4583 1544 4595
rect 1640 4701 1706 4713
rect 1640 4667 1656 4701
rect 1690 4667 1706 4701
rect 1640 4629 1706 4667
rect 1640 4595 1656 4629
rect 1690 4595 1706 4629
rect 1640 4583 1706 4595
rect 1802 4701 1868 4713
rect 1802 4667 1818 4701
rect 1852 4667 1868 4701
rect 1802 4629 1868 4667
rect 1802 4595 1818 4629
rect 1852 4595 1868 4629
rect 1802 4583 1868 4595
rect 1964 4701 2030 4713
rect 1964 4667 1980 4701
rect 2014 4667 2030 4701
rect 1964 4629 2030 4667
rect 1964 4595 1980 4629
rect 2014 4595 2030 4629
rect 1964 4583 2030 4595
rect 2126 4701 2192 4713
rect 2126 4667 2142 4701
rect 2176 4667 2192 4701
rect 2126 4629 2192 4667
rect 2126 4595 2142 4629
rect 2176 4595 2192 4629
rect 2126 4583 2192 4595
rect 2288 4701 2354 4713
rect 2288 4667 2304 4701
rect 2338 4667 2354 4701
rect 2288 4629 2354 4667
rect 2288 4595 2304 4629
rect 2338 4595 2354 4629
rect 2288 4583 2354 4595
rect 2450 4701 2516 4713
rect 2450 4667 2466 4701
rect 2500 4667 2516 4701
rect 2450 4629 2516 4667
rect 2450 4595 2466 4629
rect 2500 4595 2516 4629
rect 2450 4583 2516 4595
rect 2612 4701 2678 4713
rect 2612 4667 2628 4701
rect 2662 4667 2678 4701
rect 2612 4629 2678 4667
rect 2612 4595 2628 4629
rect 2662 4595 2678 4629
rect 2612 4583 2678 4595
rect 2774 4701 2840 4713
rect 2774 4667 2790 4701
rect 2824 4667 2840 4701
rect 2774 4629 2840 4667
rect 2774 4595 2790 4629
rect 2824 4595 2840 4629
rect 2774 4583 2840 4595
rect 2936 4701 3002 4713
rect 2936 4667 2952 4701
rect 2986 4667 3002 4701
rect 2936 4629 3002 4667
rect 2936 4595 2952 4629
rect 2986 4595 3002 4629
rect 2936 4583 3002 4595
rect 3098 4701 3164 4713
rect 3098 4667 3114 4701
rect 3148 4667 3164 4701
rect 3098 4629 3164 4667
rect 3098 4595 3114 4629
rect 3148 4595 3164 4629
rect 3098 4583 3164 4595
rect 3260 4701 3326 4713
rect 3260 4667 3276 4701
rect 3310 4667 3326 4701
rect 3260 4629 3326 4667
rect 3260 4595 3276 4629
rect 3310 4595 3326 4629
rect 3260 4583 3326 4595
rect 3422 4701 3488 4713
rect 3422 4667 3438 4701
rect 3472 4667 3488 4701
rect 3422 4629 3488 4667
rect 3422 4595 3438 4629
rect 3472 4595 3488 4629
rect 3422 4583 3488 4595
rect 3584 4701 3650 4713
rect 3584 4667 3600 4701
rect 3634 4667 3650 4701
rect 3584 4629 3650 4667
rect 3584 4595 3600 4629
rect 3634 4595 3650 4629
rect 3584 4583 3650 4595
rect 3746 4701 3812 4713
rect 3746 4667 3762 4701
rect 3796 4667 3812 4701
rect 3746 4629 3812 4667
rect 3746 4595 3762 4629
rect 3796 4595 3812 4629
rect 3746 4583 3812 4595
rect 3908 4701 3974 4713
rect 3908 4667 3924 4701
rect 3958 4667 3974 4701
rect 3908 4629 3974 4667
rect 3908 4595 3924 4629
rect 3958 4595 3974 4629
rect 3908 4583 3974 4595
rect 4070 4701 4136 4713
rect 4070 4667 4086 4701
rect 4120 4667 4136 4701
rect 4070 4629 4136 4667
rect 4070 4595 4086 4629
rect 4120 4595 4136 4629
rect 4070 4583 4136 4595
rect 344 863 410 875
rect 344 829 360 863
rect 394 829 410 863
rect 344 793 410 829
rect 344 757 360 793
rect 394 757 410 793
rect 344 745 410 757
rect 506 863 572 875
rect 506 829 522 863
rect 556 829 572 863
rect 506 793 572 829
rect 506 757 522 793
rect 556 757 572 793
rect 506 745 572 757
rect 668 863 734 875
rect 668 829 684 863
rect 718 829 734 863
rect 668 793 734 829
rect 668 757 684 793
rect 718 757 734 793
rect 668 745 734 757
rect 830 863 896 875
rect 830 829 846 863
rect 880 829 896 863
rect 830 793 896 829
rect 830 757 846 793
rect 880 757 896 793
rect 830 745 896 757
rect 992 863 1058 875
rect 992 829 1008 863
rect 1042 829 1058 863
rect 992 793 1058 829
rect 992 757 1008 793
rect 1042 757 1058 793
rect 992 745 1058 757
rect 1154 863 1220 875
rect 1154 829 1170 863
rect 1204 829 1220 863
rect 1154 793 1220 829
rect 1154 757 1170 793
rect 1204 757 1220 793
rect 1154 745 1220 757
rect 1316 863 1382 875
rect 1316 829 1332 863
rect 1366 829 1382 863
rect 1316 793 1382 829
rect 1316 757 1332 793
rect 1366 757 1382 793
rect 1316 745 1382 757
rect 1478 863 1544 875
rect 1478 829 1494 863
rect 1528 829 1544 863
rect 1478 793 1544 829
rect 1478 757 1494 793
rect 1528 757 1544 793
rect 1478 745 1544 757
rect 1640 863 1706 875
rect 1640 829 1656 863
rect 1690 829 1706 863
rect 1640 793 1706 829
rect 1640 757 1656 793
rect 1690 757 1706 793
rect 1640 745 1706 757
rect 1802 863 1868 875
rect 1802 829 1818 863
rect 1852 829 1868 863
rect 1802 793 1868 829
rect 1802 757 1818 793
rect 1852 757 1868 793
rect 1802 745 1868 757
rect 1964 863 2030 875
rect 1964 829 1980 863
rect 2014 829 2030 863
rect 1964 793 2030 829
rect 1964 757 1980 793
rect 2014 757 2030 793
rect 1964 745 2030 757
rect 2126 863 2192 875
rect 2126 829 2142 863
rect 2176 829 2192 863
rect 2126 793 2192 829
rect 2126 757 2142 793
rect 2176 757 2192 793
rect 2126 745 2192 757
rect 2288 863 2354 875
rect 2288 829 2304 863
rect 2338 829 2354 863
rect 2288 793 2354 829
rect 2288 757 2304 793
rect 2338 757 2354 793
rect 2288 745 2354 757
rect 2450 863 2516 875
rect 2450 829 2466 863
rect 2500 829 2516 863
rect 2450 793 2516 829
rect 2450 757 2466 793
rect 2500 757 2516 793
rect 2450 745 2516 757
rect 2612 863 2678 875
rect 2612 829 2628 863
rect 2662 829 2678 863
rect 2612 793 2678 829
rect 2612 757 2628 793
rect 2662 757 2678 793
rect 2612 745 2678 757
rect 2774 863 2840 875
rect 2774 829 2790 863
rect 2824 829 2840 863
rect 2774 793 2840 829
rect 2774 757 2790 793
rect 2824 757 2840 793
rect 2774 745 2840 757
rect 2936 863 3002 875
rect 2936 829 2952 863
rect 2986 829 3002 863
rect 2936 793 3002 829
rect 2936 757 2952 793
rect 2986 757 3002 793
rect 2936 745 3002 757
rect 3098 863 3164 875
rect 3098 829 3114 863
rect 3148 829 3164 863
rect 3098 793 3164 829
rect 3098 757 3114 793
rect 3148 757 3164 793
rect 3098 745 3164 757
rect 3260 863 3326 875
rect 3260 829 3276 863
rect 3310 829 3326 863
rect 3260 793 3326 829
rect 3260 757 3276 793
rect 3310 757 3326 793
rect 3260 745 3326 757
rect 3422 863 3488 875
rect 3422 829 3438 863
rect 3472 829 3488 863
rect 3422 793 3488 829
rect 3422 757 3438 793
rect 3472 757 3488 793
rect 3422 745 3488 757
rect 3584 863 3650 875
rect 3584 829 3600 863
rect 3634 829 3650 863
rect 3584 793 3650 829
rect 3584 757 3600 793
rect 3634 757 3650 793
rect 3584 745 3650 757
rect 3746 863 3812 875
rect 3746 829 3762 863
rect 3796 829 3812 863
rect 3746 793 3812 829
rect 3746 757 3762 793
rect 3796 757 3812 793
rect 3746 745 3812 757
rect 3908 863 3974 875
rect 3908 829 3924 863
rect 3958 829 3974 863
rect 3908 793 3974 829
rect 3908 757 3924 793
rect 3958 757 3974 793
rect 3908 745 3974 757
rect 4070 863 4136 875
rect 4070 829 4086 863
rect 4120 829 4136 863
rect 4070 793 4136 829
rect 4070 757 4086 793
rect 4120 757 4136 793
rect 4070 745 4136 757
rect 198 631 232 671
rect 4248 631 4282 652
rect 198 597 279 631
rect 4209 597 4282 631
rect 1327 548 2573 549
rect 1327 515 1400 548
rect 1327 481 1328 515
rect 1362 514 1400 515
rect 1434 514 1468 548
rect 1502 514 1536 548
rect 1570 514 1604 548
rect 1638 514 1672 548
rect 1706 514 1740 548
rect 1774 514 1808 548
rect 1842 514 1876 548
rect 1910 514 1944 548
rect 1978 514 2012 548
rect 2046 514 2080 548
rect 2114 514 2148 548
rect 2182 514 2216 548
rect 2250 514 2284 548
rect 2318 514 2352 548
rect 2386 514 2420 548
rect 2454 514 2488 548
rect 2522 514 2573 548
rect 1362 513 2573 514
rect 1362 481 1363 513
rect 1327 469 1363 481
rect 1327 447 1329 469
rect 1327 413 1328 447
rect 1362 413 1363 435
rect 2537 478 2573 513
rect 2537 444 2538 478
rect 2572 444 2573 478
rect 2537 431 2573 444
rect 1327 397 1363 413
rect 1632 397 1670 431
rect 1704 397 1742 431
rect 1776 397 1814 431
rect 1848 397 1886 431
rect 1920 397 1958 431
rect 1992 397 2030 431
rect 2064 397 2102 431
rect 2136 397 2174 431
rect 2208 397 2247 431
rect 2281 397 2320 431
rect 2354 397 2393 431
rect 2427 397 2466 431
rect 2500 410 2539 431
rect 2500 397 2538 410
rect 1327 379 1329 397
rect 1327 345 1328 379
rect 2537 376 2538 397
rect 2572 376 2573 397
rect 1362 345 1363 363
rect 1327 325 1363 345
rect 1327 311 1329 325
rect 1327 277 1328 311
rect 1362 277 1363 291
rect 1327 253 1363 277
rect 1327 243 1329 253
rect 1327 209 1328 243
rect 1401 361 1502 375
rect 1401 359 1468 361
rect 1435 327 1468 359
rect 1435 325 1502 327
rect 2537 342 2573 376
rect 1401 291 1502 325
rect 1638 291 1681 325
rect 1715 291 1758 325
rect 1792 291 1835 325
rect 1869 291 1912 325
rect 1946 291 1989 325
rect 2023 291 2066 325
rect 2100 291 2143 325
rect 2177 291 2220 325
rect 2254 291 2297 325
rect 2331 291 2375 325
rect 2409 291 2453 325
rect 2537 308 2538 342
rect 2572 308 2573 342
rect 1435 289 1502 291
rect 1435 257 1468 289
rect 1401 255 1468 257
rect 1401 241 1502 255
rect 2537 274 2573 308
rect 2537 240 2538 274
rect 2572 240 2573 274
rect 2537 219 2573 240
rect 1362 209 1363 219
rect 1327 181 1363 209
rect 1632 185 1670 219
rect 1704 185 1742 219
rect 1776 185 1814 219
rect 1848 185 1886 219
rect 1920 185 1958 219
rect 1992 185 2030 219
rect 2064 185 2102 219
rect 2136 185 2174 219
rect 2208 185 2247 219
rect 2281 185 2320 219
rect 2354 185 2393 219
rect 2427 185 2466 219
rect 2500 206 2539 219
rect 2500 185 2538 206
rect 1327 147 1329 181
rect 1327 103 1363 147
rect 2537 172 2538 185
rect 2572 172 2573 185
rect 2537 138 2573 172
rect 2537 104 2538 138
rect 2572 104 2573 138
rect 2537 103 2573 104
rect 1327 102 2573 103
rect 1327 68 1361 102
rect 1395 68 1429 102
rect 1463 68 1497 102
rect 1531 68 1565 102
rect 1599 68 1633 102
rect 1667 68 1701 102
rect 1735 68 1769 102
rect 1803 68 1837 102
rect 1871 68 1905 102
rect 1939 68 1973 102
rect 2007 68 2041 102
rect 2075 68 2109 102
rect 2143 68 2177 102
rect 2211 68 2245 102
rect 2279 68 2313 102
rect 2347 68 2401 102
rect 2435 68 2469 102
rect 2503 68 2573 102
rect 1327 67 2573 68
<< viali >>
rect 2142 12375 2176 12377
rect 2142 12343 2176 12375
rect 2142 12271 2176 12305
rect 2304 12375 2338 12377
rect 2304 12343 2338 12375
rect 2304 12271 2338 12305
rect 2466 12375 2500 12377
rect 2466 12343 2500 12375
rect 2466 12271 2500 12305
rect 2628 12375 2662 12377
rect 2628 12343 2662 12375
rect 2628 12271 2662 12305
rect 2790 12375 2824 12377
rect 2790 12343 2824 12375
rect 2790 12271 2824 12305
rect 2952 12375 2986 12377
rect 2952 12343 2986 12375
rect 2952 12271 2986 12305
rect 3114 12375 3148 12377
rect 3114 12343 3148 12375
rect 3114 12271 3148 12305
rect 3276 12375 3310 12377
rect 3276 12343 3310 12375
rect 3276 12271 3310 12305
rect 3438 12375 3472 12377
rect 3438 12343 3472 12375
rect 3438 12271 3472 12305
rect 3600 12375 3634 12377
rect 3600 12343 3634 12375
rect 3600 12271 3634 12305
rect 3762 12375 3796 12377
rect 3762 12343 3796 12375
rect 3762 12271 3796 12305
rect 3924 12375 3958 12377
rect 3924 12343 3958 12375
rect 3924 12271 3958 12305
rect 4086 12375 4120 12377
rect 4086 12343 4120 12375
rect 4086 12271 4120 12305
rect 1322 10208 1356 10242
rect 1322 10136 1356 10170
rect -42 8917 -33 8951
rect -33 8917 -8 8951
rect 30 8917 35 8951
rect 35 8917 64 8951
rect 102 8917 103 8951
rect 103 8917 136 8951
rect 174 8917 205 8951
rect 205 8917 208 8951
rect 246 8917 273 8951
rect 273 8917 280 8951
rect 360 8537 394 8539
rect 360 8505 394 8537
rect 360 8435 394 8467
rect 360 8433 394 8435
rect 522 8537 556 8539
rect 522 8505 556 8537
rect 522 8435 556 8467
rect 522 8433 556 8435
rect 684 8537 718 8539
rect 684 8505 718 8537
rect 684 8435 718 8467
rect 684 8433 718 8435
rect 846 8537 880 8539
rect 846 8505 880 8537
rect 846 8435 880 8467
rect 846 8433 880 8435
rect 1008 8537 1042 8539
rect 1008 8505 1042 8537
rect 1008 8435 1042 8467
rect 1008 8433 1042 8435
rect 1170 8537 1204 8539
rect 1170 8505 1204 8537
rect 1170 8435 1204 8467
rect 1170 8433 1204 8435
rect 1332 8537 1366 8539
rect 1332 8505 1366 8537
rect 1332 8435 1366 8467
rect 1332 8433 1366 8435
rect 1494 8537 1528 8539
rect 1494 8505 1528 8537
rect 1494 8435 1528 8467
rect 1494 8433 1528 8435
rect 1656 8537 1690 8539
rect 1656 8505 1690 8537
rect 1656 8435 1690 8467
rect 1656 8433 1690 8435
rect 1818 8537 1852 8539
rect 1818 8505 1852 8537
rect 1818 8435 1852 8467
rect 1818 8433 1852 8435
rect 1980 8537 2014 8539
rect 1980 8505 2014 8537
rect 1980 8435 2014 8467
rect 1980 8433 2014 8435
rect 2142 8537 2176 8539
rect 2142 8505 2176 8537
rect 2142 8435 2176 8467
rect 2142 8433 2176 8435
rect 2304 8537 2338 8539
rect 2304 8505 2338 8537
rect 2304 8435 2338 8467
rect 2304 8433 2338 8435
rect 2466 8537 2500 8539
rect 2466 8505 2500 8537
rect 2466 8435 2500 8467
rect 2466 8433 2500 8435
rect 2628 8537 2662 8539
rect 2628 8505 2662 8537
rect 2628 8435 2662 8467
rect 2628 8433 2662 8435
rect 2790 8537 2824 8539
rect 2790 8505 2824 8537
rect 2790 8435 2824 8467
rect 2790 8433 2824 8435
rect 2952 8537 2986 8539
rect 2952 8505 2986 8537
rect 2952 8435 2986 8467
rect 2952 8433 2986 8435
rect 3114 8537 3148 8539
rect 3114 8505 3148 8537
rect 3114 8435 3148 8467
rect 3114 8433 3148 8435
rect 3276 8537 3310 8539
rect 3276 8505 3310 8537
rect 3276 8435 3310 8467
rect 3276 8433 3310 8435
rect 3438 8505 3472 8539
rect 3438 8433 3472 8467
rect 3600 8505 3634 8539
rect 3600 8433 3634 8467
rect 3762 8505 3796 8539
rect 3762 8433 3796 8467
rect 3924 8505 3958 8539
rect 3924 8433 3958 8467
rect 4086 8505 4120 8539
rect 4086 8433 4120 8467
rect 360 4667 394 4701
rect 360 4595 394 4629
rect 522 4667 556 4701
rect 522 4595 556 4629
rect 684 4667 718 4701
rect 684 4595 718 4629
rect 846 4667 880 4701
rect 846 4595 880 4629
rect 1008 4667 1042 4701
rect 1008 4595 1042 4629
rect 1170 4667 1204 4701
rect 1170 4595 1204 4629
rect 1332 4667 1366 4701
rect 1332 4595 1366 4629
rect 1494 4667 1528 4701
rect 1494 4595 1528 4629
rect 1656 4667 1690 4701
rect 1656 4595 1690 4629
rect 1818 4667 1852 4701
rect 1818 4595 1852 4629
rect 1980 4667 2014 4701
rect 1980 4595 2014 4629
rect 2142 4667 2176 4701
rect 2142 4595 2176 4629
rect 2304 4667 2338 4701
rect 2304 4595 2338 4629
rect 2466 4667 2500 4701
rect 2466 4595 2500 4629
rect 2628 4667 2662 4701
rect 2628 4595 2662 4629
rect 2790 4667 2824 4701
rect 2790 4595 2824 4629
rect 2952 4667 2986 4701
rect 2952 4595 2986 4629
rect 3114 4667 3148 4701
rect 3114 4595 3148 4629
rect 3276 4667 3310 4701
rect 3276 4595 3310 4629
rect 3438 4667 3472 4701
rect 3438 4595 3472 4629
rect 3600 4667 3634 4701
rect 3600 4595 3634 4629
rect 3762 4667 3796 4701
rect 3762 4595 3796 4629
rect 3924 4667 3958 4701
rect 3924 4595 3958 4629
rect 4086 4667 4120 4701
rect 4086 4595 4120 4629
rect 360 829 394 863
rect 360 759 394 791
rect 360 757 394 759
rect 522 829 556 863
rect 522 759 556 791
rect 522 757 556 759
rect 684 829 718 863
rect 684 759 718 791
rect 684 757 718 759
rect 846 829 880 863
rect 846 759 880 791
rect 846 757 880 759
rect 1008 829 1042 863
rect 1008 759 1042 791
rect 1008 757 1042 759
rect 1170 829 1204 863
rect 1170 759 1204 791
rect 1170 757 1204 759
rect 1332 829 1366 863
rect 1332 759 1366 791
rect 1332 757 1366 759
rect 1494 829 1528 863
rect 1494 759 1528 791
rect 1494 757 1528 759
rect 1656 829 1690 863
rect 1656 759 1690 791
rect 1656 757 1690 759
rect 1818 829 1852 863
rect 1818 759 1852 791
rect 1818 757 1852 759
rect 1980 829 2014 863
rect 1980 759 2014 791
rect 1980 757 2014 759
rect 2142 829 2176 863
rect 2142 759 2176 791
rect 2142 757 2176 759
rect 2304 829 2338 863
rect 2304 759 2338 791
rect 2304 757 2338 759
rect 2466 829 2500 863
rect 2466 759 2500 791
rect 2466 757 2500 759
rect 2628 829 2662 863
rect 2628 759 2662 791
rect 2628 757 2662 759
rect 2790 829 2824 863
rect 2790 759 2824 791
rect 2790 757 2824 759
rect 2952 829 2986 863
rect 2952 759 2986 791
rect 2952 757 2986 759
rect 3114 829 3148 863
rect 3114 759 3148 791
rect 3114 757 3148 759
rect 3276 829 3310 863
rect 3276 759 3310 791
rect 3276 757 3310 759
rect 3438 829 3472 863
rect 3438 759 3472 791
rect 3438 757 3472 759
rect 3600 829 3634 863
rect 3600 759 3634 791
rect 3600 757 3634 759
rect 3762 829 3796 863
rect 3762 759 3796 791
rect 3762 757 3796 759
rect 3924 829 3958 863
rect 3924 759 3958 791
rect 3924 757 3958 759
rect 4086 829 4120 863
rect 4086 759 4120 791
rect 4086 757 4120 759
rect 1329 447 1363 469
rect 1329 435 1362 447
rect 1362 435 1363 447
rect 1598 397 1632 431
rect 1670 397 1704 431
rect 1742 397 1776 431
rect 1814 397 1848 431
rect 1886 397 1920 431
rect 1958 397 1992 431
rect 2030 397 2064 431
rect 2102 397 2136 431
rect 2174 397 2208 431
rect 2247 397 2281 431
rect 2320 397 2354 431
rect 2393 397 2427 431
rect 2466 397 2500 431
rect 2539 410 2573 431
rect 2539 397 2572 410
rect 2572 397 2573 410
rect 1329 379 1363 397
rect 1329 363 1362 379
rect 1362 363 1363 379
rect 1329 311 1363 325
rect 1329 291 1362 311
rect 1362 291 1363 311
rect 1329 243 1363 253
rect 1329 219 1362 243
rect 1362 219 1363 243
rect 1468 327 1502 361
rect 1604 291 1638 325
rect 1681 291 1715 325
rect 1758 291 1792 325
rect 1835 291 1869 325
rect 1912 291 1946 325
rect 1989 291 2023 325
rect 2066 291 2100 325
rect 2143 291 2177 325
rect 2220 291 2254 325
rect 2297 291 2331 325
rect 2375 291 2409 325
rect 2453 291 2487 325
rect 1468 255 1502 289
rect 1598 185 1632 219
rect 1670 185 1704 219
rect 1742 185 1776 219
rect 1814 185 1848 219
rect 1886 185 1920 219
rect 1958 185 1992 219
rect 2030 185 2064 219
rect 2102 185 2136 219
rect 2174 185 2208 219
rect 2247 185 2281 219
rect 2320 185 2354 219
rect 2393 185 2427 219
rect 2466 185 2500 219
rect 2539 206 2573 219
rect 2539 185 2572 206
rect 2572 185 2573 206
rect 1329 147 1363 181
<< metal1 >>
rect 1691 12730 2281 12782
rect 2333 12730 2345 12782
rect 2397 12730 2409 12782
rect 2461 12730 2473 12782
rect 2525 12730 3577 12782
rect 3629 12730 3641 12782
rect 3693 12730 3705 12782
rect 3757 12730 3769 12782
rect 3821 12730 4434 12782
rect 1691 12650 4434 12702
rect 1691 12570 2281 12622
rect 2333 12570 2345 12622
rect 2397 12570 2409 12622
rect 2461 12570 2473 12622
rect 2525 12570 3577 12622
rect 3629 12570 3641 12622
rect 3693 12570 3705 12622
rect 3757 12570 3769 12622
rect 3821 12570 4434 12622
rect 1922 12490 1928 12542
rect 1980 12490 1992 12542
rect 2044 12490 2050 12542
tri 2050 12490 2056 12496 nw
tri 4194 12490 4200 12496 ne
rect 4200 12490 4206 12542
rect 4258 12490 4270 12542
rect 4322 12490 4328 12542
tri 1794 12406 1845 12457 se
rect 1845 12411 4328 12457
rect 1845 12406 1860 12411
tri 1860 12406 1865 12411 nw
tri 1769 10328 1794 10353 se
rect 1794 10328 1840 12406
tri 1840 12386 1860 12406 nw
rect 2130 12377 2350 12383
rect 2130 12343 2142 12377
rect 2176 12343 2304 12377
rect 2338 12343 2350 12377
rect 2130 12305 2350 12343
rect 2130 12271 2142 12305
rect 2176 12271 2304 12305
rect 2338 12271 2350 12305
rect 2130 12265 2350 12271
rect 2454 12377 2674 12383
rect 2454 12343 2466 12377
rect 2500 12343 2628 12377
rect 2662 12343 2674 12377
rect 2454 12305 2674 12343
rect 2454 12271 2466 12305
rect 2500 12271 2628 12305
rect 2662 12271 2674 12305
rect 2454 12265 2674 12271
rect 2778 12377 2998 12383
rect 2778 12343 2790 12377
rect 2824 12343 2952 12377
rect 2986 12343 2998 12377
rect 2778 12305 2998 12343
rect 2778 12271 2790 12305
rect 2824 12271 2952 12305
rect 2986 12271 2998 12305
rect 2778 12265 2998 12271
rect 3102 12377 3322 12383
rect 3102 12343 3114 12377
rect 3148 12343 3276 12377
rect 3310 12343 3322 12377
rect 3102 12305 3322 12343
rect 3102 12271 3114 12305
rect 3148 12271 3276 12305
rect 3310 12271 3322 12305
rect 3102 12265 3322 12271
rect 3426 12377 3646 12383
rect 3426 12343 3438 12377
rect 3472 12343 3600 12377
rect 3634 12343 3646 12377
rect 3426 12305 3646 12343
rect 3426 12271 3438 12305
rect 3472 12271 3600 12305
rect 3634 12271 3646 12305
rect 3426 12265 3646 12271
rect 3750 12377 3970 12383
rect 3750 12343 3762 12377
rect 3796 12343 3924 12377
rect 3958 12343 3970 12377
rect 3750 12305 3970 12343
rect 3750 12271 3762 12305
rect 3796 12271 3924 12305
rect 3958 12271 3970 12305
rect 3750 12265 3970 12271
rect 4074 12377 4132 12383
rect 4074 12343 4086 12377
rect 4120 12343 4132 12377
rect 4074 12305 4132 12343
rect 4074 12271 4086 12305
rect 4120 12271 4132 12305
tri 4049 12209 4074 12234 se
rect 4074 12209 4132 12271
tri 1840 10328 1865 10353 sw
rect -547 10282 1865 10328
rect 1866 10283 1867 10327
rect 1903 10283 1904 10327
rect 1905 10303 2487 10328
tri 2487 10303 2512 10328 sw
rect 1905 10282 2512 10303
tri -225 10257 -200 10282 ne
rect -547 10220 -232 10226
rect -547 10168 -284 10220
rect -547 10156 -232 10168
rect -547 10104 -284 10156
rect -547 10092 -232 10104
rect -547 10040 -284 10092
rect -547 10034 -232 10040
tri -481 10008 -455 10034 ne
rect -455 10008 -399 10034
tri -399 10008 -373 10034 nw
rect -200 9999 -142 10282
tri -142 10257 -117 10282 nw
tri 2429 10257 2454 10282 ne
rect 1316 10248 1564 10254
rect 1316 10242 1512 10248
rect -111 10220 1138 10226
rect -59 10168 991 10220
rect -111 10156 991 10168
rect -59 10104 991 10156
rect -111 10092 991 10104
rect -59 10040 991 10092
rect 1107 10040 1138 10220
rect 1316 10208 1322 10242
rect 1356 10208 1512 10242
rect 1316 10196 1512 10208
rect 1316 10184 1564 10196
rect 1316 10170 1512 10184
rect 1316 10136 1322 10170
rect 1356 10136 1512 10170
rect 1316 10132 1512 10136
rect 1316 10124 1564 10132
rect 1638 10191 1691 10195
rect -111 10034 1138 10040
tri 31 10008 57 10034 ne
rect 57 10008 113 10034
tri 113 10008 139 10034 nw
tri 543 10008 569 10034 ne
rect 569 10008 625 10034
tri 625 10008 651 10034 nw
tri 1055 10008 1081 10034 ne
rect 1081 10008 1138 10034
tri 1081 9999 1090 10008 ne
rect 1090 9999 1138 10008
tri 1090 9951 1138 9999 ne
rect 312 9369 370 9421
rect 313 9367 369 9368
rect 824 9343 882 9395
rect 825 9341 881 9342
rect 313 9330 369 9331
rect -200 9277 -142 9302
tri -142 9277 -117 9302 sw
tri 287 9277 312 9302 se
rect 312 9277 370 9329
rect 825 9304 881 9305
tri 370 9277 395 9302 sw
tri 799 9277 824 9302 se
rect 824 9277 882 9303
tri 882 9277 907 9302 sw
tri 1217 9277 1242 9302 se
rect -200 9219 1288 9277
tri 323 9194 348 9219 ne
rect -547 9138 292 9146
rect -367 9022 -264 9138
rect -84 9022 292 9138
rect -547 9013 292 9022
rect -84 8951 292 8957
rect -84 8917 -42 8951
rect -8 8917 30 8951
rect 64 8917 102 8951
rect 136 8917 174 8951
rect 208 8917 246 8951
rect 280 8917 292 8951
rect -84 8911 292 8917
rect -84 8870 -56 8911
tri -56 8870 -15 8911 nw
rect 348 8539 406 9219
tri 406 9194 431 9219 nw
tri 1364 9146 1389 9171 se
rect 1389 9146 1441 9250
rect 462 9138 1441 9146
rect 462 9022 466 9138
rect 582 9022 991 9138
rect 1107 9022 1325 9138
rect 462 9013 1441 9022
tri 1555 8957 1592 8994 se
rect 1638 8985 1639 10191
rect 1592 8957 1639 8985
rect 1577 8911 1639 8957
tri 1949 8705 1974 8730 se
rect 1974 8705 2026 8738
rect 1964 8659 2026 8705
rect 2454 8659 2512 10282
tri 3843 8684 3888 8729 se
tri 2512 8659 2537 8684 sw
tri 3818 8659 3843 8684 se
rect 3843 8659 3888 8684
rect 2454 8601 2564 8659
rect 2565 8602 2566 8658
rect 2602 8602 2603 8658
rect 2604 8601 3888 8659
rect 348 8505 360 8539
rect 394 8505 406 8539
rect 348 8467 406 8505
rect 348 8433 360 8467
rect 394 8433 406 8467
rect 348 8427 406 8433
rect 510 8539 730 8545
rect 510 8505 522 8539
rect 556 8505 684 8539
rect 718 8505 730 8539
rect 510 8467 730 8505
rect 510 8433 522 8467
rect 556 8433 684 8467
rect 718 8433 730 8467
rect 510 8427 730 8433
rect 834 8539 1054 8545
rect 834 8505 846 8539
rect 880 8505 1008 8539
rect 1042 8505 1054 8539
rect 834 8467 1054 8505
rect 834 8433 846 8467
rect 880 8433 1008 8467
rect 1042 8433 1054 8467
rect 834 8427 1054 8433
rect 1158 8539 1378 8545
rect 1158 8505 1170 8539
rect 1204 8505 1332 8539
rect 1366 8505 1378 8539
rect 1158 8467 1378 8505
rect 1158 8433 1170 8467
rect 1204 8433 1332 8467
rect 1366 8433 1378 8467
rect 1158 8427 1378 8433
rect 1482 8539 1702 8545
rect 1482 8505 1494 8539
rect 1528 8505 1656 8539
rect 1690 8505 1702 8539
rect 1482 8467 1702 8505
rect 1482 8433 1494 8467
rect 1528 8433 1656 8467
rect 1690 8433 1702 8467
rect 1482 8427 1702 8433
rect 1806 8539 2026 8545
rect 1806 8505 1818 8539
rect 1852 8505 1980 8539
rect 2014 8505 2026 8539
rect 1806 8467 2026 8505
rect 1806 8433 1818 8467
rect 1852 8433 1980 8467
rect 2014 8433 2026 8467
rect 1806 8427 2026 8433
rect 2130 8539 2188 8545
rect 2130 8505 2142 8539
rect 2176 8505 2188 8539
rect 2130 8467 2188 8505
rect 2130 8433 2142 8467
rect 2176 8433 2188 8467
rect 2130 8427 2188 8433
rect 2292 8539 2350 8545
rect 2292 8505 2304 8539
rect 2338 8505 2350 8539
rect 2292 8467 2350 8505
rect 2292 8433 2304 8467
rect 2338 8433 2350 8467
rect 2292 8427 2350 8433
rect 2454 8539 2512 8601
tri 2512 8576 2537 8601 nw
tri 4049 8576 4074 8601 ne
rect 2454 8505 2466 8539
rect 2500 8505 2512 8539
rect 2454 8467 2512 8505
rect 2454 8433 2466 8467
rect 2500 8433 2512 8467
rect 2454 8427 2512 8433
rect 2616 8539 2674 8545
rect 2616 8505 2628 8539
rect 2662 8505 2674 8539
rect 2616 8467 2674 8505
rect 2616 8433 2628 8467
rect 2662 8433 2674 8467
rect 2616 8427 2674 8433
rect 2778 8539 2836 8545
rect 2778 8505 2790 8539
rect 2824 8505 2836 8539
rect 2778 8467 2836 8505
rect 2778 8433 2790 8467
rect 2824 8433 2836 8467
rect 2778 8427 2836 8433
rect 2940 8539 2998 8545
rect 2940 8505 2952 8539
rect 2986 8505 2998 8539
rect 2940 8467 2998 8505
rect 2940 8433 2952 8467
rect 2986 8433 2998 8467
rect 2940 8427 2998 8433
rect 3102 8539 3160 8545
rect 3102 8505 3114 8539
rect 3148 8505 3160 8539
rect 3102 8467 3160 8505
rect 3102 8433 3114 8467
rect 3148 8433 3160 8467
rect 3102 8427 3160 8433
rect 3264 8539 3322 8545
rect 3264 8505 3276 8539
rect 3310 8505 3322 8539
rect 3264 8467 3322 8505
rect 3264 8433 3276 8467
rect 3310 8433 3322 8467
rect 3264 8427 3322 8433
rect 3426 8539 3484 8545
rect 3426 8505 3438 8539
rect 3472 8505 3484 8539
rect 3426 8467 3484 8505
rect 3426 8433 3438 8467
rect 3472 8433 3484 8467
rect 3426 8427 3484 8433
rect 3588 8539 3646 8545
rect 3588 8505 3600 8539
rect 3634 8505 3646 8539
rect 3588 8467 3646 8505
rect 3588 8433 3600 8467
rect 3634 8433 3646 8467
rect 3588 8427 3646 8433
rect 3750 8539 3808 8545
rect 3750 8505 3762 8539
rect 3796 8505 3808 8539
rect 3750 8467 3808 8505
rect 3750 8433 3762 8467
rect 3796 8433 3808 8467
rect 3750 8427 3808 8433
rect 3912 8539 3970 8545
rect 3912 8505 3924 8539
rect 3958 8505 3970 8539
rect 3912 8467 3970 8505
rect 3912 8433 3924 8467
rect 3958 8433 3970 8467
rect 3912 8427 3970 8433
rect 4074 8539 4132 8601
rect 4074 8505 4086 8539
rect 4120 8505 4132 8539
rect 4074 8467 4132 8505
rect 4074 8433 4086 8467
rect 4120 8433 4132 8467
rect 4074 8427 4132 8433
rect 348 4701 406 4707
rect 348 4667 360 4701
rect 394 4667 406 4701
rect 348 4629 406 4667
rect 348 4595 360 4629
rect 394 4595 406 4629
rect 348 4589 406 4595
rect 510 4701 568 4707
rect 510 4667 522 4701
rect 556 4667 568 4701
rect 510 4629 568 4667
rect 510 4595 522 4629
rect 556 4595 568 4629
rect 510 4589 568 4595
rect 672 4701 730 4707
rect 672 4667 684 4701
rect 718 4667 730 4701
rect 672 4629 730 4667
rect 672 4595 684 4629
rect 718 4595 730 4629
rect 672 4589 730 4595
rect 834 4701 892 4707
rect 834 4667 846 4701
rect 880 4667 892 4701
rect 834 4629 892 4667
rect 834 4595 846 4629
rect 880 4595 892 4629
rect 834 4589 892 4595
rect 996 4701 1054 4707
rect 996 4667 1008 4701
rect 1042 4667 1054 4701
rect 996 4629 1054 4667
rect 996 4595 1008 4629
rect 1042 4595 1054 4629
rect 996 4589 1054 4595
rect 1158 4701 1216 4707
rect 1158 4667 1170 4701
rect 1204 4667 1216 4701
rect 1158 4629 1216 4667
rect 1158 4595 1170 4629
rect 1204 4595 1216 4629
rect 1158 4589 1216 4595
rect 1320 4701 1378 4707
rect 1320 4667 1332 4701
rect 1366 4667 1378 4701
rect 1320 4629 1378 4667
rect 1320 4595 1332 4629
rect 1366 4595 1378 4629
rect 1320 4589 1378 4595
rect 1482 4701 1540 4707
rect 1482 4667 1494 4701
rect 1528 4667 1540 4701
rect 1482 4629 1540 4667
rect 1482 4595 1494 4629
rect 1528 4595 1540 4629
rect 1482 4589 1540 4595
rect 1644 4701 1702 4707
rect 1644 4667 1656 4701
rect 1690 4667 1702 4701
rect 1644 4629 1702 4667
rect 1644 4595 1656 4629
rect 1690 4595 1702 4629
rect 1644 4589 1702 4595
rect 1806 4701 1864 4707
rect 1806 4667 1818 4701
rect 1852 4667 1864 4701
rect 1806 4629 1864 4667
rect 1806 4595 1818 4629
rect 1852 4595 1864 4629
rect 1806 4589 1864 4595
rect 1968 4701 2026 4707
rect 1968 4667 1980 4701
rect 2014 4667 2026 4701
rect 1968 4629 2026 4667
rect 1968 4595 1980 4629
rect 2014 4595 2026 4629
rect 1968 4589 2026 4595
rect 2130 4701 2188 4707
rect 2130 4667 2142 4701
rect 2176 4667 2188 4701
rect 2130 4629 2188 4667
rect 2130 4595 2142 4629
rect 2176 4595 2188 4629
rect 2130 4589 2188 4595
rect 2292 4701 2350 4707
rect 2292 4667 2304 4701
rect 2338 4667 2350 4701
rect 2292 4629 2350 4667
rect 2292 4595 2304 4629
rect 2338 4595 2350 4629
rect 2292 4589 2350 4595
rect 2454 4701 2512 4707
rect 2454 4667 2466 4701
rect 2500 4667 2512 4701
rect 2454 4629 2512 4667
rect 2454 4595 2466 4629
rect 2500 4595 2512 4629
rect 2454 4589 2512 4595
rect 2616 4701 2674 4707
rect 2616 4667 2628 4701
rect 2662 4667 2674 4701
rect 2616 4629 2674 4667
rect 2616 4595 2628 4629
rect 2662 4595 2674 4629
rect 2616 4589 2674 4595
rect 2778 4701 2836 4707
rect 2778 4667 2790 4701
rect 2824 4667 2836 4701
rect 2778 4629 2836 4667
rect 2778 4595 2790 4629
rect 2824 4595 2836 4629
rect 2778 4589 2836 4595
rect 2940 4701 2998 4707
rect 2940 4667 2952 4701
rect 2986 4667 2998 4701
rect 2940 4629 2998 4667
rect 2940 4595 2952 4629
rect 2986 4595 2998 4629
rect 2940 4589 2998 4595
rect 3102 4701 3160 4707
rect 3102 4667 3114 4701
rect 3148 4667 3160 4701
rect 3102 4629 3160 4667
rect 3102 4595 3114 4629
rect 3148 4595 3160 4629
rect 3102 4589 3160 4595
rect 3264 4701 3322 4707
rect 3264 4667 3276 4701
rect 3310 4667 3322 4701
rect 3264 4629 3322 4667
rect 3264 4595 3276 4629
rect 3310 4595 3322 4629
rect 3264 4589 3322 4595
rect 3426 4701 3484 4707
rect 3426 4667 3438 4701
rect 3472 4667 3484 4701
rect 3426 4629 3484 4667
rect 3426 4595 3438 4629
rect 3472 4595 3484 4629
rect 3426 4589 3484 4595
rect 3588 4701 3646 4707
rect 3588 4667 3600 4701
rect 3634 4667 3646 4701
rect 3588 4629 3646 4667
rect 3588 4595 3600 4629
rect 3634 4595 3646 4629
rect 3588 4589 3646 4595
rect 3750 4701 3808 4707
rect 3750 4667 3762 4701
rect 3796 4667 3808 4701
rect 3750 4629 3808 4667
rect 3750 4595 3762 4629
rect 3796 4595 3808 4629
rect 3750 4589 3808 4595
rect 3912 4701 3970 4707
rect 3912 4667 3924 4701
rect 3958 4667 3970 4701
rect 3912 4629 3970 4667
rect 3912 4595 3924 4629
rect 3958 4595 3970 4629
rect 3912 4589 3970 4595
rect 4074 4701 4132 4707
rect 4074 4667 4086 4701
rect 4120 4667 4132 4701
rect 4074 4629 4132 4667
rect 4074 4595 4086 4629
rect 4120 4595 4132 4629
rect 4074 4589 4132 4595
rect 348 863 568 869
rect 348 829 360 863
rect 394 829 522 863
rect 556 829 568 863
rect 348 791 568 829
rect 348 757 360 791
rect 394 757 522 791
rect 556 757 568 791
rect 348 751 568 757
rect 672 863 892 869
rect 672 829 684 863
rect 718 829 846 863
rect 880 829 892 863
rect 672 791 892 829
rect 672 757 684 791
rect 718 757 846 791
rect 880 757 892 791
rect 672 751 892 757
rect 996 863 1216 869
rect 996 829 1008 863
rect 1042 829 1170 863
rect 1204 829 1216 863
rect 996 791 1216 829
rect 996 757 1008 791
rect 1042 757 1170 791
rect 1204 757 1216 791
rect 996 751 1216 757
rect 1320 863 1540 869
rect 1320 829 1332 863
rect 1366 829 1494 863
rect 1528 829 1540 863
rect 1320 791 1540 829
rect 1320 757 1332 791
rect 1366 757 1494 791
rect 1528 757 1540 791
rect 1320 751 1540 757
rect 1644 863 1864 869
rect 1644 829 1656 863
rect 1690 829 1818 863
rect 1852 829 1864 863
rect 1644 791 1864 829
rect 1644 757 1656 791
rect 1690 757 1818 791
rect 1852 757 1864 791
rect 1644 751 1864 757
rect 1968 863 2188 869
rect 1968 829 1980 863
rect 2014 829 2142 863
rect 2176 829 2188 863
rect 1968 791 2188 829
rect 1968 757 1980 791
rect 2014 757 2142 791
rect 2176 757 2188 791
rect 1968 751 2188 757
rect 2292 863 2512 869
rect 2292 829 2304 863
rect 2338 829 2466 863
rect 2500 829 2512 863
rect 2292 791 2512 829
rect 2292 757 2304 791
rect 2338 757 2466 791
rect 2500 757 2512 791
rect 2292 751 2512 757
rect 2616 863 2836 869
rect 2616 829 2628 863
rect 2662 829 2790 863
rect 2824 829 2836 863
rect 2616 791 2836 829
rect 2616 757 2628 791
rect 2662 757 2790 791
rect 2824 757 2836 791
rect 2616 751 2836 757
rect 2940 863 3160 869
rect 2940 829 2952 863
rect 2986 829 3114 863
rect 3148 829 3160 863
rect 2940 791 3160 829
rect 2940 757 2952 791
rect 2986 757 3114 791
rect 3148 757 3160 791
rect 2940 751 3160 757
rect 3264 863 3484 869
rect 3264 829 3276 863
rect 3310 829 3438 863
rect 3472 829 3484 863
rect 3264 791 3484 829
rect 3264 757 3276 791
rect 3310 757 3438 791
rect 3472 757 3484 791
rect 3264 751 3484 757
rect 3588 863 3808 869
rect 3588 829 3600 863
rect 3634 829 3762 863
rect 3796 829 3808 863
rect 3588 791 3808 829
rect 3588 757 3600 791
rect 3634 757 3762 791
rect 3796 757 3808 791
rect 3588 751 3808 757
rect 3912 863 4132 869
rect 3912 829 3924 863
rect 3958 829 4086 863
rect 4120 829 4132 863
rect 3912 791 4132 829
rect 3912 757 3924 791
rect 3958 757 4086 791
rect 4120 757 4132 791
rect 3912 751 4132 757
tri 4166 662 4242 738 se
rect 4242 662 4288 670
tri 238 659 241 662 sw
tri 4163 659 4166 662 se
rect 4166 659 4288 662
rect 192 637 241 659
tri 241 637 263 659 sw
tri 4141 637 4163 659 se
rect 4163 637 4288 659
rect 192 591 267 637
rect 4213 591 4288 637
tri 1298 566 1323 591 ne
rect 1323 469 4212 591
rect 1323 435 1329 469
rect 1363 435 4212 469
rect 1323 431 4212 435
rect 1323 416 1598 431
rect 1323 397 1400 416
tri 1400 397 1419 416 nw
tri 1561 397 1580 416 ne
rect 1580 397 1598 416
rect 1632 397 1670 431
rect 1704 397 1742 431
rect 1776 397 1814 431
rect 1848 397 1886 431
rect 1920 397 1958 431
rect 1992 397 2030 431
rect 2064 397 2102 431
rect 2136 397 2174 431
rect 2208 397 2247 431
rect 2281 397 2320 431
rect 2354 397 2393 431
rect 2427 397 2466 431
rect 2500 397 2539 431
rect 2573 400 4212 431
rect 2573 397 3838 400
rect 1323 363 1329 397
rect 1363 363 1369 397
tri 1369 366 1400 397 nw
tri 1580 391 1586 397 ne
rect 1586 391 3838 397
tri 3838 391 3847 400 nw
tri 4187 391 4196 400 ne
rect 4196 391 4212 400
tri 4196 375 4212 391 ne
rect 1462 366 1564 373
rect 1323 325 1369 363
rect 1323 291 1329 325
rect 1363 291 1369 325
rect 1323 253 1369 291
rect 1323 219 1329 253
rect 1363 219 1369 253
rect 1462 361 1512 366
rect 1462 327 1468 361
rect 1502 327 1512 361
rect 1462 314 1512 327
tri 3891 363 3900 372 se
rect 1462 302 1564 314
rect 1462 289 1512 302
rect 1462 255 1468 289
rect 1502 255 1512 289
rect 1462 250 1512 255
rect 1592 325 3900 363
rect 1592 291 1604 325
rect 1638 291 1681 325
rect 1715 291 1758 325
rect 1792 291 1835 325
rect 1869 291 1912 325
rect 1946 291 1989 325
rect 2023 291 2066 325
rect 2100 291 2143 325
rect 2177 291 2220 325
rect 2254 291 2297 325
rect 2331 291 2375 325
rect 2409 291 2453 325
rect 2487 291 3900 325
rect 1592 253 3900 291
tri 1369 219 1400 250 sw
rect 1462 243 1564 250
tri 3891 244 3900 253 ne
tri 4196 225 4212 241 se
tri 1580 219 1586 225 se
rect 1586 219 3838 225
rect 1323 200 1400 219
tri 1400 200 1419 219 sw
tri 1561 200 1580 219 se
rect 1580 200 1598 219
rect 1323 185 1598 200
rect 1632 185 1670 219
rect 1704 185 1742 219
rect 1776 185 1814 219
rect 1848 185 1886 219
rect 1920 185 1958 219
rect 1992 185 2030 219
rect 2064 185 2102 219
rect 2136 185 2174 219
rect 2208 185 2247 219
rect 2281 185 2320 219
rect 2354 185 2393 219
rect 2427 185 2466 219
rect 2500 185 2539 219
rect 2573 216 3838 219
tri 3838 216 3847 225 sw
tri 4187 216 4196 225 se
rect 4196 216 4212 225
rect 2573 185 4212 216
rect 1323 181 4212 185
rect 1323 147 1329 181
rect 1363 147 4212 181
rect 1323 136 4212 147
rect 1323 108 2611 136
tri 2611 108 2639 136 nw
rect 1323 62 1382 108
tri 2565 62 2611 108 nw
<< rmetal1 >>
rect 1865 10327 1867 10328
rect 1865 10283 1866 10327
rect 1865 10282 1867 10283
rect 1903 10327 1905 10328
rect 1904 10283 1905 10327
rect 1903 10282 1905 10283
rect 312 9368 370 9369
rect 312 9367 313 9368
rect 369 9367 370 9368
rect 824 9342 882 9343
rect 824 9341 825 9342
rect 881 9341 882 9342
rect 312 9330 313 9331
rect 369 9330 370 9331
rect 312 9329 370 9330
rect 824 9304 825 9305
rect 881 9304 882 9305
rect 824 9303 882 9304
rect 2564 8658 2566 8659
rect 2564 8602 2565 8658
rect 2564 8601 2566 8602
rect 2602 8658 2604 8659
rect 2603 8602 2604 8658
rect 2602 8601 2604 8602
<< via1 >>
rect 2281 12730 2333 12782
rect 2345 12730 2397 12782
rect 2409 12730 2461 12782
rect 2473 12730 2525 12782
rect 3577 12730 3629 12782
rect 3641 12730 3693 12782
rect 3705 12730 3757 12782
rect 3769 12730 3821 12782
rect 2281 12570 2333 12622
rect 2345 12570 2397 12622
rect 2409 12570 2461 12622
rect 2473 12570 2525 12622
rect 3577 12570 3629 12622
rect 3641 12570 3693 12622
rect 3705 12570 3757 12622
rect 3769 12570 3821 12622
rect 1928 12490 1980 12542
rect 1992 12490 2044 12542
rect 4206 12490 4258 12542
rect 4270 12490 4322 12542
rect -284 10168 -232 10220
rect -284 10104 -232 10156
rect -284 10040 -232 10092
rect -111 10168 -59 10220
rect -111 10104 -59 10156
rect -111 10040 -59 10092
rect 991 10040 1107 10220
rect 1512 10196 1564 10248
rect 1512 10132 1564 10184
rect -547 9022 -367 9138
rect -264 9022 -84 9138
rect 466 9022 582 9138
rect 991 9022 1107 9138
rect 1325 9022 1441 9138
rect 1512 314 1564 366
rect 1512 250 1564 302
<< metal2 >>
rect 2268 12730 2281 12782
rect 2333 12730 2345 12782
rect 2397 12730 2409 12782
rect 2461 12730 2473 12782
rect 2525 12730 2536 12782
rect 2268 12622 2536 12730
rect 2268 12570 2281 12622
rect 2333 12570 2345 12622
rect 2397 12570 2409 12622
rect 2461 12570 2473 12622
rect 2525 12570 2536 12622
rect -570 9138 -344 10416
rect -570 9022 -547 9138
rect -367 9022 -344 9138
rect -570 9016 -344 9022
rect -288 10220 -59 10416
rect -288 10168 -284 10220
rect -232 10168 -111 10220
rect -288 10156 -59 10168
rect -288 10104 -284 10156
rect -232 10104 -111 10156
rect -288 10092 -59 10104
rect -288 10040 -284 10092
rect -232 10040 -111 10092
rect -288 9138 -59 10040
rect -288 9022 -264 9138
rect -84 9022 -59 9138
rect -288 9016 -59 9022
rect 0 0 268 10416
rect 324 9138 592 10416
rect 324 9022 466 9138
rect 582 9022 592 9138
rect 324 0 592 9022
rect 648 0 916 10416
rect 972 10220 1126 10416
rect 972 10040 991 10220
rect 1107 10040 1126 10220
rect 972 9138 1126 10040
rect 972 9022 991 9138
rect 1107 9022 1126 9138
rect 972 0 1126 9022
rect 1188 0 1240 10416
rect 1296 9138 1441 10416
rect 1494 10284 1691 10416
tri 1595 10259 1620 10284 ne
rect 1296 9022 1325 9138
rect 1296 0 1441 9022
rect 1512 10248 1564 10254
rect 1512 10184 1564 10196
rect 1512 366 1564 10132
rect 1620 8911 1691 10284
rect 1512 302 1564 314
rect 1512 0 1564 250
tri 1620 8603 1747 8730 se
rect 1747 8603 1888 12542
rect 1922 12490 1928 12542
rect 1980 12490 1992 12542
rect 2044 12490 2050 12542
tri 1922 12468 1944 12490 ne
rect 1620 0 1888 8603
rect 1944 8659 2050 12490
tri 2091 8659 2106 8674 se
rect 2106 8659 2212 12542
tri 1944 8512 2091 8659 se
rect 2091 8512 2212 8659
rect 1944 0 2212 8512
rect 2268 0 2536 12570
rect 3564 12730 3577 12782
rect 3629 12730 3641 12782
rect 3693 12730 3705 12782
rect 3757 12730 3769 12782
rect 3821 12730 3832 12782
rect 3564 12622 3832 12730
rect 3564 12570 3577 12622
rect 3629 12570 3641 12622
rect 3693 12570 3705 12622
rect 3757 12570 3769 12622
rect 3821 12570 3832 12622
rect 2592 0 2860 12542
rect 2916 0 3184 12542
rect 3240 171 3508 12542
rect 3240 136 3473 171
tri 3473 136 3508 171 nw
rect 3564 168 3832 12570
rect 3888 244 4156 12542
rect 4200 12490 4206 12542
rect 4258 12490 4270 12542
rect 4322 12490 4434 12542
tri 4200 12478 4212 12490 ne
tri 3564 136 3596 168 ne
rect 3596 136 3832 168
rect 4212 136 4434 12490
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_0
timestamp 1704896540
transform 1 0 2628 0 1 8433
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_1
timestamp 1704896540
transform 1 0 360 0 1 4595
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_2
timestamp 1704896540
transform 1 0 522 0 1 4595
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_3
timestamp 1704896540
transform 1 0 684 0 1 4595
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_4
timestamp 1704896540
transform 1 0 846 0 1 4595
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_5
timestamp 1704896540
transform 1 0 1008 0 1 4595
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_6
timestamp 1704896540
transform 1 0 1170 0 1 4595
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_7
timestamp 1704896540
transform 1 0 1332 0 1 4595
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_8
timestamp 1704896540
transform 1 0 1494 0 1 4595
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_9
timestamp 1704896540
transform 1 0 1656 0 1 4595
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_10
timestamp 1704896540
transform 1 0 1818 0 1 4595
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_11
timestamp 1704896540
transform 1 0 1980 0 1 4595
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_12
timestamp 1704896540
transform 1 0 2142 0 1 4595
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_13
timestamp 1704896540
transform 1 0 2304 0 1 4595
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_14
timestamp 1704896540
transform 1 0 2466 0 1 4595
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_15
timestamp 1704896540
transform 1 0 2628 0 1 4595
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_16
timestamp 1704896540
transform 1 0 2790 0 1 4595
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_17
timestamp 1704896540
transform 1 0 2952 0 1 4595
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_18
timestamp 1704896540
transform 1 0 3114 0 1 4595
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_19
timestamp 1704896540
transform 1 0 3276 0 1 4595
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_20
timestamp 1704896540
transform 1 0 3438 0 1 4595
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_21
timestamp 1704896540
transform 1 0 3438 0 1 12271
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_22
timestamp 1704896540
transform 1 0 3762 0 1 12271
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_23
timestamp 1704896540
transform 1 0 4086 0 1 12271
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_24
timestamp 1704896540
transform 1 0 4086 0 1 4595
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_25
timestamp 1704896540
transform 1 0 3924 0 1 4595
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_26
timestamp 1704896540
transform 1 0 3762 0 1 4595
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_27
timestamp 1704896540
transform 1 0 3600 0 1 4595
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_28
timestamp 1704896540
transform 1 0 3600 0 1 12271
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_29
timestamp 1704896540
transform 1 0 3924 0 1 12271
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_30
timestamp 1704896540
transform 1 0 4086 0 1 8433
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_31
timestamp 1704896540
transform 1 0 3924 0 1 8433
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_32
timestamp 1704896540
transform 1 0 3762 0 1 8433
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_33
timestamp 1704896540
transform 1 0 3600 0 1 8433
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_34
timestamp 1704896540
transform 1 0 3438 0 1 8433
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_35
timestamp 1704896540
transform 1 0 3600 0 1 757
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_36
timestamp 1704896540
transform 1 0 3762 0 1 757
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_37
timestamp 1704896540
transform 1 0 3924 0 1 757
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_38
timestamp 1704896540
transform 1 0 4086 0 1 757
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_39
timestamp 1704896540
transform 1 0 3438 0 1 757
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_40
timestamp 1704896540
transform 1 0 3276 0 1 757
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_41
timestamp 1704896540
transform 1 0 3114 0 1 757
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_42
timestamp 1704896540
transform 1 0 2952 0 1 757
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_43
timestamp 1704896540
transform 1 0 2790 0 1 757
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_44
timestamp 1704896540
transform 1 0 2628 0 1 757
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_45
timestamp 1704896540
transform 1 0 2466 0 1 757
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_46
timestamp 1704896540
transform 1 0 2304 0 1 757
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_47
timestamp 1704896540
transform 1 0 2142 0 1 757
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_48
timestamp 1704896540
transform 1 0 1980 0 1 757
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_49
timestamp 1704896540
transform 1 0 1818 0 1 757
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_50
timestamp 1704896540
transform 1 0 1656 0 1 757
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_51
timestamp 1704896540
transform 1 0 1494 0 1 757
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_52
timestamp 1704896540
transform 1 0 1332 0 1 757
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_53
timestamp 1704896540
transform 1 0 1170 0 1 757
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_54
timestamp 1704896540
transform 1 0 1008 0 1 757
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_55
timestamp 1704896540
transform 1 0 846 0 1 757
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_56
timestamp 1704896540
transform 1 0 684 0 1 757
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_57
timestamp 1704896540
transform 1 0 522 0 1 757
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_58
timestamp 1704896540
transform 1 0 360 0 1 757
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_59
timestamp 1704896540
transform 1 0 2142 0 1 12271
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_60
timestamp 1704896540
transform 1 0 2304 0 1 12271
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_61
timestamp 1704896540
transform 1 0 2466 0 1 12271
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_62
timestamp 1704896540
transform 1 0 2628 0 1 12271
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_63
timestamp 1704896540
transform 1 0 2790 0 1 12271
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_64
timestamp 1704896540
transform 1 0 2952 0 1 12271
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_65
timestamp 1704896540
transform 1 0 3114 0 1 12271
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_66
timestamp 1704896540
transform 1 0 3276 0 1 12271
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_67
timestamp 1704896540
transform 1 0 360 0 1 8433
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_68
timestamp 1704896540
transform 1 0 522 0 1 8433
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_69
timestamp 1704896540
transform 1 0 684 0 1 8433
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_70
timestamp 1704896540
transform 1 0 846 0 1 8433
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_71
timestamp 1704896540
transform 1 0 1008 0 1 8433
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_72
timestamp 1704896540
transform 1 0 1170 0 1 8433
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_73
timestamp 1704896540
transform 1 0 1332 0 1 8433
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_74
timestamp 1704896540
transform 1 0 1494 0 1 8433
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_75
timestamp 1704896540
transform 1 0 1656 0 1 8433
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_76
timestamp 1704896540
transform 1 0 1818 0 1 8433
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_77
timestamp 1704896540
transform 1 0 1980 0 1 8433
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_78
timestamp 1704896540
transform 1 0 2142 0 1 8433
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_79
timestamp 1704896540
transform 1 0 2304 0 1 8433
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_80
timestamp 1704896540
transform 1 0 2466 0 1 8433
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_81
timestamp 1704896540
transform 1 0 2790 0 1 8433
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_82
timestamp 1704896540
transform 1 0 2952 0 1 8433
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_83
timestamp 1704896540
transform 1 0 3114 0 1 8433
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_84
timestamp 1704896540
transform 1 0 3276 0 1 8433
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1704896540
transform 0 1 1322 -1 0 10242
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1704896540
transform 0 1 1468 1 0 255
box 0 0 1 1
use L1M1_CDNS_52468879185193  L1M1_CDNS_52468879185193_0
timestamp 1704896540
transform -1 0 280 0 -1 8951
box 0 0 1 1
use L1M1_CDNS_52468879185193  L1M1_CDNS_52468879185193_1
timestamp 1704896540
transform 0 1 1329 1 0 147
box 0 0 1 1
use L1M1_CDNS_52468879185307  L1M1_CDNS_52468879185307_0
timestamp 1704896540
transform 1 0 -376 0 1 10288
box -12 -6 1414 40
use L1M1_CDNS_52468879185316  L1M1_CDNS_52468879185316_0
timestamp 1704896540
transform 1 0 -330 0 -1 9140
box -12 -6 622 40
use L1M1_CDNS_52468879185335  L1M1_CDNS_52468879185335_0
timestamp 1704896540
transform 1 0 476 0 -1 8951
box -12 -6 1126 40
use L1M1_CDNS_52468879185381  L1M1_CDNS_52468879185381_0
timestamp 1704896540
transform 0 1 1395 1 0 9172
box -12 -6 910 40
use L1M1_CDNS_52468879185381  L1M1_CDNS_52468879185381_1
timestamp 1704896540
transform 1 0 476 0 -1 9140
box -12 -6 910 40
use L1M1_CDNS_52468879185950  L1M1_CDNS_52468879185950_0
timestamp 1704896540
transform 0 -1 4282 1 0 670
box -12 -6 11638 40
use L1M1_CDNS_52468879185952  L1M1_CDNS_52468879185952_0
timestamp 1704896540
transform 1 0 279 0 -1 631
box -12 -6 3934 40
use L1M1_CDNS_52468879185955  L1M1_CDNS_52468879185955_0
timestamp 1704896540
transform 0 -1 1282 1 0 9239
box -12 -6 982 40
use L1M1_CDNS_524688791851010  L1M1_CDNS_524688791851010_0
timestamp 1704896540
transform -1 0 4228 0 1 12502
box -12 -6 2206 40
use L1M1_CDNS_524688791851011  L1M1_CDNS_524688791851011_0
timestamp 1704896540
transform 0 1 1598 1 0 8997
box -12 -6 1198 40
use L1M1_CDNS_524688791851011  L1M1_CDNS_524688791851011_1
timestamp 1704896540
transform 1 0 1367 0 -1 548
box -12 -6 1198 40
use L1M1_CDNS_524688791851011  L1M1_CDNS_524688791851011_2
timestamp 1704896540
transform 1 0 1367 0 -1 102
box -12 -6 1198 40
use L1M1_CDNS_524688791851012  L1M1_CDNS_524688791851012_0
timestamp 1704896540
transform 0 1 1980 -1 0 10224
box -12 -6 1486 40
use L1M1_CDNS_524688791851012  L1M1_CDNS_524688791851012_1
timestamp 1704896540
transform -1 0 1952 0 -1 8699
box -12 -6 1486 40
use L1M1_CDNS_524688791851013  L1M1_CDNS_524688791851013_0
timestamp 1704896540
transform 0 -1 232 1 0 671
box -12 -6 8038 40
use L1M1_CDNS_524688791851014  L1M1_CDNS_524688791851014_0
timestamp 1704896540
transform -1 0 -154 0 1 9239
box -12 -6 46 760
use L1M1_CDNS_524688791851015  L1M1_CDNS_524688791851015_0
timestamp 1704896540
transform -1 0 614 0 -1 10209
box -12 -6 46 904
use L1M1_CDNS_524688791851015  L1M1_CDNS_524688791851015_1
timestamp 1704896540
transform -1 0 102 0 -1 10209
box -12 -6 46 904
use L1M1_CDNS_524688791851015  L1M1_CDNS_524688791851015_2
timestamp 1704896540
transform -1 0 -410 0 -1 10209
box -12 -6 46 904
use L1M1_CDNS_524688791851016  L1M1_CDNS_524688791851016_0
timestamp 1704896540
transform -1 0 870 0 -1 9993
box -12 -6 46 616
use L1M1_CDNS_524688791851016  L1M1_CDNS_524688791851016_1
timestamp 1704896540
transform -1 0 358 0 -1 9993
box -12 -6 46 616
use L1M1_CDNS_524688791851017  L1M1_CDNS_524688791851017_0
timestamp 1704896540
transform 0 -1 2014 1 0 10406
box -12 -6 1918 40
use L1M1_CDNS_524688791851018  L1M1_CDNS_524688791851018_0
timestamp 1704896540
transform -1 0 1126 0 -1 10209
box -12 -6 46 832
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1704896540
transform -1 0 2050 0 1 12490
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_1
timestamp 1704896540
transform 0 1 1512 1 0 244
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_2
timestamp 1704896540
transform 0 1 1512 1 0 10126
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_3
timestamp 1704896540
transform 1 0 4200 0 1 12490
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_0
timestamp 1704896540
transform 0 1 991 1 0 10034
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_0
timestamp 1704896540
transform 0 1 466 1 0 9016
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_1
timestamp 1704896540
transform 0 1 991 1 0 9016
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_2
timestamp 1704896540
transform 0 1 1325 1 0 9016
box 0 0 1 1
use M1M2_CDNS_52468879185200  M1M2_CDNS_52468879185200_0
timestamp 1704896540
transform 0 1 -547 1 0 9016
box 0 0 1 1
use M1M2_CDNS_52468879185200  M1M2_CDNS_52468879185200_1
timestamp 1704896540
transform 0 1 -264 1 0 9016
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_0
timestamp 1704896540
transform 0 1 -284 1 0 10034
box 0 0 1 1
use M1M2_CDNS_52468879185203  M1M2_CDNS_52468879185203_1
timestamp 1704896540
transform 0 -1 -59 1 0 10034
box 0 0 1 1
use M1M2_CDNS_52468879185208  M1M2_CDNS_52468879185208_0
timestamp 1704896540
transform 0 1 336 1 0 10034
box 0 0 192 244
use M1M2_CDNS_52468879185208  M1M2_CDNS_52468879185208_1
timestamp 1704896540
transform 0 1 12 1 0 10034
box 0 0 192 244
use M1M2_CDNS_52468879185209  M1M2_CDNS_52468879185209_0
timestamp 1704896540
transform 0 1 3888 -1 0 8729
box 0 0 128 244
use M1M2_CDNS_52468879185209  M1M2_CDNS_52468879185209_1
timestamp 1704896540
transform 0 1 3888 -1 0 12209
box 0 0 128 244
use M1M2_CDNS_52468879185209  M1M2_CDNS_52468879185209_2
timestamp 1704896540
transform 0 1 3900 1 0 244
box 0 0 128 244
use M1M2_CDNS_52468879185209  M1M2_CDNS_52468879185209_3
timestamp 1704896540
transform 0 1 12 1 0 9016
box 0 0 128 244
use M1M2_CDNS_52468879185297  M1M2_CDNS_52468879185297_0
timestamp 1704896540
transform -1 0 3827 0 1 12570
box 0 0 1 1
use M1M2_CDNS_52468879185297  M1M2_CDNS_52468879185297_1
timestamp 1704896540
transform -1 0 3827 0 1 12730
box 0 0 1 1
use M1M2_CDNS_52468879185297  M1M2_CDNS_52468879185297_2
timestamp 1704896540
transform -1 0 2531 0 1 12570
box 0 0 1 1
use M1M2_CDNS_52468879185297  M1M2_CDNS_52468879185297_3
timestamp 1704896540
transform -1 0 2531 0 1 12730
box 0 0 1 1
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_0
timestamp 1704896540
transform 0 1 -547 1 0 10034
box 0 0 192 180
use M1M2_CDNS_524688791851019  M1M2_CDNS_524688791851019_0
timestamp 1704896540
transform 0 1 1974 1 0 8700
box 0 0 1536 52
use M1M2_CDNS_524688791851020  M1M2_CDNS_524688791851020_0
timestamp 1704896540
transform 0 1 1974 1 0 10394
box 0 0 1984 52
use M1M2_CDNS_524688791851021  M1M2_CDNS_524688791851021_0
timestamp 1704896540
transform 0 1 4212 1 0 136
box 0 0 12224 116
use M1M2_CDNS_524688791851022  M1M2_CDNS_524688791851022_0
timestamp 1704896540
transform 0 -1 1691 -1 0 10191
box 0 0 1280 52
use M1M2_CDNS_524688791851023  M1M2_CDNS_524688791851023_0
timestamp 1704896540
transform 0 1 1389 1 0 9250
box 0 0 832 52
use nfet_CDNS_524688791851024  nfet_CDNS_524688791851024_0
timestamp 1704896540
transform -1 0 57 0 1 9240
box -79 -52 535 1052
use nfet_CDNS_524688791851024  nfet_CDNS_524688791851024_1
timestamp 1704896540
transform -1 0 569 0 1 9240
box -79 -52 535 1052
use nfet_CDNS_524688791851024  nfet_CDNS_524688791851024_2
timestamp 1704896540
transform -1 0 1081 0 1 9240
box -79 -52 535 1052
use nfet_CDNS_524688791851025  nfet_CDNS_524688791851025_0
timestamp 1704896540
transform -1 0 1237 0 1 9240
box -79 -52 179 1052
use pTran_CDNS_524688791851027  pTran_CDNS_524688791851027_0
timestamp 1704896540
transform 0 -1 2483 1 0 230
box -89 -36 245 1036
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_0
timestamp 1704896540
transform 0 -1 410 -1 0 809
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_1
timestamp 1704896540
transform 0 -1 572 -1 0 809
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_2
timestamp 1704896540
transform 0 -1 734 -1 0 809
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_3
timestamp 1704896540
transform 0 -1 896 -1 0 809
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_4
timestamp 1704896540
transform 0 -1 1058 -1 0 809
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_5
timestamp 1704896540
transform 0 -1 1220 -1 0 809
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_6
timestamp 1704896540
transform 0 -1 1382 -1 0 809
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_7
timestamp 1704896540
transform 0 -1 1544 -1 0 809
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_8
timestamp 1704896540
transform 0 -1 1706 -1 0 809
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_9
timestamp 1704896540
transform 0 -1 1868 -1 0 809
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_10
timestamp 1704896540
transform 0 -1 2030 -1 0 809
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_11
timestamp 1704896540
transform 0 -1 2192 -1 0 809
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_12
timestamp 1704896540
transform 0 -1 2354 -1 0 809
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_13
timestamp 1704896540
transform 0 -1 2516 -1 0 809
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_14
timestamp 1704896540
transform 0 -1 2678 -1 0 809
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_15
timestamp 1704896540
transform 0 -1 2840 -1 0 809
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_16
timestamp 1704896540
transform 0 -1 3002 -1 0 809
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_17
timestamp 1704896540
transform 0 -1 3164 -1 0 809
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_18
timestamp 1704896540
transform 0 -1 3326 -1 0 809
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_19
timestamp 1704896540
transform 0 -1 3488 -1 0 809
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_20
timestamp 1704896540
transform 0 -1 3650 -1 0 809
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_21
timestamp 1704896540
transform 0 -1 3812 -1 0 809
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_22
timestamp 1704896540
transform 0 -1 3974 -1 0 809
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_23
timestamp 1704896540
transform 0 -1 4136 -1 0 809
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_24
timestamp 1704896540
transform 0 -1 3326 -1 0 8485
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_25
timestamp 1704896540
transform 0 -1 3164 -1 0 8485
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_26
timestamp 1704896540
transform 0 -1 3002 -1 0 8485
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_27
timestamp 1704896540
transform 0 -1 2840 -1 0 8485
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_28
timestamp 1704896540
transform 0 -1 2678 -1 0 8485
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_29
timestamp 1704896540
transform 0 -1 2516 -1 0 8485
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_30
timestamp 1704896540
transform 0 -1 2354 -1 0 8485
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_31
timestamp 1704896540
transform 0 -1 2192 -1 0 8485
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_32
timestamp 1704896540
transform 0 -1 2030 -1 0 8485
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_33
timestamp 1704896540
transform 0 -1 1868 -1 0 8485
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_34
timestamp 1704896540
transform 0 -1 1706 -1 0 8485
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_35
timestamp 1704896540
transform 0 -1 1544 -1 0 8485
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_36
timestamp 1704896540
transform 0 -1 1382 -1 0 8485
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_37
timestamp 1704896540
transform 0 -1 1220 -1 0 8485
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_38
timestamp 1704896540
transform 0 -1 1058 -1 0 8485
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_39
timestamp 1704896540
transform 0 -1 896 -1 0 8485
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_40
timestamp 1704896540
transform 0 -1 734 -1 0 8485
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_41
timestamp 1704896540
transform 0 -1 572 -1 0 8485
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_42
timestamp 1704896540
transform 0 -1 410 -1 0 8485
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_43
timestamp 1704896540
transform 0 -1 3812 1 0 12325
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_44
timestamp 1704896540
transform 0 -1 3974 1 0 12325
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_45
timestamp 1704896540
transform 0 -1 3650 1 0 12325
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_46
timestamp 1704896540
transform 0 -1 734 1 0 8487
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_47
timestamp 1704896540
transform 0 -1 572 1 0 8487
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_48
timestamp 1704896540
transform 0 -1 410 1 0 8487
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_49
timestamp 1704896540
transform 0 -1 3488 1 0 12325
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_50
timestamp 1704896540
transform 0 -1 3326 1 0 8487
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_51
timestamp 1704896540
transform 0 -1 3164 1 0 8487
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_52
timestamp 1704896540
transform 0 -1 3002 1 0 8487
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_53
timestamp 1704896540
transform 0 -1 2840 1 0 8487
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_54
timestamp 1704896540
transform 0 -1 2678 1 0 8487
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_55
timestamp 1704896540
transform 0 -1 2516 1 0 8487
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_56
timestamp 1704896540
transform 0 -1 2354 1 0 8487
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_57
timestamp 1704896540
transform 0 -1 2192 1 0 8487
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_58
timestamp 1704896540
transform 0 -1 2030 1 0 8487
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_59
timestamp 1704896540
transform 0 -1 1868 1 0 8487
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_60
timestamp 1704896540
transform 0 -1 1706 1 0 8487
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_61
timestamp 1704896540
transform 0 -1 1544 1 0 8487
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_62
timestamp 1704896540
transform 0 -1 1382 1 0 8487
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_63
timestamp 1704896540
transform 0 -1 1220 1 0 8487
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_64
timestamp 1704896540
transform 0 -1 1058 1 0 8487
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_65
timestamp 1704896540
transform 0 -1 896 1 0 8487
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_66
timestamp 1704896540
transform 0 -1 2192 1 0 12325
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_67
timestamp 1704896540
transform 0 -1 2354 1 0 12325
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_68
timestamp 1704896540
transform 0 -1 2516 1 0 12325
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_69
timestamp 1704896540
transform 0 -1 2678 1 0 12325
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_70
timestamp 1704896540
transform 0 -1 2840 1 0 12325
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_71
timestamp 1704896540
transform 0 -1 3002 1 0 12325
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_72
timestamp 1704896540
transform 0 -1 3164 1 0 12325
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_73
timestamp 1704896540
transform 0 -1 3326 1 0 12325
box 0 0 1 1
use PYL1_CDNS_524688791857  PYL1_CDNS_524688791857_74
timestamp 1704896540
transform 0 -1 4136 1 0 12325
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_0
timestamp 1704896540
transform 0 1 -366 -1 0 10338
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_1
timestamp 1704896540
transform 0 1 -110 -1 0 10338
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_2
timestamp 1704896540
transform 0 1 146 -1 0 10338
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_3
timestamp 1704896540
transform 0 1 402 -1 0 10338
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_4
timestamp 1704896540
transform 0 1 658 -1 0 10338
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_5
timestamp 1704896540
transform 0 1 914 -1 0 10338
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_6
timestamp 1704896540
transform 0 1 1137 -1 0 10338
box 0 0 1 1
use PYL1_CDNS_5246887918562  PYL1_CDNS_5246887918562_7
timestamp 1704896540
transform 1 0 1385 0 1 241
box 0 0 1 1
use PYL1_CDNS_524688791851004  PYL1_CDNS_524688791851004_0
timestamp 1704896540
transform 0 1 2044 1 0 12487
box 0 0 66 2174
use PYL1_CDNS_524688791851005  PYL1_CDNS_524688791851005_0
timestamp 1704896540
transform -1 0 2030 0 -1 12470
box 0 0 66 3738
use PYL1_CDNS_524688791851006  PYL1_CDNS_524688791851006_0
timestamp 1704896540
transform 0 1 257 -1 0 8715
box 0 0 66 1698
use PYL1_CDNS_524688791851007  PYL1_CDNS_524688791851007_0
timestamp 1704896540
transform -1 0 248 0 1 671
box 0 0 66 7954
use PYL1_CDNS_524688791851008  PYL1_CDNS_524688791851008_0
timestamp 1704896540
transform -1 0 4298 0 -1 12482
box 0 0 66 11830
use PYL1_CDNS_524688791851009  PYL1_CDNS_524688791851009_0
timestamp 1704896540
transform 0 -1 4213 -1 0 647
box 0 0 66 3466
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_0
timestamp 1704896540
transform 0 -1 3488 -1 0 12273
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_1
timestamp 1704896540
transform 0 -1 3650 -1 0 12273
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_2
timestamp 1704896540
transform 0 -1 3326 -1 0 12273
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_3
timestamp 1704896540
transform 0 -1 3002 -1 0 8435
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_4
timestamp 1704896540
transform 0 -1 734 -1 0 8435
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_5
timestamp 1704896540
transform 0 -1 1058 -1 0 8435
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_6
timestamp 1704896540
transform 0 -1 2840 -1 0 4597
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_7
timestamp 1704896540
transform 0 -1 2516 -1 0 8435
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_8
timestamp 1704896540
transform 0 -1 2516 -1 0 4597
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_9
timestamp 1704896540
transform 0 -1 2840 -1 0 12273
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_10
timestamp 1704896540
transform 0 -1 2354 -1 0 4597
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_11
timestamp 1704896540
transform 0 -1 2354 -1 0 8435
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_12
timestamp 1704896540
transform 0 -1 1058 -1 0 4597
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_13
timestamp 1704896540
transform 0 -1 2192 -1 0 4597
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_14
timestamp 1704896540
transform 0 -1 2192 -1 0 8435
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_15
timestamp 1704896540
transform 0 -1 734 -1 0 4597
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_16
timestamp 1704896540
transform 0 -1 2030 -1 0 4597
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_17
timestamp 1704896540
transform 0 -1 2030 -1 0 8435
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_18
timestamp 1704896540
transform 0 -1 3002 -1 0 12273
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_19
timestamp 1704896540
transform 0 -1 1220 -1 0 8435
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_20
timestamp 1704896540
transform 0 -1 4136 -1 0 8435
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_21
timestamp 1704896540
transform 0 -1 2678 -1 0 12273
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_22
timestamp 1704896540
transform 0 -1 1220 -1 0 4597
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_23
timestamp 1704896540
transform 0 -1 3650 -1 0 4597
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_24
timestamp 1704896540
transform 0 -1 3812 -1 0 4597
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_25
timestamp 1704896540
transform 0 -1 3650 -1 0 8435
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_26
timestamp 1704896540
transform 0 -1 2840 -1 0 8435
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_27
timestamp 1704896540
transform 0 -1 3974 -1 0 4597
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_28
timestamp 1704896540
transform 0 -1 4136 -1 0 4597
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_29
timestamp 1704896540
transform 0 -1 1382 -1 0 8435
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_30
timestamp 1704896540
transform 0 -1 1382 -1 0 4597
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_31
timestamp 1704896540
transform 0 -1 4136 -1 0 12273
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_32
timestamp 1704896540
transform 0 -1 2678 -1 0 8435
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_33
timestamp 1704896540
transform 0 -1 3812 -1 0 12273
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_34
timestamp 1704896540
transform 0 -1 3974 -1 0 12273
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_35
timestamp 1704896540
transform 0 -1 3812 -1 0 8435
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_36
timestamp 1704896540
transform 0 -1 3164 -1 0 12273
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_37
timestamp 1704896540
transform 0 -1 1544 -1 0 8435
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_38
timestamp 1704896540
transform 0 -1 896 -1 0 4597
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_39
timestamp 1704896540
transform 0 -1 1544 -1 0 4597
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_40
timestamp 1704896540
transform 0 -1 3974 -1 0 8435
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_41
timestamp 1704896540
transform 0 -1 2192 -1 0 12273
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_42
timestamp 1704896540
transform 0 -1 410 -1 0 8435
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_43
timestamp 1704896540
transform 0 -1 1706 -1 0 8435
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_44
timestamp 1704896540
transform 0 -1 410 -1 0 4597
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_45
timestamp 1704896540
transform 0 -1 1706 -1 0 4597
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_46
timestamp 1704896540
transform 0 -1 1868 -1 0 8435
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_47
timestamp 1704896540
transform 0 -1 1868 -1 0 4597
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_48
timestamp 1704896540
transform 0 -1 2354 -1 0 12273
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_49
timestamp 1704896540
transform 0 -1 572 -1 0 8435
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_50
timestamp 1704896540
transform 0 -1 3488 -1 0 8435
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_51
timestamp 1704896540
transform 0 -1 572 -1 0 4597
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_52
timestamp 1704896540
transform 0 -1 3488 -1 0 4597
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_53
timestamp 1704896540
transform 0 -1 2516 -1 0 12273
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_54
timestamp 1704896540
transform 0 -1 3326 -1 0 4597
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_55
timestamp 1704896540
transform 0 -1 3326 -1 0 8435
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_56
timestamp 1704896540
transform 0 -1 3164 -1 0 4597
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_57
timestamp 1704896540
transform 0 -1 3164 -1 0 8435
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_58
timestamp 1704896540
transform 0 -1 3002 -1 0 4597
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_59
timestamp 1704896540
transform 0 -1 896 -1 0 8435
box -50 0 3786 66
use PYres_CDNS_524688791851026  PYres_CDNS_524688791851026_60
timestamp 1704896540
transform 0 -1 2678 -1 0 4597
box -50 0 3786 66
use sky130_fd_io__tk_em1o_CDNS_52468879185340  sky130_fd_io__tk_em1o_CDNS_52468879185340_0
timestamp 1704896540
transform 1 0 1813 0 1 10282
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_0
timestamp 1704896540
transform 0 -1 882 1 0 9251
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_1
timestamp 1704896540
transform 0 -1 370 1 0 9277
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_52468879185985  sky130_fd_io__tk_em1o_CDNS_52468879185985_2
timestamp 1704896540
transform 1 0 2512 0 1 8601
box 0 0 1 1
<< labels >>
flabel comment s 4422 12678 4422 12678 3 FreeSans 200 180 0 0 voutref
flabel comment s 1701 12677 1701 12677 3 FreeSans 200 0 0 0 voutref
flabel comment s 1222 10407 1222 10407 3 FreeSans 200 270 0 0 voutref
flabel comment s 1220 14 1220 14 3 FreeSans 200 90 0 0 voutref
flabel metal1 s 1691 12730 1721 12782 3 FreeSans 200 0 0 0 vgnd
port 2 nsew
flabel metal1 s 1691 12570 1721 12622 3 FreeSans 200 0 0 0 vgnd
port 2 nsew
flabel metal1 s 4399 12730 4434 12782 3 FreeSans 200 180 0 0 vgnd
port 2 nsew
flabel metal1 s 4399 12570 4434 12622 3 FreeSans 200 180 0 0 vgnd
port 2 nsew
flabel metal1 s 4287 12411 4328 12457 3 FreeSans 200 180 0 0 ngate
port 3 nsew
flabel metal1 s -547 10034 -513 10226 3 FreeSans 200 0 0 0 vgnd
port 2 nsew
flabel metal1 s -547 9013 -513 9146 3 FreeSans 200 0 0 0 vgnd
port 2 nsew
flabel metal1 s -547 10282 -513 10328 3 FreeSans 200 0 0 0 ngate
port 3 nsew
flabel metal2 s 972 0 1126 41 3 FreeSans 200 90 0 0 vgnd
port 2 nsew
flabel metal2 s 1512 0 1564 41 3 FreeSans 200 90 0 0 biasen_n
port 4 nsew
flabel metal2 s 4212 136 4434 177 3 FreeSans 200 90 0 0 vpwr_ka
port 5 nsew
flabel metal2 s 1296 0 1441 41 3 FreeSans 200 90 0 0 vgnd
port 2 nsew
flabel metal2 s 1944 0 2212 41 3 FreeSans 200 90 0 0 vgnd
port 2 nsew
flabel metal2 s 0 0 268 41 3 FreeSans 200 90 0 0 vgnd
port 2 nsew
flabel metal2 s 1620 0 1888 41 3 FreeSans 200 90 0 0 vgnd
port 2 nsew
flabel metal2 s 324 0 592 41 3 FreeSans 200 90 0 0 vgnd
port 2 nsew
flabel metal2 s 3596 136 3832 177 3 FreeSans 200 90 0 0 vgnd
port 2 nsew
flabel metal2 s 2592 0 2860 41 3 FreeSans 200 90 0 0 vgnd
port 2 nsew
flabel metal2 s 2916 0 3184 41 3 FreeSans 200 90 0 0 vgnd
port 2 nsew
flabel metal2 s 3240 136 3473 177 3 FreeSans 200 90 0 0 vgnd
port 2 nsew
flabel metal2 s 2268 0 2536 41 3 FreeSans 200 90 0 0 vgnd
port 2 nsew
<< properties >>
string GDS_END 80485516
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 80431718
string path -1.675 223.350 36.850 223.350 
<< end >>
