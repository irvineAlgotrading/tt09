magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< pwell >>
rect -76 -26 964 226
<< mvnnmos >>
rect 0 0 180 200
rect 236 0 416 200
rect 472 0 652 200
rect 708 0 888 200
<< mvndiff >>
rect -50 0 0 200
rect 416 182 472 200
rect 416 148 427 182
rect 461 148 472 182
rect 416 114 472 148
rect 416 80 427 114
rect 461 80 472 114
rect 416 46 472 80
rect 416 12 427 46
rect 461 12 472 46
rect 416 0 472 12
rect 888 0 938 200
<< mvndiffc >>
rect 427 148 461 182
rect 427 80 461 114
rect 427 12 461 46
<< poly >>
rect 0 200 180 226
rect 0 -26 180 0
rect 236 200 416 226
rect 472 200 652 226
rect 236 -26 416 0
rect 472 -26 652 0
rect 708 200 888 226
rect 708 -26 888 0
<< locali >>
rect 427 182 461 198
rect 427 114 461 148
rect 427 46 461 80
rect 427 -4 461 12
<< metal1 >>
rect -51 -16 -5 186
rect 185 -16 231 186
rect 657 -16 703 186
rect 893 -16 939 186
use DFM1sd2_CDNS_52468879185159  DFM1sd2_CDNS_52468879185159_0
timestamp 1704896540
transform 1 0 652 0 1 0
box -26 -26 82 226
use DFM1sd2_CDNS_52468879185159  DFM1sd2_CDNS_52468879185159_1
timestamp 1704896540
transform 1 0 180 0 1 0
box -26 -26 82 226
use hvDFL1sd2_CDNS_52468879185133  hvDFL1sd2_CDNS_52468879185133_0
timestamp 1704896540
transform 1 0 416 0 1 0
box 0 0 1 1
use hvDFM1sd_CDNS_52468879185147  hvDFM1sd_CDNS_52468879185147_0
timestamp 1704896540
transform -1 0 0 0 1 0
box -26 -26 79 226
use hvDFM1sd_CDNS_52468879185147  hvDFM1sd_CDNS_52468879185147_1
timestamp 1704896540
transform 1 0 888 0 1 0
box -26 -26 79 226
<< labels >>
flabel comment s -28 85 -28 85 0 FreeSans 300 0 0 0 S
flabel comment s 208 85 208 85 0 FreeSans 300 0 0 0 D
flabel comment s 444 97 444 97 0 FreeSans 300 0 0 0 S
flabel comment s 680 85 680 85 0 FreeSans 300 0 0 0 D
flabel comment s 916 85 916 85 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 86849270
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86846820
<< end >>
