magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< poly >>
rect 119 369 219 392
rect 119 335 152 369
rect 186 335 219 369
rect 119 274 219 335
rect 119 240 152 274
rect 186 240 219 274
rect 119 218 219 240
rect 275 369 375 392
rect 275 335 309 369
rect 343 335 375 369
rect 275 274 375 335
rect 275 240 309 274
rect 343 240 375 274
rect 275 218 375 240
<< polycont >>
rect 152 335 186 369
rect 152 240 186 274
rect 309 335 343 369
rect 309 240 343 274
<< locali >>
rect 74 556 108 594
rect 386 556 420 594
rect 230 472 264 510
rect 152 369 186 385
rect 152 279 186 317
rect 152 224 186 240
rect 309 369 343 385
rect 309 287 343 325
rect 309 224 343 240
rect 384 154 422 188
rect 72 24 110 58
<< viali >>
rect 74 594 108 628
rect 74 522 108 556
rect 386 594 420 628
rect 230 510 264 544
rect 386 522 420 556
rect 230 438 264 472
rect 152 335 186 351
rect 152 317 186 335
rect 152 274 186 279
rect 152 245 186 274
rect 309 335 343 359
rect 309 325 343 335
rect 309 274 343 287
rect 309 253 343 274
rect 350 154 384 188
rect 422 154 456 188
rect 38 24 72 58
rect 110 24 144 58
<< metal1 >>
rect 68 628 426 690
rect 68 594 74 628
rect 108 594 386 628
rect 420 594 426 628
rect 68 590 426 594
rect 68 556 114 590
tri 114 556 148 590 nw
tri 346 556 380 590 ne
rect 380 556 426 590
rect 68 522 74 556
rect 108 522 114 556
rect 68 510 114 522
rect 224 544 270 556
rect 224 510 230 544
rect 264 510 270 544
rect 380 522 386 556
rect 420 522 426 556
rect 224 478 270 510
tri 270 478 304 512 sw
rect 380 510 426 522
rect 224 472 426 478
rect 224 438 230 472
rect 264 438 426 472
rect 224 426 426 438
tri 346 392 380 426 ne
rect 146 351 192 363
rect 146 317 152 351
rect 186 317 192 351
rect 146 279 192 317
rect 146 245 152 279
rect 186 245 192 279
rect 146 233 192 245
rect 303 359 349 371
rect 303 325 309 359
rect 343 325 349 359
rect 303 287 349 325
rect 303 253 309 287
rect 343 253 349 287
rect 303 241 349 253
tri 346 194 380 228 se
rect 380 194 426 426
tri 426 194 460 228 sw
rect 338 188 468 194
rect 338 154 350 188
rect 384 154 422 188
rect 456 154 468 188
rect 338 148 468 154
rect 26 58 457 64
rect 26 24 38 58
rect 72 24 110 58
rect 144 24 457 58
rect 26 18 457 24
rect 68 0 457 18
use nfet_CDNS_52468879185814  nfet_CDNS_52468879185814_0
timestamp 1704896540
transform 1 0 119 0 1 36
box -82 -32 182 182
use nfet_CDNS_52468879185814  nfet_CDNS_52468879185814_1
timestamp 1704896540
transform 1 0 275 0 1 36
box -82 -32 182 182
use pfet_CDNS_52468879185725  pfet_CDNS_52468879185725_0
timestamp 1704896540
transform 1 0 275 0 -1 624
box -119 -66 219 266
use pfet_CDNS_52468879185725  pfet_CDNS_52468879185725_1
timestamp 1704896540
transform 1 0 119 0 -1 624
box -119 -66 219 266
<< properties >>
string GDS_END 25732846
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 25729942
string path 2.275 12.750 2.275 16.000 
<< end >>
