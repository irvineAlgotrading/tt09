magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< pwell >>
rect -26 -26 226 1026
<< ndiff >>
rect 0 930 60 1000
rect 140 930 200 1000
rect 0 896 11 930
rect 45 896 60 930
rect 140 896 155 930
rect 189 896 200 930
rect 0 862 60 896
rect 140 862 200 896
rect 0 828 11 862
rect 45 828 60 862
rect 140 828 155 862
rect 189 828 200 862
rect 0 794 60 828
rect 140 794 200 828
rect 0 760 11 794
rect 45 760 60 794
rect 140 760 155 794
rect 189 760 200 794
rect 0 726 60 760
rect 140 726 200 760
rect 0 692 11 726
rect 45 692 60 726
rect 140 692 155 726
rect 189 692 200 726
rect 0 658 60 692
rect 140 658 200 692
rect 0 624 11 658
rect 45 624 60 658
rect 140 624 155 658
rect 189 624 200 658
rect 0 590 60 624
rect 140 590 200 624
rect 0 556 11 590
rect 45 556 60 590
rect 140 556 155 590
rect 189 556 200 590
rect 0 522 60 556
rect 140 522 200 556
rect 0 488 11 522
rect 45 488 60 522
rect 140 488 155 522
rect 189 488 200 522
rect 0 454 60 488
rect 140 454 200 488
rect 0 420 11 454
rect 45 420 60 454
rect 140 420 155 454
rect 189 420 200 454
rect 0 386 60 420
rect 140 386 200 420
rect 0 352 11 386
rect 45 352 60 386
rect 140 352 155 386
rect 189 352 200 386
rect 0 318 60 352
rect 140 318 200 352
rect 0 284 11 318
rect 45 284 60 318
rect 140 284 155 318
rect 189 284 200 318
rect 0 250 60 284
rect 140 250 200 284
rect 0 216 11 250
rect 45 216 60 250
rect 140 216 155 250
rect 189 216 200 250
rect 0 182 60 216
rect 140 182 200 216
rect 0 148 11 182
rect 45 148 60 182
rect 140 148 155 182
rect 189 148 200 182
rect 0 114 60 148
rect 140 114 200 148
rect 0 80 11 114
rect 45 80 60 114
rect 140 80 155 114
rect 189 80 200 114
rect 0 46 60 80
rect 140 46 200 80
rect 0 12 11 46
rect 45 12 60 46
rect 140 12 155 46
rect 189 12 200 46
rect 0 0 60 12
rect 140 0 200 12
<< ndiffc >>
rect 11 896 45 930
rect 155 896 189 930
rect 11 828 45 862
rect 155 828 189 862
rect 11 760 45 794
rect 155 760 189 794
rect 11 692 45 726
rect 155 692 189 726
rect 11 624 45 658
rect 155 624 189 658
rect 11 556 45 590
rect 155 556 189 590
rect 11 488 45 522
rect 155 488 189 522
rect 11 420 45 454
rect 155 420 189 454
rect 11 352 45 386
rect 155 352 189 386
rect 11 284 45 318
rect 155 284 189 318
rect 11 216 45 250
rect 155 216 189 250
rect 11 148 45 182
rect 155 148 189 182
rect 11 80 45 114
rect 155 80 189 114
rect 11 12 45 46
rect 155 12 189 46
<< psubdiff >>
rect 60 930 140 1000
rect 60 896 83 930
rect 117 896 140 930
rect 60 862 140 896
rect 60 828 83 862
rect 117 828 140 862
rect 60 794 140 828
rect 60 760 83 794
rect 117 760 140 794
rect 60 726 140 760
rect 60 692 83 726
rect 117 692 140 726
rect 60 658 140 692
rect 60 624 83 658
rect 117 624 140 658
rect 60 590 140 624
rect 60 556 83 590
rect 117 556 140 590
rect 60 522 140 556
rect 60 488 83 522
rect 117 488 140 522
rect 60 454 140 488
rect 60 420 83 454
rect 117 420 140 454
rect 60 386 140 420
rect 60 352 83 386
rect 117 352 140 386
rect 60 318 140 352
rect 60 284 83 318
rect 117 284 140 318
rect 60 250 140 284
rect 60 216 83 250
rect 117 216 140 250
rect 60 182 140 216
rect 60 148 83 182
rect 117 148 140 182
rect 60 114 140 148
rect 60 80 83 114
rect 117 80 140 114
rect 60 46 140 80
rect 60 12 83 46
rect 117 12 140 46
rect 60 0 140 12
<< psubdiffcont >>
rect 83 896 117 930
rect 83 828 117 862
rect 83 760 117 794
rect 83 692 117 726
rect 83 624 117 658
rect 83 556 117 590
rect 83 488 117 522
rect 83 420 117 454
rect 83 352 117 386
rect 83 284 117 318
rect 83 216 117 250
rect 83 148 117 182
rect 83 80 117 114
rect 83 12 117 46
<< locali >>
rect 11 930 189 946
rect 45 896 83 930
rect 117 896 155 930
rect 11 862 189 896
rect 45 828 83 862
rect 117 828 155 862
rect 11 794 189 828
rect 45 760 83 794
rect 117 760 155 794
rect 11 726 189 760
rect 45 692 83 726
rect 117 692 155 726
rect 11 658 189 692
rect 45 624 83 658
rect 117 624 155 658
rect 11 590 189 624
rect 45 556 83 590
rect 117 556 155 590
rect 11 522 189 556
rect 45 488 83 522
rect 117 488 155 522
rect 11 454 189 488
rect 45 420 83 454
rect 117 420 155 454
rect 11 386 189 420
rect 45 352 83 386
rect 117 352 155 386
rect 11 318 189 352
rect 45 284 83 318
rect 117 284 155 318
rect 11 250 189 284
rect 45 216 83 250
rect 117 216 155 250
rect 11 182 189 216
rect 45 148 83 182
rect 117 148 155 182
rect 11 114 189 148
rect 45 80 83 114
rect 117 80 155 114
rect 11 46 189 80
rect 45 12 83 46
rect 117 12 155 46
rect 11 -4 189 12
<< properties >>
string GDS_END 42978856
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 42975588
<< end >>
