magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< metal4 >>
rect 0 35157 254 40000
rect 14746 35157 15000 40000
rect 0 14007 254 19000
rect 6904 14009 8104 14209
rect 14746 14007 15000 19000
<< metal5 >>
rect 0 35157 254 40000
rect 14746 35157 15000 40000
rect 2000 20574 12990 33596
rect 0 14007 254 18997
rect 14746 14007 15000 18997
use sky130_ef_io__minesd_pad_and_pg  sky130_ef_io__minesd_pad_and_pg_0
timestamp 1704896540
transform 1 0 -8 0 1 13
box 8 13994 15008 39987
<< labels >>
flabel metal4 s 0 35157 254 40000 3 FreeSans 1015 0 0 0 VSSIO
port 4 nsew
flabel metal4 s 14746 35157 15000 40000 3 FreeSans 1015 180 0 0 VSSIO
port 4 nsew
flabel metal4 s 6904 14009 8104 14209 0 FreeSans 1400 0 0 0 P_CORE
port 1 nsew
flabel metal5 s 2000 20574 12990 33596 0 FreeSans 3906 0 0 0 P_PAD
port 2 nsew
flabel metal5 s 14746 14007 15000 18997 3 FreeSans 1015 180 0 0 VDDIO
port 3 nsew
flabel metal5 s 0 14007 254 18997 3 FreeSans 1015 0 0 0 VDDIO
port 3 nsew
flabel metal4 s 14746 14007 15000 19000 3 FreeSans 1015 180 0 0 VDDIO
port 3 nsew
flabel metal4 s 0 14007 254 19000 3 FreeSans 1015 0 0 0 VDDIO
port 3 nsew
flabel metal5 s 0 35157 254 40000 3 FreeSans 1015 0 0 0 VSSIO
port 4 nsew
flabel metal5 s 14746 35157 15000 40000 3 FreeSans 1015 180 0 0 VSSIO
port 4 nsew
flabel metal4 s 14873 37578 14873 37578 3 FreeSans 1015 180 0 0 VSSIO
flabel metal4 s 127 37578 127 37578 3 FreeSans 1015 0 0 0 VSSIO
<< properties >>
string GDS_END 7537876
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io__analog.gds
string GDS_START 7535634
<< end >>
