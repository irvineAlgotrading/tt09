magic
tech sky130B
timestamp 1704896540
<< metal1 >>
rect 0 0 3 218
rect 189 0 192 218
<< via1 >>
rect 3 0 189 218
<< metal2 >>
rect 0 0 3 218
rect 189 0 192 218
<< properties >>
string GDS_END 86909422
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86906602
<< end >>
