magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< pwell >>
rect -79 -26 196 166
<< mvnmos >>
rect 0 0 120 140
<< mvndiff >>
rect -53 114 0 140
rect -53 80 -45 114
rect -11 80 0 114
rect -53 46 0 80
rect -53 12 -45 46
rect -11 12 0 46
rect -53 0 0 12
rect 120 0 170 140
<< mvndiffc >>
rect -45 80 -11 114
rect -45 12 -11 46
<< poly >>
rect 0 140 120 166
rect 0 -26 120 0
<< locali >>
rect -45 114 -11 130
rect -45 46 -11 80
rect -45 -4 -11 12
use DFL1sd_CDNS_5246887918531  DFL1sd_CDNS_5246887918531_0
timestamp 1704896540
transform -1 0 0 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s -28 63 -28 63 0 FreeSans 300 0 0 0 S
flabel comment s 145 70 145 70 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 4320
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 3548
<< end >>
