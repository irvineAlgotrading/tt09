magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -66 377 738 897
<< pwell >>
rect 402 217 668 283
rect 58 43 668 217
rect -26 -43 698 43
<< mvnmos >>
rect 141 107 241 191
rect 297 107 397 191
rect 485 107 585 257
<< mvpmos >>
rect 141 443 241 527
rect 283 443 383 527
rect 485 443 585 743
<< mvndiff >>
rect 428 249 485 257
rect 428 215 440 249
rect 474 215 485 249
rect 428 191 485 215
rect 84 166 141 191
rect 84 132 96 166
rect 130 132 141 166
rect 84 107 141 132
rect 241 166 297 191
rect 241 132 252 166
rect 286 132 297 166
rect 241 107 297 132
rect 397 149 485 191
rect 397 115 440 149
rect 474 115 485 149
rect 397 107 485 115
rect 585 249 642 257
rect 585 215 596 249
rect 630 215 642 249
rect 585 149 642 215
rect 585 115 596 149
rect 630 115 642 149
rect 585 107 642 115
<< mvpdiff >>
rect 428 735 485 743
rect 428 701 440 735
rect 474 701 485 735
rect 428 652 485 701
rect 428 618 440 652
rect 474 618 485 652
rect 428 568 485 618
rect 428 534 440 568
rect 474 534 485 568
rect 428 527 485 534
rect 84 502 141 527
rect 84 468 96 502
rect 130 468 141 502
rect 84 443 141 468
rect 241 443 283 527
rect 383 485 485 527
rect 383 451 440 485
rect 474 451 485 485
rect 383 443 485 451
rect 585 735 642 743
rect 585 701 596 735
rect 630 701 642 735
rect 585 652 642 701
rect 585 618 596 652
rect 630 618 642 652
rect 585 568 642 618
rect 585 534 596 568
rect 630 534 642 568
rect 585 485 642 534
rect 585 451 596 485
rect 630 451 642 485
rect 585 443 642 451
<< mvndiffc >>
rect 440 215 474 249
rect 96 132 130 166
rect 252 132 286 166
rect 440 115 474 149
rect 596 215 630 249
rect 596 115 630 149
<< mvpdiffc >>
rect 440 701 474 735
rect 440 618 474 652
rect 440 534 474 568
rect 96 468 130 502
rect 440 451 474 485
rect 596 701 630 735
rect 596 618 630 652
rect 596 534 630 568
rect 596 451 630 485
<< mvpsubdiff >>
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 672 831
<< mvpsubdiffcont >>
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
<< poly >>
rect 485 743 585 769
rect 141 527 241 553
rect 283 527 383 553
rect 141 361 241 443
rect 117 341 241 361
rect 117 307 137 341
rect 171 307 241 341
rect 117 273 241 307
rect 117 239 137 273
rect 171 239 241 273
rect 117 217 241 239
rect 283 361 383 443
rect 485 395 585 443
rect 485 361 505 395
rect 539 361 585 395
rect 283 341 397 361
rect 283 307 322 341
rect 356 307 397 341
rect 283 273 397 307
rect 283 239 322 273
rect 356 239 397 273
rect 485 257 585 361
rect 283 217 397 239
rect 141 191 241 217
rect 297 191 397 217
rect 141 81 241 107
rect 297 81 397 107
rect 485 81 585 107
<< polycont >>
rect 137 307 171 341
rect 137 239 171 273
rect 505 361 539 395
rect 322 307 356 341
rect 322 239 356 273
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 672 831
rect 166 735 560 751
rect 200 701 238 735
rect 272 701 310 735
rect 344 701 382 735
rect 416 701 440 735
rect 488 701 526 735
rect 166 652 560 701
rect 166 618 440 652
rect 474 618 560 652
rect 166 568 560 618
rect 80 502 130 535
rect 80 468 96 502
rect 80 415 130 468
rect 166 534 440 568
rect 474 534 560 568
rect 166 485 560 534
rect 166 451 440 485
rect 474 451 560 485
rect 596 735 647 751
rect 630 701 647 735
rect 596 652 647 701
rect 630 618 647 652
rect 596 568 647 618
rect 630 534 647 568
rect 596 485 647 534
rect 630 451 647 485
rect 80 395 555 415
rect 80 381 505 395
rect 121 341 187 345
rect 121 307 137 341
rect 171 307 187 341
rect 121 273 187 307
rect 121 239 137 273
rect 171 239 187 273
rect 121 235 187 239
rect 236 199 270 381
rect 489 361 505 381
rect 539 361 555 395
rect 489 345 555 361
rect 306 341 372 345
rect 306 307 322 341
rect 356 307 372 341
rect 306 273 372 307
rect 306 239 322 273
rect 356 239 372 273
rect 306 235 372 239
rect 408 249 526 265
rect 408 215 440 249
rect 474 215 526 249
rect 18 166 200 199
rect 18 132 96 166
rect 130 132 200 166
rect 18 113 200 132
rect 18 79 20 113
rect 54 79 92 113
rect 126 79 164 113
rect 198 79 200 113
rect 236 166 302 199
rect 236 132 252 166
rect 286 132 302 166
rect 236 99 302 132
rect 408 149 526 215
rect 408 115 440 149
rect 474 115 526 149
rect 408 113 526 115
rect 18 73 200 79
rect 408 79 414 113
rect 448 79 486 113
rect 520 79 526 113
rect 596 249 647 451
rect 630 215 647 249
rect 596 149 647 215
rect 630 115 647 149
rect 596 99 647 115
rect 408 73 526 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 166 701 200 735
rect 238 701 272 735
rect 310 701 344 735
rect 382 701 416 735
rect 454 701 474 735
rect 474 701 488 735
rect 526 701 560 735
rect 20 79 54 113
rect 92 79 126 113
rect 164 79 198 113
rect 414 79 448 113
rect 486 79 520 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
<< metal1 >>
rect 0 831 672 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 672 831
rect 0 791 672 797
rect 0 735 672 763
rect 0 701 166 735
rect 200 701 238 735
rect 272 701 310 735
rect 344 701 382 735
rect 416 701 454 735
rect 488 701 526 735
rect 560 701 672 735
rect 0 689 672 701
rect 0 113 672 125
rect 0 79 20 113
rect 54 79 92 113
rect 126 79 164 113
rect 198 79 414 113
rect 448 79 486 113
rect 520 79 672 113
rect 0 51 672 79
rect 0 17 672 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 672 17
rect 0 -23 672 -17
<< labels >>
rlabel comment s 0 0 0 0 4 or2_1
flabel metal1 s 0 51 672 125 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel metal1 s 0 0 672 23 0 FreeSans 340 0 0 0 VNB
port 4 nsew ground bidirectional
flabel metal1 s 0 689 672 763 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 791 672 814 0 FreeSans 340 0 0 0 VPB
port 5 nsew power bidirectional
flabel locali s 319 242 353 276 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 607 168 641 202 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 607 242 641 276 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 607 464 641 498 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 607 538 641 572 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 607 612 641 646 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 127 242 161 276 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 672 814
string GDS_END 376290
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 367608
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
<< end >>
