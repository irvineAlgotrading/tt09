magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< pwell >>
rect 18 4654 188 4742
rect 18 4632 120 4654
rect 0 3632 120 4632
rect 2632 4136 2880 4254
rect 4312 4136 4432 4632
rect 2232 4010 2352 4128
rect 1752 3876 1872 4002
rect 1552 3758 1872 3876
rect 1832 3750 1872 3758
rect 1832 3632 1952 3750
rect 0 -97 120 903
rect 1832 785 1952 903
rect 1832 777 1872 785
rect 1552 659 1872 777
rect 1752 533 1872 659
rect 2232 407 2352 525
rect 2632 281 2880 399
rect 4312 -97 4432 399
<< mvndiff >>
rect 26 4590 94 4606
rect 26 4556 34 4590
rect 68 4556 94 4590
rect 26 4540 94 4556
rect 4338 4590 4406 4606
rect 4338 4556 4364 4590
rect 4398 4556 4406 4590
rect 4338 4540 4406 4556
rect 26 4464 94 4480
rect 26 4430 34 4464
rect 68 4430 94 4464
rect 26 4414 94 4430
rect 4338 4464 4406 4480
rect 4338 4430 4364 4464
rect 4398 4430 4406 4464
rect 4338 4414 4406 4430
rect 26 4338 94 4354
rect 26 4304 34 4338
rect 68 4304 94 4338
rect 26 4288 94 4304
rect 4338 4338 4406 4354
rect 4338 4304 4364 4338
rect 4398 4304 4406 4338
rect 4338 4288 4406 4304
rect 26 4212 94 4228
rect 26 4178 34 4212
rect 68 4178 94 4212
rect 26 4162 94 4178
rect 2658 4212 2726 4228
rect 2658 4178 2684 4212
rect 2718 4178 2726 4212
rect 2658 4162 2726 4178
rect 2786 4212 2854 4228
rect 2786 4178 2794 4212
rect 2828 4178 2854 4212
rect 2786 4162 2854 4178
rect 4338 4212 4406 4228
rect 4338 4178 4364 4212
rect 4398 4178 4406 4212
rect 4338 4162 4406 4178
rect 26 4086 94 4102
rect 26 4052 34 4086
rect 68 4052 94 4086
rect 26 4036 94 4052
rect 2258 4086 2326 4102
rect 2258 4052 2284 4086
rect 2318 4052 2326 4086
rect 2258 4036 2326 4052
rect 26 3960 94 3976
rect 26 3926 34 3960
rect 68 3926 94 3960
rect 26 3910 94 3926
rect 1778 3960 1846 3976
rect 1778 3926 1804 3960
rect 1838 3926 1846 3960
rect 1778 3910 1846 3926
rect 26 3834 94 3850
rect 26 3800 34 3834
rect 68 3800 94 3834
rect 26 3784 94 3800
rect 1578 3834 1646 3850
rect 1578 3800 1604 3834
rect 1638 3800 1646 3834
rect 1578 3784 1646 3800
rect 26 3708 94 3724
rect 26 3674 34 3708
rect 68 3674 94 3708
rect 26 3658 94 3674
rect 1858 3708 1926 3724
rect 1858 3674 1884 3708
rect 1918 3674 1926 3708
rect 1858 3658 1926 3674
rect 26 861 94 877
rect 26 827 34 861
rect 68 827 94 861
rect 26 811 94 827
rect 1858 861 1926 877
rect 1858 827 1884 861
rect 1918 827 1926 861
rect 1858 811 1926 827
rect 26 735 94 751
rect 26 701 34 735
rect 68 701 94 735
rect 26 685 94 701
rect 1578 735 1646 751
rect 1578 701 1604 735
rect 1638 701 1646 735
rect 1578 685 1646 701
rect 26 609 94 625
rect 26 575 34 609
rect 68 575 94 609
rect 26 559 94 575
rect 1778 609 1846 625
rect 1778 575 1804 609
rect 1838 575 1846 609
rect 1778 559 1846 575
rect 26 483 94 499
rect 26 449 34 483
rect 68 449 94 483
rect 26 433 94 449
rect 2258 483 2326 499
rect 2258 449 2284 483
rect 2318 449 2326 483
rect 2258 433 2326 449
rect 26 357 94 373
rect 26 323 34 357
rect 68 323 94 357
rect 26 307 94 323
rect 2658 357 2726 373
rect 2658 323 2684 357
rect 2718 323 2726 357
rect 2658 307 2726 323
rect 2786 357 2854 373
rect 2786 323 2794 357
rect 2828 323 2854 357
rect 2786 307 2854 323
rect 4338 357 4406 373
rect 4338 323 4364 357
rect 4398 323 4406 357
rect 4338 307 4406 323
rect 26 231 94 247
rect 26 197 34 231
rect 68 197 94 231
rect 26 181 94 197
rect 4338 231 4406 247
rect 4338 197 4364 231
rect 4398 197 4406 231
rect 4338 181 4406 197
rect 26 105 94 121
rect 26 71 34 105
rect 68 71 94 105
rect 26 55 94 71
rect 4338 105 4406 121
rect 4338 71 4364 105
rect 4398 71 4406 105
rect 4338 55 4406 71
rect 26 -21 94 -5
rect 26 -55 34 -21
rect 68 -55 94 -21
rect 26 -71 94 -55
rect 4338 -21 4406 -5
rect 4338 -55 4364 -21
rect 4398 -55 4406 -21
rect 4338 -71 4406 -55
<< mvndiffc >>
rect 34 4556 68 4590
rect 4364 4556 4398 4590
rect 34 4430 68 4464
rect 4364 4430 4398 4464
rect 34 4304 68 4338
rect 4364 4304 4398 4338
rect 34 4178 68 4212
rect 2684 4178 2718 4212
rect 2794 4178 2828 4212
rect 4364 4178 4398 4212
rect 34 4052 68 4086
rect 2284 4052 2318 4086
rect 34 3926 68 3960
rect 1804 3926 1838 3960
rect 34 3800 68 3834
rect 1604 3800 1638 3834
rect 34 3674 68 3708
rect 1884 3674 1918 3708
rect 34 827 68 861
rect 1884 827 1918 861
rect 34 701 68 735
rect 1604 701 1638 735
rect 34 575 68 609
rect 1804 575 1838 609
rect 34 449 68 483
rect 2284 449 2318 483
rect 34 323 68 357
rect 2684 323 2718 357
rect 2794 323 2828 357
rect 4364 323 4398 357
rect 34 197 68 231
rect 4364 197 4398 231
rect 34 71 68 105
rect 4364 71 4398 105
rect 34 -55 68 -21
rect 4364 -55 4398 -21
<< locali >>
rect 34 4590 164 4606
rect 84 4556 122 4590
rect 156 4556 164 4590
rect 34 4540 164 4556
rect 4262 4593 4398 4606
rect 4262 4559 4280 4593
rect 4314 4559 4352 4593
rect 4386 4590 4398 4593
rect 4262 4556 4364 4559
rect 4262 4540 4398 4556
rect 34 4464 164 4480
rect 80 4430 118 4464
rect 152 4430 164 4464
rect 34 4414 164 4430
rect 4268 4464 4398 4480
rect 4268 4430 4280 4464
rect 4314 4430 4352 4464
rect 4268 4414 4398 4430
rect 34 4338 164 4354
rect 80 4304 118 4338
rect 152 4304 164 4338
rect 34 4288 164 4304
rect 4268 4338 4398 4354
rect 4268 4304 4280 4338
rect 4314 4304 4352 4338
rect 4268 4288 4398 4304
rect 34 4212 164 4228
rect 80 4178 118 4212
rect 152 4178 164 4212
rect 34 4162 164 4178
rect 2588 4212 2718 4228
rect 2588 4178 2600 4212
rect 2634 4178 2672 4212
rect 2588 4162 2718 4178
rect 2794 4212 2924 4228
rect 2840 4178 2878 4212
rect 2912 4178 2924 4212
rect 2794 4162 2924 4178
rect 4268 4212 4398 4228
rect 4268 4178 4280 4212
rect 4314 4178 4352 4212
rect 4268 4162 4398 4178
rect 34 4086 164 4102
rect 80 4052 118 4086
rect 152 4052 164 4086
rect 34 4036 164 4052
rect 2188 4086 2318 4102
rect 2188 4052 2200 4086
rect 2234 4052 2272 4086
rect 2188 4036 2318 4052
rect 34 3960 164 3976
rect 80 3926 118 3960
rect 152 3926 164 3960
rect 34 3910 164 3926
rect 1708 3960 1838 3976
rect 1708 3926 1720 3960
rect 1754 3926 1792 3960
rect 1708 3910 1838 3926
rect 34 3834 164 3850
rect 80 3800 118 3834
rect 152 3800 164 3834
rect 34 3784 164 3800
rect 1508 3834 1638 3850
rect 1508 3800 1520 3834
rect 1554 3800 1592 3834
rect 1508 3784 1638 3800
rect 34 3708 164 3724
rect 80 3674 118 3708
rect 152 3674 164 3708
rect 34 3658 164 3674
rect 1788 3708 1918 3724
rect 1788 3674 1800 3708
rect 1834 3674 1872 3708
rect 1788 3658 1918 3674
rect 34 861 164 877
rect 80 827 118 861
rect 152 827 164 861
rect 34 811 164 827
rect 1788 861 1918 877
rect 1788 827 1800 861
rect 1834 827 1872 861
rect 1788 811 1918 827
rect 34 735 164 751
rect 80 701 118 735
rect 152 701 164 735
rect 34 685 164 701
rect 1508 735 1638 751
rect 1508 701 1520 735
rect 1554 701 1592 735
rect 1508 685 1638 701
rect 34 609 164 625
rect 80 575 118 609
rect 152 575 164 609
rect 34 559 164 575
rect 1708 609 1838 625
rect 1708 575 1720 609
rect 1754 575 1792 609
rect 1708 559 1838 575
rect 34 483 164 499
rect 80 449 118 483
rect 152 449 164 483
rect 34 433 164 449
rect 2188 483 2318 499
rect 2188 449 2200 483
rect 2234 449 2272 483
rect 2188 433 2318 449
rect 34 357 164 373
rect 80 323 118 357
rect 152 323 164 357
rect 34 307 164 323
rect 2588 357 2718 373
rect 2588 323 2600 357
rect 2634 323 2672 357
rect 2588 307 2718 323
rect 2794 357 2924 373
rect 2840 323 2878 357
rect 2912 323 2924 357
rect 2794 307 2924 323
rect 4268 357 4398 373
rect 4268 323 4280 357
rect 4314 323 4352 357
rect 4268 307 4398 323
rect 34 231 164 247
rect 80 197 118 231
rect 152 197 164 231
rect 34 181 164 197
rect 4268 231 4398 247
rect 4268 197 4280 231
rect 4314 197 4352 231
rect 4268 181 4398 197
rect 34 105 164 121
rect 80 71 118 105
rect 152 71 164 105
rect 34 55 164 71
rect 4268 105 4398 121
rect 4268 71 4280 105
rect 4314 71 4352 105
rect 4268 55 4398 71
rect 34 -21 164 -5
rect 84 -55 122 -21
rect 156 -55 164 -21
rect 34 -71 164 -55
rect 4262 -21 4398 -5
rect 4296 -55 4334 -21
rect 4262 -71 4398 -55
<< viali >>
rect 50 4556 68 4590
rect 68 4556 84 4590
rect 122 4556 156 4590
rect 4280 4559 4314 4593
rect 4352 4590 4386 4593
rect 4352 4559 4364 4590
rect 4364 4559 4386 4590
rect 46 4430 68 4464
rect 68 4430 80 4464
rect 118 4430 152 4464
rect 4280 4430 4314 4464
rect 4352 4430 4364 4464
rect 4364 4430 4386 4464
rect 46 4304 68 4338
rect 68 4304 80 4338
rect 118 4304 152 4338
rect 4280 4304 4314 4338
rect 4352 4304 4364 4338
rect 4364 4304 4386 4338
rect 46 4178 68 4212
rect 68 4178 80 4212
rect 118 4178 152 4212
rect 2600 4178 2634 4212
rect 2672 4178 2684 4212
rect 2684 4178 2706 4212
rect 2806 4178 2828 4212
rect 2828 4178 2840 4212
rect 2878 4178 2912 4212
rect 4280 4178 4314 4212
rect 4352 4178 4364 4212
rect 4364 4178 4386 4212
rect 46 4052 68 4086
rect 68 4052 80 4086
rect 118 4052 152 4086
rect 2200 4052 2234 4086
rect 2272 4052 2284 4086
rect 2284 4052 2306 4086
rect 46 3926 68 3960
rect 68 3926 80 3960
rect 118 3926 152 3960
rect 1720 3926 1754 3960
rect 1792 3926 1804 3960
rect 1804 3926 1826 3960
rect 46 3800 68 3834
rect 68 3800 80 3834
rect 118 3800 152 3834
rect 1520 3800 1554 3834
rect 1592 3800 1604 3834
rect 1604 3800 1626 3834
rect 46 3674 68 3708
rect 68 3674 80 3708
rect 118 3674 152 3708
rect 1800 3674 1834 3708
rect 1872 3674 1884 3708
rect 1884 3674 1906 3708
rect 46 827 68 861
rect 68 827 80 861
rect 118 827 152 861
rect 1800 827 1834 861
rect 1872 827 1884 861
rect 1884 827 1906 861
rect 46 701 68 735
rect 68 701 80 735
rect 118 701 152 735
rect 1520 701 1554 735
rect 1592 701 1604 735
rect 1604 701 1626 735
rect 46 575 68 609
rect 68 575 80 609
rect 118 575 152 609
rect 1720 575 1754 609
rect 1792 575 1804 609
rect 1804 575 1826 609
rect 46 449 68 483
rect 68 449 80 483
rect 118 449 152 483
rect 2200 449 2234 483
rect 2272 449 2284 483
rect 2284 449 2306 483
rect 46 323 68 357
rect 68 323 80 357
rect 118 323 152 357
rect 2600 323 2634 357
rect 2672 323 2684 357
rect 2684 323 2706 357
rect 2806 323 2828 357
rect 2828 323 2840 357
rect 2878 323 2912 357
rect 4280 323 4314 357
rect 4352 323 4364 357
rect 4364 323 4386 357
rect 46 197 68 231
rect 68 197 80 231
rect 118 197 152 231
rect 4280 197 4314 231
rect 4352 197 4364 231
rect 4364 197 4386 231
rect 46 71 68 105
rect 68 71 80 105
rect 118 71 152 105
rect 4280 71 4314 105
rect 4352 71 4364 105
rect 4364 71 4386 105
rect 50 -55 68 -21
rect 68 -55 84 -21
rect 122 -55 156 -21
rect 4262 -55 4296 -21
rect 4334 -55 4364 -21
rect 4364 -55 4368 -21
<< metal1 >>
rect 44 4590 162 4602
rect 44 4556 50 4590
rect 84 4556 122 4590
rect 156 4556 162 4590
rect 44 4544 162 4556
rect 4274 4593 4392 4605
rect 4274 4559 4280 4593
rect 4314 4559 4352 4593
rect 4386 4559 4392 4593
rect 4274 4533 4392 4559
rect 4275 4531 4391 4532
rect 4274 4495 4392 4531
rect 4275 4494 4391 4495
tri 4257 4476 4274 4493 se
rect 4274 4476 4392 4493
rect 40 4468 158 4476
tri 158 4468 166 4476 sw
tri 4249 4468 4257 4476 se
rect 4257 4468 4392 4476
rect 40 4464 2196 4468
rect 40 4430 46 4464
rect 80 4430 118 4464
rect 152 4430 2196 4464
rect 40 4426 2196 4430
rect 2197 4427 2198 4467
rect 2234 4427 2235 4467
rect 2236 4464 4392 4468
rect 2236 4430 4280 4464
rect 4314 4430 4352 4464
rect 4386 4430 4392 4464
rect 2236 4426 4392 4430
rect 40 4418 175 4426
tri 175 4418 183 4426 nw
tri 4266 4418 4274 4426 ne
rect 4274 4418 4392 4426
rect 40 4342 158 4418
tri 158 4401 175 4418 nw
tri 158 4342 183 4367 sw
tri 4266 4342 4274 4350 se
rect 4274 4342 4392 4350
rect 40 4338 2196 4342
rect 40 4304 46 4338
rect 80 4304 118 4338
rect 152 4304 2196 4338
rect 40 4300 2196 4304
rect 2197 4301 2198 4341
rect 2234 4301 2235 4341
rect 2236 4338 4392 4342
rect 2236 4304 4280 4338
rect 4314 4304 4352 4338
rect 4386 4304 4392 4338
rect 2236 4300 4392 4304
rect 40 4292 158 4300
tri 158 4292 166 4300 nw
tri 4249 4292 4257 4300 ne
rect 4257 4292 4392 4300
tri 4257 4275 4274 4292 ne
tri 4257 4224 4274 4241 se
rect 4274 4224 4392 4292
rect 40 4216 158 4224
tri 158 4216 166 4224 sw
tri 2586 4216 2594 4224 se
rect 2594 4216 2918 4224
tri 2918 4216 2926 4224 sw
tri 4249 4216 4257 4224 se
rect 4257 4216 4392 4224
rect 40 4212 1356 4216
rect 1358 4215 1394 4216
rect 40 4178 46 4212
rect 80 4178 118 4212
rect 152 4178 1356 4212
rect 40 4174 1356 4178
rect 1357 4175 1395 4215
rect 1396 4212 3576 4216
rect 1396 4178 2600 4212
rect 2634 4178 2672 4212
rect 2706 4178 2806 4212
rect 2840 4178 2878 4212
rect 2912 4178 3576 4212
rect 1358 4174 1394 4175
rect 1396 4174 3576 4178
rect 3577 4175 3578 4215
rect 3614 4175 3615 4215
rect 3616 4212 4392 4216
rect 3616 4178 4280 4212
rect 4314 4178 4352 4212
rect 4386 4178 4392 4212
rect 3616 4174 4392 4178
rect 40 4090 158 4174
tri 158 4149 183 4174 nw
tri 2586 4166 2594 4174 ne
rect 2594 4166 2918 4174
tri 2918 4166 2926 4174 nw
tri 4266 4166 4274 4174 ne
rect 4274 4166 4392 4174
tri 158 4090 183 4115 sw
tri 2186 4090 2194 4098 se
rect 2194 4090 2312 4098
rect 40 4086 1156 4090
rect 40 4052 46 4086
rect 80 4052 118 4086
rect 152 4052 1156 4086
rect 40 4048 1156 4052
rect 1157 4049 1158 4089
rect 1194 4049 1195 4089
rect 1196 4086 2312 4090
rect 1196 4052 2200 4086
rect 2234 4052 2272 4086
rect 2306 4052 2312 4086
rect 1196 4048 2312 4052
rect 40 4040 158 4048
tri 158 4040 166 4048 nw
tri 1689 4040 1697 4048 ne
rect 1697 4040 1832 4048
tri 1697 4023 1714 4040 ne
tri 1697 3972 1714 3989 se
rect 1714 3972 1832 4040
tri 1832 4023 1857 4048 nw
tri 2186 4040 2194 4048 ne
rect 2194 4040 2312 4048
rect 40 3964 158 3972
tri 158 3964 166 3972 sw
tri 1689 3964 1697 3972 se
rect 1697 3964 1832 3972
rect 40 3960 916 3964
rect 40 3926 46 3960
rect 80 3926 118 3960
rect 152 3926 916 3960
rect 40 3922 916 3926
rect 917 3923 918 3963
rect 954 3923 955 3963
rect 956 3960 1832 3964
rect 956 3926 1720 3960
rect 1754 3926 1792 3960
rect 1826 3926 1832 3960
rect 956 3922 1832 3926
rect 40 3914 175 3922
tri 175 3914 183 3922 nw
tri 1706 3914 1714 3922 ne
rect 1714 3914 1832 3922
rect 40 3838 158 3914
tri 158 3897 175 3914 nw
tri 158 3838 183 3863 sw
tri 1506 3838 1514 3846 se
rect 1514 3838 1632 3846
rect 40 3834 816 3838
rect 40 3800 46 3834
rect 80 3800 118 3834
rect 152 3800 816 3834
rect 40 3796 816 3800
rect 817 3797 818 3837
rect 854 3797 855 3837
rect 856 3834 1632 3838
rect 856 3800 1520 3834
rect 1554 3800 1592 3834
rect 1626 3800 1632 3834
rect 856 3796 1632 3800
rect 40 3788 158 3796
tri 158 3788 166 3796 nw
tri 1489 3788 1497 3796 ne
rect 1497 3788 1632 3796
tri 1497 3771 1514 3788 ne
rect 40 3635 46 3751
rect 98 3720 104 3751
tri 1497 3720 1514 3737 se
rect 1514 3720 1632 3788
rect 98 3712 158 3720
tri 158 3712 166 3720 sw
tri 1489 3712 1497 3720 se
rect 1497 3712 1632 3720
tri 1632 3712 1657 3737 sw
tri 1786 3712 1794 3720 se
rect 1794 3712 1912 3720
rect 98 3708 956 3712
rect 958 3711 994 3712
rect 98 3699 118 3708
rect 80 3687 118 3699
rect 98 3674 118 3687
rect 152 3674 956 3708
rect 98 3670 956 3674
rect 957 3671 995 3711
rect 996 3708 1912 3712
rect 996 3674 1800 3708
rect 1834 3674 1872 3708
rect 1906 3674 1912 3708
rect 958 3670 994 3671
rect 996 3670 1912 3674
rect 98 3662 158 3670
tri 158 3662 166 3670 nw
tri 1786 3662 1794 3670 ne
rect 1794 3662 1912 3670
rect 98 3635 104 3662
rect 40 784 46 900
rect 98 873 104 900
rect 98 865 158 873
tri 158 865 166 873 sw
tri 1786 865 1794 873 se
rect 1794 865 1912 873
rect 98 861 956 865
rect 958 864 994 865
rect 98 848 118 861
rect 80 836 118 848
rect 98 827 118 836
rect 152 827 956 861
rect 98 823 956 827
rect 957 824 995 864
rect 996 861 1912 865
rect 996 827 1800 861
rect 1834 827 1872 861
rect 1906 827 1912 861
rect 958 823 994 824
rect 996 823 1912 827
rect 98 815 158 823
tri 158 815 166 823 nw
tri 1489 815 1497 823 ne
rect 1497 815 1632 823
rect 98 784 104 815
tri 1497 798 1514 815 ne
tri 1497 747 1514 764 se
rect 1514 747 1632 815
tri 1632 798 1657 823 nw
tri 1786 815 1794 823 ne
rect 1794 815 1912 823
rect 40 739 158 747
tri 158 739 166 747 sw
tri 1489 739 1497 747 se
rect 1497 739 1632 747
rect 40 735 816 739
rect 40 701 46 735
rect 80 701 118 735
rect 152 701 816 735
rect 40 697 816 701
rect 817 698 818 738
rect 854 698 855 738
rect 856 735 1632 739
rect 856 701 1520 735
rect 1554 701 1592 735
rect 1626 701 1632 735
rect 856 697 1632 701
rect 40 613 158 697
tri 158 672 183 697 nw
tri 1506 689 1514 697 ne
rect 1514 689 1632 697
tri 158 613 183 638 sw
tri 1706 613 1714 621 se
rect 1714 613 1832 621
rect 40 609 916 613
rect 40 575 46 609
rect 80 575 118 609
rect 152 575 916 609
rect 40 571 916 575
rect 917 572 918 612
rect 954 572 955 612
rect 956 609 1832 613
rect 956 575 1720 609
rect 1754 575 1792 609
rect 1826 575 1832 609
rect 956 571 1832 575
rect 40 563 158 571
tri 158 563 166 571 nw
tri 1689 563 1697 571 ne
rect 1697 563 1832 571
tri 1697 546 1714 563 ne
tri 1697 495 1714 512 se
rect 1714 495 1832 563
rect 40 487 158 495
tri 158 487 166 495 sw
tri 1689 487 1697 495 se
rect 1697 487 1832 495
tri 1832 487 1857 512 sw
tri 2186 487 2194 495 se
rect 2194 487 2312 495
rect 40 483 1156 487
rect 40 449 46 483
rect 80 449 118 483
rect 152 449 1156 483
rect 40 445 1156 449
rect 1157 446 1158 486
rect 1194 446 1195 486
rect 1196 483 2312 487
rect 1196 449 2200 483
rect 2234 449 2272 483
rect 2306 449 2312 483
rect 1196 445 2312 449
rect 40 361 158 445
tri 158 420 183 445 nw
tri 2186 437 2194 445 ne
rect 2194 437 2312 445
tri 158 361 183 386 sw
tri 2586 361 2594 369 se
rect 2594 361 2918 369
tri 2918 361 2926 369 sw
tri 4266 361 4274 369 se
rect 4274 361 4392 369
rect 40 357 1356 361
rect 1358 360 1394 361
rect 40 323 46 357
rect 80 323 118 357
rect 152 323 1356 357
rect 40 319 1356 323
rect 1357 320 1395 360
rect 1396 357 3576 361
rect 1396 323 2600 357
rect 2634 323 2672 357
rect 2706 323 2806 357
rect 2840 323 2878 357
rect 2912 323 3576 357
rect 1358 319 1394 320
rect 1396 319 3576 323
rect 3577 320 3578 360
rect 3614 320 3615 360
rect 3616 357 4392 361
rect 3616 323 4280 357
rect 4314 323 4352 357
rect 4386 323 4392 357
rect 3616 319 4392 323
rect 40 311 158 319
tri 158 311 166 319 nw
tri 2586 311 2594 319 ne
rect 2594 311 2918 319
tri 2918 311 2926 319 nw
tri 4249 311 4257 319 ne
rect 4257 311 4392 319
tri 4257 294 4274 311 ne
tri 4257 243 4274 260 se
rect 4274 243 4392 311
rect 40 235 158 243
tri 158 235 166 243 sw
tri 4249 235 4257 243 se
rect 4257 235 4392 243
rect 40 231 2196 235
rect 40 197 46 231
rect 80 197 118 231
rect 152 197 2196 231
rect 40 193 2196 197
rect 2197 194 2198 234
rect 2234 194 2235 234
rect 2236 231 4392 235
rect 2236 197 4280 231
rect 4314 197 4352 231
rect 4386 197 4392 231
rect 2236 193 4392 197
rect 40 185 175 193
tri 175 185 183 193 nw
tri 4266 185 4274 193 ne
rect 4274 185 4392 193
rect 40 109 158 185
tri 158 168 175 185 nw
tri 158 109 183 134 sw
tri 4266 109 4274 117 se
rect 4274 109 4392 117
rect 40 105 2196 109
rect 40 71 46 105
rect 80 71 118 105
rect 152 71 2196 105
rect 40 67 2196 71
rect 2197 68 2198 108
rect 2234 68 2235 108
rect 2236 105 4392 109
rect 2236 71 4280 105
rect 4314 71 4352 105
rect 4386 71 4392 105
rect 2236 67 4392 71
rect 40 59 158 67
tri 158 59 166 67 nw
tri 4266 59 4274 67 ne
rect 4274 59 4392 67
rect 44 -21 162 -9
rect 44 -55 50 -21
rect 84 -55 122 -21
rect 156 -55 162 -21
rect 44 -67 162 -55
rect 45 -69 161 -68
rect 44 -105 162 -69
rect 45 -106 161 -105
rect 44 -159 162 -107
rect 4256 -21 4374 -9
rect 4256 -55 4262 -21
rect 4296 -55 4334 -21
rect 4368 -55 4374 -21
rect 4256 -67 4374 -55
rect 4257 -69 4373 -68
rect 4256 -105 4374 -69
rect 4257 -106 4373 -105
rect 4256 -159 4374 -107
<< rmetal1 >>
rect 4274 4532 4392 4533
rect 4274 4531 4275 4532
rect 4391 4531 4392 4532
rect 4274 4494 4275 4495
rect 4391 4494 4392 4495
rect 4274 4493 4392 4494
rect 2196 4467 2198 4468
rect 2196 4427 2197 4467
rect 2196 4426 2198 4427
rect 2234 4467 2236 4468
rect 2235 4427 2236 4467
rect 2234 4426 2236 4427
rect 2196 4341 2198 4342
rect 2196 4301 2197 4341
rect 2196 4300 2198 4301
rect 2234 4341 2236 4342
rect 2235 4301 2236 4341
rect 2234 4300 2236 4301
rect 1356 4215 1358 4216
rect 1394 4215 1396 4216
rect 1356 4175 1357 4215
rect 1395 4175 1396 4215
rect 3576 4215 3578 4216
rect 1356 4174 1358 4175
rect 1394 4174 1396 4175
rect 3576 4175 3577 4215
rect 3576 4174 3578 4175
rect 3614 4215 3616 4216
rect 3615 4175 3616 4215
rect 3614 4174 3616 4175
rect 1156 4089 1158 4090
rect 1156 4049 1157 4089
rect 1156 4048 1158 4049
rect 1194 4089 1196 4090
rect 1195 4049 1196 4089
rect 1194 4048 1196 4049
rect 916 3963 918 3964
rect 916 3923 917 3963
rect 916 3922 918 3923
rect 954 3963 956 3964
rect 955 3923 956 3963
rect 954 3922 956 3923
rect 816 3837 818 3838
rect 816 3797 817 3837
rect 816 3796 818 3797
rect 854 3837 856 3838
rect 855 3797 856 3837
rect 854 3796 856 3797
rect 956 3711 958 3712
rect 994 3711 996 3712
rect 956 3671 957 3711
rect 995 3671 996 3711
rect 956 3670 958 3671
rect 994 3670 996 3671
rect 956 864 958 865
rect 994 864 996 865
rect 956 824 957 864
rect 995 824 996 864
rect 956 823 958 824
rect 994 823 996 824
rect 816 738 818 739
rect 816 698 817 738
rect 816 697 818 698
rect 854 738 856 739
rect 855 698 856 738
rect 854 697 856 698
rect 916 612 918 613
rect 916 572 917 612
rect 916 571 918 572
rect 954 612 956 613
rect 955 572 956 612
rect 954 571 956 572
rect 1156 486 1158 487
rect 1156 446 1157 486
rect 1156 445 1158 446
rect 1194 486 1196 487
rect 1195 446 1196 486
rect 1194 445 1196 446
rect 1356 360 1358 361
rect 1394 360 1396 361
rect 1356 320 1357 360
rect 1395 320 1396 360
rect 3576 360 3578 361
rect 1356 319 1358 320
rect 1394 319 1396 320
rect 3576 320 3577 360
rect 3576 319 3578 320
rect 3614 360 3616 361
rect 3615 320 3616 360
rect 3614 319 3616 320
rect 2196 234 2198 235
rect 2196 194 2197 234
rect 2196 193 2198 194
rect 2234 234 2236 235
rect 2235 194 2236 234
rect 2234 193 2236 194
rect 2196 108 2198 109
rect 2196 68 2197 108
rect 2196 67 2198 68
rect 2234 108 2236 109
rect 2235 68 2236 108
rect 2234 67 2236 68
rect 44 -68 162 -67
rect 44 -69 45 -68
rect 161 -69 162 -68
rect 44 -106 45 -105
rect 161 -106 162 -105
rect 44 -107 162 -106
rect 4256 -68 4374 -67
rect 4256 -69 4257 -68
rect 4373 -69 4374 -68
rect 4256 -106 4257 -105
rect 4373 -106 4374 -105
rect 4256 -107 4374 -106
<< via1 >>
rect 46 3708 98 3751
rect 46 3699 80 3708
rect 80 3699 98 3708
rect 46 3674 80 3687
rect 80 3674 98 3687
rect 46 3635 98 3674
rect 46 861 98 900
rect 46 848 80 861
rect 80 848 98 861
rect 46 827 80 836
rect 80 827 98 836
rect 46 784 98 827
<< metal2 >>
rect 40 3699 46 3751
rect 98 3699 104 3751
rect 40 3687 104 3699
rect 40 3635 46 3687
rect 98 3635 104 3687
rect 40 900 104 3635
rect 40 848 46 900
rect 98 848 104 900
rect 40 836 104 848
rect 40 784 46 836
rect 98 784 104 836
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_0
timestamp 1704896540
transform -1 0 4406 0 1 4166
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_1
timestamp 1704896540
transform -1 0 4406 0 1 4292
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_2
timestamp 1704896540
transform -1 0 4406 0 1 4418
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_3
timestamp 1704896540
transform -1 0 4406 0 1 4544
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_4
timestamp 1704896540
transform -1 0 2726 0 1 4166
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_5
timestamp 1704896540
transform -1 0 2326 0 1 4040
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_6
timestamp 1704896540
transform -1 0 1846 0 1 3914
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_7
timestamp 1704896540
transform -1 0 1926 0 1 3662
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_8
timestamp 1704896540
transform -1 0 1646 0 1 3788
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_9
timestamp 1704896540
transform -1 0 2726 0 1 311
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_10
timestamp 1704896540
transform -1 0 1926 0 1 815
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_11
timestamp 1704896540
transform -1 0 1646 0 1 689
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_12
timestamp 1704896540
transform -1 0 1846 0 1 563
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_13
timestamp 1704896540
transform -1 0 2326 0 1 437
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_14
timestamp 1704896540
transform -1 0 4406 0 1 311
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_15
timestamp 1704896540
transform -1 0 4406 0 1 185
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_16
timestamp 1704896540
transform -1 0 4406 0 1 59
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_17
timestamp 1704896540
transform -1 0 4406 0 1 -67
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_18
timestamp 1704896540
transform 1 0 26 0 1 4544
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_19
timestamp 1704896540
transform 1 0 2786 0 1 4166
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_20
timestamp 1704896540
transform 1 0 26 0 1 3662
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_21
timestamp 1704896540
transform 1 0 26 0 1 3788
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_22
timestamp 1704896540
transform 1 0 26 0 1 3914
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_23
timestamp 1704896540
transform 1 0 26 0 1 4040
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_24
timestamp 1704896540
transform 1 0 26 0 1 4166
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_25
timestamp 1704896540
transform 1 0 26 0 1 4292
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_26
timestamp 1704896540
transform 1 0 26 0 1 4418
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_27
timestamp 1704896540
transform 1 0 2786 0 1 311
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_28
timestamp 1704896540
transform 1 0 26 0 1 -67
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_29
timestamp 1704896540
transform 1 0 26 0 1 59
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_30
timestamp 1704896540
transform 1 0 26 0 1 185
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_31
timestamp 1704896540
transform 1 0 26 0 1 311
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_32
timestamp 1704896540
transform 1 0 26 0 1 437
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_33
timestamp 1704896540
transform 1 0 26 0 1 563
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_34
timestamp 1704896540
transform 1 0 26 0 1 689
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_35
timestamp 1704896540
transform 1 0 26 0 1 815
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_0
timestamp 1704896540
transform 0 1 2806 1 0 4178
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_1
timestamp 1704896540
transform 0 1 46 1 0 3674
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_2
timestamp 1704896540
transform 0 1 46 1 0 3800
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_3
timestamp 1704896540
transform 0 1 46 1 0 3926
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_4
timestamp 1704896540
transform 0 1 46 1 0 4052
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_5
timestamp 1704896540
transform 0 1 46 1 0 4178
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_6
timestamp 1704896540
transform 0 1 46 1 0 4304
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_7
timestamp 1704896540
transform 0 1 46 1 0 4430
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_8
timestamp 1704896540
transform 0 1 50 1 0 4556
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_9
timestamp 1704896540
transform 0 1 2806 1 0 323
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_10
timestamp 1704896540
transform 0 1 50 1 0 -55
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_11
timestamp 1704896540
transform 0 1 46 1 0 71
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_12
timestamp 1704896540
transform 0 1 46 1 0 197
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_13
timestamp 1704896540
transform 0 1 46 1 0 323
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_14
timestamp 1704896540
transform 0 1 46 1 0 449
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_15
timestamp 1704896540
transform 0 1 46 1 0 575
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_16
timestamp 1704896540
transform 0 1 46 1 0 701
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_17
timestamp 1704896540
transform 0 1 46 1 0 827
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_18
timestamp 1704896540
transform 0 -1 4386 1 0 4178
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_19
timestamp 1704896540
transform 0 -1 4386 1 0 4304
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_20
timestamp 1704896540
transform 0 -1 4386 1 0 4430
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_21
timestamp 1704896540
transform 0 -1 4386 1 0 4559
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_22
timestamp 1704896540
transform 0 -1 2706 1 0 4178
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_23
timestamp 1704896540
transform 0 -1 2306 1 0 4052
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_24
timestamp 1704896540
transform 0 -1 1826 1 0 3926
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_25
timestamp 1704896540
transform 0 -1 1626 1 0 3800
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_26
timestamp 1704896540
transform 0 -1 1906 1 0 3674
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_27
timestamp 1704896540
transform 0 -1 2706 1 0 323
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_28
timestamp 1704896540
transform 0 -1 1906 1 0 827
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_29
timestamp 1704896540
transform 0 -1 1626 1 0 701
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_30
timestamp 1704896540
transform 0 -1 1826 1 0 575
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_31
timestamp 1704896540
transform 0 -1 2306 1 0 449
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_32
timestamp 1704896540
transform 0 -1 4386 1 0 323
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_33
timestamp 1704896540
transform 0 -1 4386 1 0 197
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_34
timestamp 1704896540
transform 0 -1 4386 1 0 71
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_35
timestamp 1704896540
transform 0 -1 4368 1 0 -55
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_0
timestamp 1704896540
transform 1 0 40 0 -1 900
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_1
timestamp 1704896540
transform 1 0 40 0 1 3635
box 0 0 1 1
use nDFres_CDNS_524688791851282  nDFres_CDNS_524688791851282_0
timestamp 1704896540
transform -1 0 1816 0 -1 3724
box -68 -26 1748 92
use nDFres_CDNS_524688791851282  nDFres_CDNS_524688791851282_1
timestamp 1704896540
transform 1 0 136 0 -1 877
box -68 -26 1748 92
use nDFres_CDNS_524688791851283  nDFres_CDNS_524688791851283_0
timestamp 1704896540
transform -1 0 2216 0 -1 499
box -68 -26 2148 92
use nDFres_CDNS_524688791851283  nDFres_CDNS_524688791851283_1
timestamp 1704896540
transform 1 0 136 0 -1 4102
box -68 -26 2148 92
use nDFres_CDNS_524688791851284  nDFres_CDNS_524688791851284_0
timestamp 1704896540
transform -1 0 2616 0 -1 4228
box -68 -26 2548 92
use nDFres_CDNS_524688791851284  nDFres_CDNS_524688791851284_1
timestamp 1704896540
transform 1 0 136 0 -1 373
box -68 -26 2548 92
use nDFres_CDNS_524688791851285  nDFres_CDNS_524688791851285_0
timestamp 1704896540
transform -1 0 4296 0 -1 4480
box -68 -26 4228 92
use nDFres_CDNS_524688791851285  nDFres_CDNS_524688791851285_1
timestamp 1704896540
transform -1 0 4296 0 -1 247
box -68 -26 4228 92
use nDFres_CDNS_524688791851285  nDFres_CDNS_524688791851285_2
timestamp 1704896540
transform 1 0 136 0 -1 4354
box -68 -26 4228 92
use nDFres_CDNS_524688791851285  nDFres_CDNS_524688791851285_3
timestamp 1704896540
transform 1 0 136 0 -1 4606
box -68 -26 4228 92
use nDFres_CDNS_524688791851285  nDFres_CDNS_524688791851285_4
timestamp 1704896540
transform 1 0 136 0 -1 -5
box -68 -26 4228 92
use nDFres_CDNS_524688791851285  nDFres_CDNS_524688791851285_5
timestamp 1704896540
transform 1 0 136 0 -1 121
box -68 -26 4228 92
use nDFres_CDNS_524688791851286  nDFres_CDNS_524688791851286_0
timestamp 1704896540
transform -1 0 4296 0 -1 4228
box -68 -26 1468 92
use nDFres_CDNS_524688791851286  nDFres_CDNS_524688791851286_1
timestamp 1704896540
transform -1 0 1536 0 -1 751
box -68 -26 1468 92
use nDFres_CDNS_524688791851286  nDFres_CDNS_524688791851286_2
timestamp 1704896540
transform 1 0 136 0 -1 3850
box -68 -26 1468 92
use nDFres_CDNS_524688791851286  nDFres_CDNS_524688791851286_3
timestamp 1704896540
transform 1 0 2896 0 -1 373
box -68 -26 1468 92
use nDFres_CDNS_524688791851287  nDFres_CDNS_524688791851287_0
timestamp 1704896540
transform -1 0 1736 0 -1 3976
box -68 -26 1668 92
use nDFres_CDNS_524688791851287  nDFres_CDNS_524688791851287_1
timestamp 1704896540
transform 1 0 136 0 -1 625
box -68 -26 1668 92
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851279  sky130_fd_io__sio_tk_em1o_CDNS_524688791851279_0
timestamp 1704896540
transform -1 0 1008 0 1 3922
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851279  sky130_fd_io__sio_tk_em1o_CDNS_524688791851279_1
timestamp 1704896540
transform -1 0 3668 0 1 4174
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851279  sky130_fd_io__sio_tk_em1o_CDNS_524688791851279_2
timestamp 1704896540
transform -1 0 2288 0 1 4426
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851279  sky130_fd_io__sio_tk_em1o_CDNS_524688791851279_3
timestamp 1704896540
transform -1 0 2288 0 1 193
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851279  sky130_fd_io__sio_tk_em1o_CDNS_524688791851279_4
timestamp 1704896540
transform -1 0 1248 0 1 445
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851279  sky130_fd_io__sio_tk_em1o_CDNS_524688791851279_5
timestamp 1704896540
transform -1 0 908 0 1 697
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851279  sky130_fd_io__sio_tk_em1o_CDNS_524688791851279_6
timestamp 1704896540
transform 1 0 764 0 1 3796
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851279  sky130_fd_io__sio_tk_em1o_CDNS_524688791851279_7
timestamp 1704896540
transform 1 0 1104 0 1 4048
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851279  sky130_fd_io__sio_tk_em1o_CDNS_524688791851279_8
timestamp 1704896540
transform 1 0 2144 0 1 4300
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851279  sky130_fd_io__sio_tk_em1o_CDNS_524688791851279_9
timestamp 1704896540
transform 1 0 2144 0 1 67
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851279  sky130_fd_io__sio_tk_em1o_CDNS_524688791851279_10
timestamp 1704896540
transform 1 0 3524 0 1 319
box 0 0 1 1
use sky130_fd_io__sio_tk_em1o_CDNS_524688791851279  sky130_fd_io__sio_tk_em1o_CDNS_524688791851279_11
timestamp 1704896540
transform 1 0 864 0 1 571
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_52468879185538  sky130_fd_io__sio_tk_em1s_CDNS_52468879185538_0
timestamp 1704896540
transform 0 1 4256 -1 0 -15
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_52468879185538  sky130_fd_io__sio_tk_em1s_CDNS_52468879185538_1
timestamp 1704896540
transform 0 1 44 -1 0 -15
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_52468879185538  sky130_fd_io__sio_tk_em1s_CDNS_52468879185538_2
timestamp 1704896540
transform 0 1 4274 1 0 4441
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851278  sky130_fd_io__sio_tk_em1s_CDNS_524688791851278_0
timestamp 1704896540
transform -1 0 1048 0 1 3670
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851278  sky130_fd_io__sio_tk_em1s_CDNS_524688791851278_1
timestamp 1704896540
transform -1 0 1448 0 1 4174
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851278  sky130_fd_io__sio_tk_em1s_CDNS_524688791851278_2
timestamp 1704896540
transform 1 0 1304 0 1 319
box 0 0 1 1
use sky130_fd_io__sio_tk_em1s_CDNS_524688791851278  sky130_fd_io__sio_tk_em1s_CDNS_524688791851278_3
timestamp 1704896540
transform 1 0 904 0 1 823
box 0 0 1 1
<< labels >>
flabel metal1 s 4256 -159 4374 -107 0 FreeSans 200 90 0 0 vgnd
port 3 nsew
flabel metal1 s 4352 59 4392 117 0 FreeSans 200 0 0 0 r1
port 1 nsew
flabel metal1 s 4352 4418 4392 4476 0 FreeSans 200 0 0 0 r0
port 2 nsew
flabel metal1 s 44 -159 162 -107 0 FreeSans 200 90 0 0 vgnd
port 3 nsew
flabel mvpsubdiff s 103 4698 103 4698 0 FreeSans 200 90 0 0 vgnd
<< properties >>
string GDS_END 86234506
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86217640
<< end >>
