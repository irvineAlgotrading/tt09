magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -376 920 880 1366
rect -376 138 880 424
<< pwell >>
rect 103 1409 381 1939
rect 103 846 385 872
rect 103 702 491 846
rect 103 628 417 702
rect 35 504 417 628
rect 35 466 313 504
<< scnmos >>
rect 183 1713 213 1913
rect 271 1713 301 1913
rect 183 1435 213 1507
rect 271 1435 301 1507
rect 183 736 213 846
rect 271 736 301 846
rect 115 492 145 602
rect 203 492 233 602
rect 303 530 333 602
<< scpmos >>
rect 183 1219 213 1329
rect 271 1219 301 1329
rect 183 956 213 1066
rect 271 956 301 1066
rect 115 262 145 372
rect 203 262 233 372
rect 291 262 321 372
<< ndiff >>
rect 129 1898 183 1913
rect 129 1864 137 1898
rect 171 1864 183 1898
rect 129 1830 183 1864
rect 129 1796 137 1830
rect 171 1796 183 1830
rect 129 1762 183 1796
rect 129 1728 137 1762
rect 171 1728 183 1762
rect 129 1713 183 1728
rect 213 1898 271 1913
rect 213 1864 225 1898
rect 259 1864 271 1898
rect 213 1830 271 1864
rect 213 1796 225 1830
rect 259 1796 271 1830
rect 213 1762 271 1796
rect 213 1728 225 1762
rect 259 1728 271 1762
rect 213 1713 271 1728
rect 301 1898 355 1913
rect 301 1864 313 1898
rect 347 1864 355 1898
rect 301 1830 355 1864
rect 301 1796 313 1830
rect 347 1796 355 1830
rect 301 1762 355 1796
rect 301 1728 313 1762
rect 347 1728 355 1762
rect 301 1713 355 1728
rect 129 1489 183 1507
rect 129 1455 137 1489
rect 171 1455 183 1489
rect 129 1435 183 1455
rect 213 1489 271 1507
rect 213 1455 225 1489
rect 259 1455 271 1489
rect 213 1435 271 1455
rect 301 1489 355 1507
rect 301 1455 313 1489
rect 347 1455 355 1489
rect 301 1435 355 1455
rect 129 808 183 846
rect 129 774 137 808
rect 171 774 183 808
rect 129 736 183 774
rect 213 736 271 846
rect 301 808 359 846
rect 301 774 313 808
rect 347 774 359 808
rect 301 736 359 774
rect 61 564 115 602
rect 61 530 69 564
rect 103 530 115 564
rect 61 492 115 530
rect 145 564 203 602
rect 145 530 157 564
rect 191 530 203 564
rect 145 492 203 530
rect 233 564 303 602
rect 233 530 245 564
rect 279 530 303 564
rect 333 583 391 602
rect 333 549 345 583
rect 379 549 391 583
rect 333 530 391 549
rect 233 492 287 530
<< pdiff >>
rect 129 1291 183 1329
rect 129 1257 137 1291
rect 171 1257 183 1291
rect 129 1219 183 1257
rect 213 1291 271 1329
rect 213 1257 225 1291
rect 259 1257 271 1291
rect 213 1219 271 1257
rect 301 1291 355 1329
rect 301 1257 313 1291
rect 347 1257 355 1291
rect 301 1219 355 1257
rect 129 1028 183 1066
rect 129 994 137 1028
rect 171 994 183 1028
rect 129 956 183 994
rect 213 1028 271 1066
rect 213 994 225 1028
rect 259 994 271 1028
rect 213 956 271 994
rect 301 1028 356 1066
rect 301 994 313 1028
rect 347 994 356 1028
rect 301 956 356 994
rect 61 334 115 372
rect 61 300 69 334
rect 103 300 115 334
rect 61 262 115 300
rect 145 334 203 372
rect 145 300 157 334
rect 191 300 203 334
rect 145 262 203 300
rect 233 334 291 372
rect 233 300 245 334
rect 279 300 291 334
rect 233 262 291 300
rect 321 334 376 372
rect 321 300 333 334
rect 367 300 376 334
rect 321 262 376 300
<< ndiffc >>
rect 137 1864 171 1898
rect 137 1796 171 1830
rect 137 1728 171 1762
rect 225 1864 259 1898
rect 225 1796 259 1830
rect 225 1728 259 1762
rect 313 1864 347 1898
rect 313 1796 347 1830
rect 313 1728 347 1762
rect 137 1455 171 1489
rect 225 1455 259 1489
rect 313 1455 347 1489
rect 137 774 171 808
rect 313 774 347 808
rect 69 530 103 564
rect 157 530 191 564
rect 245 530 279 564
rect 345 549 379 583
<< pdiffc >>
rect 137 1257 171 1291
rect 225 1257 259 1291
rect 313 1257 347 1291
rect 137 994 171 1028
rect 225 994 259 1028
rect 313 994 347 1028
rect 69 300 103 334
rect 157 300 191 334
rect 245 300 279 334
rect 333 300 367 334
<< psubdiff >>
rect 229 1561 259 1595
rect 293 1561 321 1595
rect 431 790 465 820
rect 431 728 465 756
<< nsubdiff >>
rect 225 1124 259 1158
rect 293 1124 321 1158
rect 249 174 279 208
rect 313 174 341 208
<< psubdiffcont >>
rect 259 1561 293 1595
rect 431 756 465 790
<< nsubdiffcont >>
rect 259 1124 293 1158
rect 279 174 313 208
<< poly >>
rect 183 1983 409 2011
rect 183 1981 445 1983
rect 183 1913 213 1981
rect 379 1973 445 1981
rect 379 1939 395 1973
rect 429 1939 445 1973
rect 271 1913 301 1939
rect 379 1929 445 1939
rect 183 1687 213 1713
rect 271 1641 301 1713
rect 121 1631 301 1641
rect 121 1597 137 1631
rect 171 1611 301 1631
rect 171 1597 187 1611
rect 121 1585 187 1597
rect 183 1507 213 1533
rect 271 1507 301 1533
rect 183 1329 213 1435
rect 271 1329 301 1435
rect 183 1204 213 1219
rect 78 1174 213 1204
rect 271 1204 301 1219
rect 271 1174 406 1204
rect 41 1164 108 1174
rect 41 1130 57 1164
rect 91 1130 108 1164
rect 376 1164 443 1174
rect 41 1120 108 1130
rect 376 1144 393 1164
rect 377 1130 393 1144
rect 427 1130 443 1164
rect 377 1120 443 1130
rect 183 1066 213 1092
rect 271 1066 301 1092
rect 183 846 213 956
rect 271 846 301 956
rect 183 720 213 736
rect 115 690 213 720
rect 271 720 301 736
rect 271 690 399 720
rect 115 602 145 690
rect 365 680 449 690
rect 365 660 399 680
rect 375 646 399 660
rect 433 646 449 680
rect 375 636 449 646
rect 203 602 233 628
rect 303 602 333 628
rect 115 372 145 492
rect 203 476 233 492
rect 303 476 333 530
rect 203 446 333 476
rect 203 372 233 446
rect 291 372 321 446
rect 115 150 145 262
rect 101 148 145 150
rect 101 134 155 148
rect 101 100 111 134
rect 145 100 155 134
rect 203 130 233 262
rect 291 236 321 262
rect 203 100 287 130
rect 101 84 155 100
rect 255 64 287 100
rect 255 54 317 64
rect 255 20 267 54
rect 301 20 317 54
rect 255 4 317 20
<< polycont >>
rect 395 1939 429 1973
rect 137 1597 171 1631
rect 57 1130 91 1164
rect 393 1130 427 1164
rect 399 646 433 680
rect 111 100 145 134
rect 267 20 301 54
<< locali >>
rect 381 1973 429 1989
rect 137 1898 171 1913
rect 137 1830 171 1864
rect 137 1762 171 1796
rect 137 1709 171 1728
rect 225 1898 259 1927
rect 225 1830 259 1864
rect 225 1762 259 1796
rect 117 1631 171 1647
rect 117 1597 137 1631
rect 117 1580 171 1597
rect 137 1489 171 1580
rect 137 1291 171 1455
rect 225 1595 259 1728
rect 313 1898 347 1913
rect 313 1830 347 1864
rect 313 1762 347 1796
rect 313 1709 347 1728
rect 381 1939 395 1973
rect 381 1923 429 1939
rect 293 1561 309 1595
rect 225 1489 259 1561
rect 225 1433 259 1455
rect 313 1489 347 1513
rect 313 1399 347 1455
rect 381 1399 415 1923
rect 313 1365 415 1399
rect 137 1216 171 1257
rect 225 1291 259 1333
rect 57 1164 103 1180
rect 91 1130 103 1164
rect 57 1114 103 1130
rect 69 564 103 1114
rect 225 1158 259 1257
rect 313 1291 347 1365
rect 313 1216 347 1257
rect 381 1164 427 1180
rect 293 1124 309 1158
rect 381 1130 393 1164
rect 137 1028 171 1070
rect 137 918 171 994
rect 225 1028 259 1124
rect 381 1114 427 1130
rect 225 952 259 994
rect 313 1028 347 1070
rect 313 918 347 994
rect 381 918 415 1114
rect 137 884 415 918
rect 137 808 171 884
rect 137 730 171 774
rect 313 824 347 850
rect 313 808 360 824
rect 347 790 360 808
rect 394 790 471 824
rect 313 732 347 774
rect 431 740 465 756
rect 387 680 433 698
rect 387 646 399 680
rect 387 632 433 646
rect 69 444 103 530
rect 157 564 191 606
rect 157 488 191 530
rect 245 564 279 590
rect 245 488 279 530
rect 345 622 433 632
rect 345 598 421 622
rect 345 583 391 598
rect 379 578 391 583
rect 69 410 191 444
rect 345 424 379 549
rect 69 334 103 376
rect 69 208 103 300
rect 157 334 191 410
rect 333 390 379 424
rect 157 258 191 300
rect 245 334 279 376
rect 245 208 279 300
rect 333 334 367 390
rect 333 258 367 300
rect 69 174 245 208
rect 313 174 329 208
rect 245 168 279 174
rect 94 100 111 134
rect 145 100 161 134
rect 251 20 267 54
rect 301 20 317 54
<< viali >>
rect 137 1913 171 1947
rect 313 1913 347 1947
rect 225 1561 259 1595
rect 225 1124 259 1158
rect 360 790 394 824
rect 245 590 279 624
rect 245 174 279 208
rect 111 100 145 134
rect 267 20 301 54
<< metal1 >>
rect 126 1959 156 2011
rect 328 1959 358 2011
rect 125 1947 182 1959
rect 125 1913 137 1947
rect 171 1913 182 1947
rect 125 1901 182 1913
rect 302 1947 359 1959
rect 302 1913 313 1947
rect 347 1913 359 1947
rect 302 1901 359 1913
rect 213 1595 299 1601
rect 213 1561 225 1595
rect 259 1561 321 1595
rect 213 1555 299 1561
rect 213 1158 299 1164
rect 213 1124 225 1158
rect 259 1124 299 1158
rect 213 1118 299 1124
rect 334 824 420 830
rect 334 790 360 824
rect 394 790 420 824
rect 334 789 420 790
rect 347 784 420 789
rect 219 624 305 630
rect 219 590 245 624
rect 279 590 305 624
rect 219 584 305 590
rect 233 208 319 214
rect 233 174 245 208
rect 279 174 319 208
rect 233 168 319 174
rect 99 134 157 156
rect 99 100 111 134
rect 145 128 157 134
rect 145 100 500 128
rect 99 94 500 100
rect 255 54 315 60
rect 255 20 267 54
rect 301 20 315 54
rect 255 4 315 20
<< labels >>
rlabel metal1 s 126 1959 156 2011 4 BL
port 2 nsew
rlabel metal1 s 328 1959 358 2011 4 BR
port 3 nsew
rlabel metal1 s 255 4 315 60 4 DIN
port 1 nsew
rlabel metal1 s 99 94 500 128 4 EN
port 4 nsew
rlabel metal1 s 219 584 305 630 4 GND
port 6 nsew
rlabel metal1 s 334 789 420 830 4 GND
port 6 nsew
rlabel metal1 s 213 1561 321 1595 4 GND
port 6 nsew
rlabel metal1 s 233 168 319 214 4 VDD
port 5 nsew
rlabel metal1 s 213 1118 299 1164 4 VDD
port 5 nsew
rlabel metal1 s 285 32 285 32 4 din
rlabel metal1 s 141 1985 141 1985 4 bl
rlabel metal1 s 343 1985 343 1985 4 br
rlabel metal1 s 299 111 299 111 4 en
rlabel metal1 s 276 191 276 191 4 vdd
rlabel metal1 s 256 1141 256 1141 4 vdd
rlabel metal1 s 262 607 262 607 4 gnd
rlabel metal1 s 377 809 377 809 4 gnd
rlabel metal1 s 267 1578 267 1578 4 gnd
<< properties >>
string FIXED_BBOX 0 0 500 2011
string GDS_END 247866
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_2kbyte_1rw1r_32x512_8.gds
string GDS_START 234822
<< end >>
