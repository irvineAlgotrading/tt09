magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< pwell >>
rect -68 -266 2912 92
<< ndiff >>
rect -42 50 0 66
rect -42 16 -34 50
rect -42 0 0 16
rect 2843 -190 2886 -174
rect 2877 -224 2886 -190
rect 2843 -240 2886 -224
<< ndiffc >>
rect -34 16 0 50
rect 2843 -224 2877 -190
<< ndiffres >>
rect 0 0 2886 66
rect 2820 -54 2886 0
rect -42 -120 2886 -54
rect -42 -174 24 -120
rect -42 -240 2843 -174
<< locali >>
rect -34 50 0 66
rect -34 0 0 16
rect 2843 -190 2878 -174
rect 2877 -224 2878 -190
rect 2843 -240 2878 -224
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_0
timestamp 1704896540
transform 1 0 2835 0 1 -236
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_1
timestamp 1704896540
transform 1 0 -42 0 1 4
box 0 0 1 1
<< properties >>
string GDS_END 86618810
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86617686
<< end >>
