magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< obsli1 >>
rect -1208 6870 1508 7182
rect -1208 -894 -896 6870
rect 0 0 300 6000
rect -189 -651 489 -649
rect -190 -894 489 -651
rect 1196 -894 1508 6870
rect -1208 -1182 1508 -894
<< obsm1 >>
rect -1208 6700 1508 7182
rect -1208 6450 -607 6700
tri -607 6450 -357 6700 nw
tri 658 6450 908 6700 ne
rect 908 6450 1508 6700
rect -1208 -450 -709 6450
tri -709 6348 -607 6450 nw
tri -449 6374 -373 6450 se
rect -373 6374 674 6450
tri 674 6374 750 6450 sw
tri -709 -450 -607 -348 sw
rect -449 -374 750 6374
tri 908 6348 1010 6450 ne
tri -449 -386 -437 -374 ne
rect -437 -386 738 -374
tri 738 -386 750 -374 nw
tri -437 -450 -373 -386 ne
rect -373 -450 674 -386
tri 674 -450 738 -386 nw
tri 908 -450 1010 -348 se
rect 1010 -450 1508 6450
rect -1208 -700 -607 -450
tri -607 -700 -357 -450 sw
tri 658 -700 908 -450 se
rect 908 -700 1508 -450
rect -1208 -1182 1508 -700
<< obsm2 >>
rect -1208 6700 1508 7182
rect -1208 6450 -607 6700
tri -607 6450 -357 6700 nw
tri 658 6450 908 6700 ne
rect 908 6450 1508 6700
rect -1208 -450 -709 6450
tri -709 6348 -607 6450 nw
tri -449 6374 -373 6450 se
rect -373 6374 674 6450
tri 674 6374 750 6450 sw
tri -709 -450 -607 -348 sw
rect -449 -374 750 6374
tri 908 6348 1010 6450 ne
tri -449 -388 -435 -374 ne
rect -435 -388 736 -374
tri 736 -388 750 -374 nw
tri -435 -450 -373 -388 ne
rect -373 -450 674 -388
tri 674 -450 736 -388 nw
tri 908 -450 1010 -348 se
rect 1010 -450 1508 6450
rect -1208 -700 -607 -450
tri -607 -700 -357 -450 sw
tri 658 -700 908 -450 se
rect 908 -700 1508 -450
rect -1208 -1182 1508 -700
<< obsm3 >>
rect -1208 5182 1508 7182
rect -968 818 1268 5182
rect -1208 -1182 1508 818
<< properties >>
string FIXED_BBOX -1208 -1182 1508 7182
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 4406438
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 3906210
<< end >>
