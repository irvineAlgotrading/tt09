magic
tech sky130B
timestamp 1704896540
<< metal1 >>
rect 0 0 3 1146
rect 93 0 96 1146
<< via1 >>
rect 3 0 93 1146
<< metal2 >>
rect 0 0 3 1146
rect 93 0 96 1146
<< properties >>
string GDS_END 88816032
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 88808988
<< end >>
