magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect 0 3844 1126 4012
rect 0 168 168 3844
rect 958 168 1126 3844
rect 0 0 1126 168
<< pwell >>
rect 228 3698 898 3784
rect 228 314 314 3698
rect 812 314 898 3698
rect 228 228 898 314
<< mvpsubdiff >>
rect 254 3724 278 3758
rect 312 3724 351 3758
rect 385 3724 423 3758
rect 457 3724 495 3758
rect 529 3724 567 3758
rect 601 3724 701 3758
rect 735 3734 872 3758
rect 735 3724 838 3734
rect 254 3666 288 3724
rect 254 3598 288 3632
rect 254 3530 288 3564
rect 254 3462 288 3496
rect 254 3394 288 3428
rect 254 3326 288 3360
rect 254 3258 288 3292
rect 254 3190 288 3224
rect 254 3122 288 3156
rect 254 3054 288 3088
rect 254 2986 288 3020
rect 254 2918 288 2952
rect 254 2850 288 2884
rect 254 2782 288 2816
rect 254 2714 288 2748
rect 254 2646 288 2680
rect 838 3665 872 3700
rect 838 3596 872 3631
rect 838 3527 872 3562
rect 838 3458 872 3493
rect 838 3389 872 3424
rect 838 3320 872 3355
rect 838 3251 872 3286
rect 838 3182 872 3217
rect 838 3113 872 3148
rect 838 3044 872 3079
rect 838 2975 872 3010
rect 838 2906 872 2941
rect 838 2837 872 2872
rect 838 2768 872 2803
rect 838 2699 872 2734
rect 838 2630 872 2665
rect 254 2578 288 2612
rect 838 2561 872 2596
rect 254 2510 288 2544
rect 254 2442 288 2476
rect 254 2374 288 2408
rect 254 2306 288 2340
rect 254 2238 288 2272
rect 254 2170 288 2204
rect 254 2102 288 2136
rect 254 2034 288 2068
rect 254 1966 288 2000
rect 254 1898 288 1932
rect 254 1830 288 1864
rect 254 1761 288 1796
rect 254 1692 288 1727
rect 254 1623 288 1658
rect 254 1554 288 1589
rect 254 1485 288 1520
rect 838 2492 872 2527
rect 838 2423 872 2458
rect 838 2354 872 2389
rect 838 2285 872 2320
rect 838 2216 872 2251
rect 838 2148 872 2182
rect 838 2080 872 2114
rect 838 2012 872 2046
rect 838 1944 872 1978
rect 838 1876 872 1910
rect 838 1808 872 1842
rect 838 1740 872 1774
rect 838 1672 872 1706
rect 838 1604 872 1638
rect 838 1536 872 1570
rect 254 1416 288 1451
rect 838 1468 872 1502
rect 254 1347 288 1382
rect 254 1278 288 1313
rect 254 1209 288 1244
rect 254 1140 288 1175
rect 254 1071 288 1106
rect 254 1002 288 1037
rect 254 933 288 968
rect 254 864 288 899
rect 254 795 288 830
rect 254 726 288 761
rect 254 657 288 692
rect 254 588 288 623
rect 254 519 288 554
rect 254 450 288 485
rect 254 381 288 416
rect 838 1400 872 1434
rect 838 1332 872 1366
rect 838 1264 872 1298
rect 838 1196 872 1230
rect 838 1128 872 1162
rect 838 1060 872 1094
rect 838 992 872 1026
rect 838 924 872 958
rect 838 856 872 890
rect 838 788 872 822
rect 838 720 872 754
rect 838 652 872 686
rect 838 584 872 618
rect 838 516 872 550
rect 838 448 872 482
rect 254 312 288 347
rect 838 380 872 414
rect 838 288 872 346
rect 288 278 360 288
rect 254 254 360 278
rect 394 254 435 288
rect 469 254 510 288
rect 544 254 586 288
rect 620 254 662 288
rect 696 254 738 288
rect 772 254 814 288
rect 848 254 872 288
<< mvnsubdiff >>
rect 68 3911 185 3945
rect 219 3911 256 3945
rect 290 3911 327 3945
rect 361 3911 398 3945
rect 432 3911 469 3945
rect 503 3911 539 3945
rect 573 3911 609 3945
rect 643 3911 679 3945
rect 713 3911 749 3945
rect 783 3911 819 3945
rect 853 3911 889 3945
rect 923 3911 1058 3945
rect 68 3795 102 3911
rect 68 3727 102 3761
rect 68 3659 102 3693
rect 68 3591 102 3625
rect 68 3523 102 3557
rect 68 3455 102 3489
rect 68 3387 102 3421
rect 68 3319 102 3353
rect 68 3251 102 3285
rect 68 3183 102 3217
rect 68 3115 102 3149
rect 68 3047 102 3081
rect 68 2979 102 3013
rect 68 2911 102 2945
rect 68 2843 102 2877
rect 68 2775 102 2809
rect 68 2707 102 2741
rect 68 2639 102 2673
rect 68 2571 102 2605
rect 68 2503 102 2537
rect 68 2435 102 2469
rect 68 2367 102 2401
rect 68 2299 102 2333
rect 68 2231 102 2265
rect 68 2163 102 2197
rect 68 2094 102 2129
rect 68 2025 102 2060
rect 68 1956 102 1991
rect 68 1887 102 1922
rect 68 1818 102 1853
rect 68 1749 102 1784
rect 68 1680 102 1715
rect 68 1611 102 1646
rect 68 1542 102 1577
rect 68 1473 102 1508
rect 68 1404 102 1439
rect 68 1335 102 1370
rect 68 1266 102 1301
rect 68 1197 102 1232
rect 68 1128 102 1163
rect 68 1059 102 1094
rect 68 990 102 1025
rect 68 921 102 956
rect 68 852 102 887
rect 68 783 102 818
rect 68 714 102 749
rect 68 645 102 680
rect 68 576 102 611
rect 68 507 102 542
rect 68 438 102 473
rect 68 369 102 404
rect 68 300 102 335
rect 68 231 102 266
rect 68 101 102 197
rect 1024 101 1058 3911
rect 68 67 203 101
rect 237 67 277 101
rect 311 67 351 101
rect 385 67 425 101
rect 459 67 499 101
rect 533 67 573 101
rect 607 67 647 101
rect 681 67 721 101
rect 755 67 796 101
rect 830 67 871 101
rect 905 67 946 101
rect 980 67 1058 101
<< mvpsubdiffcont >>
rect 278 3724 312 3758
rect 351 3724 385 3758
rect 423 3724 457 3758
rect 495 3724 529 3758
rect 567 3724 601 3758
rect 701 3724 735 3758
rect 254 3632 288 3666
rect 254 3564 288 3598
rect 254 3496 288 3530
rect 254 3428 288 3462
rect 254 3360 288 3394
rect 254 3292 288 3326
rect 254 3224 288 3258
rect 254 3156 288 3190
rect 254 3088 288 3122
rect 254 3020 288 3054
rect 254 2952 288 2986
rect 254 2884 288 2918
rect 254 2816 288 2850
rect 254 2748 288 2782
rect 254 2680 288 2714
rect 254 2612 288 2646
rect 838 3700 872 3734
rect 838 3631 872 3665
rect 838 3562 872 3596
rect 838 3493 872 3527
rect 838 3424 872 3458
rect 838 3355 872 3389
rect 838 3286 872 3320
rect 838 3217 872 3251
rect 838 3148 872 3182
rect 838 3079 872 3113
rect 838 3010 872 3044
rect 838 2941 872 2975
rect 838 2872 872 2906
rect 838 2803 872 2837
rect 838 2734 872 2768
rect 838 2665 872 2699
rect 254 2544 288 2578
rect 838 2596 872 2630
rect 254 2476 288 2510
rect 254 2408 288 2442
rect 254 2340 288 2374
rect 254 2272 288 2306
rect 254 2204 288 2238
rect 254 2136 288 2170
rect 254 2068 288 2102
rect 254 2000 288 2034
rect 254 1932 288 1966
rect 254 1864 288 1898
rect 254 1796 288 1830
rect 254 1727 288 1761
rect 254 1658 288 1692
rect 254 1589 288 1623
rect 254 1520 288 1554
rect 838 2527 872 2561
rect 838 2458 872 2492
rect 838 2389 872 2423
rect 838 2320 872 2354
rect 838 2251 872 2285
rect 838 2182 872 2216
rect 838 2114 872 2148
rect 838 2046 872 2080
rect 838 1978 872 2012
rect 838 1910 872 1944
rect 838 1842 872 1876
rect 838 1774 872 1808
rect 838 1706 872 1740
rect 838 1638 872 1672
rect 838 1570 872 1604
rect 254 1451 288 1485
rect 838 1502 872 1536
rect 838 1434 872 1468
rect 254 1382 288 1416
rect 254 1313 288 1347
rect 254 1244 288 1278
rect 254 1175 288 1209
rect 254 1106 288 1140
rect 254 1037 288 1071
rect 254 968 288 1002
rect 254 899 288 933
rect 254 830 288 864
rect 254 761 288 795
rect 254 692 288 726
rect 254 623 288 657
rect 254 554 288 588
rect 254 485 288 519
rect 254 416 288 450
rect 838 1366 872 1400
rect 838 1298 872 1332
rect 838 1230 872 1264
rect 838 1162 872 1196
rect 838 1094 872 1128
rect 838 1026 872 1060
rect 838 958 872 992
rect 838 890 872 924
rect 838 822 872 856
rect 838 754 872 788
rect 838 686 872 720
rect 838 618 872 652
rect 838 550 872 584
rect 838 482 872 516
rect 838 414 872 448
rect 254 347 288 381
rect 838 346 872 380
rect 254 278 288 312
rect 360 254 394 288
rect 435 254 469 288
rect 510 254 544 288
rect 586 254 620 288
rect 662 254 696 288
rect 738 254 772 288
rect 814 254 848 288
<< mvnsubdiffcont >>
rect 185 3911 219 3945
rect 256 3911 290 3945
rect 327 3911 361 3945
rect 398 3911 432 3945
rect 469 3911 503 3945
rect 539 3911 573 3945
rect 609 3911 643 3945
rect 679 3911 713 3945
rect 749 3911 783 3945
rect 819 3911 853 3945
rect 889 3911 923 3945
rect 68 3761 102 3795
rect 68 3693 102 3727
rect 68 3625 102 3659
rect 68 3557 102 3591
rect 68 3489 102 3523
rect 68 3421 102 3455
rect 68 3353 102 3387
rect 68 3285 102 3319
rect 68 3217 102 3251
rect 68 3149 102 3183
rect 68 3081 102 3115
rect 68 3013 102 3047
rect 68 2945 102 2979
rect 68 2877 102 2911
rect 68 2809 102 2843
rect 68 2741 102 2775
rect 68 2673 102 2707
rect 68 2605 102 2639
rect 68 2537 102 2571
rect 68 2469 102 2503
rect 68 2401 102 2435
rect 68 2333 102 2367
rect 68 2265 102 2299
rect 68 2197 102 2231
rect 68 2129 102 2163
rect 68 2060 102 2094
rect 68 1991 102 2025
rect 68 1922 102 1956
rect 68 1853 102 1887
rect 68 1784 102 1818
rect 68 1715 102 1749
rect 68 1646 102 1680
rect 68 1577 102 1611
rect 68 1508 102 1542
rect 68 1439 102 1473
rect 68 1370 102 1404
rect 68 1301 102 1335
rect 68 1232 102 1266
rect 68 1163 102 1197
rect 68 1094 102 1128
rect 68 1025 102 1059
rect 68 956 102 990
rect 68 887 102 921
rect 68 818 102 852
rect 68 749 102 783
rect 68 680 102 714
rect 68 611 102 645
rect 68 542 102 576
rect 68 473 102 507
rect 68 404 102 438
rect 68 335 102 369
rect 68 266 102 300
rect 68 197 102 231
rect 203 67 237 101
rect 277 67 311 101
rect 351 67 385 101
rect 425 67 459 101
rect 499 67 533 101
rect 573 67 607 101
rect 647 67 681 101
rect 721 67 755 101
rect 796 67 830 101
rect 871 67 905 101
rect 946 67 980 101
<< poly >>
rect 415 2606 711 2624
rect 415 2572 444 2606
rect 478 2572 512 2606
rect 546 2572 580 2606
rect 614 2572 648 2606
rect 682 2572 711 2606
rect 415 2555 711 2572
rect 415 1485 711 1503
rect 415 1451 444 1485
rect 478 1451 512 1485
rect 546 1451 580 1485
rect 614 1451 648 1485
rect 682 1451 711 1485
rect 415 1434 711 1451
rect 428 382 698 386
rect 415 370 711 382
rect 415 336 444 370
rect 478 336 512 370
rect 546 336 580 370
rect 614 336 648 370
rect 682 336 711 370
rect 415 320 711 336
<< polycont >>
rect 444 2572 478 2606
rect 512 2572 546 2606
rect 580 2572 614 2606
rect 648 2572 682 2606
rect 444 1451 478 1485
rect 512 1451 546 1485
rect 580 1451 614 1485
rect 648 1451 682 1485
rect 444 336 478 370
rect 512 336 546 370
rect 580 336 614 370
rect 648 336 682 370
<< locali >>
rect 68 3911 185 3945
rect 219 3911 256 3945
rect 290 3911 327 3945
rect 361 3911 398 3945
rect 432 3911 469 3945
rect 503 3911 539 3945
rect 573 3911 609 3945
rect 643 3911 679 3945
rect 713 3911 749 3945
rect 783 3911 819 3945
rect 853 3911 889 3945
rect 923 3911 1058 3945
rect 68 3841 102 3911
rect 68 3795 102 3807
rect 68 3727 102 3735
rect 68 3659 102 3663
rect 68 3553 102 3557
rect 68 3481 102 3489
rect 68 3409 102 3421
rect 68 3337 102 3353
rect 68 3265 102 3285
rect 68 3193 102 3217
rect 68 3121 102 3149
rect 68 3049 102 3081
rect 68 2979 102 3013
rect 68 2911 102 2943
rect 68 2843 102 2871
rect 68 2775 102 2799
rect 68 2707 102 2726
rect 68 2639 102 2653
rect 68 2571 102 2580
rect 68 2503 102 2507
rect 68 2468 102 2469
rect 68 2395 102 2401
rect 68 2322 102 2333
rect 68 2249 102 2265
rect 68 2176 102 2197
rect 68 2103 102 2129
rect 68 2030 102 2060
rect 68 1957 102 1991
rect 68 1887 102 1922
rect 68 1818 102 1850
rect 68 1749 102 1777
rect 68 1680 102 1704
rect 68 1611 102 1631
rect 68 1542 102 1558
rect 68 1473 102 1485
rect 68 1404 102 1412
rect 68 1335 102 1339
rect 68 1300 102 1301
rect 68 1227 102 1232
rect 68 1154 102 1163
rect 68 1081 102 1094
rect 68 1008 102 1025
rect 68 935 102 956
rect 68 862 102 887
rect 68 789 102 818
rect 68 716 102 749
rect 68 645 102 680
rect 68 576 102 609
rect 68 507 102 536
rect 68 438 102 463
rect 68 369 102 390
rect 68 300 102 317
rect 254 3724 278 3758
rect 312 3724 351 3758
rect 390 3724 423 3758
rect 466 3724 495 3758
rect 542 3724 567 3758
rect 618 3724 660 3758
rect 694 3724 701 3758
rect 735 3724 736 3758
rect 770 3734 872 3758
rect 770 3724 838 3734
rect 254 3666 365 3724
rect 288 3654 365 3666
rect 838 3665 872 3700
rect 360 2631 404 3654
rect 546 3564 580 3606
rect 546 3488 580 3530
rect 546 3413 580 3454
rect 546 3338 580 3379
rect 546 3263 580 3304
rect 546 3188 580 3229
rect 546 3113 580 3154
rect 546 3038 580 3079
rect 546 2963 580 3004
rect 546 2888 580 2929
rect 546 2813 580 2854
rect 546 2738 580 2779
rect 736 3582 770 3620
rect 736 3510 770 3548
rect 736 3438 770 3476
rect 736 3366 770 3404
rect 736 3294 770 3332
rect 736 3222 770 3260
rect 736 3150 770 3188
rect 736 3078 770 3116
rect 736 3006 770 3044
rect 736 2934 770 2972
rect 736 2862 770 2900
rect 736 2790 770 2828
rect 736 2718 770 2756
rect 360 2547 394 2631
rect 472 2606 506 2628
rect 736 2646 770 2684
rect 428 2572 444 2606
rect 478 2590 512 2606
rect 506 2572 512 2590
rect 546 2572 580 2606
rect 614 2572 648 2606
rect 682 2572 698 2606
rect 736 2574 770 2612
rect 360 2108 404 2547
rect 254 2102 404 2108
rect 288 2069 404 2102
rect 288 2036 326 2069
rect 254 2035 326 2036
rect 360 2035 404 2069
rect 254 2034 404 2035
rect 288 2000 404 2034
rect 254 1998 404 2000
rect 288 1996 404 1998
rect 288 1962 326 1996
rect 360 1962 404 1996
rect 288 1932 404 1962
rect 254 1925 404 1932
rect 288 1923 404 1925
rect 288 1889 326 1923
rect 360 1889 404 1923
rect 288 1864 404 1889
rect 254 1852 404 1864
rect 288 1850 404 1852
rect 288 1816 326 1850
rect 360 1816 404 1850
rect 288 1796 404 1816
rect 254 1779 404 1796
rect 288 1777 404 1779
rect 288 1743 326 1777
rect 360 1743 404 1777
rect 288 1727 404 1743
rect 254 1706 404 1727
rect 288 1704 404 1706
rect 288 1670 326 1704
rect 360 1670 404 1704
rect 288 1658 404 1670
rect 254 1633 404 1658
rect 288 1631 404 1633
rect 288 1597 326 1631
rect 360 1597 404 1631
rect 288 1589 404 1597
rect 254 1560 404 1589
rect 546 2443 580 2485
rect 546 2367 580 2409
rect 546 2292 580 2333
rect 546 2217 580 2258
rect 546 2142 580 2183
rect 546 2067 580 2108
rect 546 1992 580 2033
rect 546 1917 580 1958
rect 546 1842 580 1883
rect 546 1767 580 1808
rect 546 1692 580 1733
rect 546 1617 580 1658
rect 736 2502 770 2540
rect 736 2430 770 2468
rect 736 2358 770 2396
rect 736 2286 770 2324
rect 736 2214 770 2252
rect 736 2142 770 2180
rect 736 2069 770 2108
rect 736 1996 770 2035
rect 736 1923 770 1962
rect 736 1850 770 1889
rect 736 1777 770 1816
rect 736 1704 770 1743
rect 736 1631 770 1670
rect 288 1558 404 1560
rect 288 1524 326 1558
rect 360 1524 404 1558
rect 736 1558 770 1597
rect 288 1520 404 1524
rect 254 1510 404 1520
rect 254 1487 394 1510
rect 288 1485 394 1487
rect 472 1485 506 1507
rect 736 1485 770 1524
rect 288 1451 326 1485
rect 360 1451 394 1485
rect 428 1451 444 1485
rect 478 1469 512 1485
rect 506 1451 512 1469
rect 546 1451 580 1485
rect 614 1451 648 1485
rect 682 1451 698 1485
rect 254 1426 394 1451
rect 254 1416 404 1426
rect 288 1412 404 1416
rect 288 1380 326 1412
rect 254 1378 326 1380
rect 360 1378 404 1412
rect 736 1412 770 1451
rect 254 1347 404 1378
rect 288 1339 404 1347
rect 288 1307 326 1339
rect 254 1305 326 1307
rect 360 1305 404 1339
rect 254 1278 404 1305
rect 288 1266 404 1278
rect 288 1234 326 1266
rect 254 1232 326 1234
rect 360 1232 404 1266
rect 254 1209 404 1232
rect 288 1193 404 1209
rect 288 1161 326 1193
rect 254 1159 326 1161
rect 360 1159 404 1193
rect 254 1140 404 1159
rect 288 1120 404 1140
rect 288 1088 326 1120
rect 254 1086 326 1088
rect 360 1086 404 1120
rect 254 1071 404 1086
rect 288 1047 404 1071
rect 288 1015 326 1047
rect 254 1013 326 1015
rect 360 1013 404 1047
rect 254 1002 404 1013
rect 288 974 404 1002
rect 288 942 326 974
rect 254 940 326 942
rect 360 940 404 974
rect 254 933 404 940
rect 288 901 404 933
rect 288 869 326 901
rect 254 867 326 869
rect 360 867 404 901
rect 254 864 404 867
rect 288 828 404 864
rect 288 796 326 828
rect 254 795 326 796
rect 288 794 326 795
rect 360 794 404 828
rect 288 761 404 794
rect 254 757 404 761
rect 288 755 404 757
rect 288 721 326 755
rect 360 721 404 755
rect 288 692 404 721
rect 254 684 404 692
rect 288 682 404 684
rect 288 648 326 682
rect 360 648 404 682
rect 288 623 404 648
rect 254 611 404 623
rect 288 609 404 611
rect 288 575 326 609
rect 360 575 404 609
rect 288 554 404 575
rect 254 538 404 554
rect 288 536 404 538
rect 288 502 326 536
rect 360 502 404 536
rect 288 485 404 502
rect 254 465 404 485
rect 288 463 404 465
rect 288 429 326 463
rect 360 462 404 463
rect 546 1322 580 1364
rect 546 1246 580 1288
rect 546 1171 580 1212
rect 546 1096 580 1137
rect 546 1021 580 1062
rect 546 946 580 987
rect 546 871 580 912
rect 546 796 580 837
rect 546 721 580 762
rect 546 646 580 687
rect 546 571 580 612
rect 546 496 580 537
rect 736 1339 770 1378
rect 736 1266 770 1305
rect 736 1193 770 1232
rect 736 1120 770 1159
rect 736 1047 770 1086
rect 736 974 770 1013
rect 736 901 770 940
rect 736 828 770 867
rect 736 755 770 794
rect 736 682 770 721
rect 736 609 770 648
rect 736 536 770 575
rect 736 463 770 502
rect 288 416 360 429
rect 254 392 360 416
rect 288 390 360 392
rect 288 356 326 390
rect 472 370 506 408
rect 736 390 770 429
rect 288 347 360 356
rect 254 312 360 347
rect 428 336 444 370
rect 506 336 512 370
rect 546 336 580 370
rect 614 336 648 370
rect 682 336 698 370
rect 838 3596 872 3620
rect 838 3527 872 3548
rect 838 3458 872 3476
rect 838 3389 872 3404
rect 838 3320 872 3332
rect 838 3251 872 3260
rect 838 3182 872 3188
rect 838 3113 872 3116
rect 838 3078 872 3079
rect 838 3006 872 3010
rect 838 2934 872 2941
rect 838 2862 872 2872
rect 838 2790 872 2803
rect 838 2718 872 2734
rect 838 2646 872 2665
rect 838 2574 872 2596
rect 838 2502 872 2527
rect 838 2430 872 2458
rect 838 2358 872 2389
rect 838 2286 872 2320
rect 838 2216 872 2251
rect 838 2148 872 2180
rect 838 2080 872 2108
rect 838 2012 872 2036
rect 838 1944 872 1964
rect 838 1876 872 1891
rect 838 1808 872 1818
rect 838 1740 872 1745
rect 838 1633 872 1638
rect 838 1560 872 1570
rect 838 1487 872 1502
rect 838 1414 872 1434
rect 838 1341 872 1366
rect 838 1268 872 1298
rect 838 1196 872 1230
rect 838 1128 872 1161
rect 838 1060 872 1088
rect 838 992 872 1015
rect 838 924 872 942
rect 838 856 872 869
rect 838 788 872 796
rect 838 720 872 723
rect 838 684 872 686
rect 838 611 872 618
rect 838 538 872 550
rect 838 465 872 482
rect 838 392 872 414
rect 288 288 360 312
rect 838 288 872 346
rect 288 278 356 288
rect 254 254 356 278
rect 394 254 432 288
rect 469 254 508 288
rect 544 254 584 288
rect 620 254 660 288
rect 696 254 736 288
rect 772 254 814 288
rect 848 254 872 288
rect 68 231 102 244
rect 68 101 102 171
rect 1024 101 1058 3911
rect 68 67 203 101
rect 237 67 277 101
rect 311 67 351 101
rect 385 67 425 101
rect 459 67 499 101
rect 533 67 573 101
rect 607 67 647 101
rect 681 67 721 101
rect 755 67 796 101
rect 830 67 871 101
rect 905 67 946 101
rect 980 67 1058 101
<< viali >>
rect 68 3807 102 3841
rect 68 3761 102 3769
rect 68 3735 102 3761
rect 68 3693 102 3697
rect 68 3663 102 3693
rect 68 3591 102 3625
rect 68 3523 102 3553
rect 68 3519 102 3523
rect 68 3455 102 3481
rect 68 3447 102 3455
rect 68 3387 102 3409
rect 68 3375 102 3387
rect 68 3319 102 3337
rect 68 3303 102 3319
rect 68 3251 102 3265
rect 68 3231 102 3251
rect 68 3183 102 3193
rect 68 3159 102 3183
rect 68 3115 102 3121
rect 68 3087 102 3115
rect 68 3047 102 3049
rect 68 3015 102 3047
rect 68 2945 102 2977
rect 68 2943 102 2945
rect 68 2877 102 2905
rect 68 2871 102 2877
rect 68 2809 102 2833
rect 68 2799 102 2809
rect 68 2741 102 2760
rect 68 2726 102 2741
rect 68 2673 102 2687
rect 68 2653 102 2673
rect 68 2605 102 2614
rect 68 2580 102 2605
rect 68 2537 102 2541
rect 68 2507 102 2537
rect 68 2435 102 2468
rect 68 2434 102 2435
rect 68 2367 102 2395
rect 68 2361 102 2367
rect 68 2299 102 2322
rect 68 2288 102 2299
rect 68 2231 102 2249
rect 68 2215 102 2231
rect 68 2163 102 2176
rect 68 2142 102 2163
rect 68 2094 102 2103
rect 68 2069 102 2094
rect 68 2025 102 2030
rect 68 1996 102 2025
rect 68 1956 102 1957
rect 68 1923 102 1956
rect 68 1853 102 1884
rect 68 1850 102 1853
rect 68 1784 102 1811
rect 68 1777 102 1784
rect 68 1715 102 1738
rect 68 1704 102 1715
rect 68 1646 102 1665
rect 68 1631 102 1646
rect 68 1577 102 1592
rect 68 1558 102 1577
rect 68 1508 102 1519
rect 68 1485 102 1508
rect 68 1439 102 1446
rect 68 1412 102 1439
rect 68 1370 102 1373
rect 68 1339 102 1370
rect 68 1266 102 1300
rect 68 1197 102 1227
rect 68 1193 102 1197
rect 68 1128 102 1154
rect 68 1120 102 1128
rect 68 1059 102 1081
rect 68 1047 102 1059
rect 68 990 102 1008
rect 68 974 102 990
rect 68 921 102 935
rect 68 901 102 921
rect 68 852 102 862
rect 68 828 102 852
rect 68 783 102 789
rect 68 755 102 783
rect 68 714 102 716
rect 68 682 102 714
rect 68 611 102 643
rect 68 609 102 611
rect 68 542 102 570
rect 68 536 102 542
rect 68 473 102 497
rect 68 463 102 473
rect 68 404 102 424
rect 68 390 102 404
rect 68 335 102 351
rect 68 317 102 335
rect 68 266 102 278
rect 68 244 102 266
rect 356 3724 385 3758
rect 385 3724 390 3758
rect 432 3724 457 3758
rect 457 3724 466 3758
rect 508 3724 529 3758
rect 529 3724 542 3758
rect 584 3724 601 3758
rect 601 3724 618 3758
rect 660 3724 694 3758
rect 736 3724 770 3758
rect 254 3632 288 3654
rect 288 3632 360 3654
rect 254 3598 360 3632
rect 254 3564 288 3598
rect 288 3564 360 3598
rect 254 3530 360 3564
rect 254 3496 288 3530
rect 288 3496 360 3530
rect 254 3462 360 3496
rect 254 3428 288 3462
rect 288 3428 360 3462
rect 254 3394 360 3428
rect 254 3360 288 3394
rect 288 3360 360 3394
rect 254 3326 360 3360
rect 254 3292 288 3326
rect 288 3292 360 3326
rect 254 3258 360 3292
rect 254 3224 288 3258
rect 288 3224 360 3258
rect 254 3190 360 3224
rect 254 3156 288 3190
rect 288 3156 360 3190
rect 254 3122 360 3156
rect 254 3088 288 3122
rect 288 3088 360 3122
rect 254 3054 360 3088
rect 254 3020 288 3054
rect 288 3020 360 3054
rect 254 2986 360 3020
rect 254 2952 288 2986
rect 288 2952 360 2986
rect 254 2918 360 2952
rect 254 2884 288 2918
rect 288 2884 360 2918
rect 254 2850 360 2884
rect 254 2816 288 2850
rect 288 2816 360 2850
rect 254 2782 360 2816
rect 254 2748 288 2782
rect 288 2748 360 2782
rect 254 2714 360 2748
rect 254 2680 288 2714
rect 288 2680 360 2714
rect 254 2646 360 2680
rect 254 2612 288 2646
rect 288 2612 360 2646
rect 546 3606 580 3640
rect 546 3530 580 3564
rect 546 3454 580 3488
rect 546 3379 580 3413
rect 546 3304 580 3338
rect 546 3229 580 3263
rect 546 3154 580 3188
rect 546 3079 580 3113
rect 546 3004 580 3038
rect 546 2929 580 2963
rect 546 2854 580 2888
rect 546 2779 580 2813
rect 546 2704 580 2738
rect 736 3620 770 3654
rect 736 3548 770 3582
rect 736 3476 770 3510
rect 736 3404 770 3438
rect 736 3332 770 3366
rect 736 3260 770 3294
rect 736 3188 770 3222
rect 736 3116 770 3150
rect 736 3044 770 3078
rect 736 2972 770 3006
rect 736 2900 770 2934
rect 736 2828 770 2862
rect 736 2756 770 2790
rect 736 2684 770 2718
rect 254 2578 360 2612
rect 254 2544 288 2578
rect 288 2544 360 2578
rect 472 2628 506 2662
rect 736 2612 770 2646
rect 472 2572 478 2590
rect 478 2572 506 2590
rect 472 2556 506 2572
rect 254 2510 360 2544
rect 254 2476 288 2510
rect 288 2476 360 2510
rect 254 2442 360 2476
rect 254 2408 288 2442
rect 288 2408 360 2442
rect 254 2374 360 2408
rect 254 2340 288 2374
rect 288 2340 360 2374
rect 254 2306 360 2340
rect 254 2272 288 2306
rect 288 2272 360 2306
rect 254 2238 360 2272
rect 254 2204 288 2238
rect 288 2204 360 2238
rect 254 2170 360 2204
rect 254 2136 288 2170
rect 288 2136 360 2170
rect 254 2108 360 2136
rect 736 2540 770 2574
rect 254 2068 288 2070
rect 254 2036 288 2068
rect 326 2035 360 2069
rect 254 1966 288 1998
rect 254 1964 288 1966
rect 326 1962 360 1996
rect 254 1898 288 1925
rect 254 1891 288 1898
rect 326 1889 360 1923
rect 254 1830 288 1852
rect 254 1818 288 1830
rect 326 1816 360 1850
rect 254 1761 288 1779
rect 254 1745 288 1761
rect 326 1743 360 1777
rect 254 1692 288 1706
rect 254 1672 288 1692
rect 326 1670 360 1704
rect 254 1623 288 1633
rect 254 1599 288 1623
rect 326 1597 360 1631
rect 546 2485 580 2519
rect 546 2409 580 2443
rect 546 2333 580 2367
rect 546 2258 580 2292
rect 546 2183 580 2217
rect 546 2108 580 2142
rect 546 2033 580 2067
rect 546 1958 580 1992
rect 546 1883 580 1917
rect 546 1808 580 1842
rect 546 1733 580 1767
rect 546 1658 580 1692
rect 546 1583 580 1617
rect 736 2468 770 2502
rect 736 2396 770 2430
rect 736 2324 770 2358
rect 736 2252 770 2286
rect 736 2180 770 2214
rect 736 2108 770 2142
rect 736 2035 770 2069
rect 736 1962 770 1996
rect 736 1889 770 1923
rect 736 1816 770 1850
rect 736 1743 770 1777
rect 736 1670 770 1704
rect 736 1597 770 1631
rect 254 1554 288 1560
rect 254 1526 288 1554
rect 326 1524 360 1558
rect 254 1485 288 1487
rect 472 1507 506 1541
rect 736 1524 770 1558
rect 254 1453 288 1485
rect 326 1451 360 1485
rect 472 1451 478 1469
rect 478 1451 506 1469
rect 736 1451 770 1485
rect 472 1435 506 1451
rect 254 1382 288 1414
rect 254 1380 288 1382
rect 326 1378 360 1412
rect 254 1313 288 1341
rect 254 1307 288 1313
rect 326 1305 360 1339
rect 254 1244 288 1268
rect 254 1234 288 1244
rect 326 1232 360 1266
rect 254 1175 288 1195
rect 254 1161 288 1175
rect 326 1159 360 1193
rect 254 1106 288 1122
rect 254 1088 288 1106
rect 326 1086 360 1120
rect 254 1037 288 1049
rect 254 1015 288 1037
rect 326 1013 360 1047
rect 254 968 288 976
rect 254 942 288 968
rect 326 940 360 974
rect 254 899 288 903
rect 254 869 288 899
rect 326 867 360 901
rect 254 796 288 830
rect 326 794 360 828
rect 254 726 288 757
rect 254 723 288 726
rect 326 721 360 755
rect 254 657 288 684
rect 254 650 288 657
rect 326 648 360 682
rect 254 588 288 611
rect 254 577 288 588
rect 326 575 360 609
rect 254 519 288 538
rect 254 504 288 519
rect 326 502 360 536
rect 254 450 288 465
rect 254 431 288 450
rect 326 429 360 463
rect 546 1364 580 1398
rect 546 1288 580 1322
rect 546 1212 580 1246
rect 546 1137 580 1171
rect 546 1062 580 1096
rect 546 987 580 1021
rect 546 912 580 946
rect 546 837 580 871
rect 546 762 580 796
rect 546 687 580 721
rect 546 612 580 646
rect 546 537 580 571
rect 546 462 580 496
rect 736 1378 770 1412
rect 736 1305 770 1339
rect 736 1232 770 1266
rect 736 1159 770 1193
rect 736 1086 770 1120
rect 736 1013 770 1047
rect 736 940 770 974
rect 736 867 770 901
rect 736 794 770 828
rect 736 721 770 755
rect 736 648 770 682
rect 736 575 770 609
rect 736 502 770 536
rect 254 381 288 392
rect 254 358 288 381
rect 326 356 360 390
rect 472 408 506 442
rect 736 429 770 463
rect 472 336 478 370
rect 478 336 506 370
rect 736 356 770 390
rect 838 3631 872 3654
rect 838 3620 872 3631
rect 838 3562 872 3582
rect 838 3548 872 3562
rect 838 3493 872 3510
rect 838 3476 872 3493
rect 838 3424 872 3438
rect 838 3404 872 3424
rect 838 3355 872 3366
rect 838 3332 872 3355
rect 838 3286 872 3294
rect 838 3260 872 3286
rect 838 3217 872 3222
rect 838 3188 872 3217
rect 838 3148 872 3150
rect 838 3116 872 3148
rect 838 3044 872 3078
rect 838 2975 872 3006
rect 838 2972 872 2975
rect 838 2906 872 2934
rect 838 2900 872 2906
rect 838 2837 872 2862
rect 838 2828 872 2837
rect 838 2768 872 2790
rect 838 2756 872 2768
rect 838 2699 872 2718
rect 838 2684 872 2699
rect 838 2630 872 2646
rect 838 2612 872 2630
rect 838 2561 872 2574
rect 838 2540 872 2561
rect 838 2492 872 2502
rect 838 2468 872 2492
rect 838 2423 872 2430
rect 838 2396 872 2423
rect 838 2354 872 2358
rect 838 2324 872 2354
rect 838 2285 872 2286
rect 838 2252 872 2285
rect 838 2182 872 2214
rect 838 2180 872 2182
rect 838 2114 872 2142
rect 838 2108 872 2114
rect 838 2046 872 2070
rect 838 2036 872 2046
rect 838 1978 872 1998
rect 838 1964 872 1978
rect 838 1910 872 1925
rect 838 1891 872 1910
rect 838 1842 872 1852
rect 838 1818 872 1842
rect 838 1774 872 1779
rect 838 1745 872 1774
rect 838 1672 872 1706
rect 838 1604 872 1633
rect 838 1599 872 1604
rect 838 1536 872 1560
rect 838 1526 872 1536
rect 838 1468 872 1487
rect 838 1453 872 1468
rect 838 1400 872 1414
rect 838 1380 872 1400
rect 838 1332 872 1341
rect 838 1307 872 1332
rect 838 1264 872 1268
rect 838 1234 872 1264
rect 838 1162 872 1195
rect 838 1161 872 1162
rect 838 1094 872 1122
rect 838 1088 872 1094
rect 838 1026 872 1049
rect 838 1015 872 1026
rect 838 958 872 976
rect 838 942 872 958
rect 838 890 872 903
rect 838 869 872 890
rect 838 822 872 830
rect 838 796 872 822
rect 838 754 872 757
rect 838 723 872 754
rect 838 652 872 684
rect 838 650 872 652
rect 838 584 872 611
rect 838 577 872 584
rect 838 516 872 538
rect 838 504 872 516
rect 838 448 872 465
rect 838 431 872 448
rect 838 380 872 392
rect 838 358 872 380
rect 356 254 360 288
rect 360 254 390 288
rect 432 254 435 288
rect 435 254 466 288
rect 508 254 510 288
rect 510 254 542 288
rect 584 254 586 288
rect 586 254 618 288
rect 660 254 662 288
rect 662 254 694 288
rect 736 254 738 288
rect 738 254 770 288
rect 68 197 102 205
rect 68 171 102 197
<< metal1 >>
rect 62 3841 108 3951
rect 62 3807 68 3841
rect 102 3807 108 3841
rect 62 3769 108 3807
rect 62 3735 68 3769
rect 102 3735 108 3769
rect 62 3697 108 3735
rect 62 3663 68 3697
rect 102 3663 108 3697
rect 62 3625 108 3663
rect 62 3591 68 3625
rect 102 3591 108 3625
rect 62 3553 108 3591
rect 62 3519 68 3553
rect 102 3519 108 3553
rect 62 3481 108 3519
rect 62 3447 68 3481
rect 102 3447 108 3481
rect 62 3409 108 3447
rect 62 3375 68 3409
rect 102 3375 108 3409
rect 62 3337 108 3375
rect 62 3303 68 3337
rect 102 3303 108 3337
rect 62 3265 108 3303
rect 62 3231 68 3265
rect 102 3231 108 3265
rect 62 3193 108 3231
rect 62 3159 68 3193
rect 102 3159 108 3193
rect 62 3121 108 3159
rect 62 3087 68 3121
rect 102 3087 108 3121
rect 62 3049 108 3087
rect 62 3015 68 3049
rect 102 3015 108 3049
rect 62 2977 108 3015
rect 62 2943 68 2977
rect 102 2943 108 2977
rect 62 2905 108 2943
rect 62 2871 68 2905
rect 102 2871 108 2905
rect 62 2833 108 2871
rect 62 2799 68 2833
rect 102 2799 108 2833
rect 62 2760 108 2799
rect 62 2726 68 2760
rect 102 2726 108 2760
rect 62 2687 108 2726
rect 62 2653 68 2687
rect 102 2653 108 2687
rect 62 2614 108 2653
rect 62 2580 68 2614
rect 102 2580 108 2614
rect 62 2541 108 2580
rect 62 2507 68 2541
rect 102 2507 108 2541
rect 62 2468 108 2507
rect 62 2434 68 2468
rect 102 2434 108 2468
rect 62 2395 108 2434
rect 62 2361 68 2395
rect 102 2361 108 2395
rect 62 2322 108 2361
rect 62 2288 68 2322
rect 102 2288 108 2322
rect 62 2249 108 2288
rect 62 2215 68 2249
rect 102 2215 108 2249
rect 62 2176 108 2215
rect 62 2142 68 2176
rect 102 2142 108 2176
rect 62 2103 108 2142
rect 62 2069 68 2103
rect 102 2069 108 2103
rect 62 2030 108 2069
rect 62 1996 68 2030
rect 102 1996 108 2030
rect 62 1957 108 1996
rect 62 1923 68 1957
rect 102 1923 108 1957
rect 62 1884 108 1923
rect 62 1850 68 1884
rect 102 1850 108 1884
rect 62 1811 108 1850
rect 62 1777 68 1811
rect 102 1777 108 1811
rect 62 1738 108 1777
rect 62 1704 68 1738
rect 102 1704 108 1738
rect 62 1665 108 1704
rect 62 1631 68 1665
rect 102 1631 108 1665
rect 62 1592 108 1631
rect 62 1558 68 1592
rect 102 1558 108 1592
rect 62 1519 108 1558
rect 62 1485 68 1519
rect 102 1485 108 1519
rect 62 1446 108 1485
rect 62 1412 68 1446
rect 102 1412 108 1446
rect 62 1373 108 1412
rect 62 1339 68 1373
rect 102 1339 108 1373
rect 62 1300 108 1339
rect 62 1266 68 1300
rect 102 1266 108 1300
rect 62 1227 108 1266
rect 62 1193 68 1227
rect 102 1193 108 1227
rect 62 1154 108 1193
rect 62 1120 68 1154
rect 102 1120 108 1154
rect 62 1081 108 1120
rect 62 1047 68 1081
rect 102 1047 108 1081
rect 62 1008 108 1047
rect 62 974 68 1008
rect 102 974 108 1008
rect 62 935 108 974
rect 62 901 68 935
rect 102 901 108 935
rect 62 862 108 901
rect 62 828 68 862
rect 102 828 108 862
rect 62 789 108 828
rect 62 755 68 789
rect 102 755 108 789
rect 62 716 108 755
rect 62 682 68 716
rect 102 682 108 716
rect 62 643 108 682
rect 62 609 68 643
rect 102 609 108 643
rect 62 570 108 609
rect 62 536 68 570
rect 102 536 108 570
rect 62 497 108 536
rect 62 463 68 497
rect 102 463 108 497
rect 62 424 108 463
rect 62 390 68 424
rect 102 390 108 424
rect 62 351 108 390
rect 62 317 68 351
rect 102 317 108 351
rect 62 278 108 317
rect 62 244 68 278
rect 102 244 108 278
rect 248 3758 878 3764
rect 248 3724 356 3758
rect 390 3724 432 3758
rect 466 3724 508 3758
rect 542 3724 584 3758
rect 618 3724 660 3758
rect 694 3724 736 3758
rect 770 3724 878 3758
rect 248 3718 878 3724
rect 248 3654 366 3718
tri 366 3682 402 3718 nw
tri 694 3682 730 3718 ne
rect 248 2108 254 3654
rect 360 2108 366 3654
rect 730 3654 878 3718
rect 248 2070 366 2108
rect 248 2036 254 2070
rect 288 2069 366 2070
rect 288 2036 326 2069
rect 248 2035 326 2036
rect 360 2035 366 2069
rect 248 1998 366 2035
rect 248 1964 254 1998
rect 288 1996 366 1998
rect 288 1964 326 1996
rect 248 1962 326 1964
rect 360 1962 366 1996
rect 248 1925 366 1962
rect 248 1891 254 1925
rect 288 1923 366 1925
rect 288 1891 326 1923
rect 248 1889 326 1891
rect 360 1889 366 1923
rect 248 1852 366 1889
rect 248 1818 254 1852
rect 288 1850 366 1852
rect 288 1818 326 1850
rect 248 1816 326 1818
rect 360 1816 366 1850
rect 248 1779 366 1816
rect 248 1745 254 1779
rect 288 1777 366 1779
rect 288 1745 326 1777
rect 248 1743 326 1745
rect 360 1743 366 1777
rect 248 1706 366 1743
rect 248 1672 254 1706
rect 288 1704 366 1706
rect 288 1672 326 1704
rect 248 1670 326 1672
rect 360 1670 366 1704
rect 248 1633 366 1670
rect 248 1599 254 1633
rect 288 1631 366 1633
rect 288 1599 326 1631
rect 248 1597 326 1599
rect 360 1597 366 1631
rect 248 1560 366 1597
rect 248 1526 254 1560
rect 288 1558 366 1560
rect 288 1526 326 1558
rect 248 1524 326 1526
rect 360 1524 366 1558
rect 248 1487 366 1524
rect 248 1453 254 1487
rect 288 1485 366 1487
rect 288 1453 326 1485
rect 248 1451 326 1453
rect 360 1451 366 1485
rect 248 1414 366 1451
rect 248 1380 254 1414
rect 288 1412 366 1414
rect 288 1380 326 1412
rect 248 1378 326 1380
rect 360 1378 366 1412
rect 248 1341 366 1378
rect 248 1307 254 1341
rect 288 1339 366 1341
rect 288 1307 326 1339
rect 248 1305 326 1307
rect 360 1305 366 1339
rect 248 1268 366 1305
rect 248 1234 254 1268
rect 288 1266 366 1268
rect 288 1234 326 1266
rect 248 1232 326 1234
rect 360 1232 366 1266
rect 248 1195 366 1232
rect 248 1161 254 1195
rect 288 1193 366 1195
rect 288 1161 326 1193
rect 248 1159 326 1161
rect 360 1159 366 1193
rect 248 1122 366 1159
rect 248 1088 254 1122
rect 288 1120 366 1122
rect 288 1088 326 1120
rect 248 1086 326 1088
rect 360 1086 366 1120
rect 248 1049 366 1086
rect 248 1015 254 1049
rect 288 1047 366 1049
rect 288 1015 326 1047
rect 248 1013 326 1015
rect 360 1013 366 1047
rect 248 976 366 1013
rect 248 942 254 976
rect 288 974 366 976
rect 288 942 326 974
rect 248 940 326 942
rect 360 940 366 974
rect 248 903 366 940
rect 248 869 254 903
rect 288 901 366 903
rect 288 869 326 901
rect 248 867 326 869
rect 360 867 366 901
rect 248 830 366 867
rect 248 796 254 830
rect 288 828 366 830
rect 288 796 326 828
rect 248 794 326 796
rect 360 794 366 828
rect 248 757 366 794
rect 248 723 254 757
rect 288 755 366 757
rect 288 723 326 755
rect 248 721 326 723
rect 360 721 366 755
rect 248 684 366 721
rect 248 650 254 684
rect 288 682 366 684
rect 288 650 326 682
rect 248 648 326 650
rect 360 648 366 682
rect 248 611 366 648
rect 248 577 254 611
rect 288 609 366 611
rect 288 577 326 609
rect 248 575 326 577
rect 360 575 366 609
rect 248 538 366 575
rect 248 504 254 538
rect 288 536 366 538
rect 288 504 326 536
rect 248 502 326 504
rect 360 502 366 536
rect 248 465 366 502
rect 248 431 254 465
rect 288 463 366 465
rect 288 431 326 463
rect 248 429 326 431
rect 360 429 366 463
rect 248 392 366 429
rect 248 358 254 392
rect 288 390 366 392
rect 288 358 326 390
rect 248 356 326 358
rect 360 356 366 390
rect 248 294 366 356
rect 466 2662 512 3645
rect 466 2628 472 2662
rect 506 2628 512 2662
rect 466 2590 512 2628
rect 466 2556 472 2590
rect 506 2556 512 2590
rect 466 1541 512 2556
rect 466 1507 472 1541
rect 506 1507 512 1541
rect 466 1469 512 1507
rect 466 1435 472 1469
rect 506 1435 512 1469
rect 466 442 512 1435
rect 540 3640 586 3652
rect 540 3606 546 3640
rect 580 3606 586 3640
rect 540 3564 586 3606
rect 540 3530 546 3564
rect 580 3530 586 3564
rect 540 3488 586 3530
rect 540 3454 546 3488
rect 580 3454 586 3488
rect 540 3413 586 3454
rect 540 3379 546 3413
rect 580 3379 586 3413
rect 540 3338 586 3379
rect 540 3304 546 3338
rect 580 3304 586 3338
rect 540 3263 586 3304
rect 540 3229 546 3263
rect 580 3229 586 3263
rect 540 3188 586 3229
rect 540 3154 546 3188
rect 580 3154 586 3188
rect 540 3113 586 3154
rect 540 3079 546 3113
rect 580 3079 586 3113
rect 540 3038 586 3079
rect 540 3004 546 3038
rect 580 3004 586 3038
rect 540 2963 586 3004
rect 540 2929 546 2963
rect 580 2929 586 2963
rect 540 2888 586 2929
rect 540 2854 546 2888
rect 580 2854 586 2888
rect 540 2813 586 2854
rect 540 2779 546 2813
rect 580 2779 586 2813
rect 540 2738 586 2779
rect 540 2704 546 2738
rect 580 2704 586 2738
rect 540 2519 586 2704
rect 540 2485 546 2519
rect 580 2485 586 2519
rect 540 2443 586 2485
rect 540 2409 546 2443
rect 580 2409 586 2443
rect 540 2367 586 2409
rect 540 2333 546 2367
rect 580 2333 586 2367
rect 540 2292 586 2333
rect 540 2258 546 2292
rect 580 2258 586 2292
rect 540 2217 586 2258
rect 540 2183 546 2217
rect 580 2183 586 2217
rect 540 2142 586 2183
rect 540 2108 546 2142
rect 580 2108 586 2142
rect 540 2067 586 2108
rect 540 2033 546 2067
rect 580 2033 586 2067
rect 540 1992 586 2033
rect 540 1958 546 1992
rect 580 1958 586 1992
rect 540 1917 586 1958
rect 540 1883 546 1917
rect 580 1883 586 1917
rect 540 1842 586 1883
rect 540 1808 546 1842
rect 580 1808 586 1842
rect 540 1767 586 1808
rect 540 1733 546 1767
rect 580 1733 586 1767
rect 540 1692 586 1733
rect 540 1658 546 1692
rect 580 1658 586 1692
rect 540 1617 586 1658
rect 540 1583 546 1617
rect 580 1583 586 1617
rect 540 1398 586 1583
rect 540 1364 546 1398
rect 580 1364 586 1398
rect 540 1322 586 1364
rect 540 1288 546 1322
rect 580 1288 586 1322
rect 540 1246 586 1288
rect 540 1212 546 1246
rect 580 1212 586 1246
rect 540 1171 586 1212
rect 540 1137 546 1171
rect 580 1137 586 1171
rect 540 1096 586 1137
rect 540 1062 546 1096
rect 580 1062 586 1096
rect 540 1021 586 1062
rect 540 987 546 1021
rect 580 987 586 1021
rect 540 946 586 987
rect 540 912 546 946
rect 580 912 586 946
rect 540 871 586 912
rect 540 837 546 871
rect 580 837 586 871
rect 540 796 586 837
rect 540 762 546 796
rect 580 762 586 796
rect 540 721 586 762
rect 540 687 546 721
rect 580 687 586 721
rect 540 646 586 687
rect 540 612 546 646
rect 580 612 586 646
rect 540 571 586 612
rect 540 537 546 571
rect 580 537 586 571
rect 540 496 586 537
rect 540 462 546 496
rect 580 462 586 496
rect 540 450 586 462
rect 730 3620 736 3654
rect 770 3620 838 3654
rect 872 3620 878 3654
rect 730 3582 878 3620
rect 730 3548 736 3582
rect 770 3548 838 3582
rect 872 3548 878 3582
rect 730 3510 878 3548
rect 730 3476 736 3510
rect 770 3476 838 3510
rect 872 3476 878 3510
rect 730 3438 878 3476
rect 730 3404 736 3438
rect 770 3404 838 3438
rect 872 3404 878 3438
rect 730 3366 878 3404
rect 730 3332 736 3366
rect 770 3332 838 3366
rect 872 3332 878 3366
rect 730 3294 878 3332
rect 730 3260 736 3294
rect 770 3260 838 3294
rect 872 3260 878 3294
rect 730 3222 878 3260
rect 730 3188 736 3222
rect 770 3188 838 3222
rect 872 3188 878 3222
rect 730 3150 878 3188
rect 730 3116 736 3150
rect 770 3116 838 3150
rect 872 3116 878 3150
rect 730 3078 878 3116
rect 730 3044 736 3078
rect 770 3044 838 3078
rect 872 3044 878 3078
rect 730 3006 878 3044
rect 730 2972 736 3006
rect 770 2972 838 3006
rect 872 2972 878 3006
rect 730 2934 878 2972
rect 730 2900 736 2934
rect 770 2900 838 2934
rect 872 2900 878 2934
rect 730 2862 878 2900
rect 730 2828 736 2862
rect 770 2828 838 2862
rect 872 2828 878 2862
rect 730 2790 878 2828
rect 730 2756 736 2790
rect 770 2756 838 2790
rect 872 2756 878 2790
rect 730 2718 878 2756
rect 730 2684 736 2718
rect 770 2684 838 2718
rect 872 2684 878 2718
rect 730 2646 878 2684
rect 730 2612 736 2646
rect 770 2612 838 2646
rect 872 2612 878 2646
rect 730 2574 878 2612
rect 730 2540 736 2574
rect 770 2540 838 2574
rect 872 2540 878 2574
rect 730 2502 878 2540
rect 730 2468 736 2502
rect 770 2468 838 2502
rect 872 2468 878 2502
rect 730 2430 878 2468
rect 730 2396 736 2430
rect 770 2396 838 2430
rect 872 2396 878 2430
rect 730 2358 878 2396
rect 730 2324 736 2358
rect 770 2324 838 2358
rect 872 2324 878 2358
rect 730 2286 878 2324
rect 730 2252 736 2286
rect 770 2252 838 2286
rect 872 2252 878 2286
rect 730 2214 878 2252
rect 730 2180 736 2214
rect 770 2180 838 2214
rect 872 2180 878 2214
rect 730 2142 878 2180
rect 730 2108 736 2142
rect 770 2108 838 2142
rect 872 2108 878 2142
rect 730 2070 878 2108
rect 730 2069 838 2070
rect 730 2035 736 2069
rect 770 2036 838 2069
rect 872 2036 878 2070
rect 770 2035 878 2036
rect 730 1998 878 2035
rect 730 1996 838 1998
rect 730 1962 736 1996
rect 770 1964 838 1996
rect 872 1964 878 1998
rect 770 1962 878 1964
rect 730 1925 878 1962
rect 730 1923 838 1925
rect 730 1889 736 1923
rect 770 1891 838 1923
rect 872 1891 878 1925
rect 770 1889 878 1891
rect 730 1852 878 1889
rect 730 1850 838 1852
rect 730 1816 736 1850
rect 770 1818 838 1850
rect 872 1818 878 1852
rect 770 1816 878 1818
rect 730 1779 878 1816
rect 730 1777 838 1779
rect 730 1743 736 1777
rect 770 1745 838 1777
rect 872 1745 878 1779
rect 770 1743 878 1745
rect 730 1706 878 1743
rect 730 1704 838 1706
rect 730 1670 736 1704
rect 770 1672 838 1704
rect 872 1672 878 1706
rect 770 1670 878 1672
rect 730 1633 878 1670
rect 730 1631 838 1633
rect 730 1597 736 1631
rect 770 1599 838 1631
rect 872 1599 878 1633
rect 770 1597 878 1599
rect 730 1560 878 1597
rect 730 1558 838 1560
rect 730 1524 736 1558
rect 770 1526 838 1558
rect 872 1526 878 1560
rect 770 1524 878 1526
rect 730 1487 878 1524
rect 730 1485 838 1487
rect 730 1451 736 1485
rect 770 1453 838 1485
rect 872 1453 878 1487
rect 770 1451 878 1453
rect 730 1414 878 1451
rect 730 1412 838 1414
rect 730 1378 736 1412
rect 770 1380 838 1412
rect 872 1380 878 1414
rect 770 1378 878 1380
rect 730 1341 878 1378
rect 730 1339 838 1341
rect 730 1305 736 1339
rect 770 1307 838 1339
rect 872 1307 878 1341
rect 770 1305 878 1307
rect 730 1268 878 1305
rect 730 1266 838 1268
rect 730 1232 736 1266
rect 770 1234 838 1266
rect 872 1234 878 1268
rect 770 1232 878 1234
rect 730 1195 878 1232
rect 730 1193 838 1195
rect 730 1159 736 1193
rect 770 1161 838 1193
rect 872 1161 878 1195
rect 770 1159 878 1161
rect 730 1122 878 1159
rect 730 1120 838 1122
rect 730 1086 736 1120
rect 770 1088 838 1120
rect 872 1088 878 1122
rect 770 1086 878 1088
rect 730 1049 878 1086
rect 730 1047 838 1049
rect 730 1013 736 1047
rect 770 1015 838 1047
rect 872 1015 878 1049
rect 770 1013 878 1015
rect 730 976 878 1013
rect 730 974 838 976
rect 730 940 736 974
rect 770 942 838 974
rect 872 942 878 976
rect 770 940 878 942
rect 730 903 878 940
rect 730 901 838 903
rect 730 867 736 901
rect 770 869 838 901
rect 872 869 878 903
rect 770 867 878 869
rect 730 830 878 867
rect 730 828 838 830
rect 730 794 736 828
rect 770 796 838 828
rect 872 796 878 830
rect 770 794 878 796
rect 730 757 878 794
rect 730 755 838 757
rect 730 721 736 755
rect 770 723 838 755
rect 872 723 878 757
rect 770 721 878 723
rect 730 684 878 721
rect 730 682 838 684
rect 730 648 736 682
rect 770 650 838 682
rect 872 650 878 684
rect 770 648 878 650
rect 730 611 878 648
rect 730 609 838 611
rect 730 575 736 609
rect 770 577 838 609
rect 872 577 878 611
rect 770 575 878 577
rect 730 538 878 575
rect 730 536 838 538
rect 730 502 736 536
rect 770 504 838 536
rect 872 504 878 538
rect 770 502 878 504
rect 730 465 878 502
rect 730 463 838 465
rect 466 408 472 442
rect 506 408 512 442
rect 466 370 512 408
rect 466 336 472 370
rect 506 336 512 370
tri 366 294 402 330 sw
rect 466 324 512 336
rect 730 429 736 463
rect 770 431 838 463
rect 872 431 878 465
rect 770 429 878 431
rect 730 392 878 429
rect 730 390 838 392
rect 730 356 736 390
rect 770 358 838 390
rect 872 358 878 392
rect 770 356 878 358
tri 724 324 730 330 se
rect 730 324 878 356
tri 694 294 724 324 se
rect 724 294 878 324
rect 248 288 878 294
rect 248 254 356 288
rect 390 254 432 288
rect 466 254 508 288
rect 542 254 584 288
rect 618 254 660 288
rect 694 254 736 288
rect 770 254 878 288
rect 248 248 878 254
rect 62 205 108 244
rect 62 171 68 205
rect 102 171 108 205
rect 62 159 108 171
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1704896540
transform 0 -1 506 1 0 336
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1704896540
transform 0 -1 506 1 0 1435
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1704896540
transform 0 -1 506 1 0 2556
box 0 0 1 1
use nfet_CDNS_52468879185993  nfet_CDNS_52468879185993_0
timestamp 1704896540
transform 1 0 415 0 -1 1408
box -79 -26 375 1026
use nfet_CDNS_52468879185993  nfet_CDNS_52468879185993_1
timestamp 1704896540
transform 1 0 415 0 -1 3650
box -79 -26 375 1026
use nfet_CDNS_52468879185993  nfet_CDNS_52468879185993_2
timestamp 1704896540
transform 1 0 415 0 -1 2529
box -79 -26 375 1026
use PYL1_CDNS_52468879185309  PYL1_CDNS_52468879185309_0
timestamp 1704896540
transform 0 1 428 -1 0 2622
box 0 0 1 1
use PYL1_CDNS_52468879185309  PYL1_CDNS_52468879185309_1
timestamp 1704896540
transform 0 1 428 -1 0 386
box 0 0 1 1
use PYL1_CDNS_52468879185309  PYL1_CDNS_52468879185309_2
timestamp 1704896540
transform 0 1 428 -1 0 1501
box 0 0 1 1
<< labels >>
flabel metal1 s 282 3613 337 3645 7 FreeSans 200 90 0 0 vgnd_io
port 1 nsew
flabel metal1 s 466 3613 512 3645 7 FreeSans 200 90 0 0 pd_h
port 2 nsew
flabel metal1 s 775 3613 830 3645 7 FreeSans 200 90 0 0 vgnd_io
port 1 nsew
flabel metal1 s 72 3904 95 3932 0 FreeSans 200 0 0 0 vcc_io
port 3 nsew
<< properties >>
string GDS_END 91990284
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 91954074
string path 3.375 98.200 24.325 98.200 
<< end >>
