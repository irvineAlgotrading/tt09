magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< pwell >>
rect 0 0 1912 39433
<< ndiff >>
rect 26 39399 86 39407
rect 26 39365 39 39399
rect 73 39365 86 39399
rect 26 39331 86 39365
rect 26 39297 39 39331
rect 73 39297 86 39331
rect 1826 39399 1886 39407
rect 1826 39365 1839 39399
rect 1873 39365 1886 39399
rect 1826 39331 1886 39365
rect 1826 39297 1839 39331
rect 1873 39297 1886 39331
<< ndiffc >>
rect 39 39365 73 39399
rect 39 39297 73 39331
rect 1839 39365 1873 39399
rect 1839 39297 1873 39331
<< ndiffres >>
rect 26 86 86 39297
rect 146 39347 326 39407
rect 146 86 206 39347
rect 26 26 206 86
rect 266 86 326 39347
rect 386 39347 566 39407
rect 386 86 446 39347
rect 266 26 446 86
rect 506 86 566 39347
rect 626 39347 806 39407
rect 626 86 686 39347
rect 506 26 686 86
rect 746 86 806 39347
rect 866 39347 1046 39407
rect 866 86 926 39347
rect 746 26 926 86
rect 986 86 1046 39347
rect 1106 39347 1286 39407
rect 1106 86 1166 39347
rect 986 26 1166 86
rect 1226 86 1286 39347
rect 1346 39347 1526 39407
rect 1346 86 1406 39347
rect 1226 26 1406 86
rect 1466 86 1526 39347
rect 1586 39347 1766 39407
rect 1586 86 1646 39347
rect 1466 26 1646 86
rect 1706 86 1766 39347
rect 1826 86 1886 39297
rect 1706 26 1886 86
<< locali >>
rect 23 39365 39 39399
rect 73 39365 89 39399
rect 23 39331 89 39365
rect 23 39297 39 39331
rect 73 39297 89 39331
rect 1823 39365 1839 39399
rect 1873 39365 1889 39399
rect 1823 39331 1889 39365
rect 1823 39297 1839 39331
rect 1873 39297 1889 39331
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_0
timestamp 1704896540
transform 0 -1 85 -1 0 39339
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_1
timestamp 1704896540
transform 0 -1 1885 -1 0 39407
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_2
timestamp 1704896540
transform 0 -1 85 -1 0 39407
box 0 0 1 1
use DFL1_CDNS_5246887918580  DFL1_CDNS_5246887918580_3
timestamp 1704896540
transform 0 -1 1885 -1 0 39339
box 0 0 1 1
<< properties >>
string GDS_END 6678188
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 6673504
<< end >>
