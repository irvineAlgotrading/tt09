magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -160 2141 4940 2309
rect -160 1386 120 2141
rect 4772 1386 4940 2141
rect -160 1320 45 1386
rect 4847 1320 4940 1386
<< pwell >>
rect -7 1172 137 1260
rect 1999 1172 2079 1260
rect 4755 1172 5069 1260
rect -7 792 79 1172
rect 4813 1014 5069 1172
rect 4813 792 4899 1014
rect -7 700 4899 792
<< psubdiff >>
rect 4940 1210 5043 1234
rect 4957 1176 4991 1210
rect 5025 1176 5043 1210
rect 4940 1139 5043 1176
rect 4957 1105 4991 1139
rect 5025 1105 5043 1139
rect 4940 1040 5043 1105
<< mvpsubdiff >>
rect 19 1200 111 1234
rect 53 1198 111 1200
rect 4781 1210 4940 1234
rect 4781 1198 4923 1210
rect 19 1132 53 1166
rect 19 1064 53 1098
rect 19 996 53 1030
rect 19 928 53 962
rect 19 860 53 894
rect 19 732 53 826
rect 4839 1176 4923 1198
rect 4839 1140 4940 1176
rect 4873 1139 4940 1140
rect 4873 1106 4923 1139
rect 4839 1105 4923 1106
rect 4839 1040 4940 1105
rect 4839 1016 4873 1040
rect 4839 944 4873 982
rect 4839 873 4873 910
rect 4839 802 4873 839
rect 4839 766 4873 768
rect 87 732 121 766
rect 155 732 189 766
rect 223 732 257 766
rect 291 732 325 766
rect 359 732 652 766
rect 686 732 741 766
rect 775 732 1175 766
rect 1209 732 1451 766
rect 1485 732 1559 766
rect 1593 732 1987 766
rect 2021 732 2055 766
rect 2089 732 2163 766
rect 2197 732 2231 766
rect 2265 732 2502 766
rect 2536 732 2570 766
rect 2604 732 2887 766
rect 2921 732 3303 766
rect 3337 732 3371 766
rect 3405 732 3439 766
rect 3473 732 3507 766
rect 3541 732 3575 766
rect 3609 732 3643 766
rect 3677 732 3711 766
rect 3745 732 3779 766
rect 3813 732 3877 766
rect 3911 732 4293 766
rect 4327 732 4597 766
rect 4631 732 4665 766
rect 4699 732 4733 766
rect 4767 732 4873 766
rect 19 726 4873 732
<< mvnsubdiff >>
rect 19 2134 53 2242
rect 87 2208 121 2242
rect 155 2208 189 2242
rect 223 2208 257 2242
rect 291 2208 325 2242
rect 359 2208 393 2242
rect 427 2208 461 2242
rect 495 2208 529 2242
rect 563 2208 597 2242
rect 631 2208 665 2242
rect 699 2208 733 2242
rect 767 2208 801 2242
rect 835 2208 869 2242
rect 903 2208 937 2242
rect 971 2208 1005 2242
rect 1039 2208 1073 2242
rect 1107 2208 1141 2242
rect 1175 2208 1209 2242
rect 1243 2208 1277 2242
rect 1311 2208 1345 2242
rect 1379 2208 1413 2242
rect 1447 2208 1481 2242
rect 1515 2208 1549 2242
rect 1583 2208 1617 2242
rect 1651 2208 1685 2242
rect 1719 2208 1753 2242
rect 1787 2208 1821 2242
rect 1855 2208 1889 2242
rect 1923 2208 1957 2242
rect 1991 2208 2025 2242
rect 2059 2208 2093 2242
rect 2127 2208 2161 2242
rect 2195 2208 2229 2242
rect 2263 2208 2297 2242
rect 2331 2208 2365 2242
rect 2399 2208 2433 2242
rect 2467 2208 2501 2242
rect 2535 2208 2569 2242
rect 2603 2208 2637 2242
rect 2671 2208 2705 2242
rect 2739 2208 2773 2242
rect 2807 2208 2841 2242
rect 2875 2208 2909 2242
rect 2943 2208 2977 2242
rect 3011 2208 3045 2242
rect 3079 2208 3113 2242
rect 3147 2208 3181 2242
rect 3215 2208 3249 2242
rect 3283 2208 3317 2242
rect 3351 2208 3385 2242
rect 3419 2208 3453 2242
rect 3487 2208 3521 2242
rect 3555 2208 3589 2242
rect 3623 2208 3657 2242
rect 3691 2208 3725 2242
rect 3759 2208 3793 2242
rect 3827 2208 3861 2242
rect 3895 2208 3929 2242
rect 3963 2208 3997 2242
rect 4031 2208 4065 2242
rect 4099 2208 4133 2242
rect 4167 2208 4201 2242
rect 4235 2208 4269 2242
rect 4303 2208 4337 2242
rect 4371 2208 4405 2242
rect 4439 2208 4473 2242
rect 4507 2208 4541 2242
rect 4575 2208 4609 2242
rect 4643 2208 4677 2242
rect 4711 2208 4745 2242
rect 4779 2208 4873 2242
rect 19 2066 53 2100
rect 19 1998 53 2032
rect 19 1930 53 1964
rect 19 1862 53 1896
rect 19 1794 53 1828
rect 19 1726 53 1760
rect 19 1658 53 1692
rect 19 1590 53 1624
rect 19 1522 53 1556
rect 19 1454 53 1488
rect 4839 2140 4873 2174
rect 4839 2072 4873 2106
rect 4839 2004 4873 2038
rect 4839 1936 4873 1970
rect 4839 1868 4873 1902
rect 4839 1800 4873 1834
rect 4839 1732 4873 1766
rect 4839 1664 4873 1698
rect 4839 1596 4873 1630
rect 4839 1528 4873 1562
rect 4839 1460 4873 1494
rect 4839 1422 4873 1426
rect 53 1420 111 1422
rect 19 1386 111 1420
rect 4781 1386 4873 1422
<< psubdiffcont >>
rect 4940 1176 4957 1210
rect 4991 1176 5025 1210
rect 4940 1105 4957 1139
rect 4991 1105 5025 1139
<< mvpsubdiffcont >>
rect 19 1166 53 1200
rect 19 1098 53 1132
rect 19 1030 53 1064
rect 19 962 53 996
rect 19 894 53 928
rect 19 826 53 860
rect 4923 1176 4940 1210
rect 4839 1106 4873 1140
rect 4923 1105 4940 1139
rect 4839 982 4873 1016
rect 4839 910 4873 944
rect 4839 839 4873 873
rect 4839 768 4873 802
rect 53 732 87 766
rect 121 732 155 766
rect 189 732 223 766
rect 257 732 291 766
rect 325 732 359 766
rect 652 732 686 766
rect 741 732 775 766
rect 1175 732 1209 766
rect 1451 732 1485 766
rect 1559 732 1593 766
rect 1987 732 2021 766
rect 2055 732 2089 766
rect 2163 732 2197 766
rect 2231 732 2265 766
rect 2502 732 2536 766
rect 2570 732 2604 766
rect 2887 732 2921 766
rect 3303 732 3337 766
rect 3371 732 3405 766
rect 3439 732 3473 766
rect 3507 732 3541 766
rect 3575 732 3609 766
rect 3643 732 3677 766
rect 3711 732 3745 766
rect 3779 732 3813 766
rect 3877 732 3911 766
rect 4293 732 4327 766
rect 4597 732 4631 766
rect 4665 732 4699 766
rect 4733 732 4767 766
<< mvnsubdiffcont >>
rect 53 2208 87 2242
rect 121 2208 155 2242
rect 189 2208 223 2242
rect 257 2208 291 2242
rect 325 2208 359 2242
rect 393 2208 427 2242
rect 461 2208 495 2242
rect 529 2208 563 2242
rect 597 2208 631 2242
rect 665 2208 699 2242
rect 733 2208 767 2242
rect 801 2208 835 2242
rect 869 2208 903 2242
rect 937 2208 971 2242
rect 1005 2208 1039 2242
rect 1073 2208 1107 2242
rect 1141 2208 1175 2242
rect 1209 2208 1243 2242
rect 1277 2208 1311 2242
rect 1345 2208 1379 2242
rect 1413 2208 1447 2242
rect 1481 2208 1515 2242
rect 1549 2208 1583 2242
rect 1617 2208 1651 2242
rect 1685 2208 1719 2242
rect 1753 2208 1787 2242
rect 1821 2208 1855 2242
rect 1889 2208 1923 2242
rect 1957 2208 1991 2242
rect 2025 2208 2059 2242
rect 2093 2208 2127 2242
rect 2161 2208 2195 2242
rect 2229 2208 2263 2242
rect 2297 2208 2331 2242
rect 2365 2208 2399 2242
rect 2433 2208 2467 2242
rect 2501 2208 2535 2242
rect 2569 2208 2603 2242
rect 2637 2208 2671 2242
rect 2705 2208 2739 2242
rect 2773 2208 2807 2242
rect 2841 2208 2875 2242
rect 2909 2208 2943 2242
rect 2977 2208 3011 2242
rect 3045 2208 3079 2242
rect 3113 2208 3147 2242
rect 3181 2208 3215 2242
rect 3249 2208 3283 2242
rect 3317 2208 3351 2242
rect 3385 2208 3419 2242
rect 3453 2208 3487 2242
rect 3521 2208 3555 2242
rect 3589 2208 3623 2242
rect 3657 2208 3691 2242
rect 3725 2208 3759 2242
rect 3793 2208 3827 2242
rect 3861 2208 3895 2242
rect 3929 2208 3963 2242
rect 3997 2208 4031 2242
rect 4065 2208 4099 2242
rect 4133 2208 4167 2242
rect 4201 2208 4235 2242
rect 4269 2208 4303 2242
rect 4337 2208 4371 2242
rect 4405 2208 4439 2242
rect 4473 2208 4507 2242
rect 4541 2208 4575 2242
rect 4609 2208 4643 2242
rect 4677 2208 4711 2242
rect 4745 2208 4779 2242
rect 19 2100 53 2134
rect 19 2032 53 2066
rect 19 1964 53 1998
rect 19 1896 53 1930
rect 19 1828 53 1862
rect 19 1760 53 1794
rect 19 1692 53 1726
rect 19 1624 53 1658
rect 19 1556 53 1590
rect 19 1488 53 1522
rect 19 1420 53 1454
rect 4839 2174 4873 2208
rect 4839 2106 4873 2140
rect 4839 2038 4873 2072
rect 4839 1970 4873 2004
rect 4839 1902 4873 1936
rect 4839 1834 4873 1868
rect 4839 1766 4873 1800
rect 4839 1698 4873 1732
rect 4839 1630 4873 1664
rect 4839 1562 4873 1596
rect 4839 1494 4873 1528
rect 4839 1426 4873 1460
<< locali >>
rect 19 2134 53 2242
rect 87 2208 121 2242
rect 155 2208 189 2242
rect 223 2208 257 2242
rect 291 2208 325 2242
rect 359 2208 393 2242
rect 427 2208 461 2242
rect 495 2208 529 2242
rect 563 2208 597 2242
rect 631 2208 665 2242
rect 699 2208 733 2242
rect 767 2208 801 2242
rect 835 2208 869 2242
rect 903 2208 937 2242
rect 971 2208 1005 2242
rect 1039 2208 1073 2242
rect 1107 2208 1141 2242
rect 1175 2208 1209 2242
rect 1243 2208 1277 2242
rect 1311 2208 1345 2242
rect 1379 2208 1413 2242
rect 1447 2208 1481 2242
rect 1515 2208 1549 2242
rect 1583 2208 1617 2242
rect 1651 2208 1685 2242
rect 1719 2208 1753 2242
rect 1787 2208 1821 2242
rect 1855 2208 1889 2242
rect 1923 2208 1957 2242
rect 1991 2208 2025 2242
rect 2059 2208 2093 2242
rect 2127 2208 2161 2242
rect 2195 2208 2229 2242
rect 2263 2208 2297 2242
rect 2331 2208 2365 2242
rect 2399 2208 2433 2242
rect 2467 2208 2501 2242
rect 2535 2208 2569 2242
rect 2603 2208 2637 2242
rect 2671 2208 2705 2242
rect 2739 2208 2773 2242
rect 2807 2208 2841 2242
rect 2875 2208 2909 2242
rect 2943 2208 2977 2242
rect 3011 2208 3045 2242
rect 3079 2208 3113 2242
rect 3147 2208 3181 2242
rect 3215 2208 3249 2242
rect 3283 2208 3317 2242
rect 3351 2208 3385 2242
rect 3419 2208 3453 2242
rect 3487 2208 3521 2242
rect 3555 2208 3589 2242
rect 3623 2208 3657 2242
rect 3691 2208 3725 2242
rect 3759 2208 3793 2242
rect 3827 2208 3861 2242
rect 3895 2208 3929 2242
rect 3963 2208 3997 2242
rect 4031 2208 4065 2242
rect 4099 2208 4133 2242
rect 4167 2208 4201 2242
rect 4235 2208 4269 2242
rect 4303 2208 4337 2242
rect 4371 2208 4405 2242
rect 4439 2208 4473 2242
rect 4507 2208 4541 2242
rect 4575 2208 4609 2242
rect 4643 2208 4677 2242
rect 4711 2208 4745 2242
rect 4779 2208 4873 2242
rect 19 2066 53 2100
rect 4839 2140 4873 2174
rect 4839 2072 4873 2106
rect 19 1998 53 2032
rect 19 1930 53 1964
rect 19 1862 53 1896
rect 19 1794 53 1828
rect 19 1726 53 1760
rect 311 1958 345 1996
rect 311 1886 345 1924
rect 311 1814 345 1852
rect 311 1742 345 1780
rect 597 1958 631 1996
rect 597 1886 631 1924
rect 597 1814 631 1852
rect 597 1742 631 1780
rect 949 1958 983 1996
rect 949 1886 983 1924
rect 949 1814 983 1852
rect 1411 1967 1445 2005
rect 1411 1895 1445 1933
rect 1411 1823 1445 1861
rect 1500 1958 1534 1996
rect 1500 1886 1534 1924
rect 1500 1814 1534 1852
rect 949 1742 983 1780
rect 2633 1967 2667 2005
rect 2633 1895 2667 1933
rect 2633 1823 2667 1861
rect 3447 1964 3481 2002
rect 3447 1892 3481 1930
rect 3447 1820 3481 1858
rect 1500 1742 1534 1780
rect 3447 1748 3481 1786
rect 3799 1958 3833 1996
rect 3799 1886 3833 1924
rect 3799 1814 3833 1852
rect 3799 1742 3833 1780
rect 4547 1958 4581 1996
rect 4547 1886 4581 1924
rect 4547 1814 4581 1852
rect 4547 1742 4581 1780
rect 4839 2004 4873 2038
rect 4839 1936 4873 1970
rect 4839 1868 4873 1902
rect 4839 1800 4873 1834
rect 4839 1732 4873 1766
rect 19 1658 53 1692
rect 19 1590 53 1624
rect 19 1522 53 1556
rect 19 1454 53 1488
rect 4839 1664 4873 1698
rect 4839 1596 4873 1630
rect 4839 1528 4873 1562
rect 4839 1460 4873 1494
rect 53 1420 135 1438
rect 19 1404 135 1420
rect 19 1366 169 1404
rect 19 1332 135 1366
rect 773 1366 807 1404
rect 1587 1366 1621 1404
rect 2001 1372 2077 1438
rect 3271 1366 3305 1404
rect 231 1290 265 1328
rect 1777 1290 1811 1328
rect 2179 1290 2213 1328
rect 2537 1290 2571 1328
rect 2919 1290 2953 1328
rect 3909 1366 3943 1404
rect 4757 1426 4839 1438
rect 4757 1372 4873 1426
rect 3095 1290 3129 1328
rect 3367 1290 3401 1328
rect 3535 1290 3569 1328
rect 3799 1290 3833 1328
rect 4085 1290 4119 1328
rect 4261 1290 4295 1328
rect 4643 1290 4677 1328
rect 19 1216 135 1248
rect 19 1200 63 1216
rect 53 1182 63 1200
rect 97 1182 135 1216
rect 2001 1182 2077 1248
rect 4757 1210 5076 1248
rect 4757 1176 4839 1210
rect 4873 1176 4921 1210
rect 4957 1176 4991 1210
rect 5027 1176 5076 1210
rect 4757 1173 5076 1176
rect 19 1136 53 1166
rect 19 1064 53 1098
rect 19 996 53 1030
rect 19 928 53 958
rect 4797 1140 5076 1173
rect 4797 1104 4839 1140
rect 4873 1139 5076 1140
rect 4873 1119 4923 1139
rect 4873 1104 4921 1119
rect 4957 1105 4991 1139
rect 5025 1119 5076 1139
rect 4797 1085 4921 1104
rect 4955 1085 4993 1105
rect 5027 1085 5076 1119
rect 4797 1040 5076 1085
rect 4797 1016 4873 1040
rect 4797 982 4839 1016
rect 4797 944 4873 982
rect 19 860 53 872
rect 19 732 53 800
rect 87 732 105 766
rect 155 732 177 766
rect 223 732 249 766
rect 291 732 321 766
rect 359 732 393 766
rect 427 732 439 766
rect 473 607 579 892
rect 753 826 931 892
rect 647 732 652 766
rect 719 732 741 766
rect 507 573 545 607
rect 473 561 579 573
rect 825 127 931 826
rect 1001 367 1107 892
rect 1209 732 1216 766
rect 1287 607 1393 892
rect 1485 732 1505 766
rect 1539 732 1559 766
rect 1321 573 1359 607
rect 1287 567 1393 573
rect 1653 447 1759 892
rect 1687 413 1725 447
rect 1653 407 1759 413
rect 1829 447 1935 892
rect 1969 732 1987 766
rect 2031 732 2055 766
rect 2103 732 2141 766
rect 2197 732 2213 766
rect 2265 732 2283 766
rect 1969 726 2283 732
rect 1863 413 1901 447
rect 1829 407 1935 413
rect 1035 333 1073 367
rect 1001 327 1107 333
rect 2319 287 2425 892
rect 2459 732 2500 766
rect 2536 732 2570 766
rect 2606 732 2651 766
rect 2685 607 2791 892
rect 2825 732 2831 766
rect 2865 732 2887 766
rect 2719 573 2757 607
rect 2685 567 2791 573
rect 2971 367 3077 892
rect 3147 447 3253 892
rect 4797 910 4839 944
rect 3711 840 3745 878
rect 3287 732 3303 766
rect 3337 732 3371 766
rect 3405 732 3439 766
rect 3473 732 3507 766
rect 3541 732 3575 766
rect 3609 732 3643 766
rect 3677 732 3711 766
rect 3745 732 3779 766
rect 3813 732 3877 766
rect 3911 732 3927 766
rect 3181 413 3219 447
rect 3147 407 3253 413
rect 3005 333 3043 367
rect 2971 321 3077 333
rect 2353 253 2391 287
rect 2319 247 2425 253
rect 859 93 897 127
rect 825 87 931 93
rect 3961 127 4067 892
rect 4137 445 4243 892
rect 4277 732 4283 766
rect 4327 732 4355 766
rect 4423 525 4529 892
rect 4797 873 4873 910
rect 4797 839 4839 873
rect 4797 802 4873 839
rect 4797 768 4839 802
rect 4797 766 4873 768
rect 4563 732 4572 766
rect 4631 732 4644 766
rect 4699 732 4716 766
rect 4767 732 4873 766
rect 4563 726 4873 732
rect 4457 491 4495 525
rect 4423 485 4529 491
rect 4171 411 4209 445
rect 4137 405 4243 411
rect 3995 93 4033 127
rect 3961 87 4067 93
<< viali >>
rect 311 1996 345 2030
rect 311 1924 345 1958
rect 311 1852 345 1886
rect 311 1780 345 1814
rect 311 1708 345 1742
rect 597 1996 631 2030
rect 597 1924 631 1958
rect 597 1852 631 1886
rect 597 1780 631 1814
rect 597 1708 631 1742
rect 949 1996 983 2030
rect 949 1924 983 1958
rect 949 1852 983 1886
rect 949 1780 983 1814
rect 1411 2005 1445 2039
rect 1411 1933 1445 1967
rect 1411 1861 1445 1895
rect 1411 1789 1445 1823
rect 1500 1996 1534 2030
rect 1500 1924 1534 1958
rect 1500 1852 1534 1886
rect 949 1708 983 1742
rect 1500 1780 1534 1814
rect 2633 2005 2667 2039
rect 2633 1933 2667 1967
rect 2633 1861 2667 1895
rect 2633 1789 2667 1823
rect 3447 2002 3481 2036
rect 3447 1930 3481 1964
rect 3447 1858 3481 1892
rect 1500 1708 1534 1742
rect 3447 1786 3481 1820
rect 3447 1714 3481 1748
rect 3799 1996 3833 2030
rect 3799 1924 3833 1958
rect 3799 1852 3833 1886
rect 3799 1780 3833 1814
rect 3799 1708 3833 1742
rect 4547 1996 4581 2030
rect 4547 1924 4581 1958
rect 4547 1852 4581 1886
rect 4547 1780 4581 1814
rect 4547 1708 4581 1742
rect 135 1404 169 1438
rect 135 1332 169 1366
rect 773 1404 807 1438
rect 231 1328 265 1362
rect 773 1332 807 1366
rect 1587 1404 1621 1438
rect 3271 1404 3305 1438
rect 1587 1332 1621 1366
rect 231 1256 265 1290
rect 1777 1328 1811 1362
rect 1777 1256 1811 1290
rect 2179 1328 2213 1362
rect 2179 1256 2213 1290
rect 2537 1328 2571 1362
rect 2537 1256 2571 1290
rect 2919 1328 2953 1362
rect 2919 1256 2953 1290
rect 3095 1328 3129 1362
rect 3271 1332 3305 1366
rect 3909 1404 3943 1438
rect 3095 1256 3129 1290
rect 3367 1328 3401 1362
rect 3367 1256 3401 1290
rect 3535 1328 3569 1362
rect 3535 1256 3569 1290
rect 3799 1328 3833 1362
rect 3909 1332 3943 1366
rect 3799 1256 3833 1290
rect 4085 1328 4119 1362
rect 4085 1256 4119 1290
rect 4261 1328 4295 1362
rect 4261 1256 4295 1290
rect 4643 1328 4677 1362
rect 4643 1256 4677 1290
rect 63 1182 97 1216
rect 135 1182 169 1216
rect 4839 1176 4873 1210
rect 4921 1176 4923 1210
rect 4923 1176 4940 1210
rect 4940 1176 4955 1210
rect 4993 1176 5025 1210
rect 5025 1176 5027 1210
rect 19 1132 53 1136
rect 19 1102 53 1132
rect 19 1030 53 1064
rect 19 962 53 992
rect 19 958 53 962
rect 4839 1106 4873 1138
rect 4839 1104 4873 1106
rect 4921 1105 4923 1119
rect 4923 1105 4940 1119
rect 4940 1105 4955 1119
rect 4993 1105 5025 1119
rect 5025 1105 5027 1119
rect 4921 1085 4955 1105
rect 4993 1085 5027 1105
rect 19 894 53 906
rect 19 872 53 894
rect 19 826 53 834
rect 19 800 53 826
rect 105 732 121 766
rect 121 732 139 766
rect 177 732 189 766
rect 189 732 211 766
rect 249 732 257 766
rect 257 732 283 766
rect 321 732 325 766
rect 325 732 355 766
rect 393 732 427 766
rect 613 732 647 766
rect 685 732 686 766
rect 686 732 719 766
rect 757 732 775 766
rect 775 732 791 766
rect 473 573 507 607
rect 545 573 579 607
rect 1144 732 1175 766
rect 1175 732 1178 766
rect 1216 732 1250 766
rect 1433 732 1451 766
rect 1451 732 1467 766
rect 1505 732 1539 766
rect 1577 732 1593 766
rect 1593 732 1611 766
rect 1287 573 1321 607
rect 1359 573 1393 607
rect 1653 413 1687 447
rect 1725 413 1759 447
rect 1997 732 2021 766
rect 2021 732 2031 766
rect 2069 732 2089 766
rect 2089 732 2103 766
rect 2141 732 2163 766
rect 2163 732 2175 766
rect 2213 732 2231 766
rect 2231 732 2247 766
rect 1829 413 1863 447
rect 1901 413 1935 447
rect 1001 333 1035 367
rect 1073 333 1107 367
rect 2500 732 2502 766
rect 2502 732 2534 766
rect 2572 732 2604 766
rect 2604 732 2606 766
rect 2831 732 2865 766
rect 2903 732 2921 766
rect 2921 732 2937 766
rect 2685 573 2719 607
rect 2757 573 2791 607
rect 3711 878 3745 912
rect 3711 806 3745 840
rect 3147 413 3181 447
rect 3219 413 3253 447
rect 2971 333 3005 367
rect 3043 333 3077 367
rect 2319 253 2353 287
rect 2391 253 2425 287
rect 825 93 859 127
rect 897 93 931 127
rect 4283 732 4293 766
rect 4293 732 4317 766
rect 4355 732 4389 766
rect 4572 732 4597 766
rect 4597 732 4606 766
rect 4644 732 4665 766
rect 4665 732 4678 766
rect 4716 732 4733 766
rect 4733 732 4750 766
rect 4423 491 4457 525
rect 4495 491 4529 525
rect 4137 411 4171 445
rect 4209 411 4243 445
rect 3961 93 3995 127
rect 4033 93 4067 127
<< metal1 >>
rect -12 2202 4878 2350
tri -13 2176 13 2202 ne
rect 13 2119 59 2202
tri 59 2176 85 2202 nw
tri 4707 2176 4733 2202 ne
rect 4832 2119 4878 2202
rect 585 2110 1796 2119
rect 585 2073 1744 2110
rect 299 2030 490 2036
rect 299 1996 311 2030
rect 345 2016 490 2030
rect 345 1996 438 2016
rect 299 1964 438 1996
rect 299 1958 490 1964
rect 299 1924 311 1958
rect 345 1952 490 1958
rect 345 1924 438 1952
rect 299 1900 438 1924
rect 299 1888 490 1900
rect 299 1886 438 1888
rect 299 1852 311 1886
rect 345 1852 438 1886
rect 299 1836 438 1852
rect 299 1824 490 1836
rect 299 1814 438 1824
rect 299 1780 311 1814
rect 345 1780 438 1814
rect 299 1772 438 1780
rect 299 1760 490 1772
rect 299 1742 438 1760
rect 299 1708 311 1742
rect 345 1708 438 1742
rect 299 1702 490 1708
rect 585 2030 643 2073
tri 643 2048 668 2073 nw
tri 1719 2048 1744 2073 ne
rect 1744 2046 1796 2058
rect 1392 2039 1457 2045
rect 585 1996 597 2030
rect 631 1996 643 2030
rect 585 1958 643 1996
rect 585 1924 597 1958
rect 631 1924 643 1958
rect 585 1886 643 1924
rect 585 1852 597 1886
rect 631 1852 643 1886
rect 585 1814 643 1852
rect 585 1780 597 1814
rect 631 1780 643 1814
rect 585 1742 643 1780
rect 585 1708 597 1742
rect 631 1708 643 1742
rect 585 1702 643 1708
rect 937 2030 995 2036
rect 937 1996 949 2030
rect 983 1996 995 2030
rect 937 1958 995 1996
rect 937 1924 949 1958
rect 983 1924 995 1958
rect 937 1886 995 1924
rect 937 1852 949 1886
rect 983 1852 995 1886
rect 937 1814 995 1852
rect 937 1780 949 1814
rect 983 1780 995 1814
rect 1392 2033 1411 2039
rect 1445 2005 1457 2039
rect 1444 1981 1457 2005
rect 1392 1969 1457 1981
rect 1444 1967 1457 1969
rect 1445 1933 1457 1967
rect 1444 1917 1457 1933
rect 1392 1905 1457 1917
rect 1444 1895 1457 1905
rect 1445 1861 1457 1895
rect 1444 1853 1457 1861
rect 1392 1841 1457 1853
rect 1444 1823 1457 1841
rect 1445 1789 1457 1823
rect 1392 1783 1457 1789
rect 1488 2030 1546 2036
rect 1488 1996 1500 2030
rect 1534 1996 1546 2030
rect 1488 1958 1546 1996
rect 1488 1924 1500 1958
rect 1534 1924 1546 1958
rect 1488 1886 1546 1924
rect 1488 1852 1500 1886
rect 1534 1852 1546 1886
rect 2558 2039 2679 2045
rect 1744 1982 1796 1994
rect 1744 1918 1796 1930
rect 1744 1860 1796 1866
rect 2143 2033 2195 2039
rect 2143 1969 2195 1981
rect 2143 1905 2195 1917
tri 2138 1852 2143 1857 se
rect 2558 2033 2633 2039
rect 2610 2005 2633 2033
rect 2667 2005 2679 2039
rect 2610 1981 2679 2005
rect 2558 1969 2679 1981
rect 2610 1967 2679 1969
rect 2610 1933 2633 1967
rect 2667 1933 2679 1967
rect 2610 1917 2679 1933
rect 2558 1905 2679 1917
rect 2143 1852 2195 1853
tri 2195 1852 2200 1857 sw
rect 2610 1895 2679 1905
rect 2610 1861 2633 1895
rect 2667 1861 2679 1895
rect 2610 1853 2679 1861
rect 1488 1814 1546 1852
tri 2118 1832 2138 1852 se
rect 2138 1841 2200 1852
rect 2138 1832 2143 1841
rect 937 1748 995 1780
rect 1488 1780 1500 1814
rect 1534 1780 1546 1814
rect 2195 1832 2200 1841
tri 2200 1832 2220 1852 sw
rect 2558 1841 2679 1853
rect 2143 1783 2195 1789
rect 2610 1823 2679 1841
rect 2610 1789 2633 1823
rect 2667 1789 2679 1823
rect 2558 1783 2679 1789
rect 3386 2036 3493 2042
rect 3386 2016 3447 2036
rect 3438 2002 3447 2016
rect 3481 2002 3493 2036
rect 3438 1964 3493 2002
rect 3386 1952 3447 1964
rect 3438 1930 3447 1952
rect 3481 1930 3493 1964
rect 3438 1900 3493 1930
rect 3386 1892 3493 1900
rect 3386 1888 3447 1892
rect 3438 1858 3447 1888
rect 3481 1858 3493 1892
rect 3438 1836 3493 1858
rect 3386 1824 3493 1836
tri 995 1748 1020 1773 sw
tri 1463 1748 1488 1773 se
rect 1488 1748 1546 1780
rect 937 1742 1546 1748
rect 937 1708 949 1742
rect 983 1708 1500 1742
rect 1534 1708 1546 1742
rect 937 1702 1546 1708
rect 3438 1820 3493 1824
rect 3438 1786 3447 1820
rect 3481 1786 3493 1820
rect 3438 1772 3493 1786
rect 3386 1760 3493 1772
rect 3438 1748 3493 1760
rect 3438 1714 3447 1748
rect 3481 1714 3493 1748
rect 3438 1708 3493 1714
rect 3386 1702 3493 1708
rect 3778 2030 3845 2036
rect 3778 2016 3799 2030
rect 3833 1996 3845 2030
rect 4535 2030 4593 2036
rect 3830 1964 3845 1996
rect 3778 1958 3845 1964
rect 3778 1952 3799 1958
rect 3833 1924 3845 1958
rect 3830 1900 3845 1924
rect 3778 1888 3845 1900
rect 3830 1886 3845 1888
rect 3833 1852 3845 1886
rect 3830 1836 3845 1852
rect 3778 1824 3845 1836
rect 3830 1814 3845 1824
rect 3833 1780 3845 1814
rect 3830 1772 3845 1780
rect 3778 1760 3845 1772
rect 3830 1742 3845 1760
rect 3833 1708 3845 1742
rect 3778 1702 3845 1708
rect 4082 2016 4134 2022
rect 4082 1952 4134 1964
rect 4082 1888 4134 1900
rect 4082 1824 4134 1836
rect 4535 1996 4547 2030
rect 4581 1996 4593 2030
rect 4535 1958 4593 1996
rect 4535 1924 4547 1958
rect 4581 1924 4593 1958
rect 4535 1886 4593 1924
rect 4535 1852 4547 1886
rect 4581 1852 4593 1886
rect 4535 1814 4593 1852
rect 4535 1780 4547 1814
rect 4581 1780 4593 1814
rect 4082 1760 4134 1772
tri 4134 1754 4159 1779 sw
tri 4510 1754 4535 1779 se
rect 4535 1754 4593 1780
rect 4134 1742 4593 1754
rect 4134 1708 4547 1742
rect 4581 1708 4593 1742
rect 4082 1702 4593 1708
tri 59 1687 71 1699 sw
tri 4721 1687 4733 1699 se
tri 0 1674 13 1687 se
rect 59 1674 71 1687
tri 71 1674 84 1687 sw
tri 4708 1674 4721 1687 se
rect 4721 1674 4733 1687
rect 0 1438 4878 1674
rect 0 1404 135 1438
rect 169 1404 773 1438
rect 807 1404 1587 1438
rect 1621 1404 3271 1438
rect 3305 1404 3909 1438
rect 3943 1404 4878 1438
rect 0 1398 4878 1404
tri 98 1373 123 1398 ne
rect 123 1366 181 1398
tri 181 1373 206 1398 nw
tri 736 1373 761 1398 ne
rect 123 1332 135 1366
rect 169 1332 181 1366
rect 123 1326 181 1332
rect 219 1362 277 1368
rect 219 1328 231 1362
rect 265 1328 277 1362
rect 219 1296 277 1328
rect 761 1366 819 1398
tri 819 1373 844 1398 nw
tri 1550 1373 1575 1398 ne
rect 761 1332 773 1366
rect 807 1332 819 1366
rect 761 1326 819 1332
rect 1575 1366 1633 1398
tri 1633 1373 1658 1398 nw
tri 3234 1373 3259 1398 ne
rect 1575 1332 1587 1366
rect 1621 1332 1633 1366
rect 1575 1326 1633 1332
rect 1765 1362 2225 1368
rect 1765 1328 1777 1362
rect 1811 1328 2179 1362
rect 2213 1328 2225 1362
tri 277 1296 302 1321 sw
rect 219 1290 409 1296
rect 219 1256 231 1290
rect 265 1256 409 1290
rect 219 1250 409 1256
rect 1765 1290 2225 1328
rect 1765 1256 1777 1290
rect 1811 1256 2179 1290
rect 2213 1256 2225 1290
rect 1765 1250 2225 1256
rect 2525 1362 3141 1368
rect 2525 1328 2537 1362
rect 2571 1328 2919 1362
rect 2953 1328 3095 1362
rect 3129 1328 3141 1362
rect 2525 1324 3141 1328
rect 3259 1366 3317 1398
tri 3317 1373 3342 1398 nw
tri 3872 1373 3897 1398 ne
rect 3259 1332 3271 1366
rect 3305 1332 3317 1366
rect 3259 1326 3317 1332
rect 3355 1362 3845 1368
rect 3355 1328 3367 1362
rect 3401 1328 3535 1362
rect 3569 1328 3799 1362
rect 3833 1328 3845 1362
rect 2525 1290 2583 1324
tri 2583 1299 2608 1324 nw
tri 2882 1299 2907 1324 ne
rect 2525 1256 2537 1290
rect 2571 1256 2583 1290
rect 2525 1250 2583 1256
rect 2907 1290 3141 1324
rect 2907 1256 2919 1290
rect 2953 1256 3095 1290
rect 3129 1256 3141 1290
rect 2907 1250 3141 1256
rect 3355 1290 3845 1328
rect 3897 1366 3955 1398
tri 3955 1373 3980 1398 nw
rect 3897 1332 3909 1366
rect 3943 1332 3955 1366
rect 3897 1326 3955 1332
rect 4073 1362 4689 1368
rect 4073 1328 4085 1362
rect 4119 1328 4261 1362
rect 4295 1328 4643 1362
rect 4677 1328 4689 1362
rect 3355 1256 3367 1290
rect 3401 1256 3535 1290
rect 3569 1256 3799 1290
rect 3833 1256 3845 1290
rect 3355 1250 3845 1256
rect 4073 1324 4689 1328
rect 4073 1290 4307 1324
tri 4307 1299 4332 1324 nw
tri 4606 1299 4631 1324 ne
rect 4073 1256 4085 1290
rect 4119 1256 4261 1290
rect 4295 1256 4307 1290
rect 4073 1250 4307 1256
rect 4631 1290 4689 1324
rect 4631 1256 4643 1290
rect 4677 1256 4689 1290
rect 4631 1250 4689 1256
rect -128 1176 -122 1228
rect -70 1176 -58 1228
rect -6 1222 0 1228
tri 0 1222 6 1228 sw
rect -6 1219 751 1222
rect -6 1216 524 1219
rect -6 1182 63 1216
rect 97 1215 135 1216
rect 169 1215 524 1216
rect -6 1176 70 1182
tri -52 1138 -14 1176 ne
rect -14 1163 70 1176
rect 122 1163 134 1215
rect 186 1163 198 1215
rect 250 1163 262 1215
rect 314 1163 326 1215
rect 378 1167 524 1215
rect 576 1167 588 1219
rect 640 1167 652 1219
rect 704 1176 751 1219
rect 842 1176 858 1219
rect 704 1167 858 1176
rect 910 1167 922 1219
rect 974 1167 986 1219
rect 1038 1167 1050 1219
rect 1102 1176 1108 1219
rect 1161 1217 5070 1222
rect 1161 1176 1500 1217
rect 1102 1167 1500 1176
rect 378 1165 1500 1167
rect 1552 1165 1564 1217
rect 1616 1165 1628 1217
rect 1680 1165 2229 1217
rect 2281 1165 2293 1217
rect 2345 1216 5070 1217
rect 2345 1165 4475 1216
rect 378 1164 4475 1165
rect 4527 1164 4539 1216
rect 4591 1164 4603 1216
rect 4655 1210 5070 1216
rect 4655 1176 4839 1210
rect 4873 1176 4921 1210
rect 4955 1176 4993 1210
rect 5027 1176 5070 1210
rect 4655 1164 5070 1176
rect 378 1163 5070 1164
rect -14 1148 5070 1163
rect -14 1138 4359 1148
tri -14 1136 -12 1138 ne
rect -12 1136 4359 1138
tri -12 1124 0 1136 ne
rect 0 1102 19 1136
rect 53 1132 4359 1136
rect 53 1102 1167 1132
rect 0 1064 1167 1102
rect 0 1030 19 1064
rect 53 1030 1167 1064
rect 0 992 1167 1030
rect 0 958 19 992
rect 53 958 1167 992
rect 0 952 1167 958
rect 1283 1126 4359 1132
rect 1283 952 1830 1126
rect 0 946 1830 952
rect 1946 1074 2470 1126
rect 2522 1074 2658 1126
rect 2710 1074 3500 1126
rect 1946 1062 3500 1074
rect 1946 1010 2470 1062
rect 2522 1010 2658 1062
rect 2710 1010 3500 1062
rect 1946 998 3500 1010
rect 1946 946 2470 998
rect 2522 946 2658 998
rect 2710 946 3500 998
rect 3616 946 3891 1126
rect 4007 946 4359 1126
rect 4454 1146 4676 1148
rect 4454 1094 4475 1146
rect 4527 1094 4539 1146
rect 4591 1094 4603 1146
rect 4655 1094 4676 1146
rect 4454 1075 4676 1094
rect 4454 1023 4475 1075
rect 4527 1023 4539 1075
rect 4591 1023 4603 1075
rect 4655 1023 4676 1075
rect 4454 1004 4676 1023
rect 4454 952 4475 1004
rect 4527 952 4539 1004
rect 4591 952 4603 1004
rect 4655 952 4676 1004
rect 4454 946 4676 952
rect 4768 1138 5070 1148
rect 4768 1104 4839 1138
rect 4873 1119 5070 1138
rect 4873 1104 4921 1119
rect 4768 1085 4921 1104
rect 4955 1085 4993 1119
rect 5027 1085 5070 1119
rect 4768 1053 5070 1085
rect 4768 946 4833 1053
tri 4833 996 4890 1053 nw
rect -130 906 59 918
rect -130 900 19 906
rect -130 720 -122 900
rect -6 872 19 900
rect 53 872 59 906
rect 3699 912 3757 918
rect 3699 878 3711 912
rect 3745 878 3757 912
rect -6 834 59 872
tri 3674 852 3699 877 se
rect 3699 852 3757 878
rect -6 800 19 834
rect 53 806 59 834
tri 59 806 73 820 sw
rect 53 800 73 806
rect -6 772 73 800
tri 73 772 107 806 sw
rect 2067 800 2073 852
rect 2125 800 2137 852
rect 2189 840 3757 852
rect 2189 806 3711 840
rect 3745 806 3757 840
rect 2189 800 3757 806
tri 4368 800 4468 900 se
rect 4468 800 4879 900
tri 4340 772 4368 800 se
rect 4368 772 4879 800
rect -6 720 70 772
rect 122 766 134 772
rect 186 766 198 772
rect 250 766 262 772
rect 314 766 326 772
rect 378 766 524 772
rect 314 732 321 766
rect 378 732 393 766
rect 427 732 524 766
rect 122 720 134 732
rect 186 720 198 732
rect 250 720 262 732
rect 314 720 326 732
rect 378 720 524 732
rect 576 720 588 772
rect 640 766 652 772
rect 704 766 858 772
rect 647 732 652 766
rect 719 732 757 766
rect 791 732 858 766
rect 640 720 652 732
rect 704 720 858 732
rect 910 720 922 772
rect 974 720 986 772
rect 1038 720 1050 772
rect 1102 766 1500 772
rect 1102 732 1144 766
rect 1178 732 1216 766
rect 1250 732 1433 766
rect 1467 732 1500 766
rect 1102 720 1500 732
rect 1552 720 1564 772
rect 1616 720 1628 772
rect 1680 766 2263 772
rect 1680 732 1997 766
rect 2031 732 2069 766
rect 2103 732 2141 766
rect 2175 732 2213 766
rect 2247 732 2263 766
rect 1680 720 2263 732
rect 2315 720 2327 772
rect 2379 766 3495 772
rect 2379 732 2500 766
rect 2534 732 2572 766
rect 2606 732 2831 766
rect 2865 732 2903 766
rect 2937 732 3495 766
rect 2379 720 3495 732
rect 3547 720 3559 772
rect 3611 720 3879 772
rect 3931 720 3943 772
rect 3995 766 4879 772
rect 3995 732 4283 766
rect 4317 732 4355 766
rect 4389 732 4572 766
rect 4606 732 4644 766
rect 4678 732 4716 766
rect 4750 732 4879 766
rect 3995 720 4879 732
tri 70 613 144 687 se
rect 144 681 3830 687
rect 144 641 3778 681
tri 144 613 172 641 nw
tri 3696 613 3724 641 ne
rect 3724 629 3778 641
rect 3724 617 3830 629
rect 3724 613 3778 617
tri 64 607 70 613 se
rect 70 607 138 613
tri 138 607 144 613 nw
tri 216 607 222 613 se
rect 222 607 3337 613
rect 0 573 104 607
tri 104 573 138 607 nw
tri 182 573 216 607 se
rect 216 573 473 607
rect 507 573 545 607
rect 579 573 1287 607
rect 1321 573 1359 607
rect 1393 573 2685 607
rect 2719 573 2757 607
rect 2791 605 3337 607
tri 3337 605 3345 613 sw
tri 3724 605 3732 613 ne
rect 3732 605 3778 613
rect 2791 573 3345 605
rect 0 559 90 573
tri 90 559 104 573 nw
tri 168 559 182 573 se
rect 182 561 3345 573
rect 182 559 222 561
tri 148 539 168 559 se
rect 168 539 222 559
tri 222 539 244 561 nw
tri 3315 539 3337 561 ne
rect 3337 539 3345 561
tri 134 525 148 539 se
rect 148 525 208 539
tri 208 525 222 539 nw
tri 3337 533 3343 539 ne
rect 3343 533 3345 539
tri 288 525 296 533 se
rect 296 525 3302 533
tri 3302 525 3310 533 sw
tri 3343 531 3345 533 ne
tri 3345 531 3419 605 sw
tri 3732 559 3778 605 ne
rect 3778 559 3830 565
tri 3345 525 3351 531 ne
rect 3351 525 4541 531
tri 100 491 134 525 se
rect 134 491 174 525
tri 174 491 208 525 nw
tri 254 491 288 525 se
rect 288 492 3310 525
tri 3310 492 3343 525 sw
tri 3351 492 3384 525 ne
rect 3384 492 4423 525
rect 288 491 3343 492
tri 3343 491 3344 492 sw
tri 3384 491 3385 492 ne
rect 3385 491 4423 492
rect 4457 491 4495 525
rect 4529 491 4541 525
tri 74 465 100 491 se
rect 100 465 148 491
tri 148 465 174 491 nw
tri 228 465 254 491 se
rect 254 481 3344 491
rect 254 465 296 481
tri 56 447 74 465 se
rect 74 447 130 465
tri 130 447 148 465 nw
tri 222 459 228 465 se
rect 228 459 296 465
tri 296 459 318 481 nw
tri 3280 459 3302 481 ne
rect 3302 459 3344 481
tri 210 447 222 459 se
rect 222 447 284 459
tri 284 447 296 459 nw
tri 3302 453 3308 459 ne
rect 3308 453 3344 459
tri 353 447 359 453 se
rect 359 447 1771 453
tri 22 413 56 447 se
rect 56 413 96 447
tri 96 413 130 447 nw
tri 176 413 210 447 se
rect 210 413 250 447
tri 250 413 284 447 nw
tri 319 413 353 447 se
rect 353 413 1653 447
rect 1687 413 1725 447
rect 1759 413 1771 447
tri 20 411 22 413 se
rect 22 411 94 413
tri 94 411 96 413 nw
tri 174 411 176 413 se
rect 176 411 248 413
tri 248 411 250 413 nw
tri 317 411 319 413 se
rect 319 411 1771 413
tri 18 409 20 411 se
rect 20 409 92 411
tri 92 409 94 411 nw
tri 172 409 174 411 se
rect 174 409 227 411
rect 0 367 50 409
tri 50 367 92 409 nw
tri 148 385 172 409 se
rect 172 390 227 409
tri 227 390 248 411 nw
tri 296 390 317 411 se
rect 317 401 1771 411
rect 1817 447 2073 453
rect 1817 413 1829 447
rect 1863 413 1901 447
rect 1935 413 2073 447
rect 1817 401 2073 413
rect 2125 401 2137 453
rect 2189 447 3265 453
tri 3308 451 3310 453 ne
rect 3310 451 3344 453
tri 3344 451 3384 491 sw
tri 3385 479 3397 491 ne
rect 3397 479 4541 491
rect 2189 413 3147 447
rect 3181 413 3219 447
rect 3253 413 3265 447
tri 3310 445 3316 451 ne
rect 3316 445 4255 451
rect 2189 401 3265 413
tri 3316 411 3350 445 ne
rect 3350 411 4137 445
rect 4171 411 4209 445
rect 4243 411 4255 445
tri 3350 401 3360 411 ne
rect 3360 401 4255 411
rect 317 390 359 401
rect 172 385 222 390
tri 222 385 227 390 nw
tri 291 385 296 390 se
rect 296 385 359 390
tri 130 367 148 385 se
rect 148 367 204 385
tri 204 367 222 385 nw
tri 285 379 291 385 se
rect 291 379 359 385
tri 359 379 381 401 nw
tri 3360 399 3362 401 ne
rect 3362 399 4255 401
tri 273 367 285 379 se
rect 285 372 352 379
tri 352 372 359 379 nw
tri 425 372 426 373 se
rect 426 372 3089 373
rect 285 367 347 372
tri 347 367 352 372 nw
tri 420 367 425 372 se
rect 425 367 3089 372
rect 0 357 40 367
tri 40 357 50 367 nw
tri 120 357 130 367 se
rect 130 357 170 367
tri 96 333 120 357 se
rect 120 333 170 357
tri 170 333 204 367 nw
tri 239 333 273 367 se
rect 273 333 313 367
tri 313 333 347 367 nw
tri 386 333 420 367 se
rect 420 333 1001 367
rect 1035 333 1073 367
rect 1107 333 2971 367
rect 3005 333 3043 367
rect 3077 333 3089 367
tri 92 329 96 333 se
rect 96 329 166 333
tri 166 329 170 333 nw
tri 235 329 239 333 se
rect 239 329 285 333
rect 0 287 124 329
tri 124 287 166 329 nw
tri 211 305 235 329 se
rect 235 305 285 329
tri 285 305 313 333 nw
tri 380 327 386 333 se
rect 386 327 3089 333
tri 358 305 380 327 se
rect 380 321 3089 327
rect 380 305 426 321
tri 193 287 211 305 se
rect 211 287 267 305
tri 267 287 285 305 nw
tri 352 299 358 305 se
rect 358 299 426 305
tri 426 299 448 321 nw
tri 340 287 352 299 se
rect 352 287 414 299
tri 414 287 426 299 nw
rect 2307 287 3157 293
rect 0 277 114 287
tri 114 277 124 287 nw
tri 183 277 193 287 se
rect 193 277 233 287
tri 159 253 183 277 se
rect 183 253 233 277
tri 233 253 267 287 nw
tri 306 253 340 287 se
rect 340 253 380 287
tri 380 253 414 287 nw
rect 2307 253 2319 287
rect 2353 253 2391 287
rect 2425 253 3157 287
tri 155 249 159 253 se
rect 159 249 229 253
tri 229 249 233 253 nw
tri 302 249 306 253 se
rect 306 249 352 253
rect 0 197 177 249
tri 177 197 229 249 nw
tri 294 241 302 249 se
rect 302 241 352 249
tri 278 225 294 241 se
rect 294 225 352 241
tri 352 225 380 253 nw
rect 2307 241 3157 253
rect 3209 241 3221 293
rect 3273 241 3279 293
tri 250 197 278 225 se
rect 278 197 296 225
tri 222 169 250 197 se
rect 250 169 296 197
tri 296 169 352 225 nw
rect 0 127 254 169
tri 254 127 296 169 nw
rect 1236 161 1242 213
rect 1294 161 1306 213
rect 1358 204 3199 213
rect 1358 161 3077 204
tri 3062 152 3071 161 ne
rect 3071 152 3077 161
rect 3129 152 3141 204
rect 3193 152 3199 204
rect 813 127 1986 133
rect 0 123 250 127
tri 250 123 254 127 nw
rect 813 93 825 127
rect 859 93 897 127
rect 931 93 1986 127
rect 813 81 1986 93
rect 2038 81 2050 133
rect 2102 127 3049 133
tri 3049 127 3055 133 sw
tri 3214 127 3220 133 se
rect 3220 127 4079 133
rect 2102 112 3055 127
tri 3055 112 3070 127 sw
tri 3199 112 3214 127 se
rect 3214 112 3961 127
rect 2102 93 3961 112
rect 3995 93 4033 127
rect 4067 93 4079 127
rect 2102 81 4079 93
<< via1 >>
rect 438 1964 490 2016
rect 438 1900 490 1952
rect 438 1836 490 1888
rect 438 1772 490 1824
rect 438 1708 490 1760
rect 1744 2058 1796 2110
rect 1392 2005 1411 2033
rect 1411 2005 1444 2033
rect 1392 1981 1444 2005
rect 1392 1967 1444 1969
rect 1392 1933 1411 1967
rect 1411 1933 1444 1967
rect 1392 1917 1444 1933
rect 1392 1895 1444 1905
rect 1392 1861 1411 1895
rect 1411 1861 1444 1895
rect 1392 1853 1444 1861
rect 1392 1823 1444 1841
rect 1392 1789 1411 1823
rect 1411 1789 1444 1823
rect 1744 1994 1796 2046
rect 1744 1930 1796 1982
rect 1744 1866 1796 1918
rect 2143 1981 2195 2033
rect 2143 1917 2195 1969
rect 2143 1853 2195 1905
rect 2558 1981 2610 2033
rect 2558 1917 2610 1969
rect 2558 1853 2610 1905
rect 2143 1789 2195 1841
rect 2558 1789 2610 1841
rect 3386 1964 3438 2016
rect 3386 1900 3438 1952
rect 3386 1836 3438 1888
rect 3386 1772 3438 1824
rect 3386 1708 3438 1760
rect 3778 1996 3799 2016
rect 3799 1996 3830 2016
rect 3778 1964 3830 1996
rect 3778 1924 3799 1952
rect 3799 1924 3830 1952
rect 3778 1900 3830 1924
rect 3778 1886 3830 1888
rect 3778 1852 3799 1886
rect 3799 1852 3830 1886
rect 3778 1836 3830 1852
rect 3778 1814 3830 1824
rect 3778 1780 3799 1814
rect 3799 1780 3830 1814
rect 3778 1772 3830 1780
rect 3778 1742 3830 1760
rect 3778 1708 3799 1742
rect 3799 1708 3830 1742
rect 4082 1964 4134 2016
rect 4082 1900 4134 1952
rect 4082 1836 4134 1888
rect 4082 1772 4134 1824
rect 4082 1708 4134 1760
rect -122 1176 -70 1228
rect -58 1176 -6 1228
rect 70 1182 97 1215
rect 97 1182 122 1215
rect 70 1163 122 1182
rect 134 1182 135 1215
rect 135 1182 169 1215
rect 169 1182 186 1215
rect 134 1163 186 1182
rect 198 1163 250 1215
rect 262 1163 314 1215
rect 326 1163 378 1215
rect 524 1167 576 1219
rect 588 1167 640 1219
rect 652 1167 704 1219
rect 858 1167 910 1219
rect 922 1167 974 1219
rect 986 1167 1038 1219
rect 1050 1167 1102 1219
rect 1500 1165 1552 1217
rect 1564 1165 1616 1217
rect 1628 1165 1680 1217
rect 2229 1165 2281 1217
rect 2293 1165 2345 1217
rect 4475 1164 4527 1216
rect 4539 1164 4591 1216
rect 4603 1164 4655 1216
rect 1167 952 1283 1132
rect 1830 946 1946 1126
rect 2470 1074 2522 1126
rect 2658 1074 2710 1126
rect 2470 1010 2522 1062
rect 2658 1010 2710 1062
rect 2470 946 2522 998
rect 2658 946 2710 998
rect 3500 946 3616 1126
rect 3891 946 4007 1126
rect 4475 1094 4527 1146
rect 4539 1094 4591 1146
rect 4603 1094 4655 1146
rect 4475 1023 4527 1075
rect 4539 1023 4591 1075
rect 4603 1023 4655 1075
rect 4475 952 4527 1004
rect 4539 952 4591 1004
rect 4603 952 4655 1004
rect -122 720 -6 900
rect 2073 800 2125 852
rect 2137 800 2189 852
rect 70 766 122 772
rect 134 766 186 772
rect 198 766 250 772
rect 262 766 314 772
rect 326 766 378 772
rect 70 732 105 766
rect 105 732 122 766
rect 134 732 139 766
rect 139 732 177 766
rect 177 732 186 766
rect 198 732 211 766
rect 211 732 249 766
rect 249 732 250 766
rect 262 732 283 766
rect 283 732 314 766
rect 326 732 355 766
rect 355 732 378 766
rect 70 720 122 732
rect 134 720 186 732
rect 198 720 250 732
rect 262 720 314 732
rect 326 720 378 732
rect 524 720 576 772
rect 588 766 640 772
rect 652 766 704 772
rect 588 732 613 766
rect 613 732 640 766
rect 652 732 685 766
rect 685 732 704 766
rect 588 720 640 732
rect 652 720 704 732
rect 858 720 910 772
rect 922 720 974 772
rect 986 720 1038 772
rect 1050 720 1102 772
rect 1500 766 1552 772
rect 1500 732 1505 766
rect 1505 732 1539 766
rect 1539 732 1552 766
rect 1500 720 1552 732
rect 1564 766 1616 772
rect 1564 732 1577 766
rect 1577 732 1611 766
rect 1611 732 1616 766
rect 1564 720 1616 732
rect 1628 720 1680 772
rect 2263 720 2315 772
rect 2327 720 2379 772
rect 3495 720 3547 772
rect 3559 720 3611 772
rect 3879 720 3931 772
rect 3943 720 3995 772
rect 3778 629 3830 681
rect 3778 565 3830 617
rect 2073 401 2125 453
rect 2137 401 2189 453
rect 3157 241 3209 293
rect 3221 241 3273 293
rect 1242 161 1294 213
rect 1306 161 1358 213
rect 3077 152 3129 204
rect 3141 152 3193 204
rect 1986 81 2038 133
rect 2050 81 2102 133
<< metal2 >>
rect -128 1176 -122 1228
rect -70 1176 -58 1228
rect -6 1176 0 1228
rect 56 1215 410 2350
rect 438 2016 490 2350
rect 438 1952 490 1964
rect 438 1888 490 1900
rect 438 1824 490 1836
rect 438 1760 490 1772
rect 438 1702 490 1708
rect 56 1163 70 1215
rect 122 1163 134 1215
rect 186 1163 198 1215
rect 250 1163 262 1215
rect 314 1163 326 1215
rect 378 1163 410 1215
rect 56 1146 410 1163
rect 518 1445 786 2350
rect 518 1219 722 1445
tri 722 1381 786 1445 nw
rect 518 1167 524 1219
rect 576 1167 588 1219
rect 640 1167 652 1219
rect 704 1167 722 1219
tri 410 1146 415 1151 sw
rect 56 1132 415 1146
tri 415 1132 429 1146 sw
rect 56 1126 429 1132
tri 429 1126 435 1132 sw
rect -128 720 -122 900
rect -6 720 0 900
rect 56 772 410 1126
tri 410 921 435 946 nw
rect 56 720 70 772
rect 122 720 134 772
rect 186 720 198 772
rect 250 720 262 772
rect 314 720 326 772
rect 378 720 410 772
rect 56 282 410 720
rect 56 0 372 282
tri 372 244 410 282 nw
rect 518 772 722 1167
rect 518 720 524 772
rect 576 720 588 772
rect 640 720 652 772
rect 704 720 722 772
rect 518 81 722 720
rect 842 1219 1110 2350
rect 842 1167 858 1219
rect 910 1167 922 1219
rect 974 1167 986 1219
rect 1038 1167 1050 1219
rect 1102 1167 1110 1219
rect 842 772 1110 1167
rect 1166 2275 1311 2350
rect 1166 1132 1284 2275
tri 1284 2248 1311 2275 nw
tri 1324 2248 1382 2306 se
rect 1382 2284 1434 2350
rect 1382 2248 1386 2284
rect 1166 952 1167 1132
rect 1283 952 1284 1132
rect 1166 946 1284 952
tri 1312 2236 1324 2248 se
rect 1324 2236 1386 2248
tri 1386 2236 1434 2284 nw
rect 842 720 858 772
rect 910 720 922 772
rect 974 720 986 772
rect 1038 720 1050 772
rect 1102 720 1110 772
rect 842 241 1110 720
tri 1110 241 1119 250 sw
rect 842 213 1119 241
tri 1119 213 1147 241 sw
tri 1287 213 1312 238 se
rect 1312 213 1364 2236
tri 1364 2214 1386 2236 nw
rect 1490 2176 1758 2350
rect 842 203 1147 213
tri 1147 203 1157 213 sw
tri 722 81 746 105 sw
rect 518 41 746 81
tri 746 41 786 81 sw
rect 518 0 786 41
rect 842 0 1157 203
rect 1236 161 1242 213
rect 1294 161 1306 213
rect 1358 161 1364 213
rect 1392 2033 1444 2039
rect 1392 1969 1444 1981
rect 1392 1905 1444 1917
rect 1392 1841 1444 1853
rect 1392 0 1444 1789
rect 1490 1217 1716 2176
tri 1716 2134 1758 2176 nw
rect 1814 2176 1918 2350
tri 1814 2166 1824 2176 ne
rect 1490 1165 1500 1217
rect 1552 1165 1564 1217
rect 1616 1165 1628 1217
rect 1680 1165 1716 1217
rect 1490 772 1716 1165
rect 1490 720 1500 772
rect 1552 720 1564 772
rect 1616 720 1628 772
rect 1680 720 1716 772
rect 1490 0 1716 720
rect 1744 2110 1796 2116
rect 1744 2046 1796 2058
rect 1744 1982 1796 1994
rect 1744 1918 1796 1930
rect 1744 0 1796 1866
rect 1824 1254 1918 2176
rect 2143 2033 2195 2039
rect 2143 1969 2195 1981
rect 2143 1905 2195 1917
rect 2143 1841 2195 1853
tri 1918 1254 1952 1288 sw
rect 1824 1126 1952 1254
rect 1824 946 1830 1126
rect 1946 946 1952 1126
rect 1824 864 1952 946
rect 1824 852 1940 864
tri 1940 852 1952 864 nw
tri 2118 852 2143 877 se
rect 2143 852 2195 1789
rect 1824 0 1918 852
tri 1918 830 1940 852 nw
rect 2067 800 2073 852
rect 2125 800 2137 852
rect 2189 800 2195 852
rect 2223 1217 2406 2350
rect 2223 1165 2229 1217
rect 2281 1165 2293 1217
rect 2345 1165 2406 1217
rect 2223 772 2406 1165
rect 2223 720 2263 772
rect 2315 720 2327 772
rect 2379 720 2406 772
rect 2067 401 2073 453
rect 2125 401 2137 453
rect 2189 401 2195 453
tri 2118 376 2143 401 ne
rect 1980 81 1986 133
rect 2038 81 2050 133
rect 2102 81 2108 133
tri 2031 56 2056 81 ne
rect 2056 0 2108 81
rect 2143 0 2195 401
rect 2223 0 2406 720
rect 2462 2077 2730 2350
rect 2762 2109 3078 2350
tri 2762 2085 2786 2109 ne
rect 2462 1126 2530 2077
tri 2530 2051 2556 2077 nw
tri 2612 2051 2638 2077 ne
rect 2462 1074 2470 1126
rect 2522 1074 2530 1126
rect 2462 1062 2530 1074
rect 2462 1010 2470 1062
rect 2522 1010 2530 1062
rect 2462 998 2530 1010
rect 2462 946 2470 998
rect 2522 946 2530 998
rect 2462 0 2530 946
rect 2558 2033 2610 2039
rect 2558 1969 2610 1981
rect 2558 1905 2610 1917
rect 2558 1841 2610 1853
rect 2558 0 2610 1789
rect 2638 1126 2730 2077
rect 2638 1074 2658 1126
rect 2710 1074 2730 1126
rect 2638 1062 2730 1074
rect 2638 1010 2658 1062
rect 2710 1010 2730 1062
rect 2638 998 2730 1010
rect 2638 946 2658 998
rect 2710 946 2730 998
rect 2638 0 2730 946
rect 2786 479 3054 2109
tri 3054 2085 3078 2109 nw
rect 3110 946 3343 2350
rect 3386 2016 3438 2350
rect 3386 1952 3438 1964
rect 3386 1888 3438 1900
rect 3386 1824 3438 1836
rect 3386 1760 3438 1772
rect 2786 0 2963 479
tri 2963 388 3054 479 nw
rect 3151 241 3157 293
rect 3209 241 3221 293
rect 3273 241 3279 293
tri 3202 216 3227 241 ne
rect 3071 152 3077 204
rect 3129 152 3141 204
rect 3193 152 3199 204
tri 3089 127 3114 152 ne
rect 3114 0 3166 152
tri 3166 127 3191 152 nw
rect 3227 0 3279 241
rect 3386 0 3438 1708
rect 3466 1126 3642 2350
rect 3466 946 3500 1126
rect 3616 946 3642 1126
rect 3466 772 3642 946
rect 3466 720 3495 772
rect 3547 720 3559 772
rect 3611 720 3642 772
rect 3466 0 3642 720
rect 3698 0 3750 2350
rect 3778 2016 3830 2022
rect 3778 1952 3830 1964
rect 3778 1888 3830 1900
rect 3778 1824 3830 1836
rect 3778 1760 3830 1772
rect 3778 681 3830 1708
rect 3778 617 3830 629
rect 3778 0 3830 565
rect 3858 1126 4026 2350
rect 3858 946 3891 1126
rect 4007 946 4026 1126
rect 3858 772 4026 946
rect 3858 720 3879 772
rect 3931 720 3943 772
rect 3995 720 4026 772
rect 3858 0 4026 720
rect 4082 2016 4134 2350
rect 4082 1952 4134 1964
rect 4082 1888 4134 1900
rect 4082 1824 4134 1836
rect 4082 1760 4134 1772
rect 4082 285 4134 1708
rect 4175 353 4398 2350
tri 4175 314 4214 353 ne
tri 4082 233 4134 285 ne
tri 4134 255 4186 307 sw
rect 4134 0 4186 255
rect 4214 0 4398 353
rect 4454 1216 4676 2350
rect 4454 1164 4475 1216
rect 4527 1164 4539 1216
rect 4591 1164 4603 1216
rect 4655 1164 4676 1216
rect 4454 1146 4676 1164
rect 4454 1094 4475 1146
rect 4527 1094 4539 1146
rect 4591 1094 4603 1146
rect 4655 1094 4676 1146
rect 4454 1075 4676 1094
rect 4454 1023 4475 1075
rect 4527 1023 4539 1075
rect 4591 1023 4603 1075
rect 4655 1023 4676 1075
rect 4454 1004 4676 1023
rect 4454 952 4475 1004
rect 4527 952 4539 1004
rect 4591 952 4603 1004
rect 4655 952 4676 1004
rect 4454 0 4676 952
rect 4732 0 5043 2350
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_0
timestamp 1704896540
transform -1 0 3129 0 1 1256
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_1
timestamp 1704896540
transform -1 0 2571 0 1 1256
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_2
timestamp 1704896540
transform -1 0 2953 0 1 1256
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_3
timestamp 1704896540
transform -1 0 3401 0 1 1256
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_4
timestamp 1704896540
transform -1 0 1811 0 1 1256
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_5
timestamp 1704896540
transform -1 0 2213 0 1 1256
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_6
timestamp 1704896540
transform 1 0 4643 0 1 1256
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_7
timestamp 1704896540
transform 1 0 4261 0 1 1256
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_8
timestamp 1704896540
transform 1 0 135 0 1 1332
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_9
timestamp 1704896540
transform 1 0 4085 0 1 1256
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_10
timestamp 1704896540
transform 1 0 1587 0 1 1332
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_11
timestamp 1704896540
transform 1 0 3271 0 1 1332
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_12
timestamp 1704896540
transform 1 0 773 0 1 1332
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_13
timestamp 1704896540
transform 1 0 231 0 1 1256
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_14
timestamp 1704896540
transform 1 0 3535 0 1 1256
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_15
timestamp 1704896540
transform 1 0 3799 0 1 1256
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_16
timestamp 1704896540
transform 1 0 3711 0 1 806
box 0 0 1 1
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_17
timestamp 1704896540
transform 1 0 3909 0 1 1332
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1704896540
transform -1 0 3077 0 -1 367
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1704896540
transform -1 0 3253 0 -1 447
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_2
timestamp 1704896540
transform -1 0 579 0 -1 607
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_3
timestamp 1704896540
transform 0 1 4839 1 0 1104
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_4
timestamp 1704896540
transform 0 -1 53 1 0 800
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_5
timestamp 1704896540
transform 1 0 3961 0 -1 127
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_6
timestamp 1704896540
transform 1 0 1287 0 -1 607
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_7
timestamp 1704896540
transform 1 0 2685 0 -1 607
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_8
timestamp 1704896540
transform 1 0 1001 0 -1 367
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_9
timestamp 1704896540
transform 1 0 2319 0 -1 287
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_10
timestamp 1704896540
transform 1 0 4423 0 -1 525
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_11
timestamp 1704896540
transform 1 0 825 0 -1 127
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_12
timestamp 1704896540
transform 1 0 4137 0 -1 445
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_13
timestamp 1704896540
transform 1 0 1653 0 -1 447
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_14
timestamp 1704896540
transform 1 0 1829 0 -1 447
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_15
timestamp 1704896540
transform 1 0 63 0 1 1182
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_16
timestamp 1704896540
transform 1 0 1144 0 1 732
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_17
timestamp 1704896540
transform 1 0 2500 0 1 732
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_18
timestamp 1704896540
transform 1 0 2831 0 1 732
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_19
timestamp 1704896540
transform 1 0 4283 0 1 732
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_0
timestamp 1704896540
transform 0 -1 53 1 0 958
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_1
timestamp 1704896540
transform 1 0 4572 0 -1 766
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_2
timestamp 1704896540
transform 1 0 1433 0 -1 766
box 0 0 1 1
use L1M1_CDNS_5246887918590  L1M1_CDNS_5246887918590_3
timestamp 1704896540
transform 1 0 613 0 -1 766
box 0 0 1 1
use L1M1_CDNS_52468879185193  L1M1_CDNS_52468879185193_0
timestamp 1704896540
transform 1 0 105 0 1 732
box 0 0 1 1
use L1M1_CDNS_52468879185196  L1M1_CDNS_52468879185196_0
timestamp 1704896540
transform -1 0 2247 0 -1 766
box 0 0 1 1
use L1M1_CDNS_52468879185316  L1M1_CDNS_52468879185316_0
timestamp 1704896540
transform 1 0 3307 0 -1 766
box -12 -6 622 40
use L1M1_CDNS_52468879185326  L1M1_CDNS_52468879185326_0
timestamp 1704896540
transform 0 1 19 1 0 1425
box -12 -6 694 40
use L1M1_CDNS_52468879185326  L1M1_CDNS_52468879185326_1
timestamp 1704896540
transform 0 -1 4872 1 0 1425
box -12 -6 694 40
use L1M1_CDNS_52468879185946  L1M1_CDNS_52468879185946_0
timestamp 1704896540
transform 1 0 691 0 1 2208
box -12 -6 4150 40
use L1M1_CDNS_524688791851057  L1M1_CDNS_524688791851057_0
timestamp 1704896540
transform 1 0 1411 0 1 1789
box 0 0 1 1
use L1M1_CDNS_524688791851057  L1M1_CDNS_524688791851057_1
timestamp 1704896540
transform 1 0 2633 0 1 1789
box 0 0 1 1
use L1M1_CDNS_524688791851072  L1M1_CDNS_524688791851072_0
timestamp 1704896540
transform 1 0 3447 0 -1 2036
box 0 0 1 1
use L1M1_CDNS_524688791851072  L1M1_CDNS_524688791851072_1
timestamp 1704896540
transform 1 0 949 0 1 1708
box 0 0 1 1
use L1M1_CDNS_524688791851072  L1M1_CDNS_524688791851072_2
timestamp 1704896540
transform 1 0 1500 0 1 1708
box 0 0 1 1
use L1M1_CDNS_524688791851072  L1M1_CDNS_524688791851072_3
timestamp 1704896540
transform 1 0 3799 0 1 1708
box 0 0 1 1
use L1M1_CDNS_524688791851072  L1M1_CDNS_524688791851072_4
timestamp 1704896540
transform 1 0 4547 0 1 1708
box 0 0 1 1
use L1M1_CDNS_524688791851072  L1M1_CDNS_524688791851072_5
timestamp 1704896540
transform 1 0 597 0 1 1708
box 0 0 1 1
use L1M1_CDNS_524688791851072  L1M1_CDNS_524688791851072_6
timestamp 1704896540
transform 1 0 311 0 1 1708
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1704896540
transform 0 -1 3830 -1 0 687
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_1
timestamp 1704896540
transform -1 0 1364 0 -1 213
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_2
timestamp 1704896540
transform 1 0 1980 0 1 81
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_3
timestamp 1704896540
transform 1 0 3151 0 1 241
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_4
timestamp 1704896540
transform 1 0 2067 0 1 401
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_5
timestamp 1704896540
transform 1 0 3071 0 1 152
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_6
timestamp 1704896540
transform 1 0 -128 0 1 1176
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_7
timestamp 1704896540
transform 1 0 2067 0 1 800
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_0
timestamp 1704896540
transform 0 1 1167 1 0 946
box 0 0 1 1
use M1M2_CDNS_52468879185200  M1M2_CDNS_52468879185200_0
timestamp 1704896540
transform -1 0 4013 0 1 946
box 0 0 1 1
use M1M2_CDNS_52468879185200  M1M2_CDNS_52468879185200_1
timestamp 1704896540
transform 1 0 1824 0 1 946
box 0 0 1 1
use M1M2_CDNS_52468879185200  M1M2_CDNS_52468879185200_2
timestamp 1704896540
transform 1 0 3494 0 1 946
box 0 0 1 1
use M1M2_CDNS_52468879185200  M1M2_CDNS_52468879185200_3
timestamp 1704896540
transform 1 0 -128 0 1 720
box 0 0 1 1
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_0
timestamp 1704896540
transform 0 -1 490 -1 0 2022
box 0 0 1 1
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_1
timestamp 1704896540
transform 0 -1 3830 1 0 1702
box 0 0 1 1
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_2
timestamp 1704896540
transform 0 -1 3438 1 0 1702
box 0 0 1 1
use M1M2_CDNS_52468879185202  M1M2_CDNS_52468879185202_3
timestamp 1704896540
transform 0 -1 4134 1 0 1702
box 0 0 1 1
use M1M2_CDNS_52468879185297  M1M2_CDNS_52468879185297_0
timestamp 1704896540
transform 0 1 1744 1 0 1860
box 0 0 1 1
use M1M2_CDNS_52468879185297  M1M2_CDNS_52468879185297_1
timestamp 1704896540
transform 0 -1 1444 1 0 1783
box 0 0 1 1
use M1M2_CDNS_52468879185297  M1M2_CDNS_52468879185297_2
timestamp 1704896540
transform 0 -1 2610 1 0 1783
box 0 0 1 1
use M1M2_CDNS_52468879185297  M1M2_CDNS_52468879185297_3
timestamp 1704896540
transform 0 -1 2195 1 0 1783
box 0 0 1 1
use M1M2_CDNS_52468879185371  M1M2_CDNS_52468879185371_0
timestamp 1704896540
transform 1 0 2464 0 1 946
box 0 0 1 1
use M1M2_CDNS_52468879185371  M1M2_CDNS_52468879185371_1
timestamp 1704896540
transform 1 0 2652 0 1 946
box 0 0 1 1
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_0
timestamp 1704896540
transform 0 1 2224 1 0 946
box 0 0 192 180
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_1
timestamp 1704896540
transform 1 0 4468 0 1 720
box 0 0 192 180
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_2
timestamp 1704896540
transform 1 0 524 0 1 946
box 0 0 192 180
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_3
timestamp 1704896540
transform 1 0 1507 0 1 946
box 0 0 192 180
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_4
timestamp 1704896540
transform 1 0 3133 0 1 946
box 0 0 192 180
use M1M2_CDNS_524688791851081  M1M2_CDNS_524688791851081_0
timestamp 1704896540
transform 1 0 848 0 1 946
box 0 0 256 180
use M1M2_CDNS_524688791851144  M1M2_CDNS_524688791851144_0
timestamp 1704896540
transform 1 0 67 0 1 946
box 0 0 384 180
use M1M2_CDNS_524688791851145  M1M2_CDNS_524688791851145_0
timestamp 1704896540
transform 1 0 4733 0 1 1398
box 0 0 128 820
use sky130_fd_io__refgen_inv_x1  sky130_fd_io__refgen_inv_x1_0
timestamp 1704896540
transform 1 0 152 0 1 805
box -107 21 267 1369
use sky130_fd_io__refgen_inv_x1  sky130_fd_io__refgen_inv_x1_1
timestamp 1704896540
transform 1 0 3640 0 1 805
box -107 21 267 1369
use sky130_fd_io__refgen_inv_x2  sky130_fd_io__refgen_inv_x2_0
timestamp 1704896540
transform 1 0 3288 0 1 805
box -107 21 459 1369
use sky130_fd_io__refgen_nand2  sky130_fd_io__refgen_nand2_0
timestamp 1704896540
transform -1 0 790 0 1 805
box -107 21 459 1369
use sky130_fd_io__refgen_nand2  sky130_fd_io__refgen_nand2_1
timestamp 1704896540
transform -1 0 1604 0 1 805
box -107 21 459 1369
use sky130_fd_io__refgen_nand2  sky130_fd_io__refgen_nand2_2
timestamp 1704896540
transform -1 0 4740 0 1 805
box -107 21 459 1369
use sky130_fd_io__refgen_nand2  sky130_fd_io__refgen_nand2_3
timestamp 1704896540
transform -1 0 3288 0 1 805
box -107 21 459 1369
use sky130_fd_io__refgen_nand2  sky130_fd_io__refgen_nand2_4
timestamp 1704896540
transform 1 0 3926 0 1 805
box -107 21 459 1369
use sky130_fd_io__refgen_nand2  sky130_fd_io__refgen_nand2_5
timestamp 1704896540
transform 1 0 790 0 1 805
box -107 21 459 1369
use sky130_fd_io__refgen_nand2  sky130_fd_io__refgen_nand2_6
timestamp 1704896540
transform 1 0 2474 0 1 805
box -107 21 459 1369
use sky130_fd_io__refgen_nor  sky130_fd_io__refgen_nor_0
timestamp 1704896540
transform -1 0 2474 0 1 805
box -107 21 487 1369
use sky130_fd_io__refgen_nor  sky130_fd_io__refgen_nor_1
timestamp 1704896540
transform 1 0 1604 0 1 805
box -107 21 487 1369
<< labels >>
flabel comment s 3013 87 3013 87 3 FreeSans 200 90 0 0 vreg_en_h_n
flabel comment s 3724 87 3724 87 3 FreeSans 200 90 0 0 vohref_0p5
flabel comment s 3138 81 3138 81 3 FreeSans 200 90 0 0 biasen_n
flabel comment s 2873 87 2873 87 3 FreeSans 200 90 0 0 vpb
flabel comment s 3722 2322 3722 2322 3 FreeSans 200 270 0 0 vohref_0p5
flabel comment s 2917 2332 2917 2332 3 FreeSans 200 270 0 0 vpb
flabel comment s 4284 30 4284 30 3 FreeSans 200 90 0 0 vpwr_ka
flabel comment s 4284 2322 4284 2322 3 FreeSans 200 270 0 0 vpwr_ka
flabel comment s 4110 2322 4110 2322 3 FreeSans 200 270 0 0 sel_vohref_0p5
flabel comment s 1407 2322 1407 2322 3 FreeSans 200 270 0 0 biasen_n
flabel metal1 s 0 197 32 249 3 FreeSans 200 0 0 0 ibuf_sel_h_n
port 2 nsew
flabel metal1 s 0 559 38 607 3 FreeSans 200 0 0 0 en_outop_h
port 3 nsew
flabel metal1 s -1 2202 35 2350 3 FreeSans 200 0 0 0 vcc_io
port 4 nsew
flabel metal1 s 0 357 34 409 3 FreeSans 200 0 0 0 ibuf_sel_h
port 5 nsew
flabel metal1 s 0 1398 36 1674 3 FreeSans 200 0 0 0 vcc_io
port 4 nsew
flabel metal1 s 0 277 34 329 3 FreeSans 200 0 0 0 vtrip_sel_h_n
port 6 nsew
flabel metal1 s 0 123 34 169 3 FreeSans 200 0 0 0 vtrip_sel_h
port 7 nsew
flabel metal1 s 780 946 792 1148 0 FreeSans 200 0 0 0 vgnd_io
port 8 nsew
flabel metal1 s 780 1398 792 1674 0 FreeSans 200 0 0 0 vcc_io
port 4 nsew
flabel metal2 s 3778 0 3830 41 3 FreeSans 200 90 0 0 en_outop_h
port 3 nsew
flabel metal2 s 438 2309 490 2350 3 FreeSans 200 270 0 0 en_inpop_h
port 9 nsew
flabel metal2 s 3227 0 3279 27 3 FreeSans 200 90 0 0 vreg_en_h
port 10 nsew
flabel metal2 s 3386 2309 3438 2350 3 FreeSans 200 270 0 0 en_outop_h_n
port 11 nsew
flabel metal2 s 4732 2309 4878 2350 3 FreeSans 200 270 0 0 vcc_io
port 4 nsew
flabel metal2 s 4732 0 4878 41 3 FreeSans 200 90 0 0 vcc_io
port 4 nsew
flabel metal2 s 4454 2309 4676 2350 3 FreeSans 200 270 0 0 vgnd_io
port 8 nsew
flabel metal2 s 3858 2309 4026 2350 3 FreeSans 200 270 0 0 vgnd_io
port 8 nsew
flabel metal2 s 3466 2309 3642 2350 3 FreeSans 200 270 0 0 vgnd_io
port 8 nsew
flabel metal2 s 2462 2309 2730 2350 3 FreeSans 200 270 0 0 vgnd_io
port 8 nsew
flabel metal2 s 2223 2309 2406 2350 3 FreeSans 200 270 0 0 vgnd_io
port 8 nsew
flabel metal2 s 1824 0 1918 41 3 FreeSans 200 90 0 0 vgnd_io
port 8 nsew
flabel metal2 s 1490 2309 1758 2350 3 FreeSans 200 270 0 0 vgnd_io
port 8 nsew
flabel metal2 s 842 2309 1110 2350 3 FreeSans 200 270 0 0 vgnd_io
port 8 nsew
flabel metal2 s 518 2309 786 2350 3 FreeSans 200 270 0 0 vgnd_io
port 8 nsew
flabel metal2 s 56 2309 410 2350 3 FreeSans 200 270 0 0 vgnd_io
port 8 nsew
flabel metal2 s 3858 0 4026 41 3 FreeSans 200 90 0 0 vgnd_io
port 8 nsew
flabel metal2 s 3466 0 3642 41 3 FreeSans 200 90 0 0 vgnd_io
port 8 nsew
flabel metal2 s 2638 0 2730 41 3 FreeSans 200 90 0 0 vgnd_io
port 8 nsew
flabel metal2 s 2462 0 2530 41 3 FreeSans 200 90 0 0 vgnd_io
port 8 nsew
flabel metal2 s 2223 0 2406 41 3 FreeSans 200 90 0 0 vgnd_io
port 8 nsew
flabel metal2 s 1814 2309 1918 2350 3 FreeSans 200 270 0 0 vgnd_io
port 8 nsew
flabel metal2 s 1490 0 1716 41 3 FreeSans 200 90 0 0 vgnd_io
port 8 nsew
flabel metal2 s 842 0 1110 41 3 FreeSans 200 90 0 0 vgnd_io
port 8 nsew
flabel metal2 s 518 0 786 41 3 FreeSans 200 90 0 0 vgnd_io
port 8 nsew
flabel metal2 s 56 0 372 41 3 FreeSans 200 90 0 0 vgnd_io
port 8 nsew
flabel metal2 s 1166 2309 1311 2350 3 FreeSans 200 270 0 0 vgnd_io
port 8 nsew
flabel metal2 s 3110 2309 3343 2350 3 FreeSans 200 270 0 0 vgnd_io
port 8 nsew
flabel metal2 s 4454 0 4676 41 3 FreeSans 200 90 0 0 vgnd_io
port 8 nsew
flabel metal2 s 3386 0 3438 41 3 FreeSans 200 90 0 0 en_outop_h_n
port 11 nsew
flabel metal2 s 2143 0 2195 34 3 FreeSans 200 90 0 0 vref_sel_h_n
port 12 nsew
flabel metal2 s 2056 0 2108 34 3 FreeSans 200 90 0 0 vref_sel_h
port 13 nsew
flabel metal2 s 4134 0 4186 30 3 FreeSans 200 90 0 0 sel_vohref_0p5
port 14 nsew
flabel metal2 s 1392 0 1444 30 3 FreeSans 200 90 0 0 sel_vohref
port 15 nsew
flabel metal2 s 2558 0 2610 30 3 FreeSans 200 90 0 0 sel_vcc_io_0p4
port 16 nsew
flabel metal2 s 1744 0 1796 30 3 FreeSans 200 90 0 0 sel_vcc_io
port 17 nsew
<< properties >>
string GDS_END 79876392
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 79840566
string path 96.825 18.650 100.475 18.650 
<< end >>
