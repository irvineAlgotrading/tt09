magic
tech sky130B
timestamp 1704896540
<< metal1 >>
rect 0 0 3 250
rect 861 0 864 250
<< via1 >>
rect 3 0 861 250
<< metal2 >>
rect 0 0 3 250
rect 861 0 864 250
<< properties >>
string GDS_END 94917242
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 94903286
<< end >>
