magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< pwell >>
rect -76 -26 9140 2026
<< mvnnmos >>
rect 0 0 400 2000
rect 456 0 856 2000
rect 912 0 1312 2000
rect 1368 0 1768 2000
rect 1824 0 2224 2000
rect 2280 0 2680 2000
rect 2736 0 3136 2000
rect 3192 0 3592 2000
rect 3648 0 4048 2000
rect 4104 0 4504 2000
rect 4560 0 4960 2000
rect 5016 0 5416 2000
rect 5472 0 5872 2000
rect 5928 0 6328 2000
rect 6384 0 6784 2000
rect 6840 0 7240 2000
rect 7296 0 7696 2000
rect 7752 0 8152 2000
rect 8208 0 8608 2000
rect 8664 0 9064 2000
<< mvndiff >>
rect -50 0 0 2000
rect 9064 0 9114 2000
<< poly >>
rect 0 2000 400 2032
rect 0 -32 400 0
rect 456 2000 856 2032
rect 456 -32 856 0
rect 912 2000 1312 2032
rect 912 -32 1312 0
rect 1368 2000 1768 2032
rect 1368 -32 1768 0
rect 1824 2000 2224 2032
rect 1824 -32 2224 0
rect 2280 2000 2680 2032
rect 2280 -32 2680 0
rect 2736 2000 3136 2032
rect 2736 -32 3136 0
rect 3192 2000 3592 2032
rect 3192 -32 3592 0
rect 3648 2000 4048 2032
rect 3648 -32 4048 0
rect 4104 2000 4504 2032
rect 4104 -32 4504 0
rect 4560 2000 4960 2032
rect 4560 -32 4960 0
rect 5016 2000 5416 2032
rect 5016 -32 5416 0
rect 5472 2000 5872 2032
rect 5472 -32 5872 0
rect 5928 2000 6328 2032
rect 5928 -32 6328 0
rect 6384 2000 6784 2032
rect 6384 -32 6784 0
rect 6840 2000 7240 2032
rect 6840 -32 7240 0
rect 7296 2000 7696 2032
rect 7296 -32 7696 0
rect 7752 2000 8152 2032
rect 7752 -32 8152 0
rect 8208 2000 8608 2032
rect 8208 -32 8608 0
rect 8664 2000 9064 2032
rect 8664 -32 9064 0
<< metal1 >>
rect -51 -16 -5 1986
rect 405 -16 451 1986
rect 861 -16 907 1986
rect 1317 -16 1363 1986
rect 1773 -16 1819 1986
rect 2229 -16 2275 1986
rect 2685 -16 2731 1986
rect 3141 -16 3187 1986
rect 3597 -16 3643 1986
rect 4053 -16 4099 1986
rect 4509 -16 4555 1986
rect 4965 -16 5011 1986
rect 5421 -16 5467 1986
rect 5877 -16 5923 1986
rect 6333 -16 6379 1986
rect 6789 -16 6835 1986
rect 7245 -16 7291 1986
rect 7701 -16 7747 1986
rect 8157 -16 8203 1986
rect 8613 -16 8659 1986
rect 9069 -16 9115 1986
use hvDFM1sd2_CDNS_5246887918552  hvDFM1sd2_CDNS_5246887918552_0
timestamp 1704896540
transform -1 0 0 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5246887918552  hvDFM1sd2_CDNS_5246887918552_1
timestamp 1704896540
transform 1 0 9064 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5246887918552  hvDFM1sd2_CDNS_5246887918552_2
timestamp 1704896540
transform 1 0 8608 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5246887918552  hvDFM1sd2_CDNS_5246887918552_3
timestamp 1704896540
transform 1 0 8152 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5246887918552  hvDFM1sd2_CDNS_5246887918552_4
timestamp 1704896540
transform 1 0 7696 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5246887918552  hvDFM1sd2_CDNS_5246887918552_5
timestamp 1704896540
transform 1 0 7240 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5246887918552  hvDFM1sd2_CDNS_5246887918552_6
timestamp 1704896540
transform 1 0 6784 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5246887918552  hvDFM1sd2_CDNS_5246887918552_7
timestamp 1704896540
transform 1 0 6328 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5246887918552  hvDFM1sd2_CDNS_5246887918552_8
timestamp 1704896540
transform 1 0 5872 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5246887918552  hvDFM1sd2_CDNS_5246887918552_9
timestamp 1704896540
transform 1 0 5416 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5246887918552  hvDFM1sd2_CDNS_5246887918552_10
timestamp 1704896540
transform 1 0 4960 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5246887918552  hvDFM1sd2_CDNS_5246887918552_11
timestamp 1704896540
transform 1 0 4504 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5246887918552  hvDFM1sd2_CDNS_5246887918552_12
timestamp 1704896540
transform 1 0 4048 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5246887918552  hvDFM1sd2_CDNS_5246887918552_13
timestamp 1704896540
transform 1 0 3592 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5246887918552  hvDFM1sd2_CDNS_5246887918552_14
timestamp 1704896540
transform 1 0 3136 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5246887918552  hvDFM1sd2_CDNS_5246887918552_15
timestamp 1704896540
transform 1 0 2680 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5246887918552  hvDFM1sd2_CDNS_5246887918552_16
timestamp 1704896540
transform 1 0 2224 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5246887918552  hvDFM1sd2_CDNS_5246887918552_17
timestamp 1704896540
transform 1 0 1768 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5246887918552  hvDFM1sd2_CDNS_5246887918552_18
timestamp 1704896540
transform 1 0 1312 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5246887918552  hvDFM1sd2_CDNS_5246887918552_19
timestamp 1704896540
transform 1 0 856 0 1 0
box -26 -26 82 2026
use hvDFM1sd2_CDNS_5246887918552  hvDFM1sd2_CDNS_5246887918552_20
timestamp 1704896540
transform 1 0 400 0 1 0
box -26 -26 82 2026
<< labels >>
flabel comment s -28 985 -28 985 0 FreeSans 300 0 0 0 S
flabel comment s 428 985 428 985 0 FreeSans 300 0 0 0 D
flabel comment s 884 985 884 985 0 FreeSans 300 0 0 0 S
flabel comment s 1340 985 1340 985 0 FreeSans 300 0 0 0 D
flabel comment s 1796 985 1796 985 0 FreeSans 300 0 0 0 S
flabel comment s 2252 985 2252 985 0 FreeSans 300 0 0 0 D
flabel comment s 2708 985 2708 985 0 FreeSans 300 0 0 0 S
flabel comment s 3164 985 3164 985 0 FreeSans 300 0 0 0 D
flabel comment s 3620 985 3620 985 0 FreeSans 300 0 0 0 S
flabel comment s 4076 985 4076 985 0 FreeSans 300 0 0 0 D
flabel comment s 4532 985 4532 985 0 FreeSans 300 0 0 0 S
flabel comment s 4988 985 4988 985 0 FreeSans 300 0 0 0 D
flabel comment s 5444 985 5444 985 0 FreeSans 300 0 0 0 S
flabel comment s 5900 985 5900 985 0 FreeSans 300 0 0 0 D
flabel comment s 6356 985 6356 985 0 FreeSans 300 0 0 0 S
flabel comment s 6812 985 6812 985 0 FreeSans 300 0 0 0 D
flabel comment s 7268 985 7268 985 0 FreeSans 300 0 0 0 S
flabel comment s 7724 985 7724 985 0 FreeSans 300 0 0 0 D
flabel comment s 8180 985 8180 985 0 FreeSans 300 0 0 0 S
flabel comment s 8636 985 8636 985 0 FreeSans 300 0 0 0 D
flabel comment s 9092 985 9092 985 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 6101782
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 6091366
<< end >>
