magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< pwell >>
rect -76 -26 179 326
<< mvnmos >>
rect 0 0 100 300
<< mvndiff >>
rect -50 0 0 300
rect 100 250 153 300
rect 100 216 111 250
rect 145 216 153 250
rect 100 182 153 216
rect 100 148 111 182
rect 145 148 153 182
rect 100 114 153 148
rect 100 80 111 114
rect 145 80 153 114
rect 100 46 153 80
rect 100 12 111 46
rect 145 12 153 46
rect 100 0 153 12
<< mvndiffc >>
rect 111 216 145 250
rect 111 148 145 182
rect 111 80 145 114
rect 111 12 145 46
<< poly >>
rect 0 300 100 326
rect 0 -26 100 0
<< locali >>
rect 111 250 145 266
rect 111 182 145 216
rect 111 114 145 148
rect 111 46 145 80
rect 111 -4 145 12
use hvDFL1sd_CDNS_52468879185376  hvDFL1sd_CDNS_52468879185376_0
timestamp 1704896540
transform 1 0 100 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s -25 150 -25 150 0 FreeSans 300 0 0 0 S
flabel comment s 128 131 128 131 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 87761148
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 87760392
<< end >>
