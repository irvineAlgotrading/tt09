magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< pwell >>
rect 894 821 918 872
<< poly >>
rect 0 1552 1716 1568
rect 0 1518 97 1552
rect 131 1518 165 1552
rect 199 1518 233 1552
rect 267 1518 301 1552
rect 335 1518 369 1552
rect 403 1518 437 1552
rect 471 1518 505 1552
rect 539 1518 573 1552
rect 607 1518 641 1552
rect 675 1518 709 1552
rect 743 1518 777 1552
rect 811 1518 897 1552
rect 931 1518 965 1552
rect 999 1518 1033 1552
rect 1067 1518 1101 1552
rect 1135 1518 1169 1552
rect 1203 1518 1237 1552
rect 1271 1518 1305 1552
rect 1339 1518 1373 1552
rect 1407 1518 1441 1552
rect 1475 1518 1509 1552
rect 1543 1518 1577 1552
rect 1611 1518 1716 1552
rect 0 1481 1716 1518
rect 0 1447 16 1481
rect 50 1447 1666 1481
rect 1700 1447 1716 1481
rect 0 1413 1716 1447
rect 0 1379 16 1413
rect 50 1379 1666 1413
rect 1700 1379 1716 1413
rect 0 1345 1716 1379
rect 0 1311 16 1345
rect 50 1311 1666 1345
rect 1700 1311 1716 1345
rect 0 1277 1716 1311
rect 0 1243 16 1277
rect 50 1243 1666 1277
rect 1700 1243 1716 1277
rect 0 1209 1716 1243
rect 0 1175 16 1209
rect 50 1175 1666 1209
rect 1700 1175 1716 1209
rect 0 1141 1716 1175
rect 0 1107 16 1141
rect 50 1107 1666 1141
rect 1700 1107 1716 1141
rect 0 1073 1716 1107
rect 0 1039 16 1073
rect 50 1039 1666 1073
rect 1700 1039 1716 1073
rect 0 1005 1716 1039
rect 0 971 16 1005
rect 50 971 1666 1005
rect 1700 971 1716 1005
rect 0 937 1716 971
rect 0 903 16 937
rect 50 903 1666 937
rect 1700 903 1716 937
rect 0 869 1716 903
rect 0 835 16 869
rect 50 835 1666 869
rect 1700 835 1716 869
rect 0 801 1716 835
rect 0 767 16 801
rect 50 767 1666 801
rect 1700 767 1716 801
rect 0 733 1716 767
rect 0 699 16 733
rect 50 699 1666 733
rect 1700 699 1716 733
rect 0 665 1716 699
rect 0 631 16 665
rect 50 631 1666 665
rect 1700 631 1716 665
rect 0 597 1716 631
rect 0 563 16 597
rect 50 563 1666 597
rect 1700 563 1716 597
rect 0 529 1716 563
rect 0 495 16 529
rect 50 495 1666 529
rect 1700 495 1716 529
rect 0 461 1716 495
rect 0 427 16 461
rect 50 427 1666 461
rect 1700 427 1716 461
rect 0 393 1716 427
rect 0 359 16 393
rect 50 359 1666 393
rect 1700 359 1716 393
rect 0 325 1716 359
rect 0 291 16 325
rect 50 291 1666 325
rect 1700 291 1716 325
rect 0 257 1716 291
rect 0 223 16 257
rect 50 223 1666 257
rect 1700 223 1716 257
rect 0 189 1716 223
rect 0 155 16 189
rect 50 155 1666 189
rect 1700 155 1716 189
rect 0 121 1716 155
rect 0 87 16 121
rect 50 87 1666 121
rect 1700 87 1716 121
rect 0 50 1716 87
rect 0 16 97 50
rect 131 16 165 50
rect 199 16 233 50
rect 267 16 301 50
rect 335 16 369 50
rect 403 16 437 50
rect 471 16 505 50
rect 539 16 573 50
rect 607 16 641 50
rect 675 16 709 50
rect 743 16 777 50
rect 811 16 897 50
rect 931 16 965 50
rect 999 16 1033 50
rect 1067 16 1101 50
rect 1135 16 1169 50
rect 1203 16 1237 50
rect 1271 16 1305 50
rect 1339 16 1373 50
rect 1407 16 1441 50
rect 1475 16 1509 50
rect 1543 16 1577 50
rect 1611 16 1716 50
rect 0 0 1716 16
<< polycont >>
rect 97 1518 131 1552
rect 165 1518 199 1552
rect 233 1518 267 1552
rect 301 1518 335 1552
rect 369 1518 403 1552
rect 437 1518 471 1552
rect 505 1518 539 1552
rect 573 1518 607 1552
rect 641 1518 675 1552
rect 709 1518 743 1552
rect 777 1518 811 1552
rect 897 1518 931 1552
rect 965 1518 999 1552
rect 1033 1518 1067 1552
rect 1101 1518 1135 1552
rect 1169 1518 1203 1552
rect 1237 1518 1271 1552
rect 1305 1518 1339 1552
rect 1373 1518 1407 1552
rect 1441 1518 1475 1552
rect 1509 1518 1543 1552
rect 1577 1518 1611 1552
rect 16 1447 50 1481
rect 1666 1447 1700 1481
rect 16 1379 50 1413
rect 1666 1379 1700 1413
rect 16 1311 50 1345
rect 1666 1311 1700 1345
rect 16 1243 50 1277
rect 1666 1243 1700 1277
rect 16 1175 50 1209
rect 1666 1175 1700 1209
rect 16 1107 50 1141
rect 1666 1107 1700 1141
rect 16 1039 50 1073
rect 1666 1039 1700 1073
rect 16 971 50 1005
rect 1666 971 1700 1005
rect 16 903 50 937
rect 1666 903 1700 937
rect 16 835 50 869
rect 1666 835 1700 869
rect 16 767 50 801
rect 1666 767 1700 801
rect 16 699 50 733
rect 1666 699 1700 733
rect 16 631 50 665
rect 1666 631 1700 665
rect 16 563 50 597
rect 1666 563 1700 597
rect 16 495 50 529
rect 1666 495 1700 529
rect 16 427 50 461
rect 1666 427 1700 461
rect 16 359 50 393
rect 1666 359 1700 393
rect 16 291 50 325
rect 1666 291 1700 325
rect 16 223 50 257
rect 1666 223 1700 257
rect 16 155 50 189
rect 1666 155 1700 189
rect 16 87 50 121
rect 1666 87 1700 121
rect 97 16 131 50
rect 165 16 199 50
rect 233 16 267 50
rect 301 16 335 50
rect 369 16 403 50
rect 437 16 471 50
rect 505 16 539 50
rect 573 16 607 50
rect 641 16 675 50
rect 709 16 743 50
rect 777 16 811 50
rect 897 16 931 50
rect 965 16 999 50
rect 1033 16 1067 50
rect 1101 16 1135 50
rect 1169 16 1203 50
rect 1237 16 1271 50
rect 1305 16 1339 50
rect 1373 16 1407 50
rect 1441 16 1475 50
rect 1509 16 1543 50
rect 1577 16 1611 50
<< locali >>
rect 0 1552 1716 1568
rect 0 1518 85 1552
rect 131 1518 157 1552
rect 199 1518 229 1552
rect 267 1518 301 1552
rect 335 1518 369 1552
rect 407 1518 437 1552
rect 479 1518 505 1552
rect 551 1518 573 1552
rect 623 1518 641 1552
rect 695 1518 709 1552
rect 767 1518 777 1552
rect 839 1518 877 1552
rect 931 1518 949 1552
rect 999 1518 1021 1552
rect 1067 1518 1093 1552
rect 1135 1518 1165 1552
rect 1203 1518 1237 1552
rect 1271 1518 1305 1552
rect 1343 1518 1373 1552
rect 1415 1518 1441 1552
rect 1487 1518 1509 1552
rect 1559 1518 1577 1552
rect 1631 1518 1716 1552
rect 0 1502 1716 1518
rect 0 1485 66 1502
rect 0 1447 16 1485
rect 50 1447 66 1485
rect 0 1413 66 1447
rect 1650 1485 1716 1502
rect 1650 1447 1666 1485
rect 1700 1447 1716 1485
rect 0 1379 16 1413
rect 50 1379 66 1413
rect 100 1415 1616 1431
rect 100 1397 841 1415
rect 0 1361 66 1379
rect 831 1381 841 1397
rect 875 1397 1616 1415
rect 1650 1413 1716 1447
rect 875 1381 885 1397
rect 0 1345 797 1361
rect 0 1307 16 1345
rect 50 1327 797 1345
rect 831 1343 885 1381
rect 1650 1379 1666 1413
rect 1700 1379 1716 1413
rect 1650 1361 1716 1379
rect 50 1307 66 1327
rect 0 1277 66 1307
rect 831 1309 841 1343
rect 875 1309 885 1343
rect 919 1345 1716 1361
rect 919 1327 1666 1345
rect 831 1291 885 1309
rect 1650 1307 1666 1327
rect 1700 1307 1716 1345
rect 0 1235 16 1277
rect 50 1235 66 1277
rect 100 1271 1616 1291
rect 100 1257 841 1271
rect 0 1221 66 1235
rect 831 1237 841 1257
rect 875 1257 1616 1271
rect 1650 1277 1716 1307
rect 875 1237 885 1257
rect 0 1209 797 1221
rect 0 1163 16 1209
rect 50 1187 797 1209
rect 831 1199 885 1237
rect 1650 1235 1666 1277
rect 1700 1235 1716 1277
rect 1650 1221 1716 1235
rect 50 1163 66 1187
rect 0 1141 66 1163
rect 831 1165 841 1199
rect 875 1165 885 1199
rect 919 1209 1716 1221
rect 919 1187 1666 1209
rect 831 1151 885 1165
rect 1650 1163 1666 1187
rect 1700 1163 1716 1209
rect 0 1091 16 1141
rect 50 1091 66 1141
rect 100 1127 1616 1151
rect 100 1117 841 1127
rect 0 1081 66 1091
rect 831 1093 841 1117
rect 875 1117 1616 1127
rect 1650 1141 1716 1163
rect 875 1093 885 1117
rect 0 1073 797 1081
rect 0 1019 16 1073
rect 50 1047 797 1073
rect 831 1055 885 1093
rect 1650 1091 1666 1141
rect 1700 1091 1716 1141
rect 1650 1081 1716 1091
rect 50 1019 66 1047
rect 0 1005 66 1019
rect 831 1021 841 1055
rect 875 1021 885 1055
rect 919 1073 1716 1081
rect 919 1047 1666 1073
rect 831 1011 885 1021
rect 1650 1019 1666 1047
rect 1700 1019 1716 1073
rect 0 947 16 1005
rect 50 947 66 1005
rect 100 983 1616 1011
rect 100 977 841 983
rect 0 941 66 947
rect 831 949 841 977
rect 875 977 1616 983
rect 1650 1005 1716 1019
rect 875 949 885 977
rect 0 937 797 941
rect 0 875 16 937
rect 50 907 797 937
rect 831 911 885 949
rect 1650 947 1666 1005
rect 1700 947 1716 1005
rect 1650 941 1716 947
rect 50 875 66 907
rect 0 869 66 875
rect 831 877 841 911
rect 875 877 885 911
rect 919 937 1716 941
rect 919 907 1666 937
rect 831 871 885 877
rect 1650 875 1666 907
rect 1700 875 1716 937
rect 0 803 16 869
rect 50 803 66 869
rect 100 837 1616 871
rect 1650 869 1716 875
rect 0 801 66 803
rect 0 767 16 801
rect 50 767 797 801
rect 0 765 66 767
rect 0 699 16 765
rect 50 699 66 765
rect 831 731 885 837
rect 1650 803 1666 869
rect 1700 803 1716 869
rect 1650 801 1716 803
rect 919 767 1666 801
rect 1700 767 1716 801
rect 1650 765 1716 767
rect 0 693 66 699
rect 100 697 1616 731
rect 1650 699 1666 765
rect 1700 699 1716 765
rect 0 631 16 693
rect 50 661 66 693
rect 831 691 885 697
rect 50 631 797 661
rect 0 627 797 631
rect 831 657 841 691
rect 875 657 885 691
rect 1650 693 1716 699
rect 1650 661 1666 693
rect 0 621 66 627
rect 0 563 16 621
rect 50 563 66 621
rect 831 619 885 657
rect 919 631 1666 661
rect 1700 631 1716 693
rect 919 627 1716 631
rect 831 591 841 619
rect 0 549 66 563
rect 100 585 841 591
rect 875 591 885 619
rect 1650 621 1716 627
rect 875 585 1616 591
rect 100 557 1616 585
rect 1650 563 1666 621
rect 1700 563 1716 621
rect 0 495 16 549
rect 50 521 66 549
rect 831 547 885 557
rect 50 495 797 521
rect 0 487 797 495
rect 831 513 841 547
rect 875 513 885 547
rect 1650 549 1716 563
rect 1650 521 1666 549
rect 0 477 66 487
rect 0 427 16 477
rect 50 427 66 477
rect 831 475 885 513
rect 919 495 1666 521
rect 1700 495 1716 549
rect 919 487 1716 495
rect 831 451 841 475
rect 0 405 66 427
rect 100 441 841 451
rect 875 451 885 475
rect 1650 477 1716 487
rect 875 441 1616 451
rect 100 417 1616 441
rect 1650 427 1666 477
rect 1700 427 1716 477
rect 0 359 16 405
rect 50 381 66 405
rect 831 403 885 417
rect 50 359 797 381
rect 0 347 797 359
rect 831 369 841 403
rect 875 369 885 403
rect 1650 405 1716 427
rect 1650 381 1666 405
rect 0 333 66 347
rect 0 291 16 333
rect 50 291 66 333
rect 831 331 885 369
rect 919 359 1666 381
rect 1700 359 1716 405
rect 919 347 1716 359
rect 831 311 841 331
rect 0 261 66 291
rect 100 297 841 311
rect 875 311 885 331
rect 1650 333 1716 347
rect 875 297 1616 311
rect 100 277 1616 297
rect 1650 291 1666 333
rect 1700 291 1716 333
rect 0 223 16 261
rect 50 241 66 261
rect 831 259 885 277
rect 50 223 797 241
rect 0 207 797 223
rect 831 225 841 259
rect 875 225 885 259
rect 1650 261 1716 291
rect 1650 241 1666 261
rect 0 189 66 207
rect 0 155 16 189
rect 50 155 66 189
rect 831 187 885 225
rect 919 223 1666 241
rect 1700 223 1716 261
rect 919 207 1716 223
rect 831 171 841 187
rect 0 121 66 155
rect 100 153 841 171
rect 875 171 885 187
rect 1650 189 1716 207
rect 875 153 1616 171
rect 100 137 1616 153
rect 1650 155 1666 189
rect 1700 155 1716 189
rect 0 83 16 121
rect 50 83 66 121
rect 0 66 66 83
rect 1650 121 1716 155
rect 1650 83 1666 121
rect 1700 83 1716 121
rect 1650 66 1716 83
rect 0 50 1716 66
rect 0 16 85 50
rect 131 16 157 50
rect 199 16 229 50
rect 267 16 301 50
rect 335 16 369 50
rect 407 16 437 50
rect 479 16 505 50
rect 551 16 573 50
rect 623 16 641 50
rect 695 16 709 50
rect 767 16 777 50
rect 839 16 877 50
rect 931 16 949 50
rect 999 16 1021 50
rect 1067 16 1093 50
rect 1135 16 1165 50
rect 1203 16 1237 50
rect 1271 16 1305 50
rect 1343 16 1373 50
rect 1415 16 1441 50
rect 1487 16 1509 50
rect 1559 16 1577 50
rect 1631 16 1716 50
rect 0 0 1716 16
<< viali >>
rect 85 1518 97 1552
rect 97 1518 119 1552
rect 157 1518 165 1552
rect 165 1518 191 1552
rect 229 1518 233 1552
rect 233 1518 263 1552
rect 301 1518 335 1552
rect 373 1518 403 1552
rect 403 1518 407 1552
rect 445 1518 471 1552
rect 471 1518 479 1552
rect 517 1518 539 1552
rect 539 1518 551 1552
rect 589 1518 607 1552
rect 607 1518 623 1552
rect 661 1518 675 1552
rect 675 1518 695 1552
rect 733 1518 743 1552
rect 743 1518 767 1552
rect 805 1518 811 1552
rect 811 1518 839 1552
rect 877 1518 897 1552
rect 897 1518 911 1552
rect 949 1518 965 1552
rect 965 1518 983 1552
rect 1021 1518 1033 1552
rect 1033 1518 1055 1552
rect 1093 1518 1101 1552
rect 1101 1518 1127 1552
rect 1165 1518 1169 1552
rect 1169 1518 1199 1552
rect 1237 1518 1271 1552
rect 1309 1518 1339 1552
rect 1339 1518 1343 1552
rect 1381 1518 1407 1552
rect 1407 1518 1415 1552
rect 1453 1518 1475 1552
rect 1475 1518 1487 1552
rect 1525 1518 1543 1552
rect 1543 1518 1559 1552
rect 1597 1518 1611 1552
rect 1611 1518 1631 1552
rect 16 1481 50 1485
rect 16 1451 50 1481
rect 1666 1481 1700 1485
rect 1666 1451 1700 1481
rect 16 1379 50 1413
rect 841 1381 875 1415
rect 16 1311 50 1341
rect 1666 1379 1700 1413
rect 16 1307 50 1311
rect 841 1309 875 1343
rect 1666 1311 1700 1341
rect 1666 1307 1700 1311
rect 16 1243 50 1269
rect 16 1235 50 1243
rect 841 1237 875 1271
rect 16 1175 50 1197
rect 1666 1243 1700 1269
rect 1666 1235 1700 1243
rect 16 1163 50 1175
rect 841 1165 875 1199
rect 1666 1175 1700 1197
rect 1666 1163 1700 1175
rect 16 1107 50 1125
rect 16 1091 50 1107
rect 841 1093 875 1127
rect 16 1039 50 1053
rect 1666 1107 1700 1125
rect 1666 1091 1700 1107
rect 16 1019 50 1039
rect 841 1021 875 1055
rect 1666 1039 1700 1053
rect 1666 1019 1700 1039
rect 16 971 50 981
rect 16 947 50 971
rect 841 949 875 983
rect 16 903 50 909
rect 1666 971 1700 981
rect 1666 947 1700 971
rect 16 875 50 903
rect 841 877 875 911
rect 1666 903 1700 909
rect 1666 875 1700 903
rect 16 835 50 837
rect 16 803 50 835
rect 16 733 50 765
rect 16 731 50 733
rect 1666 835 1700 837
rect 1666 803 1700 835
rect 1666 733 1700 765
rect 1666 731 1700 733
rect 16 665 50 693
rect 16 659 50 665
rect 841 657 875 691
rect 1666 665 1700 693
rect 16 597 50 621
rect 16 587 50 597
rect 1666 659 1700 665
rect 841 585 875 619
rect 1666 597 1700 621
rect 1666 587 1700 597
rect 16 529 50 549
rect 16 515 50 529
rect 841 513 875 547
rect 1666 529 1700 549
rect 16 461 50 477
rect 16 443 50 461
rect 1666 515 1700 529
rect 841 441 875 475
rect 1666 461 1700 477
rect 1666 443 1700 461
rect 16 393 50 405
rect 16 371 50 393
rect 841 369 875 403
rect 1666 393 1700 405
rect 16 325 50 333
rect 16 299 50 325
rect 1666 371 1700 393
rect 841 297 875 331
rect 1666 325 1700 333
rect 1666 299 1700 325
rect 16 257 50 261
rect 16 227 50 257
rect 841 225 875 259
rect 1666 257 1700 261
rect 16 155 50 189
rect 1666 227 1700 257
rect 841 153 875 187
rect 1666 155 1700 189
rect 16 87 50 117
rect 16 83 50 87
rect 1666 87 1700 117
rect 1666 83 1700 87
rect 85 16 97 50
rect 97 16 119 50
rect 157 16 165 50
rect 165 16 191 50
rect 229 16 233 50
rect 233 16 263 50
rect 301 16 335 50
rect 373 16 403 50
rect 403 16 407 50
rect 445 16 471 50
rect 471 16 479 50
rect 517 16 539 50
rect 539 16 551 50
rect 589 16 607 50
rect 607 16 623 50
rect 661 16 675 50
rect 675 16 695 50
rect 733 16 743 50
rect 743 16 767 50
rect 805 16 811 50
rect 811 16 839 50
rect 877 16 897 50
rect 897 16 911 50
rect 949 16 965 50
rect 965 16 983 50
rect 1021 16 1033 50
rect 1033 16 1055 50
rect 1093 16 1101 50
rect 1101 16 1127 50
rect 1165 16 1169 50
rect 1169 16 1199 50
rect 1237 16 1271 50
rect 1309 16 1339 50
rect 1339 16 1343 50
rect 1381 16 1407 50
rect 1407 16 1415 50
rect 1453 16 1475 50
rect 1475 16 1487 50
rect 1525 16 1543 50
rect 1543 16 1559 50
rect 1597 16 1611 50
rect 1611 16 1631 50
<< metal1 >>
rect 0 1561 1716 1568
rect 0 1552 88 1561
rect 0 1518 85 1552
rect 0 1515 88 1518
rect 0 1463 7 1515
rect 59 1509 88 1515
rect 140 1509 152 1561
rect 204 1509 216 1561
rect 268 1509 280 1561
rect 332 1552 344 1561
rect 396 1552 408 1561
rect 460 1552 472 1561
rect 524 1552 536 1561
rect 588 1552 600 1561
rect 652 1552 664 1561
rect 335 1518 344 1552
rect 407 1518 408 1552
rect 588 1518 589 1552
rect 652 1518 661 1552
rect 332 1509 344 1518
rect 396 1509 408 1518
rect 460 1509 472 1518
rect 524 1509 536 1518
rect 588 1509 600 1518
rect 652 1509 664 1518
rect 716 1509 728 1561
rect 780 1552 942 1561
rect 780 1518 805 1552
rect 839 1518 877 1552
rect 911 1518 942 1552
rect 780 1509 942 1518
rect 994 1509 1006 1561
rect 1058 1509 1070 1561
rect 1122 1552 1134 1561
rect 1186 1552 1198 1561
rect 1250 1552 1262 1561
rect 1314 1552 1326 1561
rect 1378 1552 1390 1561
rect 1442 1552 1454 1561
rect 1127 1518 1134 1552
rect 1378 1518 1381 1552
rect 1442 1518 1453 1552
rect 1122 1509 1134 1518
rect 1186 1509 1198 1518
rect 1250 1509 1262 1518
rect 1314 1509 1326 1518
rect 1378 1509 1390 1518
rect 1442 1509 1454 1518
rect 1506 1509 1518 1561
rect 1570 1509 1582 1561
rect 1634 1515 1716 1561
rect 1634 1509 1657 1515
rect 59 1502 1657 1509
rect 59 1463 66 1502
rect 0 1451 16 1463
rect 50 1451 66 1463
rect 0 1399 7 1451
rect 59 1399 66 1451
rect 0 1387 16 1399
rect 50 1387 66 1399
rect 0 1335 7 1387
rect 59 1335 66 1387
rect 0 1323 16 1335
rect 50 1323 66 1335
rect 0 1271 7 1323
rect 59 1271 66 1323
rect 0 1269 66 1271
rect 0 1259 16 1269
rect 50 1259 66 1269
rect 0 1207 7 1259
rect 59 1207 66 1259
rect 0 1197 66 1207
rect 0 1195 16 1197
rect 50 1195 66 1197
rect 0 1143 7 1195
rect 59 1143 66 1195
rect 0 1131 66 1143
rect 0 1079 7 1131
rect 59 1079 66 1131
rect 0 1067 66 1079
rect 0 1015 7 1067
rect 59 1015 66 1067
rect 0 1003 66 1015
rect 0 951 7 1003
rect 59 951 66 1003
rect 0 947 16 951
rect 50 947 66 951
rect 0 939 66 947
rect 0 887 7 939
rect 59 887 66 939
rect 0 875 16 887
rect 50 875 66 887
rect 0 837 66 875
rect 0 803 16 837
rect 50 803 66 837
rect 0 765 66 803
rect 0 731 16 765
rect 50 731 66 765
rect 0 693 66 731
rect 0 681 16 693
rect 50 681 66 693
rect 0 629 7 681
rect 59 629 66 681
rect 0 621 66 629
rect 0 617 16 621
rect 50 617 66 621
rect 0 565 7 617
rect 59 565 66 617
rect 0 553 66 565
rect 0 501 7 553
rect 59 501 66 553
rect 0 489 66 501
rect 0 437 7 489
rect 59 437 66 489
rect 0 425 66 437
rect 0 373 7 425
rect 59 373 66 425
rect 0 371 16 373
rect 50 371 66 373
rect 0 361 66 371
rect 0 309 7 361
rect 59 309 66 361
rect 0 299 16 309
rect 50 299 66 309
rect 0 297 66 299
rect 0 245 7 297
rect 59 245 66 297
rect 0 233 16 245
rect 50 233 66 245
rect 0 181 7 233
rect 59 181 66 233
rect 0 169 16 181
rect 50 169 66 181
rect 0 117 7 169
rect 59 117 66 169
rect 0 105 16 117
rect 50 105 66 117
rect 0 53 7 105
rect 59 66 66 105
rect 99 816 127 1474
rect 155 844 183 1502
rect 211 816 239 1474
rect 267 844 295 1502
rect 323 816 351 1474
rect 379 844 407 1502
rect 435 816 463 1474
rect 491 844 519 1502
rect 547 816 575 1474
rect 603 844 631 1502
rect 659 816 687 1474
rect 715 844 743 1502
rect 771 816 799 1474
rect 831 1468 885 1474
rect 831 1416 832 1468
rect 884 1416 885 1468
rect 831 1415 885 1416
rect 831 1404 841 1415
rect 875 1404 885 1415
rect 831 1352 832 1404
rect 884 1352 885 1404
rect 831 1343 885 1352
rect 831 1340 841 1343
rect 875 1340 885 1343
rect 831 1288 832 1340
rect 884 1288 885 1340
rect 831 1276 885 1288
rect 831 1224 832 1276
rect 884 1224 885 1276
rect 831 1212 885 1224
rect 831 1160 832 1212
rect 884 1160 885 1212
rect 831 1148 885 1160
rect 831 1096 832 1148
rect 884 1096 885 1148
rect 831 1093 841 1096
rect 875 1093 885 1096
rect 831 1084 885 1093
rect 831 1032 832 1084
rect 884 1032 885 1084
rect 831 1021 841 1032
rect 875 1021 885 1032
rect 831 1020 885 1021
rect 831 968 832 1020
rect 884 968 885 1020
rect 831 956 841 968
rect 875 956 885 968
rect 831 904 832 956
rect 884 904 885 956
rect 831 892 841 904
rect 875 892 885 904
rect 831 840 832 892
rect 884 840 885 892
rect 831 816 885 840
rect 917 816 945 1474
rect 973 844 1001 1502
rect 1029 816 1057 1474
rect 1085 844 1113 1502
rect 1141 816 1169 1474
rect 1197 844 1225 1502
rect 1253 816 1281 1474
rect 1309 844 1337 1502
rect 1365 816 1393 1474
rect 1421 844 1449 1502
rect 1477 816 1505 1474
rect 1533 844 1561 1502
rect 1589 816 1617 1474
rect 99 810 1617 816
rect 99 758 105 810
rect 157 758 169 810
rect 221 758 233 810
rect 285 758 297 810
rect 349 758 361 810
rect 413 758 425 810
rect 477 758 489 810
rect 541 758 553 810
rect 605 758 617 810
rect 669 758 681 810
rect 733 758 745 810
rect 797 758 919 810
rect 971 758 983 810
rect 1035 758 1047 810
rect 1099 758 1111 810
rect 1163 758 1175 810
rect 1227 758 1239 810
rect 1291 758 1303 810
rect 1355 758 1367 810
rect 1419 758 1431 810
rect 1483 758 1495 810
rect 1547 758 1559 810
rect 1611 758 1617 810
rect 99 752 1617 758
rect 99 94 127 752
rect 155 66 183 724
rect 211 94 239 752
rect 267 66 295 724
rect 323 94 351 752
rect 379 66 407 724
rect 435 94 463 752
rect 491 66 519 724
rect 547 94 575 752
rect 603 66 631 724
rect 659 94 687 752
rect 715 66 743 724
rect 771 94 799 752
rect 831 728 885 752
rect 831 676 832 728
rect 884 676 885 728
rect 831 664 841 676
rect 875 664 885 676
rect 831 612 832 664
rect 884 612 885 664
rect 831 600 841 612
rect 875 600 885 612
rect 831 548 832 600
rect 884 548 885 600
rect 831 547 885 548
rect 831 536 841 547
rect 875 536 885 547
rect 831 484 832 536
rect 884 484 885 536
rect 831 475 885 484
rect 831 472 841 475
rect 875 472 885 475
rect 831 420 832 472
rect 884 420 885 472
rect 831 408 885 420
rect 831 356 832 408
rect 884 356 885 408
rect 831 344 885 356
rect 831 292 832 344
rect 884 292 885 344
rect 831 280 885 292
rect 831 228 832 280
rect 884 228 885 280
rect 831 225 841 228
rect 875 225 885 228
rect 831 216 885 225
rect 831 164 832 216
rect 884 164 885 216
rect 831 153 841 164
rect 875 153 885 164
rect 831 152 885 153
rect 831 100 832 152
rect 884 100 885 152
rect 831 94 885 100
rect 917 94 945 752
rect 973 66 1001 724
rect 1029 94 1057 752
rect 1085 66 1113 724
rect 1141 94 1169 752
rect 1197 66 1225 724
rect 1253 94 1281 752
rect 1309 66 1337 724
rect 1365 94 1393 752
rect 1421 66 1449 724
rect 1477 94 1505 752
rect 1533 66 1561 724
rect 1589 94 1617 752
rect 1650 1463 1657 1502
rect 1709 1463 1716 1515
rect 1650 1451 1666 1463
rect 1700 1451 1716 1463
rect 1650 1399 1657 1451
rect 1709 1399 1716 1451
rect 1650 1387 1666 1399
rect 1700 1387 1716 1399
rect 1650 1335 1657 1387
rect 1709 1335 1716 1387
rect 1650 1323 1666 1335
rect 1700 1323 1716 1335
rect 1650 1271 1657 1323
rect 1709 1271 1716 1323
rect 1650 1269 1716 1271
rect 1650 1259 1666 1269
rect 1700 1259 1716 1269
rect 1650 1207 1657 1259
rect 1709 1207 1716 1259
rect 1650 1197 1716 1207
rect 1650 1195 1666 1197
rect 1700 1195 1716 1197
rect 1650 1143 1657 1195
rect 1709 1143 1716 1195
rect 1650 1131 1716 1143
rect 1650 1079 1657 1131
rect 1709 1079 1716 1131
rect 1650 1067 1716 1079
rect 1650 1015 1657 1067
rect 1709 1015 1716 1067
rect 1650 1003 1716 1015
rect 1650 951 1657 1003
rect 1709 951 1716 1003
rect 1650 947 1666 951
rect 1700 947 1716 951
rect 1650 939 1716 947
rect 1650 887 1657 939
rect 1709 887 1716 939
rect 1650 875 1666 887
rect 1700 875 1716 887
rect 1650 837 1716 875
rect 1650 803 1666 837
rect 1700 803 1716 837
rect 1650 765 1716 803
rect 1650 731 1666 765
rect 1700 731 1716 765
rect 1650 693 1716 731
rect 1650 681 1666 693
rect 1700 681 1716 693
rect 1650 629 1657 681
rect 1709 629 1716 681
rect 1650 621 1716 629
rect 1650 617 1666 621
rect 1700 617 1716 621
rect 1650 565 1657 617
rect 1709 565 1716 617
rect 1650 553 1716 565
rect 1650 501 1657 553
rect 1709 501 1716 553
rect 1650 489 1716 501
rect 1650 437 1657 489
rect 1709 437 1716 489
rect 1650 425 1716 437
rect 1650 373 1657 425
rect 1709 373 1716 425
rect 1650 371 1666 373
rect 1700 371 1716 373
rect 1650 361 1716 371
rect 1650 309 1657 361
rect 1709 309 1716 361
rect 1650 299 1666 309
rect 1700 299 1716 309
rect 1650 297 1716 299
rect 1650 245 1657 297
rect 1709 245 1716 297
rect 1650 233 1666 245
rect 1700 233 1716 245
rect 1650 181 1657 233
rect 1709 181 1716 233
rect 1650 169 1666 181
rect 1700 169 1716 181
rect 1650 117 1657 169
rect 1709 117 1716 169
rect 1650 105 1666 117
rect 1700 105 1716 117
rect 1650 66 1657 105
rect 59 59 1657 66
rect 59 53 88 59
rect 0 50 88 53
rect 0 16 85 50
rect 0 7 88 16
rect 140 7 152 59
rect 204 7 216 59
rect 268 7 280 59
rect 332 50 344 59
rect 396 50 408 59
rect 460 50 472 59
rect 524 50 536 59
rect 588 50 600 59
rect 652 50 664 59
rect 335 16 344 50
rect 407 16 408 50
rect 588 16 589 50
rect 652 16 661 50
rect 332 7 344 16
rect 396 7 408 16
rect 460 7 472 16
rect 524 7 536 16
rect 588 7 600 16
rect 652 7 664 16
rect 716 7 728 59
rect 780 50 942 59
rect 780 16 805 50
rect 839 16 877 50
rect 911 16 942 50
rect 780 7 942 16
rect 994 7 1006 59
rect 1058 7 1070 59
rect 1122 50 1134 59
rect 1186 50 1198 59
rect 1250 50 1262 59
rect 1314 50 1326 59
rect 1378 50 1390 59
rect 1442 50 1454 59
rect 1127 16 1134 50
rect 1378 16 1381 50
rect 1442 16 1453 50
rect 1122 7 1134 16
rect 1186 7 1198 16
rect 1250 7 1262 16
rect 1314 7 1326 16
rect 1378 7 1390 16
rect 1442 7 1454 16
rect 1506 7 1518 59
rect 1570 7 1582 59
rect 1634 53 1657 59
rect 1709 53 1716 105
rect 1634 7 1716 53
rect 0 0 1716 7
<< via1 >>
rect 88 1552 140 1561
rect 88 1518 119 1552
rect 119 1518 140 1552
rect 7 1485 59 1515
rect 88 1509 140 1518
rect 152 1552 204 1561
rect 152 1518 157 1552
rect 157 1518 191 1552
rect 191 1518 204 1552
rect 152 1509 204 1518
rect 216 1552 268 1561
rect 216 1518 229 1552
rect 229 1518 263 1552
rect 263 1518 268 1552
rect 216 1509 268 1518
rect 280 1552 332 1561
rect 344 1552 396 1561
rect 408 1552 460 1561
rect 472 1552 524 1561
rect 536 1552 588 1561
rect 600 1552 652 1561
rect 664 1552 716 1561
rect 280 1518 301 1552
rect 301 1518 332 1552
rect 344 1518 373 1552
rect 373 1518 396 1552
rect 408 1518 445 1552
rect 445 1518 460 1552
rect 472 1518 479 1552
rect 479 1518 517 1552
rect 517 1518 524 1552
rect 536 1518 551 1552
rect 551 1518 588 1552
rect 600 1518 623 1552
rect 623 1518 652 1552
rect 664 1518 695 1552
rect 695 1518 716 1552
rect 280 1509 332 1518
rect 344 1509 396 1518
rect 408 1509 460 1518
rect 472 1509 524 1518
rect 536 1509 588 1518
rect 600 1509 652 1518
rect 664 1509 716 1518
rect 728 1552 780 1561
rect 942 1552 994 1561
rect 728 1518 733 1552
rect 733 1518 767 1552
rect 767 1518 780 1552
rect 942 1518 949 1552
rect 949 1518 983 1552
rect 983 1518 994 1552
rect 728 1509 780 1518
rect 942 1509 994 1518
rect 1006 1552 1058 1561
rect 1006 1518 1021 1552
rect 1021 1518 1055 1552
rect 1055 1518 1058 1552
rect 1006 1509 1058 1518
rect 1070 1552 1122 1561
rect 1134 1552 1186 1561
rect 1198 1552 1250 1561
rect 1262 1552 1314 1561
rect 1326 1552 1378 1561
rect 1390 1552 1442 1561
rect 1454 1552 1506 1561
rect 1070 1518 1093 1552
rect 1093 1518 1122 1552
rect 1134 1518 1165 1552
rect 1165 1518 1186 1552
rect 1198 1518 1199 1552
rect 1199 1518 1237 1552
rect 1237 1518 1250 1552
rect 1262 1518 1271 1552
rect 1271 1518 1309 1552
rect 1309 1518 1314 1552
rect 1326 1518 1343 1552
rect 1343 1518 1378 1552
rect 1390 1518 1415 1552
rect 1415 1518 1442 1552
rect 1454 1518 1487 1552
rect 1487 1518 1506 1552
rect 1070 1509 1122 1518
rect 1134 1509 1186 1518
rect 1198 1509 1250 1518
rect 1262 1509 1314 1518
rect 1326 1509 1378 1518
rect 1390 1509 1442 1518
rect 1454 1509 1506 1518
rect 1518 1552 1570 1561
rect 1518 1518 1525 1552
rect 1525 1518 1559 1552
rect 1559 1518 1570 1552
rect 1518 1509 1570 1518
rect 1582 1552 1634 1561
rect 1582 1518 1597 1552
rect 1597 1518 1631 1552
rect 1631 1518 1634 1552
rect 1582 1509 1634 1518
rect 7 1463 16 1485
rect 16 1463 50 1485
rect 50 1463 59 1485
rect 7 1413 59 1451
rect 7 1399 16 1413
rect 16 1399 50 1413
rect 50 1399 59 1413
rect 7 1379 16 1387
rect 16 1379 50 1387
rect 50 1379 59 1387
rect 7 1341 59 1379
rect 7 1335 16 1341
rect 16 1335 50 1341
rect 50 1335 59 1341
rect 7 1307 16 1323
rect 16 1307 50 1323
rect 50 1307 59 1323
rect 7 1271 59 1307
rect 7 1235 16 1259
rect 16 1235 50 1259
rect 50 1235 59 1259
rect 7 1207 59 1235
rect 7 1163 16 1195
rect 16 1163 50 1195
rect 50 1163 59 1195
rect 7 1143 59 1163
rect 7 1125 59 1131
rect 7 1091 16 1125
rect 16 1091 50 1125
rect 50 1091 59 1125
rect 7 1079 59 1091
rect 7 1053 59 1067
rect 7 1019 16 1053
rect 16 1019 50 1053
rect 50 1019 59 1053
rect 7 1015 59 1019
rect 7 981 59 1003
rect 7 951 16 981
rect 16 951 50 981
rect 50 951 59 981
rect 7 909 59 939
rect 7 887 16 909
rect 16 887 50 909
rect 50 887 59 909
rect 7 659 16 681
rect 16 659 50 681
rect 50 659 59 681
rect 7 629 59 659
rect 7 587 16 617
rect 16 587 50 617
rect 50 587 59 617
rect 7 565 59 587
rect 7 549 59 553
rect 7 515 16 549
rect 16 515 50 549
rect 50 515 59 549
rect 7 501 59 515
rect 7 477 59 489
rect 7 443 16 477
rect 16 443 50 477
rect 50 443 59 477
rect 7 437 59 443
rect 7 405 59 425
rect 7 373 16 405
rect 16 373 50 405
rect 50 373 59 405
rect 7 333 59 361
rect 7 309 16 333
rect 16 309 50 333
rect 50 309 59 333
rect 7 261 59 297
rect 7 245 16 261
rect 16 245 50 261
rect 50 245 59 261
rect 7 227 16 233
rect 16 227 50 233
rect 50 227 59 233
rect 7 189 59 227
rect 7 181 16 189
rect 16 181 50 189
rect 50 181 59 189
rect 7 155 16 169
rect 16 155 50 169
rect 50 155 59 169
rect 7 117 59 155
rect 7 83 16 105
rect 16 83 50 105
rect 50 83 59 105
rect 7 53 59 83
rect 832 1416 884 1468
rect 832 1381 841 1404
rect 841 1381 875 1404
rect 875 1381 884 1404
rect 832 1352 884 1381
rect 832 1309 841 1340
rect 841 1309 875 1340
rect 875 1309 884 1340
rect 832 1288 884 1309
rect 832 1271 884 1276
rect 832 1237 841 1271
rect 841 1237 875 1271
rect 875 1237 884 1271
rect 832 1224 884 1237
rect 832 1199 884 1212
rect 832 1165 841 1199
rect 841 1165 875 1199
rect 875 1165 884 1199
rect 832 1160 884 1165
rect 832 1127 884 1148
rect 832 1096 841 1127
rect 841 1096 875 1127
rect 875 1096 884 1127
rect 832 1055 884 1084
rect 832 1032 841 1055
rect 841 1032 875 1055
rect 875 1032 884 1055
rect 832 983 884 1020
rect 832 968 841 983
rect 841 968 875 983
rect 875 968 884 983
rect 832 949 841 956
rect 841 949 875 956
rect 875 949 884 956
rect 832 911 884 949
rect 832 904 841 911
rect 841 904 875 911
rect 875 904 884 911
rect 832 877 841 892
rect 841 877 875 892
rect 875 877 884 892
rect 832 840 884 877
rect 105 758 157 810
rect 169 758 221 810
rect 233 758 285 810
rect 297 758 349 810
rect 361 758 413 810
rect 425 758 477 810
rect 489 758 541 810
rect 553 758 605 810
rect 617 758 669 810
rect 681 758 733 810
rect 745 758 797 810
rect 919 758 971 810
rect 983 758 1035 810
rect 1047 758 1099 810
rect 1111 758 1163 810
rect 1175 758 1227 810
rect 1239 758 1291 810
rect 1303 758 1355 810
rect 1367 758 1419 810
rect 1431 758 1483 810
rect 1495 758 1547 810
rect 1559 758 1611 810
rect 832 691 884 728
rect 832 676 841 691
rect 841 676 875 691
rect 875 676 884 691
rect 832 657 841 664
rect 841 657 875 664
rect 875 657 884 664
rect 832 619 884 657
rect 832 612 841 619
rect 841 612 875 619
rect 875 612 884 619
rect 832 585 841 600
rect 841 585 875 600
rect 875 585 884 600
rect 832 548 884 585
rect 832 513 841 536
rect 841 513 875 536
rect 875 513 884 536
rect 832 484 884 513
rect 832 441 841 472
rect 841 441 875 472
rect 875 441 884 472
rect 832 420 884 441
rect 832 403 884 408
rect 832 369 841 403
rect 841 369 875 403
rect 875 369 884 403
rect 832 356 884 369
rect 832 331 884 344
rect 832 297 841 331
rect 841 297 875 331
rect 875 297 884 331
rect 832 292 884 297
rect 832 259 884 280
rect 832 228 841 259
rect 841 228 875 259
rect 875 228 884 259
rect 832 187 884 216
rect 832 164 841 187
rect 841 164 875 187
rect 875 164 884 187
rect 832 100 884 152
rect 1657 1485 1709 1515
rect 1657 1463 1666 1485
rect 1666 1463 1700 1485
rect 1700 1463 1709 1485
rect 1657 1413 1709 1451
rect 1657 1399 1666 1413
rect 1666 1399 1700 1413
rect 1700 1399 1709 1413
rect 1657 1379 1666 1387
rect 1666 1379 1700 1387
rect 1700 1379 1709 1387
rect 1657 1341 1709 1379
rect 1657 1335 1666 1341
rect 1666 1335 1700 1341
rect 1700 1335 1709 1341
rect 1657 1307 1666 1323
rect 1666 1307 1700 1323
rect 1700 1307 1709 1323
rect 1657 1271 1709 1307
rect 1657 1235 1666 1259
rect 1666 1235 1700 1259
rect 1700 1235 1709 1259
rect 1657 1207 1709 1235
rect 1657 1163 1666 1195
rect 1666 1163 1700 1195
rect 1700 1163 1709 1195
rect 1657 1143 1709 1163
rect 1657 1125 1709 1131
rect 1657 1091 1666 1125
rect 1666 1091 1700 1125
rect 1700 1091 1709 1125
rect 1657 1079 1709 1091
rect 1657 1053 1709 1067
rect 1657 1019 1666 1053
rect 1666 1019 1700 1053
rect 1700 1019 1709 1053
rect 1657 1015 1709 1019
rect 1657 981 1709 1003
rect 1657 951 1666 981
rect 1666 951 1700 981
rect 1700 951 1709 981
rect 1657 909 1709 939
rect 1657 887 1666 909
rect 1666 887 1700 909
rect 1700 887 1709 909
rect 1657 659 1666 681
rect 1666 659 1700 681
rect 1700 659 1709 681
rect 1657 629 1709 659
rect 1657 587 1666 617
rect 1666 587 1700 617
rect 1700 587 1709 617
rect 1657 565 1709 587
rect 1657 549 1709 553
rect 1657 515 1666 549
rect 1666 515 1700 549
rect 1700 515 1709 549
rect 1657 501 1709 515
rect 1657 477 1709 489
rect 1657 443 1666 477
rect 1666 443 1700 477
rect 1700 443 1709 477
rect 1657 437 1709 443
rect 1657 405 1709 425
rect 1657 373 1666 405
rect 1666 373 1700 405
rect 1700 373 1709 405
rect 1657 333 1709 361
rect 1657 309 1666 333
rect 1666 309 1700 333
rect 1700 309 1709 333
rect 1657 261 1709 297
rect 1657 245 1666 261
rect 1666 245 1700 261
rect 1700 245 1709 261
rect 1657 227 1666 233
rect 1666 227 1700 233
rect 1700 227 1709 233
rect 1657 189 1709 227
rect 1657 181 1666 189
rect 1666 181 1700 189
rect 1700 181 1709 189
rect 1657 155 1666 169
rect 1666 155 1700 169
rect 1700 155 1709 169
rect 1657 117 1709 155
rect 1657 83 1666 105
rect 1666 83 1700 105
rect 1700 83 1709 105
rect 88 50 140 59
rect 88 16 119 50
rect 119 16 140 50
rect 88 7 140 16
rect 152 50 204 59
rect 152 16 157 50
rect 157 16 191 50
rect 191 16 204 50
rect 152 7 204 16
rect 216 50 268 59
rect 216 16 229 50
rect 229 16 263 50
rect 263 16 268 50
rect 216 7 268 16
rect 280 50 332 59
rect 344 50 396 59
rect 408 50 460 59
rect 472 50 524 59
rect 536 50 588 59
rect 600 50 652 59
rect 664 50 716 59
rect 280 16 301 50
rect 301 16 332 50
rect 344 16 373 50
rect 373 16 396 50
rect 408 16 445 50
rect 445 16 460 50
rect 472 16 479 50
rect 479 16 517 50
rect 517 16 524 50
rect 536 16 551 50
rect 551 16 588 50
rect 600 16 623 50
rect 623 16 652 50
rect 664 16 695 50
rect 695 16 716 50
rect 280 7 332 16
rect 344 7 396 16
rect 408 7 460 16
rect 472 7 524 16
rect 536 7 588 16
rect 600 7 652 16
rect 664 7 716 16
rect 728 50 780 59
rect 942 50 994 59
rect 728 16 733 50
rect 733 16 767 50
rect 767 16 780 50
rect 942 16 949 50
rect 949 16 983 50
rect 983 16 994 50
rect 728 7 780 16
rect 942 7 994 16
rect 1006 50 1058 59
rect 1006 16 1021 50
rect 1021 16 1055 50
rect 1055 16 1058 50
rect 1006 7 1058 16
rect 1070 50 1122 59
rect 1134 50 1186 59
rect 1198 50 1250 59
rect 1262 50 1314 59
rect 1326 50 1378 59
rect 1390 50 1442 59
rect 1454 50 1506 59
rect 1070 16 1093 50
rect 1093 16 1122 50
rect 1134 16 1165 50
rect 1165 16 1186 50
rect 1198 16 1199 50
rect 1199 16 1237 50
rect 1237 16 1250 50
rect 1262 16 1271 50
rect 1271 16 1309 50
rect 1309 16 1314 50
rect 1326 16 1343 50
rect 1343 16 1378 50
rect 1390 16 1415 50
rect 1415 16 1442 50
rect 1454 16 1487 50
rect 1487 16 1506 50
rect 1070 7 1122 16
rect 1134 7 1186 16
rect 1198 7 1250 16
rect 1262 7 1314 16
rect 1326 7 1378 16
rect 1390 7 1442 16
rect 1454 7 1506 16
rect 1518 50 1570 59
rect 1518 16 1525 50
rect 1525 16 1559 50
rect 1559 16 1570 50
rect 1518 7 1570 16
rect 1582 50 1634 59
rect 1657 53 1709 83
rect 1582 16 1597 50
rect 1597 16 1631 50
rect 1631 16 1634 50
rect 1582 7 1634 16
<< metal2 >>
rect 0 1561 803 1568
rect 0 1515 88 1561
rect 0 1463 7 1515
rect 59 1509 88 1515
rect 140 1509 152 1561
rect 204 1509 216 1561
rect 268 1509 280 1561
rect 332 1509 344 1561
rect 396 1509 408 1561
rect 460 1509 472 1561
rect 524 1509 536 1561
rect 588 1509 600 1561
rect 652 1509 664 1561
rect 716 1509 728 1561
rect 780 1509 803 1561
rect 59 1502 803 1509
rect 59 1463 66 1502
rect 831 1474 885 1568
rect 913 1561 1716 1568
rect 913 1509 942 1561
rect 994 1509 1006 1561
rect 1058 1509 1070 1561
rect 1122 1509 1134 1561
rect 1186 1509 1198 1561
rect 1250 1509 1262 1561
rect 1314 1509 1326 1561
rect 1378 1509 1390 1561
rect 1442 1509 1454 1561
rect 1506 1509 1518 1561
rect 1570 1509 1582 1561
rect 1634 1515 1716 1561
rect 1634 1509 1657 1515
rect 913 1502 1657 1509
rect 0 1451 66 1463
rect 0 1399 7 1451
rect 59 1418 66 1451
rect 94 1468 1622 1474
rect 94 1446 832 1468
rect 59 1399 803 1418
rect 0 1390 803 1399
rect 831 1416 832 1446
rect 884 1446 1622 1468
rect 1650 1463 1657 1502
rect 1709 1463 1716 1515
rect 1650 1451 1716 1463
rect 884 1416 885 1446
rect 1650 1418 1657 1451
rect 831 1404 885 1416
rect 0 1387 66 1390
rect 0 1335 7 1387
rect 59 1335 66 1387
rect 831 1362 832 1404
rect 0 1323 66 1335
rect 94 1352 832 1362
rect 884 1362 885 1404
rect 913 1399 1657 1418
rect 1709 1399 1716 1451
rect 913 1390 1716 1399
rect 1650 1387 1716 1390
rect 884 1352 1622 1362
rect 94 1340 1622 1352
rect 94 1334 832 1340
rect 0 1271 7 1323
rect 59 1306 66 1323
rect 59 1278 803 1306
rect 831 1288 832 1334
rect 884 1334 1622 1340
rect 1650 1335 1657 1387
rect 1709 1335 1716 1387
rect 884 1288 885 1334
rect 1650 1323 1716 1335
rect 1650 1306 1657 1323
rect 59 1271 66 1278
rect 0 1259 66 1271
rect 0 1207 7 1259
rect 59 1207 66 1259
rect 831 1276 885 1288
rect 913 1278 1657 1306
rect 831 1250 832 1276
rect 94 1224 832 1250
rect 884 1250 885 1276
rect 1650 1271 1657 1278
rect 1709 1271 1716 1323
rect 1650 1259 1716 1271
rect 884 1224 1622 1250
rect 94 1222 1622 1224
rect 0 1195 66 1207
rect 0 1143 7 1195
rect 59 1194 66 1195
rect 831 1212 885 1222
rect 59 1166 803 1194
rect 59 1143 66 1166
rect 0 1131 66 1143
rect 831 1160 832 1212
rect 884 1160 885 1212
rect 1650 1207 1657 1259
rect 1709 1207 1716 1259
rect 1650 1195 1716 1207
rect 1650 1194 1657 1195
rect 913 1166 1657 1194
rect 831 1148 885 1160
rect 831 1138 832 1148
rect 0 1079 7 1131
rect 59 1082 66 1131
rect 94 1110 832 1138
rect 831 1096 832 1110
rect 884 1138 885 1148
rect 1650 1143 1657 1166
rect 1709 1143 1716 1195
rect 884 1110 1622 1138
rect 1650 1131 1716 1143
rect 884 1096 885 1110
rect 831 1084 885 1096
rect 59 1079 803 1082
rect 0 1067 803 1079
rect 0 1015 7 1067
rect 59 1054 803 1067
rect 59 1015 66 1054
rect 831 1032 832 1084
rect 884 1032 885 1084
rect 1650 1082 1657 1131
rect 913 1079 1657 1082
rect 1709 1079 1716 1131
rect 913 1067 1716 1079
rect 913 1054 1657 1067
rect 831 1026 885 1032
rect 0 1003 66 1015
rect 0 951 7 1003
rect 59 970 66 1003
rect 94 1020 1622 1026
rect 94 998 832 1020
rect 59 951 803 970
rect 0 942 803 951
rect 831 968 832 998
rect 884 998 1622 1020
rect 1650 1015 1657 1054
rect 1709 1015 1716 1067
rect 1650 1003 1716 1015
rect 884 968 885 998
rect 1650 970 1657 1003
rect 831 956 885 968
rect 0 939 66 942
rect 0 887 7 939
rect 59 887 66 939
rect 831 914 832 956
rect 0 839 66 887
rect 94 904 832 914
rect 884 914 885 956
rect 913 951 1657 970
rect 1709 951 1716 1003
rect 913 942 1716 951
rect 1650 939 1716 942
rect 884 904 1622 914
rect 94 892 1622 904
rect 94 886 832 892
rect 831 840 832 886
rect 884 886 1622 892
rect 1650 887 1657 939
rect 1709 887 1716 939
rect 884 840 885 886
rect 831 811 885 840
rect 1650 839 1716 887
rect 0 810 1716 811
rect 0 758 105 810
rect 157 758 169 810
rect 221 758 233 810
rect 285 758 297 810
rect 349 758 361 810
rect 413 758 425 810
rect 477 758 489 810
rect 541 758 553 810
rect 605 758 617 810
rect 669 758 681 810
rect 733 758 745 810
rect 797 758 919 810
rect 971 758 983 810
rect 1035 758 1047 810
rect 1099 758 1111 810
rect 1163 758 1175 810
rect 1227 758 1239 810
rect 1291 758 1303 810
rect 1355 758 1367 810
rect 1419 758 1431 810
rect 1483 758 1495 810
rect 1547 758 1559 810
rect 1611 758 1716 810
rect 0 757 1716 758
rect 0 681 66 729
rect 831 728 885 757
rect 831 682 832 728
rect 0 629 7 681
rect 59 629 66 681
rect 94 676 832 682
rect 884 682 885 728
rect 884 676 1622 682
rect 94 664 1622 676
rect 94 654 832 664
rect 0 626 66 629
rect 0 617 803 626
rect 0 565 7 617
rect 59 598 803 617
rect 831 612 832 654
rect 884 654 1622 664
rect 1650 681 1716 729
rect 884 612 885 654
rect 1650 629 1657 681
rect 1709 629 1716 681
rect 1650 626 1716 629
rect 831 600 885 612
rect 59 565 66 598
rect 831 570 832 600
rect 0 553 66 565
rect 0 501 7 553
rect 59 514 66 553
rect 94 548 832 570
rect 884 570 885 600
rect 913 617 1716 626
rect 913 598 1657 617
rect 884 548 1622 570
rect 94 542 1622 548
rect 1650 565 1657 598
rect 1709 565 1716 617
rect 1650 553 1716 565
rect 831 536 885 542
rect 59 501 803 514
rect 0 489 803 501
rect 0 437 7 489
rect 59 486 803 489
rect 59 437 66 486
rect 831 484 832 536
rect 884 484 885 536
rect 1650 514 1657 553
rect 913 501 1657 514
rect 1709 501 1716 553
rect 913 489 1716 501
rect 913 486 1657 489
rect 831 472 885 484
rect 831 458 832 472
rect 0 425 66 437
rect 94 430 832 458
rect 0 373 7 425
rect 59 402 66 425
rect 831 420 832 430
rect 884 458 885 472
rect 884 430 1622 458
rect 1650 437 1657 486
rect 1709 437 1716 489
rect 884 420 885 430
rect 831 408 885 420
rect 59 374 803 402
rect 59 373 66 374
rect 0 361 66 373
rect 0 309 7 361
rect 59 309 66 361
rect 831 356 832 408
rect 884 356 885 408
rect 1650 425 1716 437
rect 1650 402 1657 425
rect 913 374 1657 402
rect 831 346 885 356
rect 1650 373 1657 374
rect 1709 373 1716 425
rect 1650 361 1716 373
rect 94 344 1622 346
rect 94 318 832 344
rect 0 297 66 309
rect 0 245 7 297
rect 59 290 66 297
rect 831 292 832 318
rect 884 318 1622 344
rect 884 292 885 318
rect 59 262 803 290
rect 831 280 885 292
rect 1650 309 1657 361
rect 1709 309 1716 361
rect 1650 297 1716 309
rect 1650 290 1657 297
rect 59 245 66 262
rect 0 233 66 245
rect 831 234 832 280
rect 0 181 7 233
rect 59 181 66 233
rect 94 228 832 234
rect 884 234 885 280
rect 913 262 1657 290
rect 1650 245 1657 262
rect 1709 245 1716 297
rect 884 228 1622 234
rect 94 216 1622 228
rect 94 206 832 216
rect 0 178 66 181
rect 0 169 803 178
rect 0 117 7 169
rect 59 150 803 169
rect 831 164 832 206
rect 884 206 1622 216
rect 1650 233 1716 245
rect 884 164 885 206
rect 1650 181 1657 233
rect 1709 181 1716 233
rect 1650 178 1716 181
rect 831 152 885 164
rect 59 117 66 150
rect 831 122 832 152
rect 0 105 66 117
rect 0 53 7 105
rect 59 66 66 105
rect 94 100 832 122
rect 884 122 885 152
rect 913 169 1716 178
rect 913 150 1657 169
rect 884 100 1622 122
rect 94 94 1622 100
rect 1650 117 1657 150
rect 1709 117 1716 169
rect 1650 105 1716 117
rect 59 59 803 66
rect 59 53 88 59
rect 0 7 88 53
rect 140 7 152 59
rect 204 7 216 59
rect 268 7 280 59
rect 332 7 344 59
rect 396 7 408 59
rect 460 7 472 59
rect 524 7 536 59
rect 588 7 600 59
rect 652 7 664 59
rect 716 7 728 59
rect 780 7 803 59
rect 0 0 803 7
rect 831 0 885 94
rect 1650 66 1657 105
rect 913 59 1657 66
rect 913 7 942 59
rect 994 7 1006 59
rect 1058 7 1070 59
rect 1122 7 1134 59
rect 1186 7 1198 59
rect 1250 7 1262 59
rect 1314 7 1326 59
rect 1378 7 1390 59
rect 1442 7 1454 59
rect 1506 7 1518 59
rect 1570 7 1582 59
rect 1634 53 1657 59
rect 1709 53 1716 105
rect 1634 7 1716 53
rect 913 0 1716 7
<< metal3 >>
rect 0 0 1716 1568
<< labels >>
flabel metal3 s 1189 266 1340 379 0 FreeSans 1000 0 0 0 MET3
port 4 nsew
flabel pwell s 894 821 918 872 0 FreeSans 200 0 0 0 SUB
port 3 nsew
flabel metal2 s 840 1518 878 1555 0 FreeSans 400 0 0 0 C1
port 2 nsew
flabel metal2 s 646 1533 672 1563 0 FreeSans 400 0 0 0 C0
port 1 nsew
<< properties >>
string GDS_END 216756
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 182004
string device primitive
<< end >>
