magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -89 -36 309 236
<< pmoshvt >>
rect 0 0 36 200
rect 92 0 128 200
rect 184 0 220 200
<< pdiff >>
rect -50 0 0 200
rect 36 182 92 200
rect 36 148 47 182
rect 81 148 92 182
rect 36 114 92 148
rect 36 80 47 114
rect 81 80 92 114
rect 36 46 92 80
rect 36 12 47 46
rect 81 12 92 46
rect 36 0 92 12
rect 128 182 184 200
rect 128 148 139 182
rect 173 148 184 182
rect 128 114 184 148
rect 128 80 139 114
rect 173 80 184 114
rect 128 46 184 80
rect 128 12 139 46
rect 173 12 184 46
rect 128 0 184 12
rect 220 0 270 200
<< pdiffc >>
rect 47 148 81 182
rect 47 80 81 114
rect 47 12 81 46
rect 139 148 173 182
rect 139 80 173 114
rect 139 12 173 46
<< poly >>
rect 0 200 36 226
rect 92 200 128 226
rect 184 200 220 226
rect 0 -26 36 0
rect 92 -26 128 0
rect 184 -26 220 0
<< locali >>
rect 47 182 81 198
rect 47 114 81 148
rect 47 46 81 80
rect 47 -4 81 12
rect 139 182 173 198
rect 139 114 173 148
rect 139 46 173 80
rect 139 -4 173 12
<< metal1 >>
rect -51 -16 -5 186
rect 225 -16 271 186
use hvDFL1sd2_CDNS_52468879185110  hvDFL1sd2_CDNS_52468879185110_0
timestamp 1704896540
transform 1 0 128 0 1 0
box 0 0 1 1
use hvDFL1sd2_CDNS_52468879185110  hvDFL1sd2_CDNS_52468879185110_1
timestamp 1704896540
transform 1 0 36 0 1 0
box 0 0 1 1
use hvDFM1sd_CDNS_52468879185130  hvDFM1sd_CDNS_52468879185130_0
timestamp 1704896540
transform -1 0 0 0 1 0
box -36 -36 89 236
use hvDFM1sd_CDNS_52468879185130  hvDFM1sd_CDNS_52468879185130_1
timestamp 1704896540
transform 1 0 220 0 1 0
box -36 -36 89 236
<< labels >>
flabel comment s -28 85 -28 85 0 FreeSans 300 0 0 0 S
flabel comment s 64 97 64 97 0 FreeSans 300 0 0 0 D
flabel comment s 156 97 156 97 0 FreeSans 300 0 0 0 S
flabel comment s 248 85 248 85 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 86828712
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86826758
<< end >>
