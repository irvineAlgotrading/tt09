magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 1 21 643 203
rect 29 -17 63 21
<< locali >>
rect 284 391 357 493
rect 284 357 389 391
rect 30 199 104 323
rect 145 202 248 255
rect 355 165 389 357
rect 449 199 522 323
rect 556 199 614 323
rect 355 51 441 165
rect 488 85 522 199
<< obsli1 >>
rect 0 527 644 561
rect 19 361 85 527
rect 175 323 241 493
rect 391 447 457 493
rect 423 391 457 447
rect 491 427 541 527
rect 575 391 626 493
rect 423 357 626 391
rect 175 289 316 323
rect 282 166 316 289
rect 19 17 85 165
rect 119 132 316 166
rect 119 51 153 132
rect 187 17 321 98
rect 559 17 625 165
rect 0 -17 644 17
<< metal1 >>
rect 0 496 644 592
rect 0 -48 644 48
<< labels >>
rlabel locali s 30 199 104 323 6 A1_N
port 1 nsew signal input
rlabel locali s 145 202 248 255 6 A2_N
port 2 nsew signal input
rlabel locali s 556 199 614 323 6 B1
port 3 nsew signal input
rlabel locali s 488 85 522 199 6 B2
port 4 nsew signal input
rlabel locali s 449 199 522 323 6 B2
port 4 nsew signal input
rlabel metal1 s 0 -48 644 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1 21 643 203 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 682 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 644 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 355 51 441 165 6 Y
port 9 nsew signal output
rlabel locali s 355 165 389 357 6 Y
port 9 nsew signal output
rlabel locali s 284 357 389 391 6 Y
port 9 nsew signal output
rlabel locali s 284 391 357 493 6 Y
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 644 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3937388
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3930540
<< end >>
