magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< pwell >>
rect -79 -26 112 226
<< nmos >>
rect 0 0 36 200
<< ndiff >>
rect -53 182 0 200
rect -53 148 -45 182
rect -11 148 0 182
rect -53 114 0 148
rect -53 80 -45 114
rect -11 80 0 114
rect -53 46 0 80
rect -53 12 -45 46
rect -11 12 0 46
rect -53 0 0 12
rect 36 0 86 200
<< ndiffc >>
rect -45 148 -11 182
rect -45 80 -11 114
rect -45 12 -11 46
<< poly >>
rect 0 200 36 226
rect 0 -26 36 0
<< locali >>
rect -45 182 -11 198
rect -45 114 -11 148
rect -45 46 -11 80
rect -45 -4 -11 12
<< metal1 >>
rect 41 -16 87 186
use hvDFL1sd_CDNS_52468879185132  hvDFL1sd_CDNS_52468879185132_0
timestamp 1704896540
transform -1 0 0 0 1 0
box 0 0 1 1
use hvDFM1sd_CDNS_52468879185147  hvDFM1sd_CDNS_52468879185147_0
timestamp 1704896540
transform 1 0 36 0 1 0
box -26 -26 79 226
<< labels >>
flabel comment s -28 97 -28 97 0 FreeSans 300 0 0 0 S
flabel comment s 64 85 64 85 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 86855958
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86855132
<< end >>
