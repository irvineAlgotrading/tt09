magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -122 -66 519 216
<< mvpmos >>
rect 0 0 400 150
<< mvpdiff >>
rect -56 114 0 150
rect -56 80 -45 114
rect -11 80 0 114
rect -56 46 0 80
rect -56 12 -45 46
rect -11 12 0 46
rect -56 0 0 12
rect 400 114 453 150
rect 400 80 411 114
rect 445 80 453 114
rect 400 46 453 80
rect 400 12 411 46
rect 445 12 453 46
rect 400 0 453 12
<< mvpdiffc >>
rect -45 80 -11 114
rect -45 12 -11 46
rect 411 80 445 114
rect 411 12 445 46
<< poly >>
rect 0 150 400 182
rect 0 -32 400 0
<< locali >>
rect -45 114 -11 130
rect -45 46 -11 80
rect -45 -4 -11 12
rect 411 114 445 130
rect 411 46 445 68
<< viali >>
rect 411 80 445 102
rect 411 68 445 80
rect 411 12 445 30
rect 411 -4 445 12
<< metal1 >>
rect 405 102 451 114
rect 405 68 411 102
rect 445 68 451 102
rect 405 30 451 68
rect 405 -4 411 30
rect 445 -4 451 30
rect 405 -16 451 -4
use hvDFL1sd2_CDNS_52468879185654  hvDFL1sd2_CDNS_52468879185654_0
timestamp 1704896540
transform -1 0 0 0 1 0
box 0 0 1 1
use hvDFM1sd_CDNS_52468879185172  hvDFM1sd_CDNS_52468879185172_0
timestamp 1704896540
transform 1 0 400 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s -28 63 -28 63 0 FreeSans 300 0 0 0 S
flabel comment s 428 49 428 49 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 85608810
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85607790
<< end >>
