magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect 415 600 14720 4720
<< pwell >>
rect 95 5094 249 5109
rect 95 4872 14968 5094
rect 95 525 355 4872
rect 14781 525 14968 4872
rect 95 303 14968 525
<< mvpsubdiff >>
rect 121 5021 223 5083
rect 272 4898 306 5068
rect 13600 5034 13635 5068
rect 13669 5034 13704 5068
rect 13738 5034 13773 5068
rect 13807 5034 13842 5068
rect 13876 5034 13911 5068
rect 13945 5034 13980 5068
rect 14014 5034 14049 5068
rect 14083 5034 14118 5068
rect 14152 5034 14187 5068
rect 14221 5034 14256 5068
rect 14290 5034 14325 5068
rect 14359 5034 14394 5068
rect 14428 5034 14463 5068
rect 14497 5034 14532 5068
rect 14566 5034 14601 5068
rect 14635 5034 14670 5068
rect 14704 5034 14739 5068
rect 14773 5034 14942 5068
rect 13600 5033 14942 5034
rect 13600 5000 14840 5033
rect 13600 4966 13635 5000
rect 13669 4966 13704 5000
rect 13738 4966 13773 5000
rect 13807 4966 13842 5000
rect 13876 4966 13911 5000
rect 13945 4966 13980 5000
rect 14014 4966 14049 5000
rect 14083 4966 14118 5000
rect 14152 4966 14187 5000
rect 14221 4966 14256 5000
rect 14290 4966 14325 5000
rect 14359 4966 14394 5000
rect 14428 4966 14463 5000
rect 14497 4966 14532 5000
rect 14566 4966 14601 5000
rect 14635 4966 14670 5000
rect 14704 4966 14739 5000
rect 14773 4999 14840 5000
rect 14874 4999 14942 5033
rect 14773 4966 14942 4999
rect 13600 4965 14942 4966
rect 13600 4932 14840 4965
rect 13600 4898 13635 4932
rect 13669 4898 13704 4932
rect 13738 4898 13773 4932
rect 13807 4898 13842 4932
rect 13876 4898 13911 4932
rect 13945 4898 13980 4932
rect 14014 4898 14049 4932
rect 14083 4898 14118 4932
rect 14152 4898 14187 4932
rect 14221 4898 14256 4932
rect 14290 4898 14325 4932
rect 14359 4898 14394 4932
rect 14428 4898 14463 4932
rect 14497 4898 14532 4932
rect 14566 4898 14601 4932
rect 14635 4898 14670 4932
rect 14704 4898 14739 4932
rect 14773 4898 14840 4932
rect 229 4859 329 4883
rect 229 4825 262 4859
rect 296 4825 329 4859
rect 229 4791 329 4825
rect 229 4757 262 4791
rect 296 4757 329 4791
rect 229 4723 329 4757
rect 229 4689 262 4723
rect 296 4689 329 4723
rect 229 4655 329 4689
rect 229 4621 262 4655
rect 296 4621 329 4655
rect 229 4587 329 4621
rect 229 4553 262 4587
rect 296 4553 329 4587
rect 229 4519 329 4553
rect 229 4485 262 4519
rect 296 4485 329 4519
rect 229 4451 329 4485
rect 229 4417 262 4451
rect 296 4417 329 4451
rect 229 4383 329 4417
rect 229 4349 262 4383
rect 296 4349 329 4383
rect 229 4315 329 4349
rect 229 4281 262 4315
rect 296 4281 329 4315
rect 229 4247 329 4281
rect 229 4213 262 4247
rect 296 4213 329 4247
rect 229 4179 329 4213
rect 229 4145 262 4179
rect 296 4145 329 4179
rect 229 4111 329 4145
rect 229 4077 262 4111
rect 296 4077 329 4111
rect 229 4043 329 4077
rect 229 4009 262 4043
rect 296 4009 329 4043
rect 229 3975 329 4009
rect 229 3941 262 3975
rect 296 3941 329 3975
rect 229 3907 329 3941
rect 229 3873 262 3907
rect 296 3873 329 3907
rect 229 3839 329 3873
rect 229 3805 262 3839
rect 296 3805 329 3839
rect 229 3771 329 3805
rect 229 3737 262 3771
rect 296 3737 329 3771
rect 229 3703 329 3737
rect 229 3669 262 3703
rect 296 3669 329 3703
rect 229 3635 329 3669
rect 229 3601 262 3635
rect 296 3601 329 3635
rect 229 3567 329 3601
rect 229 3533 262 3567
rect 296 3533 329 3567
rect 229 3499 329 3533
rect 229 3465 262 3499
rect 296 3465 329 3499
rect 229 3431 329 3465
rect 229 3397 262 3431
rect 296 3397 329 3431
rect 229 3363 329 3397
rect 229 3329 262 3363
rect 296 3329 329 3363
rect 229 3295 329 3329
rect 229 3261 262 3295
rect 296 3261 329 3295
rect 229 3227 329 3261
rect 229 3193 262 3227
rect 296 3193 329 3227
rect 229 3159 329 3193
rect 229 3125 262 3159
rect 296 3125 329 3159
rect 229 3091 329 3125
rect 229 3057 262 3091
rect 296 3057 329 3091
rect 229 3023 329 3057
rect 229 2989 262 3023
rect 296 2989 329 3023
rect 229 2955 329 2989
rect 229 2921 262 2955
rect 296 2921 329 2955
rect 229 2887 329 2921
rect 229 2853 262 2887
rect 296 2853 329 2887
rect 229 2819 329 2853
rect 229 2785 262 2819
rect 296 2785 329 2819
rect 229 2751 329 2785
rect 229 2717 262 2751
rect 296 2717 329 2751
rect 229 2683 329 2717
rect 229 2649 262 2683
rect 296 2649 329 2683
rect 229 2615 329 2649
rect 229 2581 262 2615
rect 296 2581 329 2615
rect 229 2547 329 2581
rect 229 2513 262 2547
rect 296 2513 329 2547
rect 229 2479 329 2513
rect 229 2445 262 2479
rect 296 2445 329 2479
rect 229 2411 329 2445
rect 229 2377 262 2411
rect 296 2377 329 2411
rect 229 2343 329 2377
rect 229 2309 262 2343
rect 296 2309 329 2343
rect 229 2275 329 2309
rect 229 2241 262 2275
rect 296 2241 329 2275
rect 229 2207 329 2241
rect 229 2173 262 2207
rect 296 2173 329 2207
rect 229 2139 329 2173
rect 229 2105 262 2139
rect 296 2105 329 2139
rect 229 2071 329 2105
rect 229 2037 262 2071
rect 296 2037 329 2071
rect 229 2003 329 2037
rect 229 1969 262 2003
rect 296 1969 329 2003
rect 229 1935 329 1969
rect 229 1901 262 1935
rect 296 1901 329 1935
rect 229 1867 329 1901
rect 229 1833 262 1867
rect 296 1833 329 1867
rect 229 1799 329 1833
rect 229 1765 262 1799
rect 296 1765 329 1799
rect 229 1731 329 1765
rect 229 1697 262 1731
rect 296 1697 329 1731
rect 229 1663 329 1697
rect 229 1629 262 1663
rect 296 1629 329 1663
rect 229 1595 329 1629
rect 229 1561 262 1595
rect 296 1561 329 1595
rect 229 1527 329 1561
rect 229 1493 262 1527
rect 296 1493 329 1527
rect 229 1459 329 1493
rect 229 1425 262 1459
rect 296 1425 329 1459
rect 229 1391 329 1425
rect 229 1357 262 1391
rect 296 1357 329 1391
rect 229 1323 329 1357
rect 229 1289 262 1323
rect 296 1289 329 1323
rect 229 1255 329 1289
rect 229 1221 262 1255
rect 296 1221 329 1255
rect 229 1187 329 1221
rect 229 1153 262 1187
rect 296 1153 329 1187
rect 229 1119 329 1153
rect 229 1085 262 1119
rect 296 1085 329 1119
rect 229 1051 329 1085
rect 229 1017 262 1051
rect 296 1017 329 1051
rect 229 983 329 1017
rect 229 949 262 983
rect 296 949 329 983
rect 229 915 329 949
rect 229 881 262 915
rect 296 881 329 915
rect 229 847 329 881
rect 229 813 262 847
rect 296 813 329 847
rect 229 779 329 813
rect 229 745 262 779
rect 296 745 329 779
rect 229 711 329 745
rect 229 677 262 711
rect 296 677 329 711
rect 229 643 329 677
rect 229 609 262 643
rect 296 609 329 643
rect 229 575 329 609
rect 229 541 262 575
rect 296 541 329 575
rect 229 514 329 541
rect 14807 499 14840 4898
rect 121 329 223 363
rect 228 465 262 499
rect 296 465 331 499
rect 365 465 400 499
rect 434 465 469 499
rect 503 465 538 499
rect 572 465 607 499
rect 641 465 676 499
rect 710 465 745 499
rect 779 465 814 499
rect 848 465 883 499
rect 917 465 952 499
rect 986 465 1021 499
rect 1055 465 1090 499
rect 1124 465 1159 499
rect 1193 465 1228 499
rect 1262 465 1297 499
rect 1331 465 1366 499
rect 1400 465 1435 499
rect 1469 465 1504 499
rect 1538 465 1573 499
rect 1607 465 1642 499
rect 1676 465 1711 499
rect 1745 465 1780 499
rect 1814 465 1849 499
rect 1883 465 1918 499
rect 1952 465 1987 499
rect 2021 465 2056 499
rect 228 431 2056 465
rect 228 397 262 431
rect 296 397 331 431
rect 365 397 400 431
rect 434 397 469 431
rect 503 397 538 431
rect 572 397 607 431
rect 641 397 676 431
rect 710 397 745 431
rect 779 397 814 431
rect 848 397 883 431
rect 917 397 952 431
rect 986 397 1021 431
rect 1055 397 1090 431
rect 1124 397 1159 431
rect 1193 397 1228 431
rect 1262 397 1297 431
rect 1331 397 1366 431
rect 1400 397 1435 431
rect 1469 397 1504 431
rect 1538 397 1573 431
rect 1607 397 1642 431
rect 1676 397 1711 431
rect 1745 397 1780 431
rect 1814 397 1849 431
rect 1883 397 1918 431
rect 1952 397 1987 431
rect 2021 397 2056 431
rect 228 363 2056 397
rect 228 329 262 363
rect 296 329 331 363
rect 365 329 400 363
rect 434 329 469 363
rect 503 329 538 363
rect 572 329 607 363
rect 641 329 676 363
rect 710 329 745 363
rect 779 329 814 363
rect 848 329 883 363
rect 917 329 952 363
rect 986 329 1021 363
rect 1055 329 1090 363
rect 1124 329 1159 363
rect 1193 329 1228 363
rect 1262 329 1297 363
rect 1331 329 1366 363
rect 1400 329 1435 363
rect 1469 329 1504 363
rect 1538 329 1573 363
rect 1607 329 1642 363
rect 1676 329 1711 363
rect 1745 329 1780 363
rect 1814 329 1849 363
rect 1883 329 1918 363
rect 1952 329 1987 363
rect 2021 329 2056 363
rect 14806 329 14942 375
<< mvnsubdiff >>
rect 482 4638 14653 4653
rect 482 4619 584 4638
rect 482 4585 497 4619
rect 531 4585 584 4619
rect 482 4570 584 4585
rect 10410 4604 10445 4638
rect 10479 4604 10514 4638
rect 10548 4604 10583 4638
rect 10617 4604 10652 4638
rect 10686 4604 10721 4638
rect 10755 4604 10790 4638
rect 10824 4604 10859 4638
rect 10893 4604 10928 4638
rect 10962 4604 10997 4638
rect 11031 4604 11066 4638
rect 11100 4604 11135 4638
rect 11169 4604 11204 4638
rect 11238 4604 11273 4638
rect 11307 4604 11342 4638
rect 11376 4604 11411 4638
rect 11445 4604 11480 4638
rect 11514 4604 11549 4638
rect 11583 4604 11618 4638
rect 11652 4604 11687 4638
rect 11721 4604 11756 4638
rect 11790 4604 11825 4638
rect 11859 4604 11894 4638
rect 11928 4604 11963 4638
rect 11997 4604 12032 4638
rect 12066 4604 12101 4638
rect 12135 4604 12170 4638
rect 12204 4604 12239 4638
rect 12273 4604 12308 4638
rect 12342 4604 12377 4638
rect 12411 4604 12446 4638
rect 12480 4604 12515 4638
rect 12549 4604 12584 4638
rect 12618 4604 12653 4638
rect 12687 4604 12722 4638
rect 12756 4604 12791 4638
rect 12825 4604 12860 4638
rect 12894 4604 12929 4638
rect 12963 4604 12998 4638
rect 13032 4604 13067 4638
rect 13101 4604 13136 4638
rect 13170 4604 13205 4638
rect 13239 4604 13274 4638
rect 13308 4604 13343 4638
rect 13377 4604 13412 4638
rect 13446 4604 13481 4638
rect 13515 4604 13550 4638
rect 13584 4604 13619 4638
rect 13653 4604 13688 4638
rect 13722 4604 13757 4638
rect 13791 4604 13826 4638
rect 13860 4604 13895 4638
rect 13929 4604 13964 4638
rect 13998 4604 14033 4638
rect 14067 4604 14102 4638
rect 14136 4604 14171 4638
rect 14205 4604 14240 4638
rect 14274 4604 14309 4638
rect 14343 4604 14378 4638
rect 14412 4604 14447 4638
rect 14481 4604 14516 4638
rect 14550 4604 14585 4638
rect 14619 4604 14653 4638
rect 10410 4570 14653 4604
rect 482 4549 565 4570
rect 482 4515 497 4549
rect 531 4536 565 4549
rect 12363 4536 12397 4570
rect 12431 4536 12466 4570
rect 12500 4536 12535 4570
rect 12569 4536 12604 4570
rect 12638 4536 12673 4570
rect 12707 4536 12742 4570
rect 12776 4536 12811 4570
rect 12845 4536 12880 4570
rect 12914 4536 12949 4570
rect 12983 4536 13018 4570
rect 13052 4536 13087 4570
rect 13121 4536 13156 4570
rect 13190 4536 13225 4570
rect 13259 4536 13294 4570
rect 13328 4536 13363 4570
rect 13397 4536 13432 4570
rect 13466 4536 13501 4570
rect 13535 4536 13570 4570
rect 13604 4536 13639 4570
rect 13673 4536 13708 4570
rect 13742 4536 13777 4570
rect 13811 4536 13846 4570
rect 13880 4536 13915 4570
rect 13949 4536 13984 4570
rect 14018 4536 14053 4570
rect 14087 4536 14122 4570
rect 14156 4536 14191 4570
rect 14225 4536 14260 4570
rect 14294 4536 14329 4570
rect 14363 4536 14398 4570
rect 14432 4536 14467 4570
rect 14501 4536 14536 4570
rect 14570 4551 14653 4570
rect 531 4515 633 4536
rect 482 4498 633 4515
rect 482 4479 565 4498
rect 482 4445 497 4479
rect 531 4464 565 4479
rect 599 4468 633 4498
rect 12363 4502 14536 4536
rect 12363 4468 12398 4502
rect 12432 4468 12467 4502
rect 12501 4468 12536 4502
rect 12570 4468 12605 4502
rect 12639 4468 12674 4502
rect 12708 4468 12743 4502
rect 12777 4468 12812 4502
rect 12846 4468 12881 4502
rect 12915 4468 12950 4502
rect 12984 4468 13019 4502
rect 13053 4468 13088 4502
rect 13122 4468 13157 4502
rect 13191 4468 13226 4502
rect 13260 4468 13295 4502
rect 13329 4468 13364 4502
rect 13398 4468 13433 4502
rect 13467 4468 13502 4502
rect 13536 4468 13571 4502
rect 13605 4468 13640 4502
rect 13674 4468 13709 4502
rect 13743 4468 13778 4502
rect 13812 4468 13847 4502
rect 13881 4468 13916 4502
rect 13950 4468 13985 4502
rect 14019 4468 14054 4502
rect 14088 4468 14123 4502
rect 14157 4468 14192 4502
rect 14226 4468 14261 4502
rect 14295 4468 14330 4502
rect 14364 4468 14399 4502
rect 14433 4468 14468 4502
rect 599 4464 14468 4468
rect 531 4453 14468 4464
rect 531 4445 682 4453
rect 482 4429 682 4445
rect 482 4426 633 4429
rect 482 4409 565 4426
rect 482 4375 497 4409
rect 531 4392 565 4409
rect 599 4395 633 4426
rect 667 4395 682 4429
rect 599 4392 682 4395
rect 531 4375 682 4392
rect 482 4356 682 4375
rect 482 4354 633 4356
rect 482 4339 565 4354
rect 482 4305 497 4339
rect 531 4320 565 4339
rect 599 4322 633 4354
rect 667 4322 682 4356
rect 599 4320 682 4322
rect 531 4305 682 4320
rect 482 4283 682 4305
rect 482 4282 633 4283
rect 482 4269 565 4282
rect 482 4235 497 4269
rect 531 4248 565 4269
rect 599 4249 633 4282
rect 667 4249 682 4283
rect 599 4248 682 4249
rect 531 4235 682 4248
rect 482 4211 682 4235
rect 482 4210 633 4211
rect 482 4199 565 4210
rect 482 4165 497 4199
rect 531 4176 565 4199
rect 599 4177 633 4210
rect 667 4177 682 4211
rect 599 4176 682 4177
rect 531 4165 682 4176
rect 482 4152 682 4165
rect 14453 4152 14468 4453
rect 482 4139 708 4152
rect 482 4138 633 4139
rect 482 4129 565 4138
rect 482 4095 497 4129
rect 531 4104 565 4129
rect 599 4105 633 4138
rect 667 4105 708 4139
rect 599 4104 708 4105
rect 531 4095 708 4104
rect 482 4067 708 4095
rect 482 4066 633 4067
rect 482 4059 565 4066
rect 482 4025 497 4059
rect 531 4032 565 4059
rect 599 4033 633 4066
rect 667 4033 708 4067
rect 599 4032 708 4033
rect 531 4025 708 4032
rect 482 3995 708 4025
rect 482 3994 633 3995
rect 482 3989 565 3994
rect 482 3955 497 3989
rect 531 3960 565 3989
rect 599 3961 633 3994
rect 667 3961 708 3995
rect 599 3960 708 3961
rect 531 3955 708 3960
rect 482 3923 708 3955
rect 482 3922 633 3923
rect 482 3920 565 3922
rect 482 3886 497 3920
rect 531 3888 565 3920
rect 599 3889 633 3922
rect 667 3889 708 3923
rect 599 3888 708 3889
rect 531 3886 708 3888
rect 482 3851 708 3886
rect 482 3817 497 3851
rect 531 3817 565 3851
rect 599 3817 633 3851
rect 667 3817 708 3851
rect 482 3749 708 3817
rect 482 3715 497 3749
rect 531 3715 565 3749
rect 599 3715 633 3749
rect 667 3715 708 3749
rect 482 3680 708 3715
rect 482 3646 497 3680
rect 531 3646 565 3680
rect 599 3646 633 3680
rect 667 3646 708 3680
rect 482 3611 708 3646
rect 482 3577 497 3611
rect 531 3577 565 3611
rect 599 3577 633 3611
rect 667 3577 708 3611
rect 482 3542 708 3577
rect 482 3508 497 3542
rect 531 3508 565 3542
rect 599 3508 633 3542
rect 667 3508 708 3542
rect 482 3473 708 3508
rect 482 3439 497 3473
rect 531 3439 565 3473
rect 599 3439 633 3473
rect 667 3439 708 3473
rect 482 3404 708 3439
rect 482 3370 497 3404
rect 531 3370 565 3404
rect 599 3370 633 3404
rect 667 3370 708 3404
rect 482 3335 708 3370
rect 482 3301 497 3335
rect 531 3301 565 3335
rect 599 3301 633 3335
rect 667 3301 708 3335
rect 482 3266 708 3301
rect 482 3232 497 3266
rect 531 3232 565 3266
rect 599 3232 633 3266
rect 667 3232 708 3266
rect 482 3197 708 3232
rect 482 3163 497 3197
rect 531 3163 565 3197
rect 599 3163 633 3197
rect 667 3163 708 3197
rect 482 3152 708 3163
rect 14427 3992 14468 4152
rect 14427 3957 14536 3992
rect 14427 3923 14468 3957
rect 14502 3924 14536 3957
rect 14502 3923 14604 3924
rect 14427 3905 14604 3923
rect 14638 3905 14653 4551
rect 14427 3889 14653 3905
rect 14427 3888 14536 3889
rect 14427 3854 14468 3888
rect 14502 3855 14536 3888
rect 14570 3871 14653 3889
rect 14570 3855 14604 3871
rect 14502 3854 14604 3855
rect 14427 3837 14604 3854
rect 14638 3837 14653 3871
rect 14427 3820 14653 3837
rect 14427 3819 14536 3820
rect 14427 3785 14468 3819
rect 14502 3786 14536 3819
rect 14570 3803 14653 3820
rect 14570 3786 14604 3803
rect 14502 3785 14604 3786
rect 14427 3769 14604 3785
rect 14638 3769 14653 3803
rect 14427 3751 14653 3769
rect 14427 3750 14536 3751
rect 14427 3716 14468 3750
rect 14502 3717 14536 3750
rect 14570 3735 14653 3751
rect 14570 3717 14604 3735
rect 14502 3716 14604 3717
rect 14427 3701 14604 3716
rect 14638 3701 14653 3735
rect 14427 3682 14653 3701
rect 14427 3681 14536 3682
rect 14427 3647 14468 3681
rect 14502 3648 14536 3681
rect 14570 3667 14653 3682
rect 14570 3648 14604 3667
rect 14502 3647 14604 3648
rect 14427 3633 14604 3647
rect 14638 3633 14653 3667
rect 14427 3613 14653 3633
rect 14427 3612 14536 3613
rect 14427 3578 14468 3612
rect 14502 3579 14536 3612
rect 14570 3599 14653 3613
rect 14570 3579 14604 3599
rect 14502 3578 14604 3579
rect 14427 3565 14604 3578
rect 14638 3565 14653 3599
rect 14427 3544 14653 3565
rect 14427 3543 14536 3544
rect 14427 3509 14468 3543
rect 14502 3510 14536 3543
rect 14570 3531 14653 3544
rect 14570 3510 14604 3531
rect 14502 3509 14604 3510
rect 14427 3497 14604 3509
rect 14638 3497 14653 3531
rect 14427 3475 14653 3497
rect 14427 3474 14536 3475
rect 14427 3440 14468 3474
rect 14502 3441 14536 3474
rect 14570 3463 14653 3475
rect 14570 3441 14604 3463
rect 14502 3440 14604 3441
rect 14427 3429 14604 3440
rect 14638 3429 14653 3463
rect 14427 3406 14653 3429
rect 14427 3405 14536 3406
rect 14427 3371 14468 3405
rect 14502 3372 14536 3405
rect 14570 3395 14653 3406
rect 14570 3372 14604 3395
rect 14502 3371 14604 3372
rect 14427 3361 14604 3371
rect 14638 3361 14653 3395
rect 14427 3337 14653 3361
rect 14427 3336 14536 3337
rect 14427 3302 14468 3336
rect 14502 3303 14536 3336
rect 14570 3327 14653 3337
rect 14570 3303 14604 3327
rect 14502 3302 14604 3303
rect 14427 3293 14604 3302
rect 14638 3293 14653 3327
rect 14427 3268 14653 3293
rect 14427 3267 14536 3268
rect 14427 3233 14468 3267
rect 14502 3234 14536 3267
rect 14570 3259 14653 3268
rect 14570 3234 14604 3259
rect 14502 3233 14604 3234
rect 14427 3225 14604 3233
rect 14638 3225 14653 3259
rect 14427 3199 14653 3225
rect 14427 3198 14536 3199
rect 14427 3164 14468 3198
rect 14502 3165 14536 3198
rect 14570 3191 14653 3199
rect 14570 3165 14604 3191
rect 14502 3164 14604 3165
rect 14427 3157 14604 3164
rect 14638 3157 14653 3191
rect 14427 3152 14653 3157
rect 482 3128 682 3152
rect 482 3094 497 3128
rect 531 3094 565 3128
rect 599 3094 633 3128
rect 667 3094 682 3128
rect 14453 3130 14653 3152
rect 14453 3129 14536 3130
rect 482 3059 682 3094
rect 482 3025 497 3059
rect 531 3025 565 3059
rect 599 3025 633 3059
rect 667 3025 682 3059
rect 482 2990 682 3025
rect 482 2956 497 2990
rect 531 2956 565 2990
rect 599 2956 633 2990
rect 667 2956 682 2990
rect 482 2921 682 2956
rect 482 2887 497 2921
rect 531 2887 565 2921
rect 599 2887 633 2921
rect 667 2887 682 2921
rect 482 2852 682 2887
rect 482 2818 497 2852
rect 531 2818 565 2852
rect 599 2818 633 2852
rect 667 2818 682 2852
rect 482 2783 682 2818
rect 482 2749 497 2783
rect 531 2749 565 2783
rect 599 2749 633 2783
rect 667 2749 682 2783
rect 482 2714 682 2749
rect 482 2680 497 2714
rect 531 2680 565 2714
rect 599 2680 633 2714
rect 667 2680 682 2714
rect 482 2645 682 2680
rect 482 2611 497 2645
rect 531 2611 565 2645
rect 599 2611 633 2645
rect 667 2611 682 2645
rect 482 2576 682 2611
rect 1541 3044 1763 3078
rect 1541 3010 1601 3044
rect 1635 3010 1669 3044
rect 1703 3010 1763 3044
rect 1541 2974 1763 3010
rect 1541 2940 1601 2974
rect 1635 2940 1669 2974
rect 1703 2940 1763 2974
rect 1541 2904 1763 2940
rect 1541 2870 1601 2904
rect 1635 2870 1669 2904
rect 1703 2870 1763 2904
rect 1541 2834 1763 2870
rect 1541 2800 1601 2834
rect 1635 2800 1669 2834
rect 1703 2800 1763 2834
rect 1541 2764 1763 2800
rect 1541 2730 1601 2764
rect 1635 2730 1669 2764
rect 1703 2730 1763 2764
rect 1541 2694 1763 2730
rect 1541 2660 1601 2694
rect 1635 2660 1669 2694
rect 1703 2660 1763 2694
rect 1541 2626 1763 2660
rect 2533 3044 2755 3078
rect 2533 3010 2593 3044
rect 2627 3010 2661 3044
rect 2695 3010 2755 3044
rect 2533 2974 2755 3010
rect 2533 2940 2593 2974
rect 2627 2940 2661 2974
rect 2695 2940 2755 2974
rect 2533 2904 2755 2940
rect 2533 2870 2593 2904
rect 2627 2870 2661 2904
rect 2695 2870 2755 2904
rect 2533 2834 2755 2870
rect 2533 2800 2593 2834
rect 2627 2800 2661 2834
rect 2695 2800 2755 2834
rect 2533 2764 2755 2800
rect 2533 2730 2593 2764
rect 2627 2730 2661 2764
rect 2695 2730 2755 2764
rect 2533 2694 2755 2730
rect 2533 2660 2593 2694
rect 2627 2660 2661 2694
rect 2695 2660 2755 2694
rect 2533 2626 2755 2660
rect 3525 3044 3747 3078
rect 3525 3010 3585 3044
rect 3619 3010 3653 3044
rect 3687 3010 3747 3044
rect 3525 2974 3747 3010
rect 3525 2940 3585 2974
rect 3619 2940 3653 2974
rect 3687 2940 3747 2974
rect 3525 2904 3747 2940
rect 3525 2870 3585 2904
rect 3619 2870 3653 2904
rect 3687 2870 3747 2904
rect 3525 2834 3747 2870
rect 3525 2800 3585 2834
rect 3619 2800 3653 2834
rect 3687 2800 3747 2834
rect 3525 2764 3747 2800
rect 3525 2730 3585 2764
rect 3619 2730 3653 2764
rect 3687 2730 3747 2764
rect 3525 2694 3747 2730
rect 3525 2660 3585 2694
rect 3619 2660 3653 2694
rect 3687 2660 3747 2694
rect 3525 2626 3747 2660
rect 4517 3044 4739 3078
rect 4517 3010 4577 3044
rect 4611 3010 4645 3044
rect 4679 3010 4739 3044
rect 4517 2974 4739 3010
rect 4517 2940 4577 2974
rect 4611 2940 4645 2974
rect 4679 2940 4739 2974
rect 4517 2904 4739 2940
rect 4517 2870 4577 2904
rect 4611 2870 4645 2904
rect 4679 2870 4739 2904
rect 4517 2834 4739 2870
rect 4517 2800 4577 2834
rect 4611 2800 4645 2834
rect 4679 2800 4739 2834
rect 4517 2764 4739 2800
rect 4517 2730 4577 2764
rect 4611 2730 4645 2764
rect 4679 2730 4739 2764
rect 4517 2694 4739 2730
rect 4517 2660 4577 2694
rect 4611 2660 4645 2694
rect 4679 2660 4739 2694
rect 4517 2626 4739 2660
rect 5509 3044 5731 3078
rect 5509 3010 5569 3044
rect 5603 3010 5637 3044
rect 5671 3010 5731 3044
rect 5509 2974 5731 3010
rect 5509 2940 5569 2974
rect 5603 2940 5637 2974
rect 5671 2940 5731 2974
rect 5509 2904 5731 2940
rect 5509 2870 5569 2904
rect 5603 2870 5637 2904
rect 5671 2870 5731 2904
rect 5509 2834 5731 2870
rect 5509 2800 5569 2834
rect 5603 2800 5637 2834
rect 5671 2800 5731 2834
rect 5509 2764 5731 2800
rect 5509 2730 5569 2764
rect 5603 2730 5637 2764
rect 5671 2730 5731 2764
rect 5509 2694 5731 2730
rect 5509 2660 5569 2694
rect 5603 2660 5637 2694
rect 5671 2660 5731 2694
rect 5509 2626 5731 2660
rect 6501 3044 6723 3078
rect 6501 3010 6561 3044
rect 6595 3010 6629 3044
rect 6663 3010 6723 3044
rect 6501 2974 6723 3010
rect 6501 2940 6561 2974
rect 6595 2940 6629 2974
rect 6663 2940 6723 2974
rect 6501 2904 6723 2940
rect 6501 2870 6561 2904
rect 6595 2870 6629 2904
rect 6663 2870 6723 2904
rect 6501 2834 6723 2870
rect 6501 2800 6561 2834
rect 6595 2800 6629 2834
rect 6663 2800 6723 2834
rect 6501 2764 6723 2800
rect 6501 2730 6561 2764
rect 6595 2730 6629 2764
rect 6663 2730 6723 2764
rect 6501 2694 6723 2730
rect 6501 2660 6561 2694
rect 6595 2660 6629 2694
rect 6663 2660 6723 2694
rect 6501 2626 6723 2660
rect 7493 3044 7715 3078
rect 7493 3010 7553 3044
rect 7587 3010 7621 3044
rect 7655 3010 7715 3044
rect 7493 2974 7715 3010
rect 7493 2940 7553 2974
rect 7587 2940 7621 2974
rect 7655 2940 7715 2974
rect 7493 2904 7715 2940
rect 7493 2870 7553 2904
rect 7587 2870 7621 2904
rect 7655 2870 7715 2904
rect 7493 2834 7715 2870
rect 7493 2800 7553 2834
rect 7587 2800 7621 2834
rect 7655 2800 7715 2834
rect 7493 2764 7715 2800
rect 7493 2730 7553 2764
rect 7587 2730 7621 2764
rect 7655 2730 7715 2764
rect 7493 2694 7715 2730
rect 7493 2660 7553 2694
rect 7587 2660 7621 2694
rect 7655 2660 7715 2694
rect 7493 2626 7715 2660
rect 8485 3044 8707 3078
rect 8485 3010 8545 3044
rect 8579 3010 8613 3044
rect 8647 3010 8707 3044
rect 8485 2974 8707 3010
rect 8485 2940 8545 2974
rect 8579 2940 8613 2974
rect 8647 2940 8707 2974
rect 8485 2904 8707 2940
rect 8485 2870 8545 2904
rect 8579 2870 8613 2904
rect 8647 2870 8707 2904
rect 8485 2834 8707 2870
rect 8485 2800 8545 2834
rect 8579 2800 8613 2834
rect 8647 2800 8707 2834
rect 8485 2764 8707 2800
rect 8485 2730 8545 2764
rect 8579 2730 8613 2764
rect 8647 2730 8707 2764
rect 8485 2694 8707 2730
rect 8485 2660 8545 2694
rect 8579 2660 8613 2694
rect 8647 2660 8707 2694
rect 8485 2626 8707 2660
rect 9477 3044 9699 3078
rect 9477 3010 9537 3044
rect 9571 3010 9605 3044
rect 9639 3010 9699 3044
rect 9477 2974 9699 3010
rect 9477 2940 9537 2974
rect 9571 2940 9605 2974
rect 9639 2940 9699 2974
rect 9477 2904 9699 2940
rect 9477 2870 9537 2904
rect 9571 2870 9605 2904
rect 9639 2870 9699 2904
rect 9477 2834 9699 2870
rect 9477 2800 9537 2834
rect 9571 2800 9605 2834
rect 9639 2800 9699 2834
rect 9477 2764 9699 2800
rect 9477 2730 9537 2764
rect 9571 2730 9605 2764
rect 9639 2730 9699 2764
rect 9477 2694 9699 2730
rect 9477 2660 9537 2694
rect 9571 2660 9605 2694
rect 9639 2660 9699 2694
rect 9477 2626 9699 2660
rect 10469 3044 10691 3078
rect 10469 3010 10529 3044
rect 10563 3010 10597 3044
rect 10631 3010 10691 3044
rect 10469 2974 10691 3010
rect 10469 2940 10529 2974
rect 10563 2940 10597 2974
rect 10631 2940 10691 2974
rect 10469 2904 10691 2940
rect 10469 2870 10529 2904
rect 10563 2870 10597 2904
rect 10631 2870 10691 2904
rect 10469 2834 10691 2870
rect 10469 2800 10529 2834
rect 10563 2800 10597 2834
rect 10631 2800 10691 2834
rect 10469 2764 10691 2800
rect 10469 2730 10529 2764
rect 10563 2730 10597 2764
rect 10631 2730 10691 2764
rect 10469 2694 10691 2730
rect 10469 2660 10529 2694
rect 10563 2660 10597 2694
rect 10631 2660 10691 2694
rect 10469 2626 10691 2660
rect 11461 3044 11683 3078
rect 11461 3010 11521 3044
rect 11555 3010 11589 3044
rect 11623 3010 11683 3044
rect 11461 2974 11683 3010
rect 11461 2940 11521 2974
rect 11555 2940 11589 2974
rect 11623 2940 11683 2974
rect 11461 2904 11683 2940
rect 11461 2870 11521 2904
rect 11555 2870 11589 2904
rect 11623 2870 11683 2904
rect 11461 2834 11683 2870
rect 11461 2800 11521 2834
rect 11555 2800 11589 2834
rect 11623 2800 11683 2834
rect 11461 2764 11683 2800
rect 11461 2730 11521 2764
rect 11555 2730 11589 2764
rect 11623 2730 11683 2764
rect 11461 2694 11683 2730
rect 11461 2660 11521 2694
rect 11555 2660 11589 2694
rect 11623 2660 11683 2694
rect 11461 2626 11683 2660
rect 12453 3044 12675 3078
rect 12453 3010 12513 3044
rect 12547 3010 12581 3044
rect 12615 3010 12675 3044
rect 12453 2974 12675 3010
rect 12453 2940 12513 2974
rect 12547 2940 12581 2974
rect 12615 2940 12675 2974
rect 12453 2904 12675 2940
rect 12453 2870 12513 2904
rect 12547 2870 12581 2904
rect 12615 2870 12675 2904
rect 12453 2834 12675 2870
rect 12453 2800 12513 2834
rect 12547 2800 12581 2834
rect 12615 2800 12675 2834
rect 12453 2764 12675 2800
rect 12453 2730 12513 2764
rect 12547 2730 12581 2764
rect 12615 2730 12675 2764
rect 12453 2694 12675 2730
rect 12453 2660 12513 2694
rect 12547 2660 12581 2694
rect 12615 2660 12675 2694
rect 12453 2626 12675 2660
rect 13445 3044 13667 3078
rect 13445 3010 13505 3044
rect 13539 3010 13573 3044
rect 13607 3010 13667 3044
rect 13445 2974 13667 3010
rect 13445 2940 13505 2974
rect 13539 2940 13573 2974
rect 13607 2940 13667 2974
rect 13445 2904 13667 2940
rect 13445 2870 13505 2904
rect 13539 2870 13573 2904
rect 13607 2870 13667 2904
rect 13445 2834 13667 2870
rect 13445 2800 13505 2834
rect 13539 2800 13573 2834
rect 13607 2800 13667 2834
rect 13445 2764 13667 2800
rect 13445 2730 13505 2764
rect 13539 2730 13573 2764
rect 13607 2730 13667 2764
rect 13445 2694 13667 2730
rect 13445 2660 13505 2694
rect 13539 2660 13573 2694
rect 13607 2660 13667 2694
rect 13445 2626 13667 2660
rect 14453 3095 14468 3129
rect 14502 3096 14536 3129
rect 14570 3123 14653 3130
rect 14570 3096 14604 3123
rect 14502 3095 14604 3096
rect 14453 3089 14604 3095
rect 14638 3089 14653 3123
rect 14453 3061 14653 3089
rect 14453 3060 14536 3061
rect 14453 3026 14468 3060
rect 14502 3027 14536 3060
rect 14570 3055 14653 3061
rect 14570 3027 14604 3055
rect 14502 3026 14604 3027
rect 14453 3021 14604 3026
rect 14638 3021 14653 3055
rect 14453 2992 14653 3021
rect 14453 2991 14536 2992
rect 14453 2957 14468 2991
rect 14502 2958 14536 2991
rect 14570 2987 14653 2992
rect 14570 2958 14604 2987
rect 14502 2957 14604 2958
rect 14453 2953 14604 2957
rect 14638 2953 14653 2987
rect 14453 2923 14653 2953
rect 14453 2922 14536 2923
rect 14453 2888 14468 2922
rect 14502 2889 14536 2922
rect 14570 2919 14653 2923
rect 14570 2889 14604 2919
rect 14502 2888 14604 2889
rect 14453 2885 14604 2888
rect 14638 2885 14653 2919
rect 14453 2854 14653 2885
rect 14453 2853 14536 2854
rect 14453 2819 14468 2853
rect 14502 2820 14536 2853
rect 14570 2851 14653 2854
rect 14570 2820 14604 2851
rect 14502 2819 14604 2820
rect 14453 2817 14604 2819
rect 14638 2817 14653 2851
rect 14453 2785 14653 2817
rect 14453 2784 14536 2785
rect 14453 2750 14468 2784
rect 14502 2751 14536 2784
rect 14570 2783 14653 2785
rect 14570 2751 14604 2783
rect 14502 2750 14604 2751
rect 14453 2749 14604 2750
rect 14638 2749 14653 2783
rect 14453 2716 14653 2749
rect 14453 2715 14536 2716
rect 14453 2681 14468 2715
rect 14502 2682 14536 2715
rect 14570 2715 14653 2716
rect 14570 2682 14604 2715
rect 14502 2681 14604 2682
rect 14638 2681 14653 2715
rect 14453 2647 14653 2681
rect 14453 2646 14536 2647
rect 14453 2612 14468 2646
rect 14502 2613 14536 2646
rect 14570 2613 14604 2647
rect 14638 2613 14653 2647
rect 14502 2612 14653 2613
rect 482 2542 497 2576
rect 531 2542 565 2576
rect 599 2542 633 2576
rect 667 2552 682 2576
rect 14453 2579 14653 2612
rect 14453 2578 14604 2579
rect 14453 2577 14536 2578
rect 14453 2552 14468 2577
rect 667 2542 708 2552
rect 482 2507 708 2542
rect 482 2473 497 2507
rect 531 2473 565 2507
rect 599 2473 633 2507
rect 667 2473 708 2507
rect 482 2438 708 2473
rect 482 2404 497 2438
rect 531 2404 565 2438
rect 599 2404 633 2438
rect 667 2404 708 2438
rect 482 2369 708 2404
rect 482 2335 497 2369
rect 531 2335 565 2369
rect 599 2335 633 2369
rect 667 2335 708 2369
rect 482 2300 708 2335
rect 482 2266 497 2300
rect 531 2266 565 2300
rect 599 2266 633 2300
rect 667 2266 708 2300
rect 482 2231 708 2266
rect 482 2197 497 2231
rect 531 2197 565 2231
rect 599 2197 633 2231
rect 667 2197 708 2231
rect 482 2163 708 2197
rect 482 2129 497 2163
rect 531 2162 708 2163
rect 531 2129 565 2162
rect 482 2128 565 2129
rect 599 2128 633 2162
rect 667 2128 708 2162
rect 482 2095 708 2128
rect 482 2061 497 2095
rect 531 2093 708 2095
rect 531 2061 565 2093
rect 482 2059 565 2061
rect 599 2059 633 2093
rect 667 2059 708 2093
rect 482 2027 708 2059
rect 482 1993 497 2027
rect 531 2024 708 2027
rect 531 1993 565 2024
rect 482 1990 565 1993
rect 599 1990 633 2024
rect 667 1990 708 2024
rect 482 1959 708 1990
rect 482 1925 497 1959
rect 531 1955 708 1959
rect 531 1925 565 1955
rect 482 1921 565 1925
rect 599 1921 633 1955
rect 667 1921 708 1955
rect 482 1891 708 1921
rect 482 1857 497 1891
rect 531 1886 708 1891
rect 531 1857 565 1886
rect 482 1852 565 1857
rect 599 1852 633 1886
rect 667 1852 708 1886
rect 482 1823 708 1852
rect 482 1789 497 1823
rect 531 1817 708 1823
rect 531 1789 565 1817
rect 482 1783 565 1789
rect 599 1783 633 1817
rect 667 1783 708 1817
rect 482 1755 708 1783
rect 482 1721 497 1755
rect 531 1748 708 1755
rect 531 1721 565 1748
rect 482 1714 565 1721
rect 599 1714 633 1748
rect 667 1714 708 1748
rect 482 1687 708 1714
rect 482 1653 497 1687
rect 531 1679 708 1687
rect 531 1653 565 1679
rect 482 1645 565 1653
rect 599 1645 633 1679
rect 667 1645 708 1679
rect 482 1619 708 1645
rect 482 1585 497 1619
rect 531 1610 708 1619
rect 531 1585 565 1610
rect 482 1576 565 1585
rect 599 1576 633 1610
rect 667 1576 708 1610
rect 482 1552 708 1576
rect 14427 2543 14468 2552
rect 14502 2544 14536 2577
rect 14570 2545 14604 2578
rect 14638 2545 14653 2579
rect 14570 2544 14653 2545
rect 14502 2543 14653 2544
rect 14427 2511 14653 2543
rect 14427 2509 14604 2511
rect 14427 2508 14536 2509
rect 14427 2474 14468 2508
rect 14502 2475 14536 2508
rect 14570 2477 14604 2509
rect 14638 2477 14653 2511
rect 14570 2475 14653 2477
rect 14502 2474 14653 2475
rect 14427 2443 14653 2474
rect 14427 2440 14604 2443
rect 14427 2439 14536 2440
rect 14427 2405 14468 2439
rect 14502 2406 14536 2439
rect 14570 2409 14604 2440
rect 14638 2409 14653 2443
rect 14570 2406 14653 2409
rect 14502 2405 14653 2406
rect 14427 2375 14653 2405
rect 14427 2371 14604 2375
rect 14427 2370 14536 2371
rect 14427 2336 14468 2370
rect 14502 2337 14536 2370
rect 14570 2341 14604 2371
rect 14638 2341 14653 2375
rect 14570 2337 14653 2341
rect 14502 2336 14653 2337
rect 14427 2307 14653 2336
rect 14427 2302 14604 2307
rect 14427 2301 14536 2302
rect 14427 2267 14468 2301
rect 14502 2268 14536 2301
rect 14570 2273 14604 2302
rect 14638 2273 14653 2307
rect 14570 2268 14653 2273
rect 14502 2267 14653 2268
rect 14427 2239 14653 2267
rect 14427 2233 14604 2239
rect 14427 2232 14536 2233
rect 14427 2198 14468 2232
rect 14502 2199 14536 2232
rect 14570 2205 14604 2233
rect 14638 2205 14653 2239
rect 14570 2199 14653 2205
rect 14502 2198 14653 2199
rect 14427 2171 14653 2198
rect 14427 2164 14604 2171
rect 14427 2163 14536 2164
rect 14427 2129 14468 2163
rect 14502 2130 14536 2163
rect 14570 2137 14604 2164
rect 14638 2137 14653 2171
rect 14570 2130 14653 2137
rect 14502 2129 14653 2130
rect 14427 2103 14653 2129
rect 14427 2095 14604 2103
rect 14427 2094 14536 2095
rect 14427 2060 14468 2094
rect 14502 2061 14536 2094
rect 14570 2069 14604 2095
rect 14638 2069 14653 2103
rect 14570 2061 14653 2069
rect 14502 2060 14653 2061
rect 14427 2035 14653 2060
rect 14427 2026 14604 2035
rect 14427 2025 14536 2026
rect 14427 1991 14468 2025
rect 14502 1992 14536 2025
rect 14570 2001 14604 2026
rect 14638 2001 14653 2035
rect 14570 1992 14653 2001
rect 14502 1991 14653 1992
rect 14427 1967 14653 1991
rect 14427 1957 14604 1967
rect 14427 1956 14536 1957
rect 14427 1922 14468 1956
rect 14502 1923 14536 1956
rect 14570 1933 14604 1957
rect 14638 1933 14653 1967
rect 14570 1923 14653 1933
rect 14502 1922 14653 1923
rect 14427 1899 14653 1922
rect 14427 1888 14604 1899
rect 14427 1887 14536 1888
rect 14427 1853 14468 1887
rect 14502 1854 14536 1887
rect 14570 1865 14604 1888
rect 14638 1865 14653 1899
rect 14570 1854 14653 1865
rect 14502 1853 14653 1854
rect 14427 1831 14653 1853
rect 14427 1819 14604 1831
rect 14427 1818 14536 1819
rect 14427 1784 14468 1818
rect 14502 1785 14536 1818
rect 14570 1797 14604 1819
rect 14638 1797 14653 1831
rect 14570 1785 14653 1797
rect 14502 1784 14653 1785
rect 14427 1763 14653 1784
rect 14427 1750 14604 1763
rect 14427 1749 14536 1750
rect 14427 1715 14468 1749
rect 14502 1716 14536 1749
rect 14570 1729 14604 1750
rect 14638 1729 14653 1763
rect 14570 1716 14653 1729
rect 14502 1715 14653 1716
rect 14427 1695 14653 1715
rect 14427 1681 14604 1695
rect 14427 1680 14536 1681
rect 14427 1646 14468 1680
rect 14502 1647 14536 1680
rect 14570 1661 14604 1681
rect 14638 1661 14653 1695
rect 14570 1647 14653 1661
rect 14502 1646 14653 1647
rect 14427 1627 14653 1646
rect 14427 1612 14604 1627
rect 14427 1611 14536 1612
rect 14427 1577 14468 1611
rect 14502 1578 14536 1611
rect 14570 1593 14604 1612
rect 14638 1593 14653 1627
rect 14570 1578 14653 1593
rect 14502 1577 14653 1578
rect 14427 1559 14653 1577
rect 14427 1552 14604 1559
rect 482 1551 682 1552
rect 482 1517 497 1551
rect 531 1541 682 1551
rect 531 1517 565 1541
rect 482 1507 565 1517
rect 599 1507 633 1541
rect 667 1507 682 1541
rect 14453 1543 14604 1552
rect 14453 1542 14536 1543
rect 482 1483 682 1507
rect 482 1449 497 1483
rect 531 1472 682 1483
rect 531 1449 565 1472
rect 482 1438 565 1449
rect 599 1438 633 1472
rect 667 1438 682 1472
rect 482 1415 682 1438
rect 482 1381 497 1415
rect 531 1403 682 1415
rect 531 1381 565 1403
rect 482 1369 565 1381
rect 599 1369 633 1403
rect 667 1369 682 1403
rect 14453 1508 14468 1542
rect 14502 1509 14536 1542
rect 14570 1525 14604 1543
rect 14638 1525 14653 1559
rect 14570 1509 14653 1525
rect 14502 1508 14653 1509
rect 14453 1491 14653 1508
rect 14453 1474 14604 1491
rect 14453 1473 14536 1474
rect 14453 1439 14468 1473
rect 14502 1440 14536 1473
rect 14570 1457 14604 1474
rect 14638 1457 14653 1491
rect 14570 1440 14653 1457
rect 14502 1439 14653 1440
rect 14453 1423 14653 1439
rect 14453 1405 14604 1423
rect 14453 1404 14536 1405
rect 482 1347 682 1369
rect 482 1313 497 1347
rect 531 1334 682 1347
rect 531 1313 565 1334
rect 482 1300 565 1313
rect 599 1300 633 1334
rect 667 1300 682 1334
rect 482 1279 682 1300
rect 482 1245 497 1279
rect 531 1265 682 1279
rect 531 1245 565 1265
rect 482 1231 565 1245
rect 599 1231 633 1265
rect 667 1231 682 1265
rect 482 1211 682 1231
rect 482 1177 497 1211
rect 531 1196 682 1211
rect 531 1177 565 1196
rect 482 1162 565 1177
rect 599 1162 633 1196
rect 667 1162 682 1196
rect 482 1143 682 1162
rect 482 1109 497 1143
rect 531 1127 682 1143
rect 531 1109 565 1127
rect 482 1093 565 1109
rect 599 1093 633 1127
rect 667 1093 682 1127
rect 482 1075 682 1093
rect 482 1041 497 1075
rect 531 1058 682 1075
rect 531 1041 565 1058
rect 482 1024 565 1041
rect 599 1024 633 1058
rect 667 1024 682 1058
rect 482 1007 682 1024
rect 482 973 497 1007
rect 531 989 682 1007
rect 531 973 565 989
rect 482 955 565 973
rect 599 955 633 989
rect 667 955 682 989
rect 482 939 682 955
rect 482 769 497 939
rect 531 920 682 939
rect 667 867 682 920
rect 14453 1370 14468 1404
rect 14502 1371 14536 1404
rect 14570 1389 14604 1405
rect 14638 1389 14653 1423
rect 14570 1371 14653 1389
rect 14502 1370 14653 1371
rect 14453 1355 14653 1370
rect 14453 1336 14604 1355
rect 14453 1335 14536 1336
rect 14453 1301 14468 1335
rect 14502 1302 14536 1335
rect 14570 1321 14604 1336
rect 14638 1321 14653 1355
rect 14570 1302 14653 1321
rect 14502 1301 14653 1302
rect 14453 1287 14653 1301
rect 14453 1267 14604 1287
rect 14453 1266 14536 1267
rect 14453 1232 14468 1266
rect 14502 1233 14536 1266
rect 14570 1253 14604 1267
rect 14638 1253 14653 1287
rect 14570 1233 14653 1253
rect 14502 1232 14653 1233
rect 14453 1218 14653 1232
rect 14453 1198 14604 1218
rect 14453 1197 14536 1198
rect 14453 1163 14468 1197
rect 14502 1164 14536 1197
rect 14570 1184 14604 1198
rect 14638 1184 14653 1218
rect 14570 1164 14653 1184
rect 14502 1163 14653 1164
rect 14453 1149 14653 1163
rect 14453 1129 14604 1149
rect 14453 1128 14536 1129
rect 14453 1094 14468 1128
rect 14502 1095 14536 1128
rect 14570 1115 14604 1129
rect 14638 1115 14653 1149
rect 14570 1095 14653 1115
rect 14502 1094 14653 1095
rect 14453 1080 14653 1094
rect 14453 1060 14604 1080
rect 14453 1059 14536 1060
rect 14453 1025 14468 1059
rect 14502 1026 14536 1059
rect 14570 1046 14604 1060
rect 14638 1046 14653 1080
rect 14570 1026 14653 1046
rect 14502 1025 14653 1026
rect 14453 1011 14653 1025
rect 14453 991 14604 1011
rect 14453 990 14536 991
rect 14453 956 14468 990
rect 14502 957 14536 990
rect 14570 977 14604 991
rect 14638 977 14653 1011
rect 14570 957 14653 977
rect 14502 956 14653 957
rect 14453 942 14653 956
rect 14453 922 14604 942
rect 14453 921 14536 922
rect 14453 887 14468 921
rect 14502 888 14536 921
rect 14570 908 14604 922
rect 14638 908 14653 942
rect 14570 888 14653 908
rect 14502 887 14653 888
rect 14453 873 14653 887
rect 14453 867 14604 873
rect 667 853 14604 867
rect 667 852 14536 853
rect 667 818 702 852
rect 736 818 771 852
rect 805 818 840 852
rect 874 818 909 852
rect 943 818 978 852
rect 1012 818 1047 852
rect 1081 818 1116 852
rect 1150 818 1185 852
rect 1219 818 1254 852
rect 1288 818 1323 852
rect 1357 818 1392 852
rect 1426 818 1461 852
rect 1495 818 1530 852
rect 1564 818 1599 852
rect 1633 818 1668 852
rect 1702 818 1737 852
rect 1771 818 1806 852
rect 1840 818 1875 852
rect 1909 818 1944 852
rect 1978 818 2013 852
rect 2047 818 2082 852
rect 2116 818 2151 852
rect 2185 818 2220 852
rect 2254 818 2289 852
rect 2323 818 2358 852
rect 2392 818 2427 852
rect 2461 818 2496 852
rect 2530 818 2565 852
rect 2599 818 2634 852
rect 2668 818 2703 852
rect 2737 818 2772 852
rect 599 784 2772 818
rect 14502 819 14536 852
rect 14570 839 14604 853
rect 14638 839 14653 873
rect 14570 819 14653 839
rect 14502 804 14653 819
rect 14502 784 14604 804
rect 482 750 565 769
rect 599 750 634 784
rect 668 750 703 784
rect 737 750 772 784
rect 806 750 841 784
rect 875 750 910 784
rect 944 750 979 784
rect 1013 750 1048 784
rect 1082 750 1117 784
rect 1151 750 1186 784
rect 1220 750 1255 784
rect 1289 750 1324 784
rect 1358 750 1393 784
rect 1427 750 1462 784
rect 1496 750 1531 784
rect 1565 750 1600 784
rect 1634 750 1669 784
rect 1703 750 1738 784
rect 1772 750 1807 784
rect 1841 750 1876 784
rect 1910 750 1945 784
rect 1979 750 2014 784
rect 2048 750 2083 784
rect 2117 750 2152 784
rect 2186 750 2221 784
rect 2255 750 2290 784
rect 2324 750 2359 784
rect 2393 750 2428 784
rect 2462 750 2497 784
rect 2531 750 2566 784
rect 2600 750 2635 784
rect 2669 750 2704 784
rect 2738 750 2772 784
rect 14570 770 14604 784
rect 14638 770 14653 804
rect 14570 750 14653 770
rect 482 716 4725 750
rect 482 682 516 716
rect 550 682 585 716
rect 619 682 654 716
rect 688 682 723 716
rect 757 682 792 716
rect 826 682 861 716
rect 895 682 930 716
rect 964 682 999 716
rect 1033 682 1068 716
rect 1102 682 1137 716
rect 1171 682 1206 716
rect 1240 682 1275 716
rect 1309 682 1344 716
rect 1378 682 1413 716
rect 1447 682 1482 716
rect 1516 682 1551 716
rect 1585 682 1620 716
rect 1654 682 1689 716
rect 1723 682 1758 716
rect 1792 682 1827 716
rect 1861 682 1896 716
rect 1930 682 1965 716
rect 1999 682 2034 716
rect 2068 682 2103 716
rect 2137 682 2172 716
rect 2206 682 2241 716
rect 2275 682 2310 716
rect 2344 682 2379 716
rect 2413 682 2448 716
rect 2482 682 2517 716
rect 2551 682 2586 716
rect 2620 682 2655 716
rect 2689 682 2724 716
rect 2758 682 2793 716
rect 2827 682 2862 716
rect 2896 682 2931 716
rect 2965 682 3000 716
rect 3034 682 3069 716
rect 3103 682 3138 716
rect 3172 682 3207 716
rect 3241 682 3276 716
rect 3310 682 3345 716
rect 3379 682 3414 716
rect 3448 682 3483 716
rect 3517 682 3552 716
rect 3586 682 3621 716
rect 3655 682 3690 716
rect 3724 682 3759 716
rect 3793 682 3828 716
rect 3862 682 3897 716
rect 3931 682 3966 716
rect 4000 682 4035 716
rect 4069 682 4104 716
rect 4138 682 4173 716
rect 4207 682 4242 716
rect 4276 682 4311 716
rect 4345 682 4380 716
rect 4414 682 4449 716
rect 4483 682 4518 716
rect 4552 682 4587 716
rect 4621 682 4656 716
rect 4690 682 4725 716
rect 14551 735 14653 750
rect 14551 701 14604 735
rect 14638 701 14653 735
rect 14551 682 14653 701
rect 482 667 14653 682
<< mvpsubdiffcont >>
rect 121 363 223 5021
rect 306 4898 13600 5068
rect 13635 5034 13669 5068
rect 13704 5034 13738 5068
rect 13773 5034 13807 5068
rect 13842 5034 13876 5068
rect 13911 5034 13945 5068
rect 13980 5034 14014 5068
rect 14049 5034 14083 5068
rect 14118 5034 14152 5068
rect 14187 5034 14221 5068
rect 14256 5034 14290 5068
rect 14325 5034 14359 5068
rect 14394 5034 14428 5068
rect 14463 5034 14497 5068
rect 14532 5034 14566 5068
rect 14601 5034 14635 5068
rect 14670 5034 14704 5068
rect 14739 5034 14773 5068
rect 13635 4966 13669 5000
rect 13704 4966 13738 5000
rect 13773 4966 13807 5000
rect 13842 4966 13876 5000
rect 13911 4966 13945 5000
rect 13980 4966 14014 5000
rect 14049 4966 14083 5000
rect 14118 4966 14152 5000
rect 14187 4966 14221 5000
rect 14256 4966 14290 5000
rect 14325 4966 14359 5000
rect 14394 4966 14428 5000
rect 14463 4966 14497 5000
rect 14532 4966 14566 5000
rect 14601 4966 14635 5000
rect 14670 4966 14704 5000
rect 14739 4966 14773 5000
rect 14840 4999 14874 5033
rect 13635 4898 13669 4932
rect 13704 4898 13738 4932
rect 13773 4898 13807 4932
rect 13842 4898 13876 4932
rect 13911 4898 13945 4932
rect 13980 4898 14014 4932
rect 14049 4898 14083 4932
rect 14118 4898 14152 4932
rect 14187 4898 14221 4932
rect 14256 4898 14290 4932
rect 14325 4898 14359 4932
rect 14394 4898 14428 4932
rect 14463 4898 14497 4932
rect 14532 4898 14566 4932
rect 14601 4898 14635 4932
rect 14670 4898 14704 4932
rect 14739 4898 14773 4932
rect 262 4825 296 4859
rect 262 4757 296 4791
rect 262 4689 296 4723
rect 262 4621 296 4655
rect 262 4553 296 4587
rect 262 4485 296 4519
rect 262 4417 296 4451
rect 262 4349 296 4383
rect 262 4281 296 4315
rect 262 4213 296 4247
rect 262 4145 296 4179
rect 262 4077 296 4111
rect 262 4009 296 4043
rect 262 3941 296 3975
rect 262 3873 296 3907
rect 262 3805 296 3839
rect 262 3737 296 3771
rect 262 3669 296 3703
rect 262 3601 296 3635
rect 262 3533 296 3567
rect 262 3465 296 3499
rect 262 3397 296 3431
rect 262 3329 296 3363
rect 262 3261 296 3295
rect 262 3193 296 3227
rect 262 3125 296 3159
rect 262 3057 296 3091
rect 262 2989 296 3023
rect 262 2921 296 2955
rect 262 2853 296 2887
rect 262 2785 296 2819
rect 262 2717 296 2751
rect 262 2649 296 2683
rect 262 2581 296 2615
rect 262 2513 296 2547
rect 262 2445 296 2479
rect 262 2377 296 2411
rect 262 2309 296 2343
rect 262 2241 296 2275
rect 262 2173 296 2207
rect 262 2105 296 2139
rect 262 2037 296 2071
rect 262 1969 296 2003
rect 262 1901 296 1935
rect 262 1833 296 1867
rect 262 1765 296 1799
rect 262 1697 296 1731
rect 262 1629 296 1663
rect 262 1561 296 1595
rect 262 1493 296 1527
rect 262 1425 296 1459
rect 262 1357 296 1391
rect 262 1289 296 1323
rect 262 1221 296 1255
rect 262 1153 296 1187
rect 262 1085 296 1119
rect 262 1017 296 1051
rect 262 949 296 983
rect 262 881 296 915
rect 262 813 296 847
rect 262 745 296 779
rect 262 677 296 711
rect 262 609 296 643
rect 262 541 296 575
rect 14840 499 14942 4965
rect 262 465 296 499
rect 331 465 365 499
rect 400 465 434 499
rect 469 465 503 499
rect 538 465 572 499
rect 607 465 641 499
rect 676 465 710 499
rect 745 465 779 499
rect 814 465 848 499
rect 883 465 917 499
rect 952 465 986 499
rect 1021 465 1055 499
rect 1090 465 1124 499
rect 1159 465 1193 499
rect 1228 465 1262 499
rect 1297 465 1331 499
rect 1366 465 1400 499
rect 1435 465 1469 499
rect 1504 465 1538 499
rect 1573 465 1607 499
rect 1642 465 1676 499
rect 1711 465 1745 499
rect 1780 465 1814 499
rect 1849 465 1883 499
rect 1918 465 1952 499
rect 1987 465 2021 499
rect 262 397 296 431
rect 331 397 365 431
rect 400 397 434 431
rect 469 397 503 431
rect 538 397 572 431
rect 607 397 641 431
rect 676 397 710 431
rect 745 397 779 431
rect 814 397 848 431
rect 883 397 917 431
rect 952 397 986 431
rect 1021 397 1055 431
rect 1090 397 1124 431
rect 1159 397 1193 431
rect 1228 397 1262 431
rect 1297 397 1331 431
rect 1366 397 1400 431
rect 1435 397 1469 431
rect 1504 397 1538 431
rect 1573 397 1607 431
rect 1642 397 1676 431
rect 1711 397 1745 431
rect 1780 397 1814 431
rect 1849 397 1883 431
rect 1918 397 1952 431
rect 1987 397 2021 431
rect 2056 375 14942 499
rect 262 329 296 363
rect 331 329 365 363
rect 400 329 434 363
rect 469 329 503 363
rect 538 329 572 363
rect 607 329 641 363
rect 676 329 710 363
rect 745 329 779 363
rect 814 329 848 363
rect 883 329 917 363
rect 952 329 986 363
rect 1021 329 1055 363
rect 1090 329 1124 363
rect 1159 329 1193 363
rect 1228 329 1262 363
rect 1297 329 1331 363
rect 1366 329 1400 363
rect 1435 329 1469 363
rect 1504 329 1538 363
rect 1573 329 1607 363
rect 1642 329 1676 363
rect 1711 329 1745 363
rect 1780 329 1814 363
rect 1849 329 1883 363
rect 1918 329 1952 363
rect 1987 329 2021 363
rect 2056 329 14806 375
<< mvnsubdiffcont >>
rect 497 4585 531 4619
rect 584 4570 10410 4638
rect 10445 4604 10479 4638
rect 10514 4604 10548 4638
rect 10583 4604 10617 4638
rect 10652 4604 10686 4638
rect 10721 4604 10755 4638
rect 10790 4604 10824 4638
rect 10859 4604 10893 4638
rect 10928 4604 10962 4638
rect 10997 4604 11031 4638
rect 11066 4604 11100 4638
rect 11135 4604 11169 4638
rect 11204 4604 11238 4638
rect 11273 4604 11307 4638
rect 11342 4604 11376 4638
rect 11411 4604 11445 4638
rect 11480 4604 11514 4638
rect 11549 4604 11583 4638
rect 11618 4604 11652 4638
rect 11687 4604 11721 4638
rect 11756 4604 11790 4638
rect 11825 4604 11859 4638
rect 11894 4604 11928 4638
rect 11963 4604 11997 4638
rect 12032 4604 12066 4638
rect 12101 4604 12135 4638
rect 12170 4604 12204 4638
rect 12239 4604 12273 4638
rect 12308 4604 12342 4638
rect 12377 4604 12411 4638
rect 12446 4604 12480 4638
rect 12515 4604 12549 4638
rect 12584 4604 12618 4638
rect 12653 4604 12687 4638
rect 12722 4604 12756 4638
rect 12791 4604 12825 4638
rect 12860 4604 12894 4638
rect 12929 4604 12963 4638
rect 12998 4604 13032 4638
rect 13067 4604 13101 4638
rect 13136 4604 13170 4638
rect 13205 4604 13239 4638
rect 13274 4604 13308 4638
rect 13343 4604 13377 4638
rect 13412 4604 13446 4638
rect 13481 4604 13515 4638
rect 13550 4604 13584 4638
rect 13619 4604 13653 4638
rect 13688 4604 13722 4638
rect 13757 4604 13791 4638
rect 13826 4604 13860 4638
rect 13895 4604 13929 4638
rect 13964 4604 13998 4638
rect 14033 4604 14067 4638
rect 14102 4604 14136 4638
rect 14171 4604 14205 4638
rect 14240 4604 14274 4638
rect 14309 4604 14343 4638
rect 14378 4604 14412 4638
rect 14447 4604 14481 4638
rect 14516 4604 14550 4638
rect 14585 4604 14619 4638
rect 497 4515 531 4549
rect 565 4536 12363 4570
rect 12397 4536 12431 4570
rect 12466 4536 12500 4570
rect 12535 4536 12569 4570
rect 12604 4536 12638 4570
rect 12673 4536 12707 4570
rect 12742 4536 12776 4570
rect 12811 4536 12845 4570
rect 12880 4536 12914 4570
rect 12949 4536 12983 4570
rect 13018 4536 13052 4570
rect 13087 4536 13121 4570
rect 13156 4536 13190 4570
rect 13225 4536 13259 4570
rect 13294 4536 13328 4570
rect 13363 4536 13397 4570
rect 13432 4536 13466 4570
rect 13501 4536 13535 4570
rect 13570 4536 13604 4570
rect 13639 4536 13673 4570
rect 13708 4536 13742 4570
rect 13777 4536 13811 4570
rect 13846 4536 13880 4570
rect 13915 4536 13949 4570
rect 13984 4536 14018 4570
rect 14053 4536 14087 4570
rect 14122 4536 14156 4570
rect 14191 4536 14225 4570
rect 14260 4536 14294 4570
rect 14329 4536 14363 4570
rect 14398 4536 14432 4570
rect 14467 4536 14501 4570
rect 14536 4551 14570 4570
rect 497 4445 531 4479
rect 565 4464 599 4498
rect 633 4468 12363 4536
rect 14536 4502 14638 4551
rect 12398 4468 12432 4502
rect 12467 4468 12501 4502
rect 12536 4468 12570 4502
rect 12605 4468 12639 4502
rect 12674 4468 12708 4502
rect 12743 4468 12777 4502
rect 12812 4468 12846 4502
rect 12881 4468 12915 4502
rect 12950 4468 12984 4502
rect 13019 4468 13053 4502
rect 13088 4468 13122 4502
rect 13157 4468 13191 4502
rect 13226 4468 13260 4502
rect 13295 4468 13329 4502
rect 13364 4468 13398 4502
rect 13433 4468 13467 4502
rect 13502 4468 13536 4502
rect 13571 4468 13605 4502
rect 13640 4468 13674 4502
rect 13709 4468 13743 4502
rect 13778 4468 13812 4502
rect 13847 4468 13881 4502
rect 13916 4468 13950 4502
rect 13985 4468 14019 4502
rect 14054 4468 14088 4502
rect 14123 4468 14157 4502
rect 14192 4468 14226 4502
rect 14261 4468 14295 4502
rect 14330 4468 14364 4502
rect 14399 4468 14433 4502
rect 497 4375 531 4409
rect 565 4392 599 4426
rect 633 4395 667 4429
rect 497 4305 531 4339
rect 565 4320 599 4354
rect 633 4322 667 4356
rect 497 4235 531 4269
rect 565 4248 599 4282
rect 633 4249 667 4283
rect 497 4165 531 4199
rect 565 4176 599 4210
rect 633 4177 667 4211
rect 497 4095 531 4129
rect 565 4104 599 4138
rect 633 4105 667 4139
rect 497 4025 531 4059
rect 565 4032 599 4066
rect 633 4033 667 4067
rect 497 3955 531 3989
rect 565 3960 599 3994
rect 633 3961 667 3995
rect 497 3886 531 3920
rect 565 3888 599 3922
rect 633 3889 667 3923
rect 497 3817 531 3851
rect 565 3817 599 3851
rect 633 3817 667 3851
rect 497 3715 531 3749
rect 565 3715 599 3749
rect 633 3715 667 3749
rect 497 3646 531 3680
rect 565 3646 599 3680
rect 633 3646 667 3680
rect 497 3577 531 3611
rect 565 3577 599 3611
rect 633 3577 667 3611
rect 497 3508 531 3542
rect 565 3508 599 3542
rect 633 3508 667 3542
rect 497 3439 531 3473
rect 565 3439 599 3473
rect 633 3439 667 3473
rect 497 3370 531 3404
rect 565 3370 599 3404
rect 633 3370 667 3404
rect 497 3301 531 3335
rect 565 3301 599 3335
rect 633 3301 667 3335
rect 497 3232 531 3266
rect 565 3232 599 3266
rect 633 3232 667 3266
rect 497 3163 531 3197
rect 565 3163 599 3197
rect 633 3163 667 3197
rect 14468 3992 14638 4502
rect 14468 3923 14502 3957
rect 14536 3924 14638 3992
rect 14604 3905 14638 3924
rect 14468 3854 14502 3888
rect 14536 3855 14570 3889
rect 14604 3837 14638 3871
rect 14468 3785 14502 3819
rect 14536 3786 14570 3820
rect 14604 3769 14638 3803
rect 14468 3716 14502 3750
rect 14536 3717 14570 3751
rect 14604 3701 14638 3735
rect 14468 3647 14502 3681
rect 14536 3648 14570 3682
rect 14604 3633 14638 3667
rect 14468 3578 14502 3612
rect 14536 3579 14570 3613
rect 14604 3565 14638 3599
rect 14468 3509 14502 3543
rect 14536 3510 14570 3544
rect 14604 3497 14638 3531
rect 14468 3440 14502 3474
rect 14536 3441 14570 3475
rect 14604 3429 14638 3463
rect 14468 3371 14502 3405
rect 14536 3372 14570 3406
rect 14604 3361 14638 3395
rect 14468 3302 14502 3336
rect 14536 3303 14570 3337
rect 14604 3293 14638 3327
rect 14468 3233 14502 3267
rect 14536 3234 14570 3268
rect 14604 3225 14638 3259
rect 14468 3164 14502 3198
rect 14536 3165 14570 3199
rect 14604 3157 14638 3191
rect 497 3094 531 3128
rect 565 3094 599 3128
rect 633 3094 667 3128
rect 497 3025 531 3059
rect 565 3025 599 3059
rect 633 3025 667 3059
rect 497 2956 531 2990
rect 565 2956 599 2990
rect 633 2956 667 2990
rect 497 2887 531 2921
rect 565 2887 599 2921
rect 633 2887 667 2921
rect 497 2818 531 2852
rect 565 2818 599 2852
rect 633 2818 667 2852
rect 497 2749 531 2783
rect 565 2749 599 2783
rect 633 2749 667 2783
rect 497 2680 531 2714
rect 565 2680 599 2714
rect 633 2680 667 2714
rect 497 2611 531 2645
rect 565 2611 599 2645
rect 633 2611 667 2645
rect 1601 3010 1635 3044
rect 1669 3010 1703 3044
rect 1601 2940 1635 2974
rect 1669 2940 1703 2974
rect 1601 2870 1635 2904
rect 1669 2870 1703 2904
rect 1601 2800 1635 2834
rect 1669 2800 1703 2834
rect 1601 2730 1635 2764
rect 1669 2730 1703 2764
rect 1601 2660 1635 2694
rect 1669 2660 1703 2694
rect 2593 3010 2627 3044
rect 2661 3010 2695 3044
rect 2593 2940 2627 2974
rect 2661 2940 2695 2974
rect 2593 2870 2627 2904
rect 2661 2870 2695 2904
rect 2593 2800 2627 2834
rect 2661 2800 2695 2834
rect 2593 2730 2627 2764
rect 2661 2730 2695 2764
rect 2593 2660 2627 2694
rect 2661 2660 2695 2694
rect 3585 3010 3619 3044
rect 3653 3010 3687 3044
rect 3585 2940 3619 2974
rect 3653 2940 3687 2974
rect 3585 2870 3619 2904
rect 3653 2870 3687 2904
rect 3585 2800 3619 2834
rect 3653 2800 3687 2834
rect 3585 2730 3619 2764
rect 3653 2730 3687 2764
rect 3585 2660 3619 2694
rect 3653 2660 3687 2694
rect 4577 3010 4611 3044
rect 4645 3010 4679 3044
rect 4577 2940 4611 2974
rect 4645 2940 4679 2974
rect 4577 2870 4611 2904
rect 4645 2870 4679 2904
rect 4577 2800 4611 2834
rect 4645 2800 4679 2834
rect 4577 2730 4611 2764
rect 4645 2730 4679 2764
rect 4577 2660 4611 2694
rect 4645 2660 4679 2694
rect 5569 3010 5603 3044
rect 5637 3010 5671 3044
rect 5569 2940 5603 2974
rect 5637 2940 5671 2974
rect 5569 2870 5603 2904
rect 5637 2870 5671 2904
rect 5569 2800 5603 2834
rect 5637 2800 5671 2834
rect 5569 2730 5603 2764
rect 5637 2730 5671 2764
rect 5569 2660 5603 2694
rect 5637 2660 5671 2694
rect 6561 3010 6595 3044
rect 6629 3010 6663 3044
rect 6561 2940 6595 2974
rect 6629 2940 6663 2974
rect 6561 2870 6595 2904
rect 6629 2870 6663 2904
rect 6561 2800 6595 2834
rect 6629 2800 6663 2834
rect 6561 2730 6595 2764
rect 6629 2730 6663 2764
rect 6561 2660 6595 2694
rect 6629 2660 6663 2694
rect 7553 3010 7587 3044
rect 7621 3010 7655 3044
rect 7553 2940 7587 2974
rect 7621 2940 7655 2974
rect 7553 2870 7587 2904
rect 7621 2870 7655 2904
rect 7553 2800 7587 2834
rect 7621 2800 7655 2834
rect 7553 2730 7587 2764
rect 7621 2730 7655 2764
rect 7553 2660 7587 2694
rect 7621 2660 7655 2694
rect 8545 3010 8579 3044
rect 8613 3010 8647 3044
rect 8545 2940 8579 2974
rect 8613 2940 8647 2974
rect 8545 2870 8579 2904
rect 8613 2870 8647 2904
rect 8545 2800 8579 2834
rect 8613 2800 8647 2834
rect 8545 2730 8579 2764
rect 8613 2730 8647 2764
rect 8545 2660 8579 2694
rect 8613 2660 8647 2694
rect 9537 3010 9571 3044
rect 9605 3010 9639 3044
rect 9537 2940 9571 2974
rect 9605 2940 9639 2974
rect 9537 2870 9571 2904
rect 9605 2870 9639 2904
rect 9537 2800 9571 2834
rect 9605 2800 9639 2834
rect 9537 2730 9571 2764
rect 9605 2730 9639 2764
rect 9537 2660 9571 2694
rect 9605 2660 9639 2694
rect 10529 3010 10563 3044
rect 10597 3010 10631 3044
rect 10529 2940 10563 2974
rect 10597 2940 10631 2974
rect 10529 2870 10563 2904
rect 10597 2870 10631 2904
rect 10529 2800 10563 2834
rect 10597 2800 10631 2834
rect 10529 2730 10563 2764
rect 10597 2730 10631 2764
rect 10529 2660 10563 2694
rect 10597 2660 10631 2694
rect 11521 3010 11555 3044
rect 11589 3010 11623 3044
rect 11521 2940 11555 2974
rect 11589 2940 11623 2974
rect 11521 2870 11555 2904
rect 11589 2870 11623 2904
rect 11521 2800 11555 2834
rect 11589 2800 11623 2834
rect 11521 2730 11555 2764
rect 11589 2730 11623 2764
rect 11521 2660 11555 2694
rect 11589 2660 11623 2694
rect 12513 3010 12547 3044
rect 12581 3010 12615 3044
rect 12513 2940 12547 2974
rect 12581 2940 12615 2974
rect 12513 2870 12547 2904
rect 12581 2870 12615 2904
rect 12513 2800 12547 2834
rect 12581 2800 12615 2834
rect 12513 2730 12547 2764
rect 12581 2730 12615 2764
rect 12513 2660 12547 2694
rect 12581 2660 12615 2694
rect 13505 3010 13539 3044
rect 13573 3010 13607 3044
rect 13505 2940 13539 2974
rect 13573 2940 13607 2974
rect 13505 2870 13539 2904
rect 13573 2870 13607 2904
rect 13505 2800 13539 2834
rect 13573 2800 13607 2834
rect 13505 2730 13539 2764
rect 13573 2730 13607 2764
rect 13505 2660 13539 2694
rect 13573 2660 13607 2694
rect 14468 3095 14502 3129
rect 14536 3096 14570 3130
rect 14604 3089 14638 3123
rect 14468 3026 14502 3060
rect 14536 3027 14570 3061
rect 14604 3021 14638 3055
rect 14468 2957 14502 2991
rect 14536 2958 14570 2992
rect 14604 2953 14638 2987
rect 14468 2888 14502 2922
rect 14536 2889 14570 2923
rect 14604 2885 14638 2919
rect 14468 2819 14502 2853
rect 14536 2820 14570 2854
rect 14604 2817 14638 2851
rect 14468 2750 14502 2784
rect 14536 2751 14570 2785
rect 14604 2749 14638 2783
rect 14468 2681 14502 2715
rect 14536 2682 14570 2716
rect 14604 2681 14638 2715
rect 14468 2612 14502 2646
rect 14536 2613 14570 2647
rect 14604 2613 14638 2647
rect 497 2542 531 2576
rect 565 2542 599 2576
rect 633 2542 667 2576
rect 497 2473 531 2507
rect 565 2473 599 2507
rect 633 2473 667 2507
rect 497 2404 531 2438
rect 565 2404 599 2438
rect 633 2404 667 2438
rect 497 2335 531 2369
rect 565 2335 599 2369
rect 633 2335 667 2369
rect 497 2266 531 2300
rect 565 2266 599 2300
rect 633 2266 667 2300
rect 497 2197 531 2231
rect 565 2197 599 2231
rect 633 2197 667 2231
rect 497 2129 531 2163
rect 565 2128 599 2162
rect 633 2128 667 2162
rect 497 2061 531 2095
rect 565 2059 599 2093
rect 633 2059 667 2093
rect 497 1993 531 2027
rect 565 1990 599 2024
rect 633 1990 667 2024
rect 497 1925 531 1959
rect 565 1921 599 1955
rect 633 1921 667 1955
rect 497 1857 531 1891
rect 565 1852 599 1886
rect 633 1852 667 1886
rect 497 1789 531 1823
rect 565 1783 599 1817
rect 633 1783 667 1817
rect 497 1721 531 1755
rect 565 1714 599 1748
rect 633 1714 667 1748
rect 497 1653 531 1687
rect 565 1645 599 1679
rect 633 1645 667 1679
rect 497 1585 531 1619
rect 565 1576 599 1610
rect 633 1576 667 1610
rect 14468 2543 14502 2577
rect 14536 2544 14570 2578
rect 14604 2545 14638 2579
rect 14468 2474 14502 2508
rect 14536 2475 14570 2509
rect 14604 2477 14638 2511
rect 14468 2405 14502 2439
rect 14536 2406 14570 2440
rect 14604 2409 14638 2443
rect 14468 2336 14502 2370
rect 14536 2337 14570 2371
rect 14604 2341 14638 2375
rect 14468 2267 14502 2301
rect 14536 2268 14570 2302
rect 14604 2273 14638 2307
rect 14468 2198 14502 2232
rect 14536 2199 14570 2233
rect 14604 2205 14638 2239
rect 14468 2129 14502 2163
rect 14536 2130 14570 2164
rect 14604 2137 14638 2171
rect 14468 2060 14502 2094
rect 14536 2061 14570 2095
rect 14604 2069 14638 2103
rect 14468 1991 14502 2025
rect 14536 1992 14570 2026
rect 14604 2001 14638 2035
rect 14468 1922 14502 1956
rect 14536 1923 14570 1957
rect 14604 1933 14638 1967
rect 14468 1853 14502 1887
rect 14536 1854 14570 1888
rect 14604 1865 14638 1899
rect 14468 1784 14502 1818
rect 14536 1785 14570 1819
rect 14604 1797 14638 1831
rect 14468 1715 14502 1749
rect 14536 1716 14570 1750
rect 14604 1729 14638 1763
rect 14468 1646 14502 1680
rect 14536 1647 14570 1681
rect 14604 1661 14638 1695
rect 14468 1577 14502 1611
rect 14536 1578 14570 1612
rect 14604 1593 14638 1627
rect 497 1517 531 1551
rect 565 1507 599 1541
rect 633 1507 667 1541
rect 497 1449 531 1483
rect 565 1438 599 1472
rect 633 1438 667 1472
rect 497 1381 531 1415
rect 565 1369 599 1403
rect 633 1369 667 1403
rect 14468 1508 14502 1542
rect 14536 1509 14570 1543
rect 14604 1525 14638 1559
rect 14468 1439 14502 1473
rect 14536 1440 14570 1474
rect 14604 1457 14638 1491
rect 497 1313 531 1347
rect 565 1300 599 1334
rect 633 1300 667 1334
rect 497 1245 531 1279
rect 565 1231 599 1265
rect 633 1231 667 1265
rect 497 1177 531 1211
rect 565 1162 599 1196
rect 633 1162 667 1196
rect 497 1109 531 1143
rect 565 1093 599 1127
rect 633 1093 667 1127
rect 497 1041 531 1075
rect 565 1024 599 1058
rect 633 1024 667 1058
rect 497 973 531 1007
rect 565 955 599 989
rect 633 955 667 989
rect 497 920 531 939
rect 497 818 667 920
rect 14468 1370 14502 1404
rect 14536 1371 14570 1405
rect 14604 1389 14638 1423
rect 14468 1301 14502 1335
rect 14536 1302 14570 1336
rect 14604 1321 14638 1355
rect 14468 1232 14502 1266
rect 14536 1233 14570 1267
rect 14604 1253 14638 1287
rect 14468 1163 14502 1197
rect 14536 1164 14570 1198
rect 14604 1184 14638 1218
rect 14468 1094 14502 1128
rect 14536 1095 14570 1129
rect 14604 1115 14638 1149
rect 14468 1025 14502 1059
rect 14536 1026 14570 1060
rect 14604 1046 14638 1080
rect 14468 956 14502 990
rect 14536 957 14570 991
rect 14604 977 14638 1011
rect 14468 887 14502 921
rect 14536 888 14570 922
rect 14604 908 14638 942
rect 702 818 736 852
rect 771 818 805 852
rect 840 818 874 852
rect 909 818 943 852
rect 978 818 1012 852
rect 1047 818 1081 852
rect 1116 818 1150 852
rect 1185 818 1219 852
rect 1254 818 1288 852
rect 1323 818 1357 852
rect 1392 818 1426 852
rect 1461 818 1495 852
rect 1530 818 1564 852
rect 1599 818 1633 852
rect 1668 818 1702 852
rect 1737 818 1771 852
rect 1806 818 1840 852
rect 1875 818 1909 852
rect 1944 818 1978 852
rect 2013 818 2047 852
rect 2082 818 2116 852
rect 2151 818 2185 852
rect 2220 818 2254 852
rect 2289 818 2323 852
rect 2358 818 2392 852
rect 2427 818 2461 852
rect 2496 818 2530 852
rect 2565 818 2599 852
rect 2634 818 2668 852
rect 2703 818 2737 852
rect 497 769 599 818
rect 2772 784 14502 852
rect 14536 819 14570 853
rect 14604 839 14638 873
rect 565 750 599 769
rect 634 750 668 784
rect 703 750 737 784
rect 772 750 806 784
rect 841 750 875 784
rect 910 750 944 784
rect 979 750 1013 784
rect 1048 750 1082 784
rect 1117 750 1151 784
rect 1186 750 1220 784
rect 1255 750 1289 784
rect 1324 750 1358 784
rect 1393 750 1427 784
rect 1462 750 1496 784
rect 1531 750 1565 784
rect 1600 750 1634 784
rect 1669 750 1703 784
rect 1738 750 1772 784
rect 1807 750 1841 784
rect 1876 750 1910 784
rect 1945 750 1979 784
rect 2014 750 2048 784
rect 2083 750 2117 784
rect 2152 750 2186 784
rect 2221 750 2255 784
rect 2290 750 2324 784
rect 2359 750 2393 784
rect 2428 750 2462 784
rect 2497 750 2531 784
rect 2566 750 2600 784
rect 2635 750 2669 784
rect 2704 750 2738 784
rect 2772 750 14570 784
rect 14604 770 14638 804
rect 516 682 550 716
rect 585 682 619 716
rect 654 682 688 716
rect 723 682 757 716
rect 792 682 826 716
rect 861 682 895 716
rect 930 682 964 716
rect 999 682 1033 716
rect 1068 682 1102 716
rect 1137 682 1171 716
rect 1206 682 1240 716
rect 1275 682 1309 716
rect 1344 682 1378 716
rect 1413 682 1447 716
rect 1482 682 1516 716
rect 1551 682 1585 716
rect 1620 682 1654 716
rect 1689 682 1723 716
rect 1758 682 1792 716
rect 1827 682 1861 716
rect 1896 682 1930 716
rect 1965 682 1999 716
rect 2034 682 2068 716
rect 2103 682 2137 716
rect 2172 682 2206 716
rect 2241 682 2275 716
rect 2310 682 2344 716
rect 2379 682 2413 716
rect 2448 682 2482 716
rect 2517 682 2551 716
rect 2586 682 2620 716
rect 2655 682 2689 716
rect 2724 682 2758 716
rect 2793 682 2827 716
rect 2862 682 2896 716
rect 2931 682 2965 716
rect 3000 682 3034 716
rect 3069 682 3103 716
rect 3138 682 3172 716
rect 3207 682 3241 716
rect 3276 682 3310 716
rect 3345 682 3379 716
rect 3414 682 3448 716
rect 3483 682 3517 716
rect 3552 682 3586 716
rect 3621 682 3655 716
rect 3690 682 3724 716
rect 3759 682 3793 716
rect 3828 682 3862 716
rect 3897 682 3931 716
rect 3966 682 4000 716
rect 4035 682 4069 716
rect 4104 682 4138 716
rect 4173 682 4207 716
rect 4242 682 4276 716
rect 4311 682 4345 716
rect 4380 682 4414 716
rect 4449 682 4483 716
rect 4518 682 4552 716
rect 4587 682 4621 716
rect 4656 682 4690 716
rect 4725 682 14551 750
rect 14604 701 14638 735
<< poly >>
rect 881 4308 1001 4324
rect 881 4274 924 4308
rect 958 4274 1001 4308
rect 881 4234 1001 4274
rect 881 4200 924 4234
rect 958 4200 1001 4234
rect 881 4184 1001 4200
rect 1311 4308 1431 4324
rect 1311 4274 1354 4308
rect 1388 4274 1431 4308
rect 1311 4234 1431 4274
rect 1311 4200 1354 4234
rect 1388 4200 1431 4234
rect 1311 4184 1431 4200
rect 1873 4308 1993 4324
rect 1873 4274 1916 4308
rect 1950 4274 1993 4308
rect 1873 4234 1993 4274
rect 1873 4200 1916 4234
rect 1950 4200 1993 4234
rect 1873 4184 1993 4200
rect 2303 4308 2423 4324
rect 2303 4274 2346 4308
rect 2380 4274 2423 4308
rect 2303 4234 2423 4274
rect 2303 4200 2346 4234
rect 2380 4200 2423 4234
rect 2303 4184 2423 4200
rect 2865 4308 2985 4324
rect 2865 4274 2908 4308
rect 2942 4274 2985 4308
rect 2865 4234 2985 4274
rect 2865 4200 2908 4234
rect 2942 4200 2985 4234
rect 2865 4184 2985 4200
rect 3295 4308 3415 4324
rect 3295 4274 3338 4308
rect 3372 4274 3415 4308
rect 3295 4234 3415 4274
rect 3295 4200 3338 4234
rect 3372 4200 3415 4234
rect 3295 4184 3415 4200
rect 3857 4308 3977 4324
rect 3857 4274 3900 4308
rect 3934 4274 3977 4308
rect 3857 4234 3977 4274
rect 3857 4200 3900 4234
rect 3934 4200 3977 4234
rect 3857 4184 3977 4200
rect 4287 4308 4407 4324
rect 4287 4274 4330 4308
rect 4364 4274 4407 4308
rect 4287 4234 4407 4274
rect 4287 4200 4330 4234
rect 4364 4200 4407 4234
rect 4287 4184 4407 4200
rect 4849 4308 4969 4324
rect 4849 4274 4892 4308
rect 4926 4274 4969 4308
rect 4849 4234 4969 4274
rect 4849 4200 4892 4234
rect 4926 4200 4969 4234
rect 4849 4184 4969 4200
rect 5279 4308 5399 4324
rect 5279 4274 5322 4308
rect 5356 4274 5399 4308
rect 5279 4234 5399 4274
rect 5279 4200 5322 4234
rect 5356 4200 5399 4234
rect 5279 4184 5399 4200
rect 5841 4308 5961 4324
rect 5841 4274 5884 4308
rect 5918 4274 5961 4308
rect 5841 4234 5961 4274
rect 5841 4200 5884 4234
rect 5918 4200 5961 4234
rect 5841 4184 5961 4200
rect 6271 4308 6391 4324
rect 6271 4274 6314 4308
rect 6348 4274 6391 4308
rect 6271 4234 6391 4274
rect 6271 4200 6314 4234
rect 6348 4200 6391 4234
rect 6271 4184 6391 4200
rect 6833 4308 6953 4324
rect 6833 4274 6876 4308
rect 6910 4274 6953 4308
rect 6833 4234 6953 4274
rect 6833 4200 6876 4234
rect 6910 4200 6953 4234
rect 6833 4184 6953 4200
rect 7263 4308 7383 4324
rect 7263 4274 7306 4308
rect 7340 4274 7383 4308
rect 7263 4234 7383 4274
rect 7263 4200 7306 4234
rect 7340 4200 7383 4234
rect 7263 4184 7383 4200
rect 7825 4308 7945 4324
rect 7825 4274 7868 4308
rect 7902 4274 7945 4308
rect 7825 4234 7945 4274
rect 7825 4200 7868 4234
rect 7902 4200 7945 4234
rect 7825 4184 7945 4200
rect 8255 4308 8375 4324
rect 8255 4274 8298 4308
rect 8332 4274 8375 4308
rect 8255 4234 8375 4274
rect 8255 4200 8298 4234
rect 8332 4200 8375 4234
rect 8255 4184 8375 4200
rect 8817 4308 8937 4324
rect 8817 4274 8860 4308
rect 8894 4274 8937 4308
rect 8817 4234 8937 4274
rect 8817 4200 8860 4234
rect 8894 4200 8937 4234
rect 8817 4184 8937 4200
rect 9247 4308 9367 4324
rect 9247 4274 9290 4308
rect 9324 4274 9367 4308
rect 9247 4234 9367 4274
rect 9247 4200 9290 4234
rect 9324 4200 9367 4234
rect 9247 4184 9367 4200
rect 9809 4308 9929 4324
rect 9809 4274 9852 4308
rect 9886 4274 9929 4308
rect 9809 4234 9929 4274
rect 9809 4200 9852 4234
rect 9886 4200 9929 4234
rect 9809 4184 9929 4200
rect 10239 4308 10359 4324
rect 10239 4274 10282 4308
rect 10316 4274 10359 4308
rect 10239 4234 10359 4274
rect 10239 4200 10282 4234
rect 10316 4200 10359 4234
rect 10239 4184 10359 4200
rect 10801 4308 10921 4324
rect 10801 4274 10844 4308
rect 10878 4274 10921 4308
rect 10801 4234 10921 4274
rect 10801 4200 10844 4234
rect 10878 4200 10921 4234
rect 10801 4184 10921 4200
rect 11231 4308 11351 4324
rect 11231 4274 11274 4308
rect 11308 4274 11351 4308
rect 11231 4234 11351 4274
rect 11231 4200 11274 4234
rect 11308 4200 11351 4234
rect 11231 4184 11351 4200
rect 11793 4308 11913 4324
rect 11793 4274 11836 4308
rect 11870 4274 11913 4308
rect 11793 4234 11913 4274
rect 11793 4200 11836 4234
rect 11870 4200 11913 4234
rect 11793 4184 11913 4200
rect 12223 4308 12343 4324
rect 12223 4274 12266 4308
rect 12300 4274 12343 4308
rect 12223 4234 12343 4274
rect 12223 4200 12266 4234
rect 12300 4200 12343 4234
rect 12223 4184 12343 4200
rect 12785 4308 12905 4324
rect 12785 4274 12828 4308
rect 12862 4274 12905 4308
rect 12785 4234 12905 4274
rect 12785 4200 12828 4234
rect 12862 4200 12905 4234
rect 12785 4184 12905 4200
rect 13215 4308 13335 4324
rect 13215 4274 13258 4308
rect 13292 4274 13335 4308
rect 13215 4234 13335 4274
rect 13215 4200 13258 4234
rect 13292 4200 13335 4234
rect 13215 4184 13335 4200
rect 13777 4308 13897 4324
rect 13777 4274 13820 4308
rect 13854 4274 13897 4308
rect 13777 4234 13897 4274
rect 13777 4200 13820 4234
rect 13854 4200 13897 4234
rect 13777 4184 13897 4200
rect 14135 4308 14255 4324
rect 14135 4274 14178 4308
rect 14212 4274 14255 4308
rect 14135 4234 14255 4274
rect 14135 4200 14178 4234
rect 14212 4200 14255 4234
rect 14135 4184 14255 4200
rect 881 3104 1001 3120
rect 881 3070 924 3104
rect 958 3070 1001 3104
rect 881 3026 1001 3070
rect 881 2992 924 3026
rect 958 2992 1001 3026
rect 881 2948 1001 2992
rect 881 2914 924 2948
rect 958 2914 1001 2948
rect 881 2870 1001 2914
rect 881 2836 924 2870
rect 958 2836 1001 2870
rect 881 2792 1001 2836
rect 881 2758 924 2792
rect 958 2758 1001 2792
rect 881 2713 1001 2758
rect 881 2679 924 2713
rect 958 2679 1001 2713
rect 881 2634 1001 2679
rect 881 2600 924 2634
rect 958 2600 1001 2634
rect 881 2584 1001 2600
rect 1311 3104 1431 3120
rect 1311 3070 1354 3104
rect 1388 3070 1431 3104
rect 1873 3104 1993 3120
rect 1311 3026 1431 3070
rect 1311 2992 1354 3026
rect 1388 2992 1431 3026
rect 1311 2948 1431 2992
rect 1311 2914 1354 2948
rect 1388 2914 1431 2948
rect 1311 2870 1431 2914
rect 1311 2836 1354 2870
rect 1388 2836 1431 2870
rect 1311 2792 1431 2836
rect 1311 2758 1354 2792
rect 1388 2758 1431 2792
rect 1311 2713 1431 2758
rect 1311 2679 1354 2713
rect 1388 2679 1431 2713
rect 1311 2634 1431 2679
rect 1311 2600 1354 2634
rect 1388 2600 1431 2634
rect 1873 3070 1916 3104
rect 1950 3070 1993 3104
rect 1873 3026 1993 3070
rect 1873 2992 1916 3026
rect 1950 2992 1993 3026
rect 1873 2948 1993 2992
rect 1873 2914 1916 2948
rect 1950 2914 1993 2948
rect 1873 2870 1993 2914
rect 1873 2836 1916 2870
rect 1950 2836 1993 2870
rect 1873 2792 1993 2836
rect 1873 2758 1916 2792
rect 1950 2758 1993 2792
rect 1873 2713 1993 2758
rect 1873 2679 1916 2713
rect 1950 2679 1993 2713
rect 1873 2634 1993 2679
rect 1311 2584 1431 2600
rect 1873 2600 1916 2634
rect 1950 2600 1993 2634
rect 1873 2584 1993 2600
rect 2303 3104 2423 3120
rect 2303 3070 2346 3104
rect 2380 3070 2423 3104
rect 2865 3104 2985 3120
rect 2303 3026 2423 3070
rect 2303 2992 2346 3026
rect 2380 2992 2423 3026
rect 2303 2948 2423 2992
rect 2303 2914 2346 2948
rect 2380 2914 2423 2948
rect 2303 2870 2423 2914
rect 2303 2836 2346 2870
rect 2380 2836 2423 2870
rect 2303 2792 2423 2836
rect 2303 2758 2346 2792
rect 2380 2758 2423 2792
rect 2303 2713 2423 2758
rect 2303 2679 2346 2713
rect 2380 2679 2423 2713
rect 2303 2634 2423 2679
rect 2303 2600 2346 2634
rect 2380 2600 2423 2634
rect 2865 3070 2908 3104
rect 2942 3070 2985 3104
rect 2865 3026 2985 3070
rect 2865 2992 2908 3026
rect 2942 2992 2985 3026
rect 2865 2948 2985 2992
rect 2865 2914 2908 2948
rect 2942 2914 2985 2948
rect 2865 2870 2985 2914
rect 2865 2836 2908 2870
rect 2942 2836 2985 2870
rect 2865 2792 2985 2836
rect 2865 2758 2908 2792
rect 2942 2758 2985 2792
rect 2865 2713 2985 2758
rect 2865 2679 2908 2713
rect 2942 2679 2985 2713
rect 2865 2634 2985 2679
rect 2303 2584 2423 2600
rect 2865 2600 2908 2634
rect 2942 2600 2985 2634
rect 2865 2584 2985 2600
rect 3295 3104 3415 3120
rect 3295 3070 3338 3104
rect 3372 3070 3415 3104
rect 3857 3104 3977 3120
rect 3295 3026 3415 3070
rect 3295 2992 3338 3026
rect 3372 2992 3415 3026
rect 3295 2948 3415 2992
rect 3295 2914 3338 2948
rect 3372 2914 3415 2948
rect 3295 2870 3415 2914
rect 3295 2836 3338 2870
rect 3372 2836 3415 2870
rect 3295 2792 3415 2836
rect 3295 2758 3338 2792
rect 3372 2758 3415 2792
rect 3295 2713 3415 2758
rect 3295 2679 3338 2713
rect 3372 2679 3415 2713
rect 3295 2634 3415 2679
rect 3295 2600 3338 2634
rect 3372 2600 3415 2634
rect 3857 3070 3900 3104
rect 3934 3070 3977 3104
rect 3857 3026 3977 3070
rect 3857 2992 3900 3026
rect 3934 2992 3977 3026
rect 3857 2948 3977 2992
rect 3857 2914 3900 2948
rect 3934 2914 3977 2948
rect 3857 2870 3977 2914
rect 3857 2836 3900 2870
rect 3934 2836 3977 2870
rect 3857 2792 3977 2836
rect 3857 2758 3900 2792
rect 3934 2758 3977 2792
rect 3857 2713 3977 2758
rect 3857 2679 3900 2713
rect 3934 2679 3977 2713
rect 3857 2634 3977 2679
rect 3295 2584 3415 2600
rect 3857 2600 3900 2634
rect 3934 2600 3977 2634
rect 3857 2584 3977 2600
rect 4287 3104 4407 3120
rect 4287 3070 4330 3104
rect 4364 3070 4407 3104
rect 4849 3104 4969 3120
rect 4287 3026 4407 3070
rect 4287 2992 4330 3026
rect 4364 2992 4407 3026
rect 4287 2948 4407 2992
rect 4287 2914 4330 2948
rect 4364 2914 4407 2948
rect 4287 2870 4407 2914
rect 4287 2836 4330 2870
rect 4364 2836 4407 2870
rect 4287 2792 4407 2836
rect 4287 2758 4330 2792
rect 4364 2758 4407 2792
rect 4287 2713 4407 2758
rect 4287 2679 4330 2713
rect 4364 2679 4407 2713
rect 4287 2634 4407 2679
rect 4287 2600 4330 2634
rect 4364 2600 4407 2634
rect 4849 3070 4892 3104
rect 4926 3070 4969 3104
rect 4849 3026 4969 3070
rect 4849 2992 4892 3026
rect 4926 2992 4969 3026
rect 4849 2948 4969 2992
rect 4849 2914 4892 2948
rect 4926 2914 4969 2948
rect 4849 2870 4969 2914
rect 4849 2836 4892 2870
rect 4926 2836 4969 2870
rect 4849 2792 4969 2836
rect 4849 2758 4892 2792
rect 4926 2758 4969 2792
rect 4849 2713 4969 2758
rect 4849 2679 4892 2713
rect 4926 2679 4969 2713
rect 4849 2634 4969 2679
rect 4287 2584 4407 2600
rect 4849 2600 4892 2634
rect 4926 2600 4969 2634
rect 4849 2584 4969 2600
rect 5279 3104 5399 3120
rect 5279 3070 5322 3104
rect 5356 3070 5399 3104
rect 5841 3104 5961 3120
rect 5279 3026 5399 3070
rect 5279 2992 5322 3026
rect 5356 2992 5399 3026
rect 5279 2948 5399 2992
rect 5279 2914 5322 2948
rect 5356 2914 5399 2948
rect 5279 2870 5399 2914
rect 5279 2836 5322 2870
rect 5356 2836 5399 2870
rect 5279 2792 5399 2836
rect 5279 2758 5322 2792
rect 5356 2758 5399 2792
rect 5279 2713 5399 2758
rect 5279 2679 5322 2713
rect 5356 2679 5399 2713
rect 5279 2634 5399 2679
rect 5279 2600 5322 2634
rect 5356 2600 5399 2634
rect 5841 3070 5884 3104
rect 5918 3070 5961 3104
rect 5841 3026 5961 3070
rect 5841 2992 5884 3026
rect 5918 2992 5961 3026
rect 5841 2948 5961 2992
rect 5841 2914 5884 2948
rect 5918 2914 5961 2948
rect 5841 2870 5961 2914
rect 5841 2836 5884 2870
rect 5918 2836 5961 2870
rect 5841 2792 5961 2836
rect 5841 2758 5884 2792
rect 5918 2758 5961 2792
rect 5841 2713 5961 2758
rect 5841 2679 5884 2713
rect 5918 2679 5961 2713
rect 5841 2634 5961 2679
rect 5279 2584 5399 2600
rect 5841 2600 5884 2634
rect 5918 2600 5961 2634
rect 5841 2584 5961 2600
rect 6271 3104 6391 3120
rect 6271 3070 6314 3104
rect 6348 3070 6391 3104
rect 6833 3104 6953 3120
rect 6271 3026 6391 3070
rect 6271 2992 6314 3026
rect 6348 2992 6391 3026
rect 6271 2948 6391 2992
rect 6271 2914 6314 2948
rect 6348 2914 6391 2948
rect 6271 2870 6391 2914
rect 6271 2836 6314 2870
rect 6348 2836 6391 2870
rect 6271 2792 6391 2836
rect 6271 2758 6314 2792
rect 6348 2758 6391 2792
rect 6271 2713 6391 2758
rect 6271 2679 6314 2713
rect 6348 2679 6391 2713
rect 6271 2634 6391 2679
rect 6271 2600 6314 2634
rect 6348 2600 6391 2634
rect 6833 3070 6876 3104
rect 6910 3070 6953 3104
rect 6833 3026 6953 3070
rect 6833 2992 6876 3026
rect 6910 2992 6953 3026
rect 6833 2948 6953 2992
rect 6833 2914 6876 2948
rect 6910 2914 6953 2948
rect 6833 2870 6953 2914
rect 6833 2836 6876 2870
rect 6910 2836 6953 2870
rect 6833 2792 6953 2836
rect 6833 2758 6876 2792
rect 6910 2758 6953 2792
rect 6833 2713 6953 2758
rect 6833 2679 6876 2713
rect 6910 2679 6953 2713
rect 6833 2634 6953 2679
rect 6271 2584 6391 2600
rect 6833 2600 6876 2634
rect 6910 2600 6953 2634
rect 6833 2584 6953 2600
rect 7263 3104 7383 3120
rect 7263 3070 7306 3104
rect 7340 3070 7383 3104
rect 7825 3104 7945 3120
rect 7263 3026 7383 3070
rect 7263 2992 7306 3026
rect 7340 2992 7383 3026
rect 7263 2948 7383 2992
rect 7263 2914 7306 2948
rect 7340 2914 7383 2948
rect 7263 2870 7383 2914
rect 7263 2836 7306 2870
rect 7340 2836 7383 2870
rect 7263 2792 7383 2836
rect 7263 2758 7306 2792
rect 7340 2758 7383 2792
rect 7263 2713 7383 2758
rect 7263 2679 7306 2713
rect 7340 2679 7383 2713
rect 7263 2634 7383 2679
rect 7263 2600 7306 2634
rect 7340 2600 7383 2634
rect 7825 3070 7868 3104
rect 7902 3070 7945 3104
rect 7825 3026 7945 3070
rect 7825 2992 7868 3026
rect 7902 2992 7945 3026
rect 7825 2948 7945 2992
rect 7825 2914 7868 2948
rect 7902 2914 7945 2948
rect 7825 2870 7945 2914
rect 7825 2836 7868 2870
rect 7902 2836 7945 2870
rect 7825 2792 7945 2836
rect 7825 2758 7868 2792
rect 7902 2758 7945 2792
rect 7825 2713 7945 2758
rect 7825 2679 7868 2713
rect 7902 2679 7945 2713
rect 7825 2634 7945 2679
rect 7263 2584 7383 2600
rect 7825 2600 7868 2634
rect 7902 2600 7945 2634
rect 7825 2584 7945 2600
rect 8255 3104 8375 3120
rect 8255 3070 8298 3104
rect 8332 3070 8375 3104
rect 8817 3104 8937 3120
rect 8255 3026 8375 3070
rect 8255 2992 8298 3026
rect 8332 2992 8375 3026
rect 8255 2948 8375 2992
rect 8255 2914 8298 2948
rect 8332 2914 8375 2948
rect 8255 2870 8375 2914
rect 8255 2836 8298 2870
rect 8332 2836 8375 2870
rect 8255 2792 8375 2836
rect 8255 2758 8298 2792
rect 8332 2758 8375 2792
rect 8255 2713 8375 2758
rect 8255 2679 8298 2713
rect 8332 2679 8375 2713
rect 8255 2634 8375 2679
rect 8255 2600 8298 2634
rect 8332 2600 8375 2634
rect 8817 3070 8860 3104
rect 8894 3070 8937 3104
rect 8817 3026 8937 3070
rect 8817 2992 8860 3026
rect 8894 2992 8937 3026
rect 8817 2948 8937 2992
rect 8817 2914 8860 2948
rect 8894 2914 8937 2948
rect 8817 2870 8937 2914
rect 8817 2836 8860 2870
rect 8894 2836 8937 2870
rect 8817 2792 8937 2836
rect 8817 2758 8860 2792
rect 8894 2758 8937 2792
rect 8817 2713 8937 2758
rect 8817 2679 8860 2713
rect 8894 2679 8937 2713
rect 8817 2634 8937 2679
rect 8255 2584 8375 2600
rect 8817 2600 8860 2634
rect 8894 2600 8937 2634
rect 8817 2584 8937 2600
rect 9247 3104 9367 3120
rect 9247 3070 9290 3104
rect 9324 3070 9367 3104
rect 9809 3104 9929 3120
rect 9247 3026 9367 3070
rect 9247 2992 9290 3026
rect 9324 2992 9367 3026
rect 9247 2948 9367 2992
rect 9247 2914 9290 2948
rect 9324 2914 9367 2948
rect 9247 2870 9367 2914
rect 9247 2836 9290 2870
rect 9324 2836 9367 2870
rect 9247 2792 9367 2836
rect 9247 2758 9290 2792
rect 9324 2758 9367 2792
rect 9247 2713 9367 2758
rect 9247 2679 9290 2713
rect 9324 2679 9367 2713
rect 9247 2634 9367 2679
rect 9247 2600 9290 2634
rect 9324 2600 9367 2634
rect 9809 3070 9852 3104
rect 9886 3070 9929 3104
rect 9809 3026 9929 3070
rect 9809 2992 9852 3026
rect 9886 2992 9929 3026
rect 9809 2948 9929 2992
rect 9809 2914 9852 2948
rect 9886 2914 9929 2948
rect 9809 2870 9929 2914
rect 9809 2836 9852 2870
rect 9886 2836 9929 2870
rect 9809 2792 9929 2836
rect 9809 2758 9852 2792
rect 9886 2758 9929 2792
rect 9809 2713 9929 2758
rect 9809 2679 9852 2713
rect 9886 2679 9929 2713
rect 9809 2634 9929 2679
rect 9247 2584 9367 2600
rect 9809 2600 9852 2634
rect 9886 2600 9929 2634
rect 9809 2584 9929 2600
rect 10239 3104 10359 3120
rect 10239 3070 10282 3104
rect 10316 3070 10359 3104
rect 10801 3104 10921 3120
rect 10239 3026 10359 3070
rect 10239 2992 10282 3026
rect 10316 2992 10359 3026
rect 10239 2948 10359 2992
rect 10239 2914 10282 2948
rect 10316 2914 10359 2948
rect 10239 2870 10359 2914
rect 10239 2836 10282 2870
rect 10316 2836 10359 2870
rect 10239 2792 10359 2836
rect 10239 2758 10282 2792
rect 10316 2758 10359 2792
rect 10239 2713 10359 2758
rect 10239 2679 10282 2713
rect 10316 2679 10359 2713
rect 10239 2634 10359 2679
rect 10239 2600 10282 2634
rect 10316 2600 10359 2634
rect 10801 3070 10844 3104
rect 10878 3070 10921 3104
rect 10801 3026 10921 3070
rect 10801 2992 10844 3026
rect 10878 2992 10921 3026
rect 10801 2948 10921 2992
rect 10801 2914 10844 2948
rect 10878 2914 10921 2948
rect 10801 2870 10921 2914
rect 10801 2836 10844 2870
rect 10878 2836 10921 2870
rect 10801 2792 10921 2836
rect 10801 2758 10844 2792
rect 10878 2758 10921 2792
rect 10801 2713 10921 2758
rect 10801 2679 10844 2713
rect 10878 2679 10921 2713
rect 10801 2634 10921 2679
rect 10239 2584 10359 2600
rect 10801 2600 10844 2634
rect 10878 2600 10921 2634
rect 10801 2584 10921 2600
rect 11231 3104 11351 3120
rect 11231 3070 11274 3104
rect 11308 3070 11351 3104
rect 11793 3104 11913 3120
rect 11231 3026 11351 3070
rect 11231 2992 11274 3026
rect 11308 2992 11351 3026
rect 11231 2948 11351 2992
rect 11231 2914 11274 2948
rect 11308 2914 11351 2948
rect 11231 2870 11351 2914
rect 11231 2836 11274 2870
rect 11308 2836 11351 2870
rect 11231 2792 11351 2836
rect 11231 2758 11274 2792
rect 11308 2758 11351 2792
rect 11231 2713 11351 2758
rect 11231 2679 11274 2713
rect 11308 2679 11351 2713
rect 11231 2634 11351 2679
rect 11231 2600 11274 2634
rect 11308 2600 11351 2634
rect 11793 3070 11836 3104
rect 11870 3070 11913 3104
rect 11793 3026 11913 3070
rect 11793 2992 11836 3026
rect 11870 2992 11913 3026
rect 11793 2948 11913 2992
rect 11793 2914 11836 2948
rect 11870 2914 11913 2948
rect 11793 2870 11913 2914
rect 11793 2836 11836 2870
rect 11870 2836 11913 2870
rect 11793 2792 11913 2836
rect 11793 2758 11836 2792
rect 11870 2758 11913 2792
rect 11793 2713 11913 2758
rect 11793 2679 11836 2713
rect 11870 2679 11913 2713
rect 11793 2634 11913 2679
rect 11231 2584 11351 2600
rect 11793 2600 11836 2634
rect 11870 2600 11913 2634
rect 11793 2584 11913 2600
rect 12223 3104 12343 3120
rect 12223 3070 12266 3104
rect 12300 3070 12343 3104
rect 12785 3104 12905 3120
rect 12223 3026 12343 3070
rect 12223 2992 12266 3026
rect 12300 2992 12343 3026
rect 12223 2948 12343 2992
rect 12223 2914 12266 2948
rect 12300 2914 12343 2948
rect 12223 2870 12343 2914
rect 12223 2836 12266 2870
rect 12300 2836 12343 2870
rect 12223 2792 12343 2836
rect 12223 2758 12266 2792
rect 12300 2758 12343 2792
rect 12223 2713 12343 2758
rect 12223 2679 12266 2713
rect 12300 2679 12343 2713
rect 12223 2634 12343 2679
rect 12223 2600 12266 2634
rect 12300 2600 12343 2634
rect 12785 3070 12828 3104
rect 12862 3070 12905 3104
rect 12785 3026 12905 3070
rect 12785 2992 12828 3026
rect 12862 2992 12905 3026
rect 12785 2948 12905 2992
rect 12785 2914 12828 2948
rect 12862 2914 12905 2948
rect 12785 2870 12905 2914
rect 12785 2836 12828 2870
rect 12862 2836 12905 2870
rect 12785 2792 12905 2836
rect 12785 2758 12828 2792
rect 12862 2758 12905 2792
rect 12785 2713 12905 2758
rect 12785 2679 12828 2713
rect 12862 2679 12905 2713
rect 12785 2634 12905 2679
rect 12223 2584 12343 2600
rect 12785 2600 12828 2634
rect 12862 2600 12905 2634
rect 12785 2584 12905 2600
rect 13215 3104 13335 3120
rect 13215 3070 13258 3104
rect 13292 3070 13335 3104
rect 13777 3104 13897 3120
rect 13215 3026 13335 3070
rect 13215 2992 13258 3026
rect 13292 2992 13335 3026
rect 13215 2948 13335 2992
rect 13215 2914 13258 2948
rect 13292 2914 13335 2948
rect 13215 2870 13335 2914
rect 13215 2836 13258 2870
rect 13292 2836 13335 2870
rect 13215 2792 13335 2836
rect 13215 2758 13258 2792
rect 13292 2758 13335 2792
rect 13215 2713 13335 2758
rect 13215 2679 13258 2713
rect 13292 2679 13335 2713
rect 13215 2634 13335 2679
rect 13215 2600 13258 2634
rect 13292 2600 13335 2634
rect 13777 3070 13820 3104
rect 13854 3070 13897 3104
rect 13777 3026 13897 3070
rect 13777 2992 13820 3026
rect 13854 2992 13897 3026
rect 13777 2948 13897 2992
rect 13777 2914 13820 2948
rect 13854 2914 13897 2948
rect 13777 2870 13897 2914
rect 13777 2836 13820 2870
rect 13854 2836 13897 2870
rect 13777 2792 13897 2836
rect 13777 2758 13820 2792
rect 13854 2758 13897 2792
rect 13777 2713 13897 2758
rect 13777 2679 13820 2713
rect 13854 2679 13897 2713
rect 13777 2634 13897 2679
rect 13215 2584 13335 2600
rect 13777 2600 13820 2634
rect 13854 2600 13897 2634
rect 13777 2584 13897 2600
rect 14135 3104 14255 3120
rect 14135 3070 14178 3104
rect 14212 3070 14255 3104
rect 14135 3026 14255 3070
rect 14135 2992 14178 3026
rect 14212 2992 14255 3026
rect 14135 2948 14255 2992
rect 14135 2914 14178 2948
rect 14212 2914 14255 2948
rect 14135 2870 14255 2914
rect 14135 2836 14178 2870
rect 14212 2836 14255 2870
rect 14135 2792 14255 2836
rect 14135 2758 14178 2792
rect 14212 2758 14255 2792
rect 14135 2713 14255 2758
rect 14135 2679 14178 2713
rect 14212 2679 14255 2713
rect 14135 2634 14255 2679
rect 14135 2600 14178 2634
rect 14212 2600 14255 2634
rect 14135 2584 14255 2600
rect 881 1504 1001 1520
rect 881 1470 924 1504
rect 958 1470 1001 1504
rect 881 1430 1001 1470
rect 881 1396 924 1430
rect 958 1396 1001 1430
rect 881 1380 1001 1396
rect 1311 1504 1431 1520
rect 1311 1470 1354 1504
rect 1388 1470 1431 1504
rect 1311 1430 1431 1470
rect 1311 1396 1354 1430
rect 1388 1396 1431 1430
rect 1311 1380 1431 1396
rect 1873 1504 1993 1520
rect 1873 1470 1916 1504
rect 1950 1470 1993 1504
rect 1873 1430 1993 1470
rect 1873 1396 1916 1430
rect 1950 1396 1993 1430
rect 1873 1380 1993 1396
rect 2303 1504 2423 1520
rect 2303 1470 2346 1504
rect 2380 1470 2423 1504
rect 2303 1430 2423 1470
rect 2303 1396 2346 1430
rect 2380 1396 2423 1430
rect 2303 1380 2423 1396
rect 2865 1504 2985 1520
rect 2865 1470 2908 1504
rect 2942 1470 2985 1504
rect 2865 1430 2985 1470
rect 2865 1396 2908 1430
rect 2942 1396 2985 1430
rect 2865 1380 2985 1396
rect 3295 1504 3415 1520
rect 3295 1470 3338 1504
rect 3372 1470 3415 1504
rect 3295 1430 3415 1470
rect 3295 1396 3338 1430
rect 3372 1396 3415 1430
rect 3295 1380 3415 1396
rect 3857 1504 3977 1520
rect 3857 1470 3900 1504
rect 3934 1470 3977 1504
rect 3857 1430 3977 1470
rect 3857 1396 3900 1430
rect 3934 1396 3977 1430
rect 3857 1380 3977 1396
rect 4287 1504 4407 1520
rect 4287 1470 4330 1504
rect 4364 1470 4407 1504
rect 4287 1430 4407 1470
rect 4287 1396 4330 1430
rect 4364 1396 4407 1430
rect 4287 1380 4407 1396
rect 4849 1504 4969 1520
rect 4849 1470 4892 1504
rect 4926 1470 4969 1504
rect 4849 1430 4969 1470
rect 4849 1396 4892 1430
rect 4926 1396 4969 1430
rect 4849 1380 4969 1396
rect 5279 1504 5399 1520
rect 5279 1470 5322 1504
rect 5356 1470 5399 1504
rect 5279 1430 5399 1470
rect 5279 1396 5322 1430
rect 5356 1396 5399 1430
rect 5279 1380 5399 1396
rect 5841 1504 5961 1520
rect 5841 1470 5884 1504
rect 5918 1470 5961 1504
rect 5841 1430 5961 1470
rect 5841 1396 5884 1430
rect 5918 1396 5961 1430
rect 5841 1380 5961 1396
rect 6271 1504 6391 1520
rect 6271 1470 6314 1504
rect 6348 1470 6391 1504
rect 6271 1430 6391 1470
rect 6271 1396 6314 1430
rect 6348 1396 6391 1430
rect 6271 1380 6391 1396
rect 6833 1504 6953 1520
rect 6833 1470 6876 1504
rect 6910 1470 6953 1504
rect 6833 1430 6953 1470
rect 6833 1396 6876 1430
rect 6910 1396 6953 1430
rect 6833 1380 6953 1396
rect 7263 1504 7383 1520
rect 7263 1470 7306 1504
rect 7340 1470 7383 1504
rect 7263 1430 7383 1470
rect 7263 1396 7306 1430
rect 7340 1396 7383 1430
rect 7263 1380 7383 1396
rect 7825 1504 7945 1520
rect 7825 1470 7868 1504
rect 7902 1470 7945 1504
rect 7825 1430 7945 1470
rect 7825 1396 7868 1430
rect 7902 1396 7945 1430
rect 7825 1380 7945 1396
rect 8255 1504 8375 1520
rect 8255 1470 8298 1504
rect 8332 1470 8375 1504
rect 8255 1430 8375 1470
rect 8255 1396 8298 1430
rect 8332 1396 8375 1430
rect 8255 1380 8375 1396
rect 8817 1504 8937 1520
rect 8817 1470 8860 1504
rect 8894 1470 8937 1504
rect 8817 1430 8937 1470
rect 8817 1396 8860 1430
rect 8894 1396 8937 1430
rect 8817 1380 8937 1396
rect 9247 1504 9367 1520
rect 9247 1470 9290 1504
rect 9324 1470 9367 1504
rect 9247 1430 9367 1470
rect 9247 1396 9290 1430
rect 9324 1396 9367 1430
rect 9247 1380 9367 1396
rect 9809 1504 9929 1520
rect 9809 1470 9852 1504
rect 9886 1470 9929 1504
rect 9809 1430 9929 1470
rect 9809 1396 9852 1430
rect 9886 1396 9929 1430
rect 9809 1380 9929 1396
rect 10239 1504 10359 1520
rect 10239 1470 10282 1504
rect 10316 1470 10359 1504
rect 10239 1430 10359 1470
rect 10239 1396 10282 1430
rect 10316 1396 10359 1430
rect 10239 1380 10359 1396
rect 10801 1504 10921 1520
rect 10801 1470 10844 1504
rect 10878 1470 10921 1504
rect 10801 1430 10921 1470
rect 10801 1396 10844 1430
rect 10878 1396 10921 1430
rect 10801 1380 10921 1396
rect 11231 1504 11351 1520
rect 11231 1470 11274 1504
rect 11308 1470 11351 1504
rect 11231 1430 11351 1470
rect 11231 1396 11274 1430
rect 11308 1396 11351 1430
rect 11231 1380 11351 1396
rect 11793 1504 11913 1520
rect 11793 1470 11836 1504
rect 11870 1470 11913 1504
rect 11793 1430 11913 1470
rect 11793 1396 11836 1430
rect 11870 1396 11913 1430
rect 11793 1380 11913 1396
rect 12223 1504 12343 1520
rect 12223 1470 12266 1504
rect 12300 1470 12343 1504
rect 12223 1430 12343 1470
rect 12223 1396 12266 1430
rect 12300 1396 12343 1430
rect 12223 1380 12343 1396
rect 12785 1504 12905 1520
rect 12785 1470 12828 1504
rect 12862 1470 12905 1504
rect 12785 1430 12905 1470
rect 12785 1396 12828 1430
rect 12862 1396 12905 1430
rect 12785 1380 12905 1396
rect 13215 1504 13335 1520
rect 13215 1470 13258 1504
rect 13292 1470 13335 1504
rect 13215 1430 13335 1470
rect 13215 1396 13258 1430
rect 13292 1396 13335 1430
rect 13215 1380 13335 1396
rect 13777 1504 13897 1520
rect 13777 1470 13820 1504
rect 13854 1470 13897 1504
rect 13777 1430 13897 1470
rect 13777 1396 13820 1430
rect 13854 1396 13897 1430
rect 13777 1380 13897 1396
rect 14135 1504 14255 1520
rect 14135 1470 14178 1504
rect 14212 1470 14255 1504
rect 14135 1430 14255 1470
rect 14135 1396 14178 1430
rect 14212 1396 14255 1430
rect 14135 1380 14255 1396
<< polycont >>
rect 924 4274 958 4308
rect 924 4200 958 4234
rect 1354 4274 1388 4308
rect 1354 4200 1388 4234
rect 1916 4274 1950 4308
rect 1916 4200 1950 4234
rect 2346 4274 2380 4308
rect 2346 4200 2380 4234
rect 2908 4274 2942 4308
rect 2908 4200 2942 4234
rect 3338 4274 3372 4308
rect 3338 4200 3372 4234
rect 3900 4274 3934 4308
rect 3900 4200 3934 4234
rect 4330 4274 4364 4308
rect 4330 4200 4364 4234
rect 4892 4274 4926 4308
rect 4892 4200 4926 4234
rect 5322 4274 5356 4308
rect 5322 4200 5356 4234
rect 5884 4274 5918 4308
rect 5884 4200 5918 4234
rect 6314 4274 6348 4308
rect 6314 4200 6348 4234
rect 6876 4274 6910 4308
rect 6876 4200 6910 4234
rect 7306 4274 7340 4308
rect 7306 4200 7340 4234
rect 7868 4274 7902 4308
rect 7868 4200 7902 4234
rect 8298 4274 8332 4308
rect 8298 4200 8332 4234
rect 8860 4274 8894 4308
rect 8860 4200 8894 4234
rect 9290 4274 9324 4308
rect 9290 4200 9324 4234
rect 9852 4274 9886 4308
rect 9852 4200 9886 4234
rect 10282 4274 10316 4308
rect 10282 4200 10316 4234
rect 10844 4274 10878 4308
rect 10844 4200 10878 4234
rect 11274 4274 11308 4308
rect 11274 4200 11308 4234
rect 11836 4274 11870 4308
rect 11836 4200 11870 4234
rect 12266 4274 12300 4308
rect 12266 4200 12300 4234
rect 12828 4274 12862 4308
rect 12828 4200 12862 4234
rect 13258 4274 13292 4308
rect 13258 4200 13292 4234
rect 13820 4274 13854 4308
rect 13820 4200 13854 4234
rect 14178 4274 14212 4308
rect 14178 4200 14212 4234
rect 924 3070 958 3104
rect 924 2992 958 3026
rect 924 2914 958 2948
rect 924 2836 958 2870
rect 924 2758 958 2792
rect 924 2679 958 2713
rect 924 2600 958 2634
rect 1354 3070 1388 3104
rect 1354 2992 1388 3026
rect 1354 2914 1388 2948
rect 1354 2836 1388 2870
rect 1354 2758 1388 2792
rect 1354 2679 1388 2713
rect 1354 2600 1388 2634
rect 1916 3070 1950 3104
rect 1916 2992 1950 3026
rect 1916 2914 1950 2948
rect 1916 2836 1950 2870
rect 1916 2758 1950 2792
rect 1916 2679 1950 2713
rect 1916 2600 1950 2634
rect 2346 3070 2380 3104
rect 2346 2992 2380 3026
rect 2346 2914 2380 2948
rect 2346 2836 2380 2870
rect 2346 2758 2380 2792
rect 2346 2679 2380 2713
rect 2346 2600 2380 2634
rect 2908 3070 2942 3104
rect 2908 2992 2942 3026
rect 2908 2914 2942 2948
rect 2908 2836 2942 2870
rect 2908 2758 2942 2792
rect 2908 2679 2942 2713
rect 2908 2600 2942 2634
rect 3338 3070 3372 3104
rect 3338 2992 3372 3026
rect 3338 2914 3372 2948
rect 3338 2836 3372 2870
rect 3338 2758 3372 2792
rect 3338 2679 3372 2713
rect 3338 2600 3372 2634
rect 3900 3070 3934 3104
rect 3900 2992 3934 3026
rect 3900 2914 3934 2948
rect 3900 2836 3934 2870
rect 3900 2758 3934 2792
rect 3900 2679 3934 2713
rect 3900 2600 3934 2634
rect 4330 3070 4364 3104
rect 4330 2992 4364 3026
rect 4330 2914 4364 2948
rect 4330 2836 4364 2870
rect 4330 2758 4364 2792
rect 4330 2679 4364 2713
rect 4330 2600 4364 2634
rect 4892 3070 4926 3104
rect 4892 2992 4926 3026
rect 4892 2914 4926 2948
rect 4892 2836 4926 2870
rect 4892 2758 4926 2792
rect 4892 2679 4926 2713
rect 4892 2600 4926 2634
rect 5322 3070 5356 3104
rect 5322 2992 5356 3026
rect 5322 2914 5356 2948
rect 5322 2836 5356 2870
rect 5322 2758 5356 2792
rect 5322 2679 5356 2713
rect 5322 2600 5356 2634
rect 5884 3070 5918 3104
rect 5884 2992 5918 3026
rect 5884 2914 5918 2948
rect 5884 2836 5918 2870
rect 5884 2758 5918 2792
rect 5884 2679 5918 2713
rect 5884 2600 5918 2634
rect 6314 3070 6348 3104
rect 6314 2992 6348 3026
rect 6314 2914 6348 2948
rect 6314 2836 6348 2870
rect 6314 2758 6348 2792
rect 6314 2679 6348 2713
rect 6314 2600 6348 2634
rect 6876 3070 6910 3104
rect 6876 2992 6910 3026
rect 6876 2914 6910 2948
rect 6876 2836 6910 2870
rect 6876 2758 6910 2792
rect 6876 2679 6910 2713
rect 6876 2600 6910 2634
rect 7306 3070 7340 3104
rect 7306 2992 7340 3026
rect 7306 2914 7340 2948
rect 7306 2836 7340 2870
rect 7306 2758 7340 2792
rect 7306 2679 7340 2713
rect 7306 2600 7340 2634
rect 7868 3070 7902 3104
rect 7868 2992 7902 3026
rect 7868 2914 7902 2948
rect 7868 2836 7902 2870
rect 7868 2758 7902 2792
rect 7868 2679 7902 2713
rect 7868 2600 7902 2634
rect 8298 3070 8332 3104
rect 8298 2992 8332 3026
rect 8298 2914 8332 2948
rect 8298 2836 8332 2870
rect 8298 2758 8332 2792
rect 8298 2679 8332 2713
rect 8298 2600 8332 2634
rect 8860 3070 8894 3104
rect 8860 2992 8894 3026
rect 8860 2914 8894 2948
rect 8860 2836 8894 2870
rect 8860 2758 8894 2792
rect 8860 2679 8894 2713
rect 8860 2600 8894 2634
rect 9290 3070 9324 3104
rect 9290 2992 9324 3026
rect 9290 2914 9324 2948
rect 9290 2836 9324 2870
rect 9290 2758 9324 2792
rect 9290 2679 9324 2713
rect 9290 2600 9324 2634
rect 9852 3070 9886 3104
rect 9852 2992 9886 3026
rect 9852 2914 9886 2948
rect 9852 2836 9886 2870
rect 9852 2758 9886 2792
rect 9852 2679 9886 2713
rect 9852 2600 9886 2634
rect 10282 3070 10316 3104
rect 10282 2992 10316 3026
rect 10282 2914 10316 2948
rect 10282 2836 10316 2870
rect 10282 2758 10316 2792
rect 10282 2679 10316 2713
rect 10282 2600 10316 2634
rect 10844 3070 10878 3104
rect 10844 2992 10878 3026
rect 10844 2914 10878 2948
rect 10844 2836 10878 2870
rect 10844 2758 10878 2792
rect 10844 2679 10878 2713
rect 10844 2600 10878 2634
rect 11274 3070 11308 3104
rect 11274 2992 11308 3026
rect 11274 2914 11308 2948
rect 11274 2836 11308 2870
rect 11274 2758 11308 2792
rect 11274 2679 11308 2713
rect 11274 2600 11308 2634
rect 11836 3070 11870 3104
rect 11836 2992 11870 3026
rect 11836 2914 11870 2948
rect 11836 2836 11870 2870
rect 11836 2758 11870 2792
rect 11836 2679 11870 2713
rect 11836 2600 11870 2634
rect 12266 3070 12300 3104
rect 12266 2992 12300 3026
rect 12266 2914 12300 2948
rect 12266 2836 12300 2870
rect 12266 2758 12300 2792
rect 12266 2679 12300 2713
rect 12266 2600 12300 2634
rect 12828 3070 12862 3104
rect 12828 2992 12862 3026
rect 12828 2914 12862 2948
rect 12828 2836 12862 2870
rect 12828 2758 12862 2792
rect 12828 2679 12862 2713
rect 12828 2600 12862 2634
rect 13258 3070 13292 3104
rect 13258 2992 13292 3026
rect 13258 2914 13292 2948
rect 13258 2836 13292 2870
rect 13258 2758 13292 2792
rect 13258 2679 13292 2713
rect 13258 2600 13292 2634
rect 13820 3070 13854 3104
rect 13820 2992 13854 3026
rect 13820 2914 13854 2948
rect 13820 2836 13854 2870
rect 13820 2758 13854 2792
rect 13820 2679 13854 2713
rect 13820 2600 13854 2634
rect 14178 3070 14212 3104
rect 14178 2992 14212 3026
rect 14178 2914 14212 2948
rect 14178 2836 14212 2870
rect 14178 2758 14212 2792
rect 14178 2679 14212 2713
rect 14178 2600 14212 2634
rect 924 1470 958 1504
rect 924 1396 958 1430
rect 1354 1470 1388 1504
rect 1354 1396 1388 1430
rect 1916 1470 1950 1504
rect 1916 1396 1950 1430
rect 2346 1470 2380 1504
rect 2346 1396 2380 1430
rect 2908 1470 2942 1504
rect 2908 1396 2942 1430
rect 3338 1470 3372 1504
rect 3338 1396 3372 1430
rect 3900 1470 3934 1504
rect 3900 1396 3934 1430
rect 4330 1470 4364 1504
rect 4330 1396 4364 1430
rect 4892 1470 4926 1504
rect 4892 1396 4926 1430
rect 5322 1470 5356 1504
rect 5322 1396 5356 1430
rect 5884 1470 5918 1504
rect 5884 1396 5918 1430
rect 6314 1470 6348 1504
rect 6314 1396 6348 1430
rect 6876 1470 6910 1504
rect 6876 1396 6910 1430
rect 7306 1470 7340 1504
rect 7306 1396 7340 1430
rect 7868 1470 7902 1504
rect 7868 1396 7902 1430
rect 8298 1470 8332 1504
rect 8298 1396 8332 1430
rect 8860 1470 8894 1504
rect 8860 1396 8894 1430
rect 9290 1470 9324 1504
rect 9290 1396 9324 1430
rect 9852 1470 9886 1504
rect 9852 1396 9886 1430
rect 10282 1470 10316 1504
rect 10282 1396 10316 1430
rect 10844 1470 10878 1504
rect 10844 1396 10878 1430
rect 11274 1470 11308 1504
rect 11274 1396 11308 1430
rect 11836 1470 11870 1504
rect 11836 1396 11870 1430
rect 12266 1470 12300 1504
rect 12266 1396 12300 1430
rect 12828 1470 12862 1504
rect 12828 1396 12862 1430
rect 13258 1470 13292 1504
rect 13258 1396 13292 1430
rect 13820 1470 13854 1504
rect 13820 1396 13854 1430
rect 14178 1470 14212 1504
rect 14178 1396 14212 1430
<< locali >>
rect 36 5111 15051 5118
rect 36 5083 361 5111
rect 121 5021 223 5083
rect 329 5077 361 5083
rect 395 5077 434 5111
rect 468 5077 507 5111
rect 541 5077 580 5111
rect 614 5077 653 5111
rect 687 5077 726 5111
rect 760 5077 799 5111
rect 833 5077 872 5111
rect 906 5077 945 5111
rect 979 5077 1018 5111
rect 1052 5077 1091 5111
rect 1125 5077 1164 5111
rect 1198 5077 1237 5111
rect 1271 5077 1310 5111
rect 1344 5077 1383 5111
rect 1417 5077 1456 5111
rect 1490 5077 1529 5111
rect 1563 5077 1602 5111
rect 1636 5077 1675 5111
rect 1709 5077 1748 5111
rect 1782 5077 1821 5111
rect 1855 5077 1894 5111
rect 1928 5077 1967 5111
rect 2001 5077 2040 5111
rect 2074 5077 2113 5111
rect 2147 5077 2186 5111
rect 2220 5077 2259 5111
rect 2293 5077 2332 5111
rect 2366 5077 2405 5111
rect 2439 5077 2478 5111
rect 2512 5077 2551 5111
rect 2585 5077 2624 5111
rect 2658 5077 2697 5111
rect 2731 5077 2770 5111
rect 2804 5077 2843 5111
rect 2877 5077 2916 5111
rect 2950 5077 2989 5111
rect 3023 5077 3062 5111
rect 3096 5077 3135 5111
rect 3169 5077 3208 5111
rect 3242 5077 3281 5111
rect 3315 5077 3354 5111
rect 3388 5077 3427 5111
rect 3461 5077 3500 5111
rect 3534 5077 3573 5111
rect 3607 5077 3646 5111
rect 3680 5077 3719 5111
rect 3753 5077 3792 5111
rect 3826 5077 3865 5111
rect 3899 5077 3938 5111
rect 3972 5077 4011 5111
rect 4045 5077 4084 5111
rect 4118 5077 4157 5111
rect 4191 5077 4229 5111
rect 4263 5077 4301 5111
rect 4335 5077 4373 5111
rect 4407 5077 4445 5111
rect 4479 5077 4517 5111
rect 4551 5077 4589 5111
rect 4623 5077 4661 5111
rect 4695 5077 4733 5111
rect 4767 5077 4805 5111
rect 4839 5077 4877 5111
rect 4911 5077 4949 5111
rect 4983 5077 5021 5111
rect 5055 5077 5093 5111
rect 5127 5077 5165 5111
rect 5199 5077 5237 5111
rect 5271 5077 5309 5111
rect 5343 5077 5381 5111
rect 5415 5077 5453 5111
rect 5487 5077 5525 5111
rect 5559 5077 5597 5111
rect 5631 5077 5669 5111
rect 5703 5077 5741 5111
rect 5775 5077 5813 5111
rect 5847 5077 5885 5111
rect 5919 5077 5957 5111
rect 5991 5077 6029 5111
rect 6063 5077 6101 5111
rect 6135 5077 6173 5111
rect 6207 5077 6245 5111
rect 6279 5077 6317 5111
rect 6351 5077 6389 5111
rect 6423 5077 6461 5111
rect 6495 5077 6533 5111
rect 6567 5077 6605 5111
rect 6639 5077 6677 5111
rect 6711 5077 6749 5111
rect 6783 5077 6821 5111
rect 6855 5077 6893 5111
rect 6927 5077 6965 5111
rect 6999 5077 7037 5111
rect 7071 5077 7109 5111
rect 7143 5077 7181 5111
rect 7215 5077 7253 5111
rect 7287 5077 7325 5111
rect 7359 5077 7397 5111
rect 7431 5077 7469 5111
rect 7503 5077 7541 5111
rect 7575 5077 7613 5111
rect 7647 5077 7685 5111
rect 7719 5077 7757 5111
rect 7791 5077 7829 5111
rect 7863 5077 7901 5111
rect 7935 5077 7973 5111
rect 8007 5077 8045 5111
rect 8079 5077 8117 5111
rect 8151 5077 8189 5111
rect 8223 5077 8261 5111
rect 8295 5077 8333 5111
rect 8367 5077 8405 5111
rect 8439 5077 8477 5111
rect 8511 5077 8549 5111
rect 8583 5077 8621 5111
rect 8655 5077 8693 5111
rect 8727 5077 8765 5111
rect 8799 5077 8837 5111
rect 8871 5077 8909 5111
rect 8943 5077 8981 5111
rect 9015 5077 9053 5111
rect 9087 5077 9125 5111
rect 9159 5077 9197 5111
rect 9231 5077 9269 5111
rect 9303 5077 9341 5111
rect 9375 5077 9413 5111
rect 9447 5077 9485 5111
rect 9519 5077 9557 5111
rect 9591 5077 9629 5111
rect 9663 5077 9701 5111
rect 9735 5077 9773 5111
rect 9807 5077 9845 5111
rect 9879 5077 9917 5111
rect 9951 5077 9989 5111
rect 10023 5077 10061 5111
rect 10095 5077 10133 5111
rect 10167 5077 10205 5111
rect 10239 5077 10277 5111
rect 10311 5077 10349 5111
rect 10383 5077 10421 5111
rect 10455 5077 10493 5111
rect 10527 5077 10565 5111
rect 10599 5077 10637 5111
rect 10671 5077 10709 5111
rect 10743 5077 10781 5111
rect 10815 5077 10853 5111
rect 10887 5077 10925 5111
rect 10959 5077 10997 5111
rect 11031 5077 11069 5111
rect 11103 5077 11141 5111
rect 11175 5077 11213 5111
rect 11247 5077 11285 5111
rect 11319 5077 11357 5111
rect 11391 5077 11429 5111
rect 11463 5077 11501 5111
rect 11535 5077 11573 5111
rect 11607 5077 11645 5111
rect 11679 5077 11717 5111
rect 11751 5077 11789 5111
rect 11823 5077 11861 5111
rect 11895 5077 11933 5111
rect 11967 5077 12005 5111
rect 12039 5077 12077 5111
rect 12111 5077 12149 5111
rect 12183 5077 12221 5111
rect 12255 5077 12293 5111
rect 12327 5077 12365 5111
rect 12399 5077 12437 5111
rect 12471 5077 12509 5111
rect 12543 5077 12581 5111
rect 12615 5077 12653 5111
rect 12687 5077 12725 5111
rect 12759 5077 12797 5111
rect 12831 5077 12869 5111
rect 12903 5077 12941 5111
rect 12975 5077 13013 5111
rect 13047 5077 13085 5111
rect 13119 5077 13157 5111
rect 13191 5077 13229 5111
rect 13263 5077 13301 5111
rect 13335 5077 13373 5111
rect 13407 5077 13445 5111
rect 13479 5077 13517 5111
rect 13551 5077 13589 5111
rect 13623 5077 13661 5111
rect 13695 5077 13733 5111
rect 13767 5077 13805 5111
rect 13839 5077 13877 5111
rect 13911 5077 13949 5111
rect 13983 5077 14021 5111
rect 14055 5077 14093 5111
rect 14127 5077 14165 5111
rect 14199 5077 14237 5111
rect 14271 5077 14309 5111
rect 14343 5077 14381 5111
rect 14415 5077 14453 5111
rect 14487 5077 14525 5111
rect 14559 5077 14597 5111
rect 14631 5077 14669 5111
rect 14703 5077 14741 5111
rect 14775 5083 15051 5111
rect 14775 5077 14807 5083
rect 329 5068 14807 5077
rect 272 5029 306 5068
rect 13600 5035 13635 5068
rect 13669 5035 13704 5068
rect 13738 5035 13773 5068
rect 13807 5035 13842 5068
rect 267 4995 269 5029
rect 303 4995 306 5029
rect 13623 5034 13635 5035
rect 13695 5034 13704 5035
rect 13767 5034 13773 5035
rect 13839 5034 13842 5035
rect 13876 5035 13911 5068
rect 13876 5034 13877 5035
rect 13623 5001 13661 5034
rect 13695 5001 13733 5034
rect 13767 5001 13805 5034
rect 13839 5001 13877 5034
rect 13945 5035 13980 5068
rect 14014 5035 14049 5068
rect 14083 5035 14118 5068
rect 14152 5035 14187 5068
rect 14221 5035 14256 5068
rect 14290 5035 14325 5068
rect 14359 5035 14394 5068
rect 14428 5035 14463 5068
rect 14497 5035 14532 5068
rect 14566 5035 14601 5068
rect 14635 5035 14670 5068
rect 13945 5034 13949 5035
rect 14014 5034 14021 5035
rect 14083 5034 14093 5035
rect 14152 5034 14165 5035
rect 14221 5034 14237 5035
rect 14290 5034 14309 5035
rect 14359 5034 14381 5035
rect 14428 5034 14453 5035
rect 14497 5034 14525 5035
rect 14566 5034 14597 5035
rect 14635 5034 14669 5035
rect 14704 5034 14739 5068
rect 14773 5057 14807 5068
rect 14773 5035 14907 5057
rect 13911 5001 13949 5034
rect 13983 5001 14021 5034
rect 14055 5001 14093 5034
rect 14127 5001 14165 5034
rect 14199 5001 14237 5034
rect 14271 5001 14309 5034
rect 14343 5001 14381 5034
rect 14415 5001 14453 5034
rect 14487 5001 14525 5034
rect 14559 5001 14597 5034
rect 14631 5001 14669 5034
rect 14703 5001 14741 5034
rect 14775 5033 14907 5035
rect 14775 5030 14840 5033
rect 14775 5001 14832 5030
rect 267 4956 306 4995
rect 13600 5000 14832 5001
rect 13600 4966 13635 5000
rect 13669 4966 13704 5000
rect 13738 4966 13773 5000
rect 13807 4966 13842 5000
rect 13876 4966 13911 5000
rect 13945 4966 13980 5000
rect 14014 4966 14049 5000
rect 14083 4966 14118 5000
rect 14152 4966 14187 5000
rect 14221 4966 14256 5000
rect 14290 4966 14325 5000
rect 14359 4966 14394 5000
rect 14428 4966 14463 5000
rect 14497 4966 14532 5000
rect 14566 4966 14601 5000
rect 14635 4966 14670 5000
rect 14704 4966 14739 5000
rect 14773 4996 14832 5000
rect 14874 5021 14907 5033
rect 14927 5021 15051 5083
rect 14874 4999 15051 5021
rect 14866 4996 15051 4999
rect 14773 4966 15051 4996
rect 13600 4965 15051 4966
rect 13600 4959 14840 4965
rect 267 4922 269 4956
rect 303 4922 306 4956
rect 13623 4932 13661 4959
rect 13695 4932 13733 4959
rect 13767 4932 13805 4959
rect 13839 4932 13877 4959
rect 13623 4925 13635 4932
rect 13695 4925 13704 4932
rect 13767 4925 13773 4932
rect 13839 4925 13842 4932
rect 267 4898 306 4922
rect 13600 4898 13635 4925
rect 13669 4898 13704 4925
rect 13738 4898 13773 4925
rect 13807 4898 13842 4925
rect 13876 4925 13877 4932
rect 13911 4932 13949 4959
rect 13983 4932 14021 4959
rect 14055 4932 14093 4959
rect 14127 4932 14165 4959
rect 14199 4932 14237 4959
rect 14271 4932 14309 4959
rect 14343 4932 14381 4959
rect 14415 4932 14453 4959
rect 14487 4932 14525 4959
rect 14559 4932 14597 4959
rect 14631 4932 14669 4959
rect 14703 4932 14741 4959
rect 14775 4958 14840 4959
rect 13876 4898 13911 4925
rect 13945 4925 13949 4932
rect 14014 4925 14021 4932
rect 14083 4925 14093 4932
rect 14152 4925 14165 4932
rect 14221 4925 14237 4932
rect 14290 4925 14309 4932
rect 14359 4925 14381 4932
rect 14428 4925 14453 4932
rect 14497 4925 14525 4932
rect 14566 4925 14597 4932
rect 14635 4925 14669 4932
rect 13945 4898 13980 4925
rect 14014 4898 14049 4925
rect 14083 4898 14118 4925
rect 14152 4898 14187 4925
rect 14221 4898 14256 4925
rect 14290 4898 14325 4925
rect 14359 4898 14394 4925
rect 14428 4898 14463 4925
rect 14497 4898 14532 4925
rect 14566 4898 14601 4925
rect 14635 4898 14670 4925
rect 14704 4898 14739 4932
rect 14775 4925 14832 4958
rect 14773 4924 14832 4925
rect 14773 4898 14840 4924
rect 267 4883 305 4898
rect 14807 4886 14840 4898
rect 229 4859 269 4883
rect 229 4825 262 4859
rect 303 4849 329 4883
rect 296 4825 329 4849
rect 229 4810 329 4825
rect 229 4791 269 4810
rect 229 4757 262 4791
rect 303 4776 329 4810
rect 296 4757 329 4776
rect 229 4737 329 4757
rect 229 4723 269 4737
rect 229 4689 262 4723
rect 303 4703 329 4737
rect 296 4689 329 4703
rect 229 4664 329 4689
rect 229 4655 269 4664
rect 229 4621 262 4655
rect 303 4630 329 4664
rect 14807 4852 14832 4886
rect 14807 4814 14840 4852
rect 14807 4780 14832 4814
rect 14807 4742 14840 4780
rect 14807 4708 14832 4742
rect 14807 4670 14840 4708
rect 296 4621 329 4630
rect 229 4591 329 4621
rect 229 4587 269 4591
rect 229 4553 262 4587
rect 303 4557 329 4591
rect 296 4553 329 4557
rect 229 4519 329 4553
rect 229 4485 262 4519
rect 296 4518 329 4519
rect 229 4484 269 4485
rect 303 4484 329 4518
rect 229 4451 329 4484
rect 229 4417 262 4451
rect 296 4445 329 4451
rect 229 4411 269 4417
rect 303 4411 329 4445
rect 229 4383 329 4411
rect 229 4349 262 4383
rect 296 4372 329 4383
rect 229 4338 269 4349
rect 303 4338 329 4372
rect 229 4315 329 4338
rect 229 4281 262 4315
rect 296 4299 329 4315
rect 229 4265 269 4281
rect 303 4265 329 4299
rect 229 4247 329 4265
rect 229 4213 262 4247
rect 296 4226 329 4247
rect 229 4192 269 4213
rect 303 4192 329 4226
rect 229 4179 329 4192
rect 229 4145 262 4179
rect 296 4153 329 4179
rect 229 4119 269 4145
rect 303 4119 329 4153
rect 229 4111 329 4119
rect 229 4077 262 4111
rect 296 4080 329 4111
rect 229 4046 269 4077
rect 303 4046 329 4080
rect 229 4043 329 4046
rect 229 4009 262 4043
rect 296 4009 329 4043
rect 229 4007 329 4009
rect 229 3975 269 4007
rect 229 3941 262 3975
rect 303 3973 329 4007
rect 296 3941 329 3973
rect 229 3934 329 3941
rect 229 3907 269 3934
rect 229 3873 262 3907
rect 303 3900 329 3934
rect 296 3873 329 3900
rect 229 3861 329 3873
rect 229 3839 269 3861
rect 229 3805 262 3839
rect 303 3827 329 3861
rect 296 3805 329 3827
rect 229 3788 329 3805
rect 229 3771 269 3788
rect 229 3737 262 3771
rect 303 3754 329 3788
rect 296 3737 329 3754
rect 229 3715 329 3737
rect 229 3703 269 3715
rect 229 3669 262 3703
rect 303 3681 329 3715
rect 296 3669 329 3681
rect 229 3642 329 3669
rect 229 3635 269 3642
rect 229 3601 262 3635
rect 303 3608 329 3642
rect 296 3601 329 3608
rect 229 3569 329 3601
rect 229 3567 269 3569
rect 229 3533 262 3567
rect 303 3535 329 3569
rect 296 3533 329 3535
rect 229 3499 329 3533
rect 229 3465 262 3499
rect 296 3496 329 3499
rect 229 3462 269 3465
rect 303 3462 329 3496
rect 229 3431 329 3462
rect 229 3397 262 3431
rect 296 3423 329 3431
rect 229 3389 269 3397
rect 303 3389 329 3423
rect 229 3363 329 3389
rect 229 3329 262 3363
rect 296 3350 329 3363
rect 229 3316 269 3329
rect 303 3316 329 3350
rect 229 3295 329 3316
rect 229 3261 262 3295
rect 296 3277 329 3295
rect 229 3243 269 3261
rect 303 3243 329 3277
rect 229 3227 329 3243
rect 229 3193 262 3227
rect 296 3204 329 3227
rect 229 3170 269 3193
rect 303 3170 329 3204
rect 229 3159 329 3170
rect 229 3125 262 3159
rect 296 3131 329 3159
rect 229 3097 269 3125
rect 303 3097 329 3131
rect 229 3091 329 3097
rect 229 3057 262 3091
rect 296 3058 329 3091
rect 229 3024 269 3057
rect 303 3024 329 3058
rect 229 3023 329 3024
rect 229 2989 262 3023
rect 296 2989 329 3023
rect 229 2985 329 2989
rect 229 2955 269 2985
rect 229 2921 262 2955
rect 303 2951 329 2985
rect 296 2921 329 2951
rect 229 2912 329 2921
rect 229 2887 269 2912
rect 229 2853 262 2887
rect 303 2878 329 2912
rect 296 2853 329 2878
rect 229 2839 329 2853
rect 229 2819 269 2839
rect 229 2785 262 2819
rect 303 2805 329 2839
rect 296 2785 329 2805
rect 229 2766 329 2785
rect 229 2751 269 2766
rect 229 2717 262 2751
rect 303 2732 329 2766
rect 296 2717 329 2732
rect 229 2693 329 2717
rect 229 2683 269 2693
rect 229 2649 262 2683
rect 303 2659 329 2693
rect 296 2649 329 2659
rect 229 2620 329 2649
rect 229 2615 269 2620
rect 229 2581 262 2615
rect 303 2586 329 2620
rect 296 2581 329 2586
rect 229 2547 329 2581
rect 229 2513 262 2547
rect 303 2513 329 2547
rect 229 2479 329 2513
rect 229 2445 262 2479
rect 296 2474 329 2479
rect 229 2440 269 2445
rect 303 2440 329 2474
rect 229 2411 329 2440
rect 229 2377 262 2411
rect 296 2401 329 2411
rect 229 2367 269 2377
rect 303 2367 329 2401
rect 229 2343 329 2367
rect 229 2309 262 2343
rect 296 2328 329 2343
rect 229 2294 269 2309
rect 303 2294 329 2328
rect 229 2275 329 2294
rect 229 2241 262 2275
rect 296 2255 329 2275
rect 229 2221 269 2241
rect 303 2221 329 2255
rect 229 2207 329 2221
rect 229 2173 262 2207
rect 296 2182 329 2207
rect 229 2148 269 2173
rect 303 2148 329 2182
rect 229 2139 329 2148
rect 229 2105 262 2139
rect 296 2109 329 2139
rect 229 2075 269 2105
rect 303 2075 329 2109
rect 229 2071 329 2075
rect 229 2037 262 2071
rect 296 2037 329 2071
rect 229 2036 329 2037
rect 229 2003 269 2036
rect 229 1969 262 2003
rect 303 2002 329 2036
rect 296 1969 329 2002
rect 229 1963 329 1969
rect 229 1935 269 1963
rect 229 1901 262 1935
rect 303 1929 329 1963
rect 296 1901 329 1929
rect 229 1890 329 1901
rect 229 1867 269 1890
rect 229 1833 262 1867
rect 303 1856 329 1890
rect 296 1833 329 1856
rect 229 1817 329 1833
rect 229 1799 269 1817
rect 229 1765 262 1799
rect 303 1783 329 1817
rect 296 1765 329 1783
rect 229 1744 329 1765
rect 229 1731 269 1744
rect 229 1697 262 1731
rect 303 1710 329 1744
rect 296 1697 329 1710
rect 229 1671 329 1697
rect 229 1663 269 1671
rect 229 1629 262 1663
rect 303 1637 329 1671
rect 296 1629 329 1637
rect 229 1598 329 1629
rect 229 1595 269 1598
rect 229 1561 262 1595
rect 303 1564 329 1598
rect 296 1561 329 1564
rect 229 1527 329 1561
rect 229 1493 262 1527
rect 296 1525 329 1527
rect 229 1491 269 1493
rect 303 1491 329 1525
rect 229 1459 329 1491
rect 229 1425 262 1459
rect 296 1452 329 1459
rect 229 1418 269 1425
rect 303 1418 329 1452
rect 229 1391 329 1418
rect 229 1357 262 1391
rect 296 1379 329 1391
rect 229 1345 269 1357
rect 303 1345 329 1379
rect 229 1323 329 1345
rect 229 1289 262 1323
rect 296 1306 329 1323
rect 229 1272 269 1289
rect 303 1272 329 1306
rect 229 1255 329 1272
rect 229 1221 262 1255
rect 296 1233 329 1255
rect 229 1199 269 1221
rect 303 1199 329 1233
rect 229 1187 329 1199
rect 229 1153 262 1187
rect 296 1159 329 1187
rect 229 1125 269 1153
rect 303 1125 329 1159
rect 229 1119 329 1125
rect 229 1085 262 1119
rect 296 1085 329 1119
rect 229 1051 269 1085
rect 303 1051 329 1085
rect 229 1017 262 1051
rect 296 1017 329 1051
rect 229 1011 329 1017
rect 229 983 269 1011
rect 229 949 262 983
rect 303 977 329 1011
rect 296 949 329 977
rect 229 937 329 949
rect 229 915 269 937
rect 229 881 262 915
rect 303 903 329 937
rect 296 881 329 903
rect 229 863 329 881
rect 229 847 269 863
rect 229 813 262 847
rect 303 829 329 863
rect 296 813 329 829
rect 229 789 329 813
rect 229 779 269 789
rect 229 745 262 779
rect 303 755 329 789
rect 296 745 329 755
rect 229 715 329 745
rect 229 711 269 715
rect 229 677 262 711
rect 303 681 329 715
rect 296 677 329 681
rect 229 643 329 677
rect 482 4638 14653 4653
rect 482 4619 584 4638
rect 482 4585 497 4619
rect 531 4585 584 4619
rect 10410 4606 10445 4638
rect 10479 4606 10514 4638
rect 10548 4606 10583 4638
rect 10617 4606 10652 4638
rect 10686 4606 10721 4638
rect 10755 4606 10790 4638
rect 10824 4606 10859 4638
rect 10893 4606 10928 4638
rect 10962 4606 10997 4638
rect 11031 4606 11066 4638
rect 11100 4606 11135 4638
rect 11169 4606 11204 4638
rect 11238 4606 11273 4638
rect 11307 4606 11342 4638
rect 11376 4606 11411 4638
rect 11445 4606 11480 4638
rect 11514 4606 11549 4638
rect 11583 4606 11618 4638
rect 11652 4606 11687 4638
rect 11721 4606 11756 4638
rect 11790 4606 11825 4638
rect 11859 4606 11894 4638
rect 11928 4606 11963 4638
rect 11997 4606 12032 4638
rect 12066 4606 12101 4638
rect 12135 4606 12170 4638
rect 12204 4606 12239 4638
rect 12273 4606 12308 4638
rect 12342 4606 12377 4638
rect 12411 4606 12446 4638
rect 12480 4606 12515 4638
rect 12549 4606 12584 4638
rect 12618 4606 12653 4638
rect 12687 4606 12722 4638
rect 12756 4606 12791 4638
rect 12825 4606 12860 4638
rect 12894 4606 12929 4638
rect 12963 4606 12998 4638
rect 13032 4606 13067 4638
rect 13101 4606 13136 4638
rect 13170 4606 13205 4638
rect 13239 4606 13274 4638
rect 13308 4606 13343 4638
rect 13377 4606 13412 4638
rect 13446 4606 13481 4638
rect 13515 4606 13550 4638
rect 13584 4606 13619 4638
rect 13653 4606 13688 4638
rect 13722 4606 13757 4638
rect 13791 4606 13826 4638
rect 13860 4606 13895 4638
rect 13929 4606 13964 4638
rect 13998 4606 14033 4638
rect 14067 4606 14102 4638
rect 14136 4606 14171 4638
rect 14205 4606 14240 4638
rect 14274 4606 14309 4638
rect 14343 4606 14378 4638
rect 14412 4606 14447 4638
rect 482 4570 584 4585
rect 14207 4604 14240 4606
rect 14280 4604 14309 4606
rect 14353 4604 14378 4606
rect 14426 4604 14447 4606
rect 14481 4604 14516 4638
rect 14550 4604 14585 4638
rect 14619 4604 14653 4638
rect 14207 4572 14246 4604
rect 14280 4572 14319 4604
rect 14353 4572 14392 4604
rect 14426 4572 14653 4604
rect 14207 4570 14653 4572
rect 482 4549 565 4570
rect 482 4515 497 4549
rect 531 4536 565 4549
rect 531 4515 633 4536
rect 482 4498 633 4515
rect 14225 4536 14260 4570
rect 14294 4536 14329 4570
rect 14363 4536 14398 4570
rect 14432 4536 14467 4570
rect 14501 4536 14536 4570
rect 14570 4551 14653 4570
rect 14207 4534 14536 4536
rect 14207 4502 14246 4534
rect 14280 4502 14319 4534
rect 14353 4502 14392 4534
rect 14426 4502 14536 4534
rect 14226 4500 14246 4502
rect 14295 4500 14319 4502
rect 14364 4500 14392 4502
rect 482 4479 565 4498
rect 482 4445 497 4479
rect 531 4464 565 4479
rect 599 4468 633 4498
rect 12363 4468 12398 4500
rect 12432 4468 12467 4500
rect 12501 4468 12536 4500
rect 12570 4468 12605 4500
rect 12639 4468 12674 4500
rect 12708 4468 12743 4500
rect 12777 4468 12812 4500
rect 12846 4468 12881 4500
rect 12915 4468 12950 4500
rect 12984 4468 13019 4500
rect 13053 4468 13088 4500
rect 13122 4468 13157 4500
rect 13191 4468 13226 4500
rect 13260 4468 13295 4500
rect 13329 4468 13364 4500
rect 13398 4468 13433 4500
rect 13467 4468 13502 4500
rect 13536 4468 13571 4500
rect 13605 4468 13640 4500
rect 13674 4468 13709 4500
rect 13743 4468 13778 4500
rect 13812 4468 13847 4500
rect 13881 4468 13916 4500
rect 13950 4468 13985 4500
rect 14019 4468 14054 4500
rect 14088 4468 14123 4500
rect 14157 4468 14192 4500
rect 14226 4468 14261 4500
rect 14295 4468 14330 4500
rect 14364 4468 14399 4500
rect 14433 4468 14468 4502
rect 599 4464 14468 4468
rect 531 4456 14468 4464
rect 531 4445 674 4456
rect 708 4453 14428 4456
rect 708 4445 780 4453
rect 482 4429 674 4445
rect 482 4426 633 4429
rect 482 4409 529 4426
rect 482 4375 497 4409
rect 563 4392 565 4426
rect 599 4392 601 4426
rect 667 4395 674 4429
rect 635 4392 674 4395
rect 531 4375 674 4392
rect 482 4356 674 4375
rect 482 4354 633 4356
rect 482 4351 565 4354
rect 482 4339 529 4351
rect 482 4305 497 4339
rect 563 4320 565 4351
rect 599 4351 633 4354
rect 599 4320 601 4351
rect 667 4322 674 4356
rect 563 4317 601 4320
rect 635 4317 674 4322
rect 531 4305 674 4317
rect 482 4283 674 4305
rect 482 4282 633 4283
rect 482 4276 565 4282
rect 482 4269 529 4276
rect 482 4235 497 4269
rect 563 4248 565 4276
rect 599 4276 633 4282
rect 599 4248 601 4276
rect 667 4249 674 4283
rect 563 4242 601 4248
rect 635 4242 674 4249
rect 531 4235 674 4242
rect 482 4211 674 4235
rect 482 4210 633 4211
rect 482 4201 565 4210
rect 482 4199 529 4201
rect 482 4165 497 4199
rect 563 4176 565 4201
rect 599 4201 633 4210
rect 599 4176 601 4201
rect 667 4177 674 4211
rect 563 4167 601 4176
rect 635 4167 674 4177
rect 531 4165 674 4167
rect 482 4139 674 4165
rect 482 4138 633 4139
rect 482 4129 565 4138
rect 482 4095 497 4129
rect 531 4126 565 4129
rect 563 4104 565 4126
rect 599 4126 633 4138
rect 599 4104 601 4126
rect 667 4105 674 4139
rect 482 4092 529 4095
rect 563 4092 601 4104
rect 635 4092 674 4105
rect 482 4067 674 4092
rect 482 4066 633 4067
rect 482 4059 565 4066
rect 482 4025 497 4059
rect 531 4052 565 4059
rect 563 4032 565 4052
rect 599 4052 633 4066
rect 599 4032 601 4052
rect 667 4033 674 4067
rect 482 4018 529 4025
rect 563 4018 601 4032
rect 635 4018 674 4033
rect 482 3995 674 4018
rect 482 3994 633 3995
rect 482 3989 565 3994
rect 482 3955 497 3989
rect 531 3978 565 3989
rect 563 3960 565 3978
rect 599 3978 633 3994
rect 599 3960 601 3978
rect 667 3961 674 3995
rect 482 3944 529 3955
rect 563 3944 601 3960
rect 635 3944 674 3961
rect 482 3923 674 3944
rect 482 3922 633 3923
rect 482 3920 565 3922
rect 482 3886 497 3920
rect 531 3904 565 3920
rect 563 3888 565 3904
rect 599 3904 633 3922
rect 599 3888 601 3904
rect 667 3889 674 3923
rect 482 3870 529 3886
rect 563 3870 601 3888
rect 635 3870 674 3889
rect 482 3851 674 3870
rect 482 3817 497 3851
rect 531 3817 565 3851
rect 599 3817 633 3851
rect 667 3817 674 3851
rect 482 3794 674 3817
rect 482 3760 529 3794
rect 563 3760 601 3794
rect 635 3760 674 3794
rect 482 3749 674 3760
rect 482 3715 497 3749
rect 531 3720 565 3749
rect 563 3715 565 3720
rect 599 3720 633 3749
rect 599 3715 601 3720
rect 667 3715 674 3749
rect 482 3686 529 3715
rect 563 3686 601 3715
rect 635 3686 674 3715
rect 482 3680 674 3686
rect 482 3646 497 3680
rect 531 3646 565 3680
rect 599 3646 633 3680
rect 667 3646 674 3680
rect 482 3612 529 3646
rect 563 3612 601 3646
rect 635 3612 674 3646
rect 482 3611 674 3612
rect 482 3577 497 3611
rect 531 3577 565 3611
rect 599 3577 633 3611
rect 667 3577 674 3611
rect 482 3572 674 3577
rect 482 3542 529 3572
rect 563 3542 601 3572
rect 635 3542 674 3572
rect 482 3508 497 3542
rect 563 3538 565 3542
rect 531 3508 565 3538
rect 599 3538 601 3542
rect 599 3508 633 3538
rect 667 3508 674 3542
rect 482 3498 674 3508
rect 482 3473 529 3498
rect 563 3473 601 3498
rect 635 3473 674 3498
rect 482 3439 497 3473
rect 563 3464 565 3473
rect 531 3439 565 3464
rect 599 3464 601 3473
rect 599 3439 633 3464
rect 667 3439 674 3473
rect 482 3424 674 3439
rect 482 3404 529 3424
rect 563 3404 601 3424
rect 635 3404 674 3424
rect 482 3370 497 3404
rect 563 3390 565 3404
rect 531 3370 565 3390
rect 599 3390 601 3404
rect 599 3370 633 3390
rect 667 3370 674 3404
rect 482 3350 674 3370
rect 482 3335 529 3350
rect 563 3335 601 3350
rect 635 3335 674 3350
rect 482 3301 497 3335
rect 563 3316 565 3335
rect 531 3301 565 3316
rect 599 3316 601 3335
rect 599 3301 633 3316
rect 667 3301 674 3335
rect 482 3276 674 3301
rect 482 3266 529 3276
rect 563 3266 601 3276
rect 635 3266 674 3276
rect 482 3232 497 3266
rect 563 3242 565 3266
rect 531 3232 565 3242
rect 599 3242 601 3266
rect 599 3232 633 3242
rect 667 3232 674 3266
rect 482 3202 674 3232
rect 482 3197 529 3202
rect 563 3197 601 3202
rect 635 3197 674 3202
rect 482 3163 497 3197
rect 563 3168 565 3197
rect 531 3163 565 3168
rect 599 3168 601 3197
rect 599 3163 633 3168
rect 667 3163 674 3197
rect 482 3128 674 3163
rect 482 3094 497 3128
rect 563 3094 565 3128
rect 599 3094 601 3128
rect 667 3094 674 3128
rect 482 3059 674 3094
rect 482 3025 497 3059
rect 531 3054 565 3059
rect 563 3025 565 3054
rect 599 3054 633 3059
rect 599 3025 601 3054
rect 667 3025 674 3059
rect 482 3020 529 3025
rect 563 3020 601 3025
rect 635 3020 674 3025
rect 482 2990 674 3020
rect 482 2956 497 2990
rect 531 2980 565 2990
rect 563 2956 565 2980
rect 599 2980 633 2990
rect 599 2956 601 2980
rect 667 2956 674 2990
rect 482 2946 529 2956
rect 563 2946 601 2956
rect 635 2946 674 2956
rect 482 2921 674 2946
rect 482 2887 497 2921
rect 531 2906 565 2921
rect 563 2887 565 2906
rect 599 2906 633 2921
rect 599 2887 601 2906
rect 667 2887 674 2921
rect 482 2872 529 2887
rect 563 2872 601 2887
rect 635 2872 674 2887
rect 482 2852 674 2872
rect 482 2818 497 2852
rect 531 2832 565 2852
rect 563 2818 565 2832
rect 599 2832 633 2852
rect 599 2818 601 2832
rect 667 2818 674 2852
rect 482 2798 529 2818
rect 563 2798 601 2818
rect 635 2798 674 2818
rect 482 2783 674 2798
rect 482 2749 497 2783
rect 531 2758 565 2783
rect 563 2749 565 2758
rect 599 2758 633 2783
rect 599 2749 601 2758
rect 667 2749 674 2783
rect 482 2724 529 2749
rect 563 2724 601 2749
rect 635 2724 674 2749
rect 482 2714 674 2724
rect 482 2680 497 2714
rect 531 2684 565 2714
rect 563 2680 565 2684
rect 599 2684 633 2714
rect 599 2680 601 2684
rect 667 2680 674 2714
rect 482 2650 529 2680
rect 563 2650 601 2680
rect 635 2650 674 2680
rect 482 2645 674 2650
rect 482 2611 497 2645
rect 531 2611 565 2645
rect 599 2611 633 2645
rect 667 2611 674 2645
rect 482 2610 674 2611
rect 482 2576 529 2610
rect 563 2576 601 2610
rect 635 2576 674 2610
rect 482 2542 497 2576
rect 531 2542 565 2576
rect 599 2542 633 2576
rect 667 2542 674 2576
rect 482 2536 674 2542
rect 482 2507 529 2536
rect 563 2507 601 2536
rect 635 2507 674 2536
rect 482 2473 497 2507
rect 563 2502 565 2507
rect 531 2473 565 2502
rect 599 2502 601 2507
rect 599 2473 633 2502
rect 667 2473 674 2507
rect 482 2462 674 2473
rect 482 2438 529 2462
rect 563 2438 601 2462
rect 635 2438 674 2462
rect 482 2404 497 2438
rect 563 2428 565 2438
rect 531 2404 565 2428
rect 599 2428 601 2438
rect 599 2404 633 2428
rect 667 2404 674 2438
rect 482 2389 674 2404
rect 482 2369 529 2389
rect 563 2369 601 2389
rect 635 2369 674 2389
rect 482 2335 497 2369
rect 563 2355 565 2369
rect 531 2335 565 2355
rect 599 2355 601 2369
rect 599 2335 633 2355
rect 667 2335 674 2369
rect 482 2316 674 2335
rect 482 2300 529 2316
rect 563 2300 601 2316
rect 635 2300 674 2316
rect 482 2266 497 2300
rect 563 2282 565 2300
rect 531 2266 565 2282
rect 599 2282 601 2300
rect 599 2266 633 2282
rect 667 2266 674 2300
rect 482 2243 674 2266
rect 482 2231 529 2243
rect 563 2231 601 2243
rect 635 2231 674 2243
rect 482 2197 497 2231
rect 563 2209 565 2231
rect 531 2197 565 2209
rect 599 2209 601 2231
rect 599 2197 633 2209
rect 667 2197 674 2231
rect 482 2170 674 2197
rect 482 2163 529 2170
rect 482 2129 497 2163
rect 563 2162 601 2170
rect 635 2162 674 2170
rect 563 2136 565 2162
rect 531 2129 565 2136
rect 482 2128 565 2129
rect 599 2136 601 2162
rect 599 2128 633 2136
rect 667 2128 674 2162
rect 482 2097 674 2128
rect 482 2095 529 2097
rect 482 2061 497 2095
rect 563 2093 601 2097
rect 635 2093 674 2097
rect 563 2063 565 2093
rect 531 2061 565 2063
rect 482 2059 565 2061
rect 599 2063 601 2093
rect 599 2059 633 2063
rect 667 2059 674 2093
rect 482 2027 674 2059
rect 482 1993 497 2027
rect 531 2024 674 2027
rect 482 1990 529 1993
rect 563 1990 565 2024
rect 599 1990 601 2024
rect 667 1990 674 2024
rect 482 1959 674 1990
rect 482 1925 497 1959
rect 531 1955 674 1959
rect 531 1951 565 1955
rect 482 1917 529 1925
rect 563 1921 565 1951
rect 599 1951 633 1955
rect 599 1921 601 1951
rect 667 1921 674 1955
rect 563 1917 601 1921
rect 635 1917 674 1921
rect 482 1891 674 1917
rect 482 1857 497 1891
rect 531 1886 674 1891
rect 531 1878 565 1886
rect 482 1844 529 1857
rect 563 1852 565 1878
rect 599 1878 633 1886
rect 599 1852 601 1878
rect 667 1852 674 1886
rect 563 1844 601 1852
rect 635 1844 674 1852
rect 482 1823 674 1844
rect 482 1789 497 1823
rect 531 1817 674 1823
rect 531 1805 565 1817
rect 482 1771 529 1789
rect 563 1783 565 1805
rect 599 1805 633 1817
rect 599 1783 601 1805
rect 667 1783 674 1817
rect 563 1771 601 1783
rect 635 1771 674 1783
rect 482 1755 674 1771
rect 482 1721 497 1755
rect 531 1748 674 1755
rect 531 1732 565 1748
rect 482 1698 529 1721
rect 563 1714 565 1732
rect 599 1732 633 1748
rect 599 1714 601 1732
rect 667 1714 674 1748
rect 563 1698 601 1714
rect 635 1698 674 1714
rect 482 1687 674 1698
rect 482 1653 497 1687
rect 531 1679 674 1687
rect 531 1659 565 1679
rect 482 1625 529 1653
rect 563 1645 565 1659
rect 599 1659 633 1679
rect 599 1645 601 1659
rect 667 1645 674 1679
rect 563 1625 601 1645
rect 635 1625 674 1645
rect 482 1619 674 1625
rect 482 1585 497 1619
rect 531 1610 674 1619
rect 531 1586 565 1610
rect 482 1552 529 1585
rect 563 1576 565 1586
rect 599 1586 633 1610
rect 599 1576 601 1586
rect 667 1576 674 1610
rect 563 1552 601 1576
rect 635 1552 674 1576
rect 482 1551 674 1552
rect 482 1517 497 1551
rect 531 1541 674 1551
rect 531 1517 565 1541
rect 482 1513 565 1517
rect 482 1483 529 1513
rect 563 1507 565 1513
rect 599 1513 633 1541
rect 599 1507 601 1513
rect 667 1507 674 1541
rect 482 1449 497 1483
rect 563 1479 601 1507
rect 635 1479 674 1507
rect 531 1472 674 1479
rect 531 1449 565 1472
rect 482 1440 565 1449
rect 482 1415 529 1440
rect 563 1438 565 1440
rect 599 1440 633 1472
rect 599 1438 601 1440
rect 667 1438 674 1472
rect 482 1381 497 1415
rect 563 1406 601 1438
rect 635 1406 674 1438
rect 531 1403 674 1406
rect 531 1381 565 1403
rect 482 1369 565 1381
rect 599 1369 633 1403
rect 667 1369 674 1403
rect 482 1367 674 1369
rect 482 1347 529 1367
rect 482 1313 497 1347
rect 563 1334 601 1367
rect 635 1334 674 1367
rect 563 1333 565 1334
rect 531 1313 565 1333
rect 482 1300 565 1313
rect 599 1333 601 1334
rect 599 1300 633 1333
rect 667 1300 674 1334
rect 482 1294 674 1300
rect 482 1279 529 1294
rect 482 1245 497 1279
rect 563 1265 601 1294
rect 635 1265 674 1294
rect 563 1260 565 1265
rect 531 1245 565 1260
rect 482 1231 565 1245
rect 599 1260 601 1265
rect 599 1231 633 1260
rect 667 1231 674 1265
rect 482 1221 674 1231
rect 482 1211 529 1221
rect 482 1177 497 1211
rect 563 1196 601 1221
rect 635 1196 674 1221
rect 563 1187 565 1196
rect 531 1177 565 1187
rect 482 1162 565 1177
rect 599 1187 601 1196
rect 599 1162 633 1187
rect 667 1162 674 1196
rect 482 1148 674 1162
rect 482 1143 529 1148
rect 482 1109 497 1143
rect 563 1127 601 1148
rect 635 1127 674 1148
rect 563 1114 565 1127
rect 531 1109 565 1114
rect 482 1093 565 1109
rect 599 1114 601 1127
rect 599 1093 633 1114
rect 667 1093 674 1127
rect 482 1075 674 1093
rect 482 1041 497 1075
rect 563 1058 601 1075
rect 635 1058 674 1075
rect 563 1041 565 1058
rect 482 1024 565 1041
rect 599 1041 601 1058
rect 599 1024 633 1041
rect 667 1024 674 1058
rect 482 1007 674 1024
rect 482 973 497 1007
rect 531 1002 674 1007
rect 563 989 601 1002
rect 635 989 674 1002
rect 482 968 529 973
rect 563 968 565 989
rect 482 955 565 968
rect 599 968 601 989
rect 599 955 633 968
rect 667 955 674 989
rect 482 939 674 955
rect 482 769 497 939
rect 531 929 674 939
rect 563 920 601 929
rect 635 920 674 929
rect 667 894 674 920
rect 14356 4432 14428 4453
rect 14390 4398 14428 4432
rect 14462 4426 14468 4456
rect 14356 4359 14428 4398
rect 14390 4325 14428 4359
rect 881 4308 1001 4324
rect 881 4274 924 4308
rect 958 4274 1001 4308
rect 881 4234 1001 4274
rect 881 4200 924 4234
rect 958 4200 1001 4234
rect 881 3104 1001 4200
rect 1311 4308 1431 4324
rect 1311 4274 1354 4308
rect 1388 4274 1431 4308
rect 1311 4234 1431 4274
rect 1311 4200 1354 4234
rect 1388 4200 1431 4234
rect 881 3070 924 3104
rect 958 3070 1001 3104
rect 881 3026 1001 3070
rect 881 2992 924 3026
rect 958 2992 1001 3026
rect 881 2948 1001 2992
rect 881 2914 924 2948
rect 958 2914 1001 2948
rect 881 2870 1001 2914
rect 881 2836 924 2870
rect 958 2836 1001 2870
rect 881 2792 1001 2836
rect 881 2758 924 2792
rect 958 2758 1001 2792
rect 881 2713 1001 2758
rect 881 2679 924 2713
rect 958 2679 1001 2713
rect 881 2634 1001 2679
rect 881 2600 924 2634
rect 958 2600 1001 2634
rect 881 1504 1001 2600
rect 1066 4064 1067 4098
rect 1101 4064 1139 4098
rect 1173 4064 1211 4098
rect 1245 4064 1246 4098
rect 1066 4025 1246 4064
rect 1066 3991 1067 4025
rect 1101 3991 1139 4025
rect 1173 3991 1211 4025
rect 1245 3991 1246 4025
rect 1066 3952 1246 3991
rect 1066 3918 1067 3952
rect 1101 3918 1139 3952
rect 1173 3918 1211 3952
rect 1245 3918 1246 3952
rect 1066 3879 1246 3918
rect 1066 3845 1067 3879
rect 1101 3845 1139 3879
rect 1173 3845 1211 3879
rect 1245 3845 1246 3879
rect 1066 3806 1246 3845
rect 1066 3772 1067 3806
rect 1101 3772 1139 3806
rect 1173 3772 1211 3806
rect 1245 3772 1246 3806
rect 1066 3733 1246 3772
rect 1066 3699 1067 3733
rect 1101 3699 1139 3733
rect 1173 3699 1211 3733
rect 1245 3699 1246 3733
rect 1066 3660 1246 3699
rect 1066 3626 1067 3660
rect 1101 3626 1139 3660
rect 1173 3626 1211 3660
rect 1245 3626 1246 3660
rect 1066 3587 1246 3626
rect 1066 3553 1067 3587
rect 1101 3553 1139 3587
rect 1173 3553 1211 3587
rect 1245 3553 1246 3587
rect 1066 3514 1246 3553
rect 1066 3480 1067 3514
rect 1101 3480 1139 3514
rect 1173 3480 1211 3514
rect 1245 3480 1246 3514
rect 1066 3441 1246 3480
rect 1066 3407 1067 3441
rect 1101 3407 1139 3441
rect 1173 3407 1211 3441
rect 1245 3407 1246 3441
rect 1066 3368 1246 3407
rect 1066 3334 1067 3368
rect 1101 3334 1139 3368
rect 1173 3334 1211 3368
rect 1245 3334 1246 3368
rect 1066 3295 1246 3334
rect 1066 3261 1067 3295
rect 1101 3261 1139 3295
rect 1173 3261 1211 3295
rect 1245 3261 1246 3295
rect 1066 3222 1246 3261
rect 1066 3188 1067 3222
rect 1101 3188 1139 3222
rect 1173 3188 1211 3222
rect 1245 3188 1246 3222
rect 1066 3149 1246 3188
rect 1066 3115 1067 3149
rect 1101 3115 1139 3149
rect 1173 3115 1211 3149
rect 1245 3115 1246 3149
rect 1066 3076 1246 3115
rect 1066 3042 1067 3076
rect 1101 3042 1139 3076
rect 1173 3042 1211 3076
rect 1245 3042 1246 3076
rect 1066 3003 1246 3042
rect 1066 2969 1067 3003
rect 1101 2969 1139 3003
rect 1173 2969 1211 3003
rect 1245 2969 1246 3003
rect 1066 2930 1246 2969
rect 1066 2896 1067 2930
rect 1101 2896 1139 2930
rect 1173 2896 1211 2930
rect 1245 2896 1246 2930
rect 1066 2857 1246 2896
rect 1066 2823 1067 2857
rect 1101 2823 1139 2857
rect 1173 2823 1211 2857
rect 1245 2823 1246 2857
rect 1066 2784 1246 2823
rect 1066 2750 1067 2784
rect 1101 2750 1139 2784
rect 1173 2750 1211 2784
rect 1245 2750 1246 2784
rect 1066 2711 1246 2750
rect 1066 2677 1067 2711
rect 1101 2677 1139 2711
rect 1173 2677 1211 2711
rect 1245 2677 1246 2711
rect 1066 2638 1246 2677
rect 1066 2604 1067 2638
rect 1101 2604 1139 2638
rect 1173 2604 1211 2638
rect 1245 2604 1246 2638
rect 1066 2565 1246 2604
rect 1066 2531 1067 2565
rect 1101 2531 1139 2565
rect 1173 2531 1211 2565
rect 1245 2531 1246 2565
rect 1066 2492 1246 2531
rect 1066 2458 1067 2492
rect 1101 2458 1139 2492
rect 1173 2458 1211 2492
rect 1245 2458 1246 2492
rect 1066 2419 1246 2458
rect 1066 2385 1067 2419
rect 1101 2385 1139 2419
rect 1173 2385 1211 2419
rect 1245 2385 1246 2419
rect 1066 2346 1246 2385
rect 1066 2312 1067 2346
rect 1101 2312 1139 2346
rect 1173 2312 1211 2346
rect 1245 2312 1246 2346
rect 1066 2273 1246 2312
rect 1066 2239 1067 2273
rect 1101 2239 1139 2273
rect 1173 2239 1211 2273
rect 1245 2239 1246 2273
rect 1066 2200 1246 2239
rect 1066 2166 1067 2200
rect 1101 2166 1139 2200
rect 1173 2166 1211 2200
rect 1245 2166 1246 2200
rect 1066 2126 1246 2166
rect 1066 2092 1067 2126
rect 1101 2092 1139 2126
rect 1173 2092 1211 2126
rect 1245 2092 1246 2126
rect 1066 2052 1246 2092
rect 1066 2018 1067 2052
rect 1101 2018 1139 2052
rect 1173 2018 1211 2052
rect 1245 2018 1246 2052
rect 1066 1978 1246 2018
rect 1066 1944 1067 1978
rect 1101 1944 1139 1978
rect 1173 1944 1211 1978
rect 1245 1944 1246 1978
rect 1066 1904 1246 1944
rect 1066 1870 1067 1904
rect 1101 1870 1139 1904
rect 1173 1870 1211 1904
rect 1245 1870 1246 1904
rect 1066 1830 1246 1870
rect 1066 1796 1067 1830
rect 1101 1796 1139 1830
rect 1173 1796 1211 1830
rect 1245 1796 1246 1830
rect 1066 1756 1246 1796
rect 1066 1722 1067 1756
rect 1101 1722 1139 1756
rect 1173 1722 1211 1756
rect 1245 1722 1246 1756
rect 1066 1682 1246 1722
rect 1066 1648 1067 1682
rect 1101 1648 1139 1682
rect 1173 1648 1211 1682
rect 1245 1648 1246 1682
rect 1066 1608 1246 1648
rect 1066 1574 1067 1608
rect 1101 1574 1139 1608
rect 1173 1574 1211 1608
rect 1245 1574 1246 1608
rect 1066 1548 1246 1574
rect 1311 3104 1431 4200
rect 1873 4308 1993 4324
rect 1873 4274 1916 4308
rect 1950 4274 1993 4308
rect 1873 4234 1993 4274
rect 1873 4200 1916 4234
rect 1950 4200 1993 4234
rect 1311 3070 1354 3104
rect 1388 3070 1431 3104
rect 1311 3026 1431 3070
rect 1311 2992 1354 3026
rect 1388 2992 1431 3026
rect 1311 2948 1431 2992
rect 1311 2914 1354 2948
rect 1388 2914 1431 2948
rect 1311 2870 1431 2914
rect 1311 2836 1354 2870
rect 1388 2836 1431 2870
rect 1311 2792 1431 2836
rect 1311 2758 1354 2792
rect 1388 2758 1431 2792
rect 1311 2713 1431 2758
rect 1311 2679 1354 2713
rect 1388 2679 1431 2713
rect 1311 2634 1431 2679
rect 1311 2600 1354 2634
rect 1388 2600 1431 2634
rect 881 1470 924 1504
rect 958 1470 1001 1504
rect 881 1430 1001 1470
rect 881 1396 924 1430
rect 958 1396 1001 1430
rect 881 1250 1001 1396
rect 881 1216 924 1250
rect 958 1216 1001 1250
rect 881 1178 1001 1216
rect 881 1144 924 1178
rect 958 1144 1001 1178
rect 1311 1504 1431 2600
rect 1533 4092 1771 4104
rect 1533 4058 1563 4092
rect 1597 4058 1707 4092
rect 1741 4058 1771 4092
rect 1533 4020 1771 4058
rect 1533 3986 1563 4020
rect 1597 3986 1707 4020
rect 1741 3986 1771 4020
rect 1533 3948 1771 3986
rect 1533 3914 1563 3948
rect 1597 3914 1707 3948
rect 1741 3914 1771 3948
rect 1533 3876 1771 3914
rect 1533 3842 1563 3876
rect 1597 3842 1707 3876
rect 1741 3842 1771 3876
rect 1533 3804 1771 3842
rect 1533 3770 1563 3804
rect 1597 3770 1707 3804
rect 1741 3770 1771 3804
rect 1533 3732 1771 3770
rect 1533 3698 1563 3732
rect 1597 3698 1707 3732
rect 1741 3698 1771 3732
rect 1533 3660 1771 3698
rect 1533 3626 1563 3660
rect 1597 3626 1707 3660
rect 1741 3626 1771 3660
rect 1533 3588 1771 3626
rect 1533 3554 1563 3588
rect 1597 3554 1707 3588
rect 1741 3554 1771 3588
rect 1533 3516 1771 3554
rect 1533 3482 1563 3516
rect 1597 3482 1707 3516
rect 1741 3482 1771 3516
rect 1533 3444 1771 3482
rect 1533 3410 1563 3444
rect 1597 3410 1707 3444
rect 1741 3410 1771 3444
rect 1533 3372 1771 3410
rect 1533 3338 1563 3372
rect 1597 3338 1707 3372
rect 1741 3338 1771 3372
rect 1533 3300 1771 3338
rect 1533 3266 1563 3300
rect 1597 3266 1707 3300
rect 1741 3266 1771 3300
rect 1533 3228 1771 3266
rect 1533 3194 1563 3228
rect 1597 3194 1707 3228
rect 1741 3194 1771 3228
rect 1533 3108 1771 3194
rect 1533 3074 1563 3108
rect 1597 3074 1635 3108
rect 1669 3074 1707 3108
rect 1741 3074 1771 3108
rect 1533 3044 1771 3074
rect 1533 3028 1601 3044
rect 1533 2994 1563 3028
rect 1597 3010 1601 3028
rect 1635 3028 1669 3044
rect 1597 2994 1635 3010
rect 1703 3028 1771 3044
rect 1703 3010 1707 3028
rect 1669 2994 1707 3010
rect 1741 2994 1771 3028
rect 1533 2974 1771 2994
rect 1533 2948 1601 2974
rect 1533 2914 1563 2948
rect 1597 2940 1601 2948
rect 1635 2948 1669 2974
rect 1597 2914 1635 2940
rect 1703 2948 1771 2974
rect 1703 2940 1707 2948
rect 1669 2914 1707 2940
rect 1741 2914 1771 2948
rect 1533 2904 1771 2914
rect 1533 2870 1601 2904
rect 1635 2870 1669 2904
rect 1703 2870 1771 2904
rect 1533 2868 1771 2870
rect 1533 2834 1563 2868
rect 1597 2834 1635 2868
rect 1669 2834 1707 2868
rect 1741 2834 1771 2868
rect 1533 2800 1601 2834
rect 1635 2800 1669 2834
rect 1703 2800 1771 2834
rect 1533 2788 1771 2800
rect 1533 2754 1563 2788
rect 1597 2764 1635 2788
rect 1597 2754 1601 2764
rect 1533 2730 1601 2754
rect 1669 2764 1707 2788
rect 1635 2730 1669 2754
rect 1703 2754 1707 2764
rect 1741 2754 1771 2788
rect 1703 2730 1771 2754
rect 1533 2708 1771 2730
rect 1533 2674 1563 2708
rect 1597 2694 1635 2708
rect 1597 2674 1601 2694
rect 1533 2660 1601 2674
rect 1669 2694 1707 2708
rect 1635 2660 1669 2674
rect 1703 2674 1707 2694
rect 1741 2674 1771 2708
rect 1703 2660 1771 2674
rect 1533 2628 1771 2660
rect 1533 2594 1563 2628
rect 1597 2594 1635 2628
rect 1669 2594 1707 2628
rect 1741 2594 1771 2628
rect 1533 2518 1771 2594
rect 1533 2484 1563 2518
rect 1597 2484 1707 2518
rect 1741 2484 1771 2518
rect 1533 2446 1771 2484
rect 1533 2412 1563 2446
rect 1597 2412 1707 2446
rect 1741 2412 1771 2446
rect 1533 2374 1771 2412
rect 1533 2340 1563 2374
rect 1597 2340 1707 2374
rect 1741 2340 1771 2374
rect 1533 2302 1771 2340
rect 1533 2268 1563 2302
rect 1597 2268 1707 2302
rect 1741 2268 1771 2302
rect 1533 2230 1771 2268
rect 1533 2196 1563 2230
rect 1597 2196 1707 2230
rect 1741 2196 1771 2230
rect 1533 2158 1771 2196
rect 1533 2124 1563 2158
rect 1597 2124 1707 2158
rect 1741 2124 1771 2158
rect 1533 2086 1771 2124
rect 1533 2052 1563 2086
rect 1597 2052 1707 2086
rect 1741 2052 1771 2086
rect 1533 2014 1771 2052
rect 1533 1980 1563 2014
rect 1597 1980 1707 2014
rect 1741 1980 1771 2014
rect 1533 1942 1771 1980
rect 1533 1908 1563 1942
rect 1597 1908 1707 1942
rect 1741 1908 1771 1942
rect 1533 1870 1771 1908
rect 1533 1836 1563 1870
rect 1597 1836 1707 1870
rect 1741 1836 1771 1870
rect 1533 1798 1771 1836
rect 1533 1764 1563 1798
rect 1597 1764 1707 1798
rect 1741 1764 1771 1798
rect 1533 1726 1771 1764
rect 1533 1692 1563 1726
rect 1597 1692 1707 1726
rect 1741 1692 1771 1726
rect 1533 1654 1771 1692
rect 1533 1620 1563 1654
rect 1597 1620 1707 1654
rect 1741 1620 1771 1654
rect 1533 1536 1771 1620
rect 1873 3104 1993 4200
rect 2303 4308 2423 4324
rect 2303 4274 2346 4308
rect 2380 4274 2423 4308
rect 2303 4234 2423 4274
rect 2303 4200 2346 4234
rect 2380 4200 2423 4234
rect 1873 3070 1916 3104
rect 1950 3070 1993 3104
rect 1873 3026 1993 3070
rect 1873 2992 1916 3026
rect 1950 2992 1993 3026
rect 1873 2948 1993 2992
rect 1873 2914 1916 2948
rect 1950 2914 1993 2948
rect 1873 2870 1993 2914
rect 1873 2836 1916 2870
rect 1950 2836 1993 2870
rect 1873 2792 1993 2836
rect 1873 2758 1916 2792
rect 1950 2758 1993 2792
rect 1873 2713 1993 2758
rect 1873 2679 1916 2713
rect 1950 2679 1993 2713
rect 1873 2634 1993 2679
rect 1873 2600 1916 2634
rect 1950 2600 1993 2634
rect 1311 1470 1354 1504
rect 1388 1470 1431 1504
rect 1311 1430 1431 1470
rect 1311 1396 1354 1430
rect 1388 1396 1431 1430
rect 1311 1250 1431 1396
rect 1311 1144 1318 1250
rect 1424 1144 1431 1250
rect 1873 1504 1993 2600
rect 2058 4064 2059 4098
rect 2093 4064 2131 4098
rect 2165 4064 2203 4098
rect 2237 4064 2238 4098
rect 2058 4025 2238 4064
rect 2058 3991 2059 4025
rect 2093 3991 2131 4025
rect 2165 3991 2203 4025
rect 2237 3991 2238 4025
rect 2058 3952 2238 3991
rect 2058 3918 2059 3952
rect 2093 3918 2131 3952
rect 2165 3918 2203 3952
rect 2237 3918 2238 3952
rect 2058 3879 2238 3918
rect 2058 3845 2059 3879
rect 2093 3845 2131 3879
rect 2165 3845 2203 3879
rect 2237 3845 2238 3879
rect 2058 3806 2238 3845
rect 2058 3772 2059 3806
rect 2093 3772 2131 3806
rect 2165 3772 2203 3806
rect 2237 3772 2238 3806
rect 2058 3733 2238 3772
rect 2058 3699 2059 3733
rect 2093 3699 2131 3733
rect 2165 3699 2203 3733
rect 2237 3699 2238 3733
rect 2058 3660 2238 3699
rect 2058 3626 2059 3660
rect 2093 3626 2131 3660
rect 2165 3626 2203 3660
rect 2237 3626 2238 3660
rect 2058 3587 2238 3626
rect 2058 3553 2059 3587
rect 2093 3553 2131 3587
rect 2165 3553 2203 3587
rect 2237 3553 2238 3587
rect 2058 3514 2238 3553
rect 2058 3480 2059 3514
rect 2093 3480 2131 3514
rect 2165 3480 2203 3514
rect 2237 3480 2238 3514
rect 2058 3441 2238 3480
rect 2058 3407 2059 3441
rect 2093 3407 2131 3441
rect 2165 3407 2203 3441
rect 2237 3407 2238 3441
rect 2058 3368 2238 3407
rect 2058 3334 2059 3368
rect 2093 3334 2131 3368
rect 2165 3334 2203 3368
rect 2237 3334 2238 3368
rect 2058 3295 2238 3334
rect 2058 3261 2059 3295
rect 2093 3261 2131 3295
rect 2165 3261 2203 3295
rect 2237 3261 2238 3295
rect 2058 3222 2238 3261
rect 2058 3188 2059 3222
rect 2093 3188 2131 3222
rect 2165 3188 2203 3222
rect 2237 3188 2238 3222
rect 2058 3149 2238 3188
rect 2058 3115 2059 3149
rect 2093 3115 2131 3149
rect 2165 3115 2203 3149
rect 2237 3115 2238 3149
rect 2058 3076 2238 3115
rect 2058 3042 2059 3076
rect 2093 3042 2131 3076
rect 2165 3042 2203 3076
rect 2237 3042 2238 3076
rect 2058 3003 2238 3042
rect 2058 2969 2059 3003
rect 2093 2969 2131 3003
rect 2165 2969 2203 3003
rect 2237 2969 2238 3003
rect 2058 2930 2238 2969
rect 2058 2896 2059 2930
rect 2093 2896 2131 2930
rect 2165 2896 2203 2930
rect 2237 2896 2238 2930
rect 2058 2857 2238 2896
rect 2058 2823 2059 2857
rect 2093 2823 2131 2857
rect 2165 2823 2203 2857
rect 2237 2823 2238 2857
rect 2058 2784 2238 2823
rect 2058 2750 2059 2784
rect 2093 2750 2131 2784
rect 2165 2750 2203 2784
rect 2237 2750 2238 2784
rect 2058 2711 2238 2750
rect 2058 2677 2059 2711
rect 2093 2677 2131 2711
rect 2165 2677 2203 2711
rect 2237 2677 2238 2711
rect 2058 2638 2238 2677
rect 2058 2604 2059 2638
rect 2093 2604 2131 2638
rect 2165 2604 2203 2638
rect 2237 2604 2238 2638
rect 2058 2565 2238 2604
rect 2058 2531 2059 2565
rect 2093 2531 2131 2565
rect 2165 2531 2203 2565
rect 2237 2531 2238 2565
rect 2058 2492 2238 2531
rect 2058 2458 2059 2492
rect 2093 2458 2131 2492
rect 2165 2458 2203 2492
rect 2237 2458 2238 2492
rect 2058 2419 2238 2458
rect 2058 2385 2059 2419
rect 2093 2385 2131 2419
rect 2165 2385 2203 2419
rect 2237 2385 2238 2419
rect 2058 2346 2238 2385
rect 2058 2312 2059 2346
rect 2093 2312 2131 2346
rect 2165 2312 2203 2346
rect 2237 2312 2238 2346
rect 2058 2273 2238 2312
rect 2058 2239 2059 2273
rect 2093 2239 2131 2273
rect 2165 2239 2203 2273
rect 2237 2239 2238 2273
rect 2058 2200 2238 2239
rect 2058 2166 2059 2200
rect 2093 2166 2131 2200
rect 2165 2166 2203 2200
rect 2237 2166 2238 2200
rect 2058 2126 2238 2166
rect 2058 2092 2059 2126
rect 2093 2092 2131 2126
rect 2165 2092 2203 2126
rect 2237 2092 2238 2126
rect 2058 2052 2238 2092
rect 2058 2018 2059 2052
rect 2093 2018 2131 2052
rect 2165 2018 2203 2052
rect 2237 2018 2238 2052
rect 2058 1978 2238 2018
rect 2058 1944 2059 1978
rect 2093 1944 2131 1978
rect 2165 1944 2203 1978
rect 2237 1944 2238 1978
rect 2058 1904 2238 1944
rect 2058 1870 2059 1904
rect 2093 1870 2131 1904
rect 2165 1870 2203 1904
rect 2237 1870 2238 1904
rect 2058 1830 2238 1870
rect 2058 1796 2059 1830
rect 2093 1796 2131 1830
rect 2165 1796 2203 1830
rect 2237 1796 2238 1830
rect 2058 1756 2238 1796
rect 2058 1722 2059 1756
rect 2093 1722 2131 1756
rect 2165 1722 2203 1756
rect 2237 1722 2238 1756
rect 2058 1682 2238 1722
rect 2058 1648 2059 1682
rect 2093 1648 2131 1682
rect 2165 1648 2203 1682
rect 2237 1648 2238 1682
rect 2058 1608 2238 1648
rect 2058 1574 2059 1608
rect 2093 1574 2131 1608
rect 2165 1574 2203 1608
rect 2237 1574 2238 1608
rect 2058 1548 2238 1574
rect 2303 3104 2423 4200
rect 2865 4308 2985 4324
rect 2865 4274 2908 4308
rect 2942 4274 2985 4308
rect 2865 4234 2985 4274
rect 2865 4200 2908 4234
rect 2942 4200 2985 4234
rect 2303 3070 2346 3104
rect 2380 3070 2423 3104
rect 2303 3026 2423 3070
rect 2303 2992 2346 3026
rect 2380 2992 2423 3026
rect 2303 2948 2423 2992
rect 2303 2914 2346 2948
rect 2380 2914 2423 2948
rect 2303 2870 2423 2914
rect 2303 2836 2346 2870
rect 2380 2836 2423 2870
rect 2303 2792 2423 2836
rect 2303 2758 2346 2792
rect 2380 2758 2423 2792
rect 2303 2713 2423 2758
rect 2303 2679 2346 2713
rect 2380 2679 2423 2713
rect 2303 2634 2423 2679
rect 2303 2600 2346 2634
rect 2380 2600 2423 2634
rect 1873 1470 1916 1504
rect 1950 1470 1993 1504
rect 1873 1430 1993 1470
rect 1873 1396 1916 1430
rect 1950 1396 1993 1430
rect 1873 1250 1993 1396
rect 1873 1144 1880 1250
rect 1986 1144 1993 1250
rect 2303 1504 2423 2600
rect 2525 4092 2763 4104
rect 2525 4058 2555 4092
rect 2589 4058 2699 4092
rect 2733 4058 2763 4092
rect 2525 4020 2763 4058
rect 2525 3986 2555 4020
rect 2589 3986 2699 4020
rect 2733 3986 2763 4020
rect 2525 3948 2763 3986
rect 2525 3914 2555 3948
rect 2589 3914 2699 3948
rect 2733 3914 2763 3948
rect 2525 3876 2763 3914
rect 2525 3842 2555 3876
rect 2589 3842 2699 3876
rect 2733 3842 2763 3876
rect 2525 3804 2763 3842
rect 2525 3770 2555 3804
rect 2589 3770 2699 3804
rect 2733 3770 2763 3804
rect 2525 3732 2763 3770
rect 2525 3698 2555 3732
rect 2589 3698 2699 3732
rect 2733 3698 2763 3732
rect 2525 3660 2763 3698
rect 2525 3626 2555 3660
rect 2589 3626 2699 3660
rect 2733 3626 2763 3660
rect 2525 3588 2763 3626
rect 2525 3554 2555 3588
rect 2589 3554 2699 3588
rect 2733 3554 2763 3588
rect 2525 3516 2763 3554
rect 2525 3482 2555 3516
rect 2589 3482 2699 3516
rect 2733 3482 2763 3516
rect 2525 3444 2763 3482
rect 2525 3410 2555 3444
rect 2589 3410 2699 3444
rect 2733 3410 2763 3444
rect 2525 3372 2763 3410
rect 2525 3338 2555 3372
rect 2589 3338 2699 3372
rect 2733 3338 2763 3372
rect 2525 3300 2763 3338
rect 2525 3266 2555 3300
rect 2589 3266 2699 3300
rect 2733 3266 2763 3300
rect 2525 3228 2763 3266
rect 2525 3194 2555 3228
rect 2589 3194 2699 3228
rect 2733 3194 2763 3228
rect 2525 3108 2763 3194
rect 2525 3074 2555 3108
rect 2589 3074 2627 3108
rect 2661 3074 2699 3108
rect 2733 3074 2763 3108
rect 2525 3044 2763 3074
rect 2525 3028 2593 3044
rect 2525 2994 2555 3028
rect 2589 3010 2593 3028
rect 2627 3028 2661 3044
rect 2589 2994 2627 3010
rect 2695 3028 2763 3044
rect 2695 3010 2699 3028
rect 2661 2994 2699 3010
rect 2733 2994 2763 3028
rect 2525 2974 2763 2994
rect 2525 2948 2593 2974
rect 2525 2914 2555 2948
rect 2589 2940 2593 2948
rect 2627 2948 2661 2974
rect 2589 2914 2627 2940
rect 2695 2948 2763 2974
rect 2695 2940 2699 2948
rect 2661 2914 2699 2940
rect 2733 2914 2763 2948
rect 2525 2904 2763 2914
rect 2525 2870 2593 2904
rect 2627 2870 2661 2904
rect 2695 2870 2763 2904
rect 2525 2868 2763 2870
rect 2525 2834 2555 2868
rect 2589 2834 2627 2868
rect 2661 2834 2699 2868
rect 2733 2834 2763 2868
rect 2525 2800 2593 2834
rect 2627 2800 2661 2834
rect 2695 2800 2763 2834
rect 2525 2788 2763 2800
rect 2525 2754 2555 2788
rect 2589 2764 2627 2788
rect 2589 2754 2593 2764
rect 2525 2730 2593 2754
rect 2661 2764 2699 2788
rect 2627 2730 2661 2754
rect 2695 2754 2699 2764
rect 2733 2754 2763 2788
rect 2695 2730 2763 2754
rect 2525 2708 2763 2730
rect 2525 2674 2555 2708
rect 2589 2694 2627 2708
rect 2589 2674 2593 2694
rect 2525 2660 2593 2674
rect 2661 2694 2699 2708
rect 2627 2660 2661 2674
rect 2695 2674 2699 2694
rect 2733 2674 2763 2708
rect 2695 2660 2763 2674
rect 2525 2628 2763 2660
rect 2525 2594 2555 2628
rect 2589 2594 2627 2628
rect 2661 2594 2699 2628
rect 2733 2594 2763 2628
rect 2525 2518 2763 2594
rect 2525 2484 2555 2518
rect 2589 2484 2699 2518
rect 2733 2484 2763 2518
rect 2525 2446 2763 2484
rect 2525 2412 2555 2446
rect 2589 2412 2699 2446
rect 2733 2412 2763 2446
rect 2525 2374 2763 2412
rect 2525 2340 2555 2374
rect 2589 2340 2699 2374
rect 2733 2340 2763 2374
rect 2525 2302 2763 2340
rect 2525 2268 2555 2302
rect 2589 2268 2699 2302
rect 2733 2268 2763 2302
rect 2525 2230 2763 2268
rect 2525 2196 2555 2230
rect 2589 2196 2699 2230
rect 2733 2196 2763 2230
rect 2525 2158 2763 2196
rect 2525 2124 2555 2158
rect 2589 2124 2699 2158
rect 2733 2124 2763 2158
rect 2525 2086 2763 2124
rect 2525 2052 2555 2086
rect 2589 2052 2699 2086
rect 2733 2052 2763 2086
rect 2525 2014 2763 2052
rect 2525 1980 2555 2014
rect 2589 1980 2699 2014
rect 2733 1980 2763 2014
rect 2525 1942 2763 1980
rect 2525 1908 2555 1942
rect 2589 1908 2699 1942
rect 2733 1908 2763 1942
rect 2525 1870 2763 1908
rect 2525 1836 2555 1870
rect 2589 1836 2699 1870
rect 2733 1836 2763 1870
rect 2525 1798 2763 1836
rect 2525 1764 2555 1798
rect 2589 1764 2699 1798
rect 2733 1764 2763 1798
rect 2525 1726 2763 1764
rect 2525 1692 2555 1726
rect 2589 1692 2699 1726
rect 2733 1692 2763 1726
rect 2525 1654 2763 1692
rect 2525 1620 2555 1654
rect 2589 1620 2699 1654
rect 2733 1620 2763 1654
rect 2525 1536 2763 1620
rect 2865 3104 2985 4200
rect 3295 4308 3415 4324
rect 3295 4274 3338 4308
rect 3372 4274 3415 4308
rect 3295 4234 3415 4274
rect 3295 4200 3338 4234
rect 3372 4200 3415 4234
rect 2865 3070 2908 3104
rect 2942 3070 2985 3104
rect 2865 3026 2985 3070
rect 2865 2992 2908 3026
rect 2942 2992 2985 3026
rect 2865 2948 2985 2992
rect 2865 2914 2908 2948
rect 2942 2914 2985 2948
rect 2865 2870 2985 2914
rect 2865 2836 2908 2870
rect 2942 2836 2985 2870
rect 2865 2792 2985 2836
rect 2865 2758 2908 2792
rect 2942 2758 2985 2792
rect 2865 2713 2985 2758
rect 2865 2679 2908 2713
rect 2942 2679 2985 2713
rect 2865 2634 2985 2679
rect 2865 2600 2908 2634
rect 2942 2600 2985 2634
rect 2303 1470 2346 1504
rect 2380 1470 2423 1504
rect 2303 1430 2423 1470
rect 2303 1396 2346 1430
rect 2380 1396 2423 1430
rect 2303 1250 2423 1396
rect 2303 1144 2310 1250
rect 2416 1144 2423 1250
rect 2865 1504 2985 2600
rect 3050 4064 3051 4098
rect 3085 4064 3123 4098
rect 3157 4064 3195 4098
rect 3229 4064 3230 4098
rect 3050 4025 3230 4064
rect 3050 3991 3051 4025
rect 3085 3991 3123 4025
rect 3157 3991 3195 4025
rect 3229 3991 3230 4025
rect 3050 3952 3230 3991
rect 3050 3918 3051 3952
rect 3085 3918 3123 3952
rect 3157 3918 3195 3952
rect 3229 3918 3230 3952
rect 3050 3879 3230 3918
rect 3050 3845 3051 3879
rect 3085 3845 3123 3879
rect 3157 3845 3195 3879
rect 3229 3845 3230 3879
rect 3050 3806 3230 3845
rect 3050 3772 3051 3806
rect 3085 3772 3123 3806
rect 3157 3772 3195 3806
rect 3229 3772 3230 3806
rect 3050 3733 3230 3772
rect 3050 3699 3051 3733
rect 3085 3699 3123 3733
rect 3157 3699 3195 3733
rect 3229 3699 3230 3733
rect 3050 3660 3230 3699
rect 3050 3626 3051 3660
rect 3085 3626 3123 3660
rect 3157 3626 3195 3660
rect 3229 3626 3230 3660
rect 3050 3587 3230 3626
rect 3050 3553 3051 3587
rect 3085 3553 3123 3587
rect 3157 3553 3195 3587
rect 3229 3553 3230 3587
rect 3050 3514 3230 3553
rect 3050 3480 3051 3514
rect 3085 3480 3123 3514
rect 3157 3480 3195 3514
rect 3229 3480 3230 3514
rect 3050 3441 3230 3480
rect 3050 3407 3051 3441
rect 3085 3407 3123 3441
rect 3157 3407 3195 3441
rect 3229 3407 3230 3441
rect 3050 3368 3230 3407
rect 3050 3334 3051 3368
rect 3085 3334 3123 3368
rect 3157 3334 3195 3368
rect 3229 3334 3230 3368
rect 3050 3295 3230 3334
rect 3050 3261 3051 3295
rect 3085 3261 3123 3295
rect 3157 3261 3195 3295
rect 3229 3261 3230 3295
rect 3050 3222 3230 3261
rect 3050 3188 3051 3222
rect 3085 3188 3123 3222
rect 3157 3188 3195 3222
rect 3229 3188 3230 3222
rect 3050 3149 3230 3188
rect 3050 3115 3051 3149
rect 3085 3115 3123 3149
rect 3157 3115 3195 3149
rect 3229 3115 3230 3149
rect 3050 3076 3230 3115
rect 3050 3042 3051 3076
rect 3085 3042 3123 3076
rect 3157 3042 3195 3076
rect 3229 3042 3230 3076
rect 3050 3003 3230 3042
rect 3050 2969 3051 3003
rect 3085 2969 3123 3003
rect 3157 2969 3195 3003
rect 3229 2969 3230 3003
rect 3050 2930 3230 2969
rect 3050 2896 3051 2930
rect 3085 2896 3123 2930
rect 3157 2896 3195 2930
rect 3229 2896 3230 2930
rect 3050 2857 3230 2896
rect 3050 2823 3051 2857
rect 3085 2823 3123 2857
rect 3157 2823 3195 2857
rect 3229 2823 3230 2857
rect 3050 2784 3230 2823
rect 3050 2750 3051 2784
rect 3085 2750 3123 2784
rect 3157 2750 3195 2784
rect 3229 2750 3230 2784
rect 3050 2711 3230 2750
rect 3050 2677 3051 2711
rect 3085 2677 3123 2711
rect 3157 2677 3195 2711
rect 3229 2677 3230 2711
rect 3050 2638 3230 2677
rect 3050 2604 3051 2638
rect 3085 2604 3123 2638
rect 3157 2604 3195 2638
rect 3229 2604 3230 2638
rect 3050 2565 3230 2604
rect 3050 2531 3051 2565
rect 3085 2531 3123 2565
rect 3157 2531 3195 2565
rect 3229 2531 3230 2565
rect 3050 2492 3230 2531
rect 3050 2458 3051 2492
rect 3085 2458 3123 2492
rect 3157 2458 3195 2492
rect 3229 2458 3230 2492
rect 3050 2419 3230 2458
rect 3050 2385 3051 2419
rect 3085 2385 3123 2419
rect 3157 2385 3195 2419
rect 3229 2385 3230 2419
rect 3050 2346 3230 2385
rect 3050 2312 3051 2346
rect 3085 2312 3123 2346
rect 3157 2312 3195 2346
rect 3229 2312 3230 2346
rect 3050 2273 3230 2312
rect 3050 2239 3051 2273
rect 3085 2239 3123 2273
rect 3157 2239 3195 2273
rect 3229 2239 3230 2273
rect 3050 2200 3230 2239
rect 3050 2166 3051 2200
rect 3085 2166 3123 2200
rect 3157 2166 3195 2200
rect 3229 2166 3230 2200
rect 3050 2126 3230 2166
rect 3050 2092 3051 2126
rect 3085 2092 3123 2126
rect 3157 2092 3195 2126
rect 3229 2092 3230 2126
rect 3050 2052 3230 2092
rect 3050 2018 3051 2052
rect 3085 2018 3123 2052
rect 3157 2018 3195 2052
rect 3229 2018 3230 2052
rect 3050 1978 3230 2018
rect 3050 1944 3051 1978
rect 3085 1944 3123 1978
rect 3157 1944 3195 1978
rect 3229 1944 3230 1978
rect 3050 1904 3230 1944
rect 3050 1870 3051 1904
rect 3085 1870 3123 1904
rect 3157 1870 3195 1904
rect 3229 1870 3230 1904
rect 3050 1830 3230 1870
rect 3050 1796 3051 1830
rect 3085 1796 3123 1830
rect 3157 1796 3195 1830
rect 3229 1796 3230 1830
rect 3050 1756 3230 1796
rect 3050 1722 3051 1756
rect 3085 1722 3123 1756
rect 3157 1722 3195 1756
rect 3229 1722 3230 1756
rect 3050 1682 3230 1722
rect 3050 1648 3051 1682
rect 3085 1648 3123 1682
rect 3157 1648 3195 1682
rect 3229 1648 3230 1682
rect 3050 1608 3230 1648
rect 3050 1574 3051 1608
rect 3085 1574 3123 1608
rect 3157 1574 3195 1608
rect 3229 1574 3230 1608
rect 3050 1548 3230 1574
rect 3295 3104 3415 4200
rect 3857 4308 3977 4324
rect 3857 4274 3900 4308
rect 3934 4274 3977 4308
rect 3857 4234 3977 4274
rect 3857 4200 3900 4234
rect 3934 4200 3977 4234
rect 3295 3070 3338 3104
rect 3372 3070 3415 3104
rect 3295 3026 3415 3070
rect 3295 2992 3338 3026
rect 3372 2992 3415 3026
rect 3295 2948 3415 2992
rect 3295 2914 3338 2948
rect 3372 2914 3415 2948
rect 3295 2870 3415 2914
rect 3295 2836 3338 2870
rect 3372 2836 3415 2870
rect 3295 2792 3415 2836
rect 3295 2758 3338 2792
rect 3372 2758 3415 2792
rect 3295 2713 3415 2758
rect 3295 2679 3338 2713
rect 3372 2679 3415 2713
rect 3295 2634 3415 2679
rect 3295 2600 3338 2634
rect 3372 2600 3415 2634
rect 2865 1470 2908 1504
rect 2942 1470 2985 1504
rect 2865 1430 2985 1470
rect 2865 1396 2908 1430
rect 2942 1396 2985 1430
rect 2865 1250 2985 1396
rect 2865 1144 2872 1250
rect 2978 1144 2985 1250
rect 3295 1504 3415 2600
rect 3517 4092 3755 4104
rect 3517 4058 3547 4092
rect 3581 4058 3691 4092
rect 3725 4058 3755 4092
rect 3517 4020 3755 4058
rect 3517 3986 3547 4020
rect 3581 3986 3691 4020
rect 3725 3986 3755 4020
rect 3517 3948 3755 3986
rect 3517 3914 3547 3948
rect 3581 3914 3691 3948
rect 3725 3914 3755 3948
rect 3517 3876 3755 3914
rect 3517 3842 3547 3876
rect 3581 3842 3691 3876
rect 3725 3842 3755 3876
rect 3517 3804 3755 3842
rect 3517 3770 3547 3804
rect 3581 3770 3691 3804
rect 3725 3770 3755 3804
rect 3517 3732 3755 3770
rect 3517 3698 3547 3732
rect 3581 3698 3691 3732
rect 3725 3698 3755 3732
rect 3517 3660 3755 3698
rect 3517 3626 3547 3660
rect 3581 3626 3691 3660
rect 3725 3626 3755 3660
rect 3517 3588 3755 3626
rect 3517 3554 3547 3588
rect 3581 3554 3691 3588
rect 3725 3554 3755 3588
rect 3517 3516 3755 3554
rect 3517 3482 3547 3516
rect 3581 3482 3691 3516
rect 3725 3482 3755 3516
rect 3517 3444 3755 3482
rect 3517 3410 3547 3444
rect 3581 3410 3691 3444
rect 3725 3410 3755 3444
rect 3517 3372 3755 3410
rect 3517 3338 3547 3372
rect 3581 3338 3691 3372
rect 3725 3338 3755 3372
rect 3517 3300 3755 3338
rect 3517 3266 3547 3300
rect 3581 3266 3691 3300
rect 3725 3266 3755 3300
rect 3517 3228 3755 3266
rect 3517 3194 3547 3228
rect 3581 3194 3691 3228
rect 3725 3194 3755 3228
rect 3517 3108 3755 3194
rect 3517 3074 3547 3108
rect 3581 3074 3619 3108
rect 3653 3074 3691 3108
rect 3725 3074 3755 3108
rect 3517 3044 3755 3074
rect 3517 3028 3585 3044
rect 3517 2994 3547 3028
rect 3581 3010 3585 3028
rect 3619 3028 3653 3044
rect 3581 2994 3619 3010
rect 3687 3028 3755 3044
rect 3687 3010 3691 3028
rect 3653 2994 3691 3010
rect 3725 2994 3755 3028
rect 3517 2974 3755 2994
rect 3517 2948 3585 2974
rect 3517 2914 3547 2948
rect 3581 2940 3585 2948
rect 3619 2948 3653 2974
rect 3581 2914 3619 2940
rect 3687 2948 3755 2974
rect 3687 2940 3691 2948
rect 3653 2914 3691 2940
rect 3725 2914 3755 2948
rect 3517 2904 3755 2914
rect 3517 2870 3585 2904
rect 3619 2870 3653 2904
rect 3687 2870 3755 2904
rect 3517 2868 3755 2870
rect 3517 2834 3547 2868
rect 3581 2834 3619 2868
rect 3653 2834 3691 2868
rect 3725 2834 3755 2868
rect 3517 2800 3585 2834
rect 3619 2800 3653 2834
rect 3687 2800 3755 2834
rect 3517 2788 3755 2800
rect 3517 2754 3547 2788
rect 3581 2764 3619 2788
rect 3581 2754 3585 2764
rect 3517 2730 3585 2754
rect 3653 2764 3691 2788
rect 3619 2730 3653 2754
rect 3687 2754 3691 2764
rect 3725 2754 3755 2788
rect 3687 2730 3755 2754
rect 3517 2708 3755 2730
rect 3517 2674 3547 2708
rect 3581 2694 3619 2708
rect 3581 2674 3585 2694
rect 3517 2660 3585 2674
rect 3653 2694 3691 2708
rect 3619 2660 3653 2674
rect 3687 2674 3691 2694
rect 3725 2674 3755 2708
rect 3687 2660 3755 2674
rect 3517 2628 3755 2660
rect 3517 2594 3547 2628
rect 3581 2594 3619 2628
rect 3653 2594 3691 2628
rect 3725 2594 3755 2628
rect 3517 2518 3755 2594
rect 3517 2484 3547 2518
rect 3581 2484 3691 2518
rect 3725 2484 3755 2518
rect 3517 2446 3755 2484
rect 3517 2412 3547 2446
rect 3581 2412 3691 2446
rect 3725 2412 3755 2446
rect 3517 2374 3755 2412
rect 3517 2340 3547 2374
rect 3581 2340 3691 2374
rect 3725 2340 3755 2374
rect 3517 2302 3755 2340
rect 3517 2268 3547 2302
rect 3581 2268 3691 2302
rect 3725 2268 3755 2302
rect 3517 2230 3755 2268
rect 3517 2196 3547 2230
rect 3581 2196 3691 2230
rect 3725 2196 3755 2230
rect 3517 2158 3755 2196
rect 3517 2124 3547 2158
rect 3581 2124 3691 2158
rect 3725 2124 3755 2158
rect 3517 2086 3755 2124
rect 3517 2052 3547 2086
rect 3581 2052 3691 2086
rect 3725 2052 3755 2086
rect 3517 2014 3755 2052
rect 3517 1980 3547 2014
rect 3581 1980 3691 2014
rect 3725 1980 3755 2014
rect 3517 1942 3755 1980
rect 3517 1908 3547 1942
rect 3581 1908 3691 1942
rect 3725 1908 3755 1942
rect 3517 1870 3755 1908
rect 3517 1836 3547 1870
rect 3581 1836 3691 1870
rect 3725 1836 3755 1870
rect 3517 1798 3755 1836
rect 3517 1764 3547 1798
rect 3581 1764 3691 1798
rect 3725 1764 3755 1798
rect 3517 1726 3755 1764
rect 3517 1692 3547 1726
rect 3581 1692 3691 1726
rect 3725 1692 3755 1726
rect 3517 1654 3755 1692
rect 3517 1620 3547 1654
rect 3581 1620 3691 1654
rect 3725 1620 3755 1654
rect 3517 1536 3755 1620
rect 3857 3104 3977 4200
rect 4287 4308 4407 4324
rect 4287 4274 4330 4308
rect 4364 4274 4407 4308
rect 4287 4234 4407 4274
rect 4287 4200 4330 4234
rect 4364 4200 4407 4234
rect 3857 3070 3900 3104
rect 3934 3070 3977 3104
rect 3857 3026 3977 3070
rect 3857 2992 3900 3026
rect 3934 2992 3977 3026
rect 3857 2948 3977 2992
rect 3857 2914 3900 2948
rect 3934 2914 3977 2948
rect 3857 2870 3977 2914
rect 3857 2836 3900 2870
rect 3934 2836 3977 2870
rect 3857 2792 3977 2836
rect 3857 2758 3900 2792
rect 3934 2758 3977 2792
rect 3857 2713 3977 2758
rect 3857 2679 3900 2713
rect 3934 2679 3977 2713
rect 3857 2634 3977 2679
rect 3857 2600 3900 2634
rect 3934 2600 3977 2634
rect 3295 1470 3338 1504
rect 3372 1470 3415 1504
rect 3295 1430 3415 1470
rect 3295 1396 3338 1430
rect 3372 1396 3415 1430
rect 3295 1250 3415 1396
rect 3295 1144 3302 1250
rect 3408 1144 3415 1250
rect 3857 1504 3977 2600
rect 4042 4064 4043 4098
rect 4077 4064 4115 4098
rect 4149 4064 4187 4098
rect 4221 4064 4222 4098
rect 4042 4025 4222 4064
rect 4042 3991 4043 4025
rect 4077 3991 4115 4025
rect 4149 3991 4187 4025
rect 4221 3991 4222 4025
rect 4042 3952 4222 3991
rect 4042 3918 4043 3952
rect 4077 3918 4115 3952
rect 4149 3918 4187 3952
rect 4221 3918 4222 3952
rect 4042 3879 4222 3918
rect 4042 3845 4043 3879
rect 4077 3845 4115 3879
rect 4149 3845 4187 3879
rect 4221 3845 4222 3879
rect 4042 3806 4222 3845
rect 4042 3772 4043 3806
rect 4077 3772 4115 3806
rect 4149 3772 4187 3806
rect 4221 3772 4222 3806
rect 4042 3733 4222 3772
rect 4042 3699 4043 3733
rect 4077 3699 4115 3733
rect 4149 3699 4187 3733
rect 4221 3699 4222 3733
rect 4042 3660 4222 3699
rect 4042 3626 4043 3660
rect 4077 3626 4115 3660
rect 4149 3626 4187 3660
rect 4221 3626 4222 3660
rect 4042 3587 4222 3626
rect 4042 3553 4043 3587
rect 4077 3553 4115 3587
rect 4149 3553 4187 3587
rect 4221 3553 4222 3587
rect 4042 3514 4222 3553
rect 4042 3480 4043 3514
rect 4077 3480 4115 3514
rect 4149 3480 4187 3514
rect 4221 3480 4222 3514
rect 4042 3441 4222 3480
rect 4042 3407 4043 3441
rect 4077 3407 4115 3441
rect 4149 3407 4187 3441
rect 4221 3407 4222 3441
rect 4042 3368 4222 3407
rect 4042 3334 4043 3368
rect 4077 3334 4115 3368
rect 4149 3334 4187 3368
rect 4221 3334 4222 3368
rect 4042 3295 4222 3334
rect 4042 3261 4043 3295
rect 4077 3261 4115 3295
rect 4149 3261 4187 3295
rect 4221 3261 4222 3295
rect 4042 3222 4222 3261
rect 4042 3188 4043 3222
rect 4077 3188 4115 3222
rect 4149 3188 4187 3222
rect 4221 3188 4222 3222
rect 4042 3149 4222 3188
rect 4042 3115 4043 3149
rect 4077 3115 4115 3149
rect 4149 3115 4187 3149
rect 4221 3115 4222 3149
rect 4042 3076 4222 3115
rect 4042 3042 4043 3076
rect 4077 3042 4115 3076
rect 4149 3042 4187 3076
rect 4221 3042 4222 3076
rect 4042 3003 4222 3042
rect 4042 2969 4043 3003
rect 4077 2969 4115 3003
rect 4149 2969 4187 3003
rect 4221 2969 4222 3003
rect 4042 2930 4222 2969
rect 4042 2896 4043 2930
rect 4077 2896 4115 2930
rect 4149 2896 4187 2930
rect 4221 2896 4222 2930
rect 4042 2857 4222 2896
rect 4042 2823 4043 2857
rect 4077 2823 4115 2857
rect 4149 2823 4187 2857
rect 4221 2823 4222 2857
rect 4042 2784 4222 2823
rect 4042 2750 4043 2784
rect 4077 2750 4115 2784
rect 4149 2750 4187 2784
rect 4221 2750 4222 2784
rect 4042 2711 4222 2750
rect 4042 2677 4043 2711
rect 4077 2677 4115 2711
rect 4149 2677 4187 2711
rect 4221 2677 4222 2711
rect 4042 2638 4222 2677
rect 4042 2604 4043 2638
rect 4077 2604 4115 2638
rect 4149 2604 4187 2638
rect 4221 2604 4222 2638
rect 4042 2565 4222 2604
rect 4042 2531 4043 2565
rect 4077 2531 4115 2565
rect 4149 2531 4187 2565
rect 4221 2531 4222 2565
rect 4042 2492 4222 2531
rect 4042 2458 4043 2492
rect 4077 2458 4115 2492
rect 4149 2458 4187 2492
rect 4221 2458 4222 2492
rect 4042 2419 4222 2458
rect 4042 2385 4043 2419
rect 4077 2385 4115 2419
rect 4149 2385 4187 2419
rect 4221 2385 4222 2419
rect 4042 2346 4222 2385
rect 4042 2312 4043 2346
rect 4077 2312 4115 2346
rect 4149 2312 4187 2346
rect 4221 2312 4222 2346
rect 4042 2273 4222 2312
rect 4042 2239 4043 2273
rect 4077 2239 4115 2273
rect 4149 2239 4187 2273
rect 4221 2239 4222 2273
rect 4042 2200 4222 2239
rect 4042 2166 4043 2200
rect 4077 2166 4115 2200
rect 4149 2166 4187 2200
rect 4221 2166 4222 2200
rect 4042 2126 4222 2166
rect 4042 2092 4043 2126
rect 4077 2092 4115 2126
rect 4149 2092 4187 2126
rect 4221 2092 4222 2126
rect 4042 2052 4222 2092
rect 4042 2018 4043 2052
rect 4077 2018 4115 2052
rect 4149 2018 4187 2052
rect 4221 2018 4222 2052
rect 4042 1978 4222 2018
rect 4042 1944 4043 1978
rect 4077 1944 4115 1978
rect 4149 1944 4187 1978
rect 4221 1944 4222 1978
rect 4042 1904 4222 1944
rect 4042 1870 4043 1904
rect 4077 1870 4115 1904
rect 4149 1870 4187 1904
rect 4221 1870 4222 1904
rect 4042 1830 4222 1870
rect 4042 1796 4043 1830
rect 4077 1796 4115 1830
rect 4149 1796 4187 1830
rect 4221 1796 4222 1830
rect 4042 1756 4222 1796
rect 4042 1722 4043 1756
rect 4077 1722 4115 1756
rect 4149 1722 4187 1756
rect 4221 1722 4222 1756
rect 4042 1682 4222 1722
rect 4042 1648 4043 1682
rect 4077 1648 4115 1682
rect 4149 1648 4187 1682
rect 4221 1648 4222 1682
rect 4042 1608 4222 1648
rect 4042 1574 4043 1608
rect 4077 1574 4115 1608
rect 4149 1574 4187 1608
rect 4221 1574 4222 1608
rect 4042 1548 4222 1574
rect 4287 3104 4407 4200
rect 4849 4308 4969 4324
rect 4849 4274 4892 4308
rect 4926 4274 4969 4308
rect 4849 4234 4969 4274
rect 4849 4200 4892 4234
rect 4926 4200 4969 4234
rect 4287 3070 4330 3104
rect 4364 3070 4407 3104
rect 4287 3026 4407 3070
rect 4287 2992 4330 3026
rect 4364 2992 4407 3026
rect 4287 2948 4407 2992
rect 4287 2914 4330 2948
rect 4364 2914 4407 2948
rect 4287 2870 4407 2914
rect 4287 2836 4330 2870
rect 4364 2836 4407 2870
rect 4287 2792 4407 2836
rect 4287 2758 4330 2792
rect 4364 2758 4407 2792
rect 4287 2713 4407 2758
rect 4287 2679 4330 2713
rect 4364 2679 4407 2713
rect 4287 2634 4407 2679
rect 4287 2600 4330 2634
rect 4364 2600 4407 2634
rect 3857 1470 3900 1504
rect 3934 1470 3977 1504
rect 3857 1430 3977 1470
rect 3857 1396 3900 1430
rect 3934 1396 3977 1430
rect 3857 1250 3977 1396
rect 3857 1144 3864 1250
rect 3970 1144 3977 1250
rect 4287 1504 4407 2600
rect 4509 4092 4747 4104
rect 4509 4058 4539 4092
rect 4573 4058 4683 4092
rect 4717 4058 4747 4092
rect 4509 4020 4747 4058
rect 4509 3986 4539 4020
rect 4573 3986 4683 4020
rect 4717 3986 4747 4020
rect 4509 3948 4747 3986
rect 4509 3914 4539 3948
rect 4573 3914 4683 3948
rect 4717 3914 4747 3948
rect 4509 3876 4747 3914
rect 4509 3842 4539 3876
rect 4573 3842 4683 3876
rect 4717 3842 4747 3876
rect 4509 3804 4747 3842
rect 4509 3770 4539 3804
rect 4573 3770 4683 3804
rect 4717 3770 4747 3804
rect 4509 3732 4747 3770
rect 4509 3698 4539 3732
rect 4573 3698 4683 3732
rect 4717 3698 4747 3732
rect 4509 3660 4747 3698
rect 4509 3626 4539 3660
rect 4573 3626 4683 3660
rect 4717 3626 4747 3660
rect 4509 3588 4747 3626
rect 4509 3554 4539 3588
rect 4573 3554 4683 3588
rect 4717 3554 4747 3588
rect 4509 3516 4747 3554
rect 4509 3482 4539 3516
rect 4573 3482 4683 3516
rect 4717 3482 4747 3516
rect 4509 3444 4747 3482
rect 4509 3410 4539 3444
rect 4573 3410 4683 3444
rect 4717 3410 4747 3444
rect 4509 3372 4747 3410
rect 4509 3338 4539 3372
rect 4573 3338 4683 3372
rect 4717 3338 4747 3372
rect 4509 3300 4747 3338
rect 4509 3266 4539 3300
rect 4573 3266 4683 3300
rect 4717 3266 4747 3300
rect 4509 3228 4747 3266
rect 4509 3194 4539 3228
rect 4573 3194 4683 3228
rect 4717 3194 4747 3228
rect 4509 3108 4747 3194
rect 4509 3074 4539 3108
rect 4573 3074 4611 3108
rect 4645 3074 4683 3108
rect 4717 3074 4747 3108
rect 4509 3044 4747 3074
rect 4509 3028 4577 3044
rect 4509 2994 4539 3028
rect 4573 3010 4577 3028
rect 4611 3028 4645 3044
rect 4573 2994 4611 3010
rect 4679 3028 4747 3044
rect 4679 3010 4683 3028
rect 4645 2994 4683 3010
rect 4717 2994 4747 3028
rect 4509 2974 4747 2994
rect 4509 2948 4577 2974
rect 4509 2914 4539 2948
rect 4573 2940 4577 2948
rect 4611 2948 4645 2974
rect 4573 2914 4611 2940
rect 4679 2948 4747 2974
rect 4679 2940 4683 2948
rect 4645 2914 4683 2940
rect 4717 2914 4747 2948
rect 4509 2904 4747 2914
rect 4509 2870 4577 2904
rect 4611 2870 4645 2904
rect 4679 2870 4747 2904
rect 4509 2868 4747 2870
rect 4509 2834 4539 2868
rect 4573 2834 4611 2868
rect 4645 2834 4683 2868
rect 4717 2834 4747 2868
rect 4509 2800 4577 2834
rect 4611 2800 4645 2834
rect 4679 2800 4747 2834
rect 4509 2788 4747 2800
rect 4509 2754 4539 2788
rect 4573 2764 4611 2788
rect 4573 2754 4577 2764
rect 4509 2730 4577 2754
rect 4645 2764 4683 2788
rect 4611 2730 4645 2754
rect 4679 2754 4683 2764
rect 4717 2754 4747 2788
rect 4679 2730 4747 2754
rect 4509 2708 4747 2730
rect 4509 2674 4539 2708
rect 4573 2694 4611 2708
rect 4573 2674 4577 2694
rect 4509 2660 4577 2674
rect 4645 2694 4683 2708
rect 4611 2660 4645 2674
rect 4679 2674 4683 2694
rect 4717 2674 4747 2708
rect 4679 2660 4747 2674
rect 4509 2628 4747 2660
rect 4509 2594 4539 2628
rect 4573 2594 4611 2628
rect 4645 2594 4683 2628
rect 4717 2594 4747 2628
rect 4509 2518 4747 2594
rect 4509 2484 4539 2518
rect 4573 2484 4683 2518
rect 4717 2484 4747 2518
rect 4509 2446 4747 2484
rect 4509 2412 4539 2446
rect 4573 2412 4683 2446
rect 4717 2412 4747 2446
rect 4509 2374 4747 2412
rect 4509 2340 4539 2374
rect 4573 2340 4683 2374
rect 4717 2340 4747 2374
rect 4509 2302 4747 2340
rect 4509 2268 4539 2302
rect 4573 2268 4683 2302
rect 4717 2268 4747 2302
rect 4509 2230 4747 2268
rect 4509 2196 4539 2230
rect 4573 2196 4683 2230
rect 4717 2196 4747 2230
rect 4509 2158 4747 2196
rect 4509 2124 4539 2158
rect 4573 2124 4683 2158
rect 4717 2124 4747 2158
rect 4509 2086 4747 2124
rect 4509 2052 4539 2086
rect 4573 2052 4683 2086
rect 4717 2052 4747 2086
rect 4509 2014 4747 2052
rect 4509 1980 4539 2014
rect 4573 1980 4683 2014
rect 4717 1980 4747 2014
rect 4509 1942 4747 1980
rect 4509 1908 4539 1942
rect 4573 1908 4683 1942
rect 4717 1908 4747 1942
rect 4509 1870 4747 1908
rect 4509 1836 4539 1870
rect 4573 1836 4683 1870
rect 4717 1836 4747 1870
rect 4509 1798 4747 1836
rect 4509 1764 4539 1798
rect 4573 1764 4683 1798
rect 4717 1764 4747 1798
rect 4509 1726 4747 1764
rect 4509 1692 4539 1726
rect 4573 1692 4683 1726
rect 4717 1692 4747 1726
rect 4509 1654 4747 1692
rect 4509 1620 4539 1654
rect 4573 1620 4683 1654
rect 4717 1620 4747 1654
rect 4509 1536 4747 1620
rect 4849 3104 4969 4200
rect 5279 4308 5399 4324
rect 5279 4274 5322 4308
rect 5356 4274 5399 4308
rect 5279 4234 5399 4274
rect 5279 4200 5322 4234
rect 5356 4200 5399 4234
rect 4849 3070 4892 3104
rect 4926 3070 4969 3104
rect 4849 3026 4969 3070
rect 4849 2992 4892 3026
rect 4926 2992 4969 3026
rect 4849 2948 4969 2992
rect 4849 2914 4892 2948
rect 4926 2914 4969 2948
rect 4849 2870 4969 2914
rect 4849 2836 4892 2870
rect 4926 2836 4969 2870
rect 4849 2792 4969 2836
rect 4849 2758 4892 2792
rect 4926 2758 4969 2792
rect 4849 2713 4969 2758
rect 4849 2679 4892 2713
rect 4926 2679 4969 2713
rect 4849 2634 4969 2679
rect 4849 2600 4892 2634
rect 4926 2600 4969 2634
rect 4287 1470 4330 1504
rect 4364 1470 4407 1504
rect 4287 1430 4407 1470
rect 4287 1396 4330 1430
rect 4364 1396 4407 1430
rect 4287 1250 4407 1396
rect 4287 1144 4294 1250
rect 4400 1144 4407 1250
rect 4849 1504 4969 2600
rect 5034 4064 5035 4098
rect 5069 4064 5107 4098
rect 5141 4064 5179 4098
rect 5213 4064 5214 4098
rect 5034 4025 5214 4064
rect 5034 3991 5035 4025
rect 5069 3991 5107 4025
rect 5141 3991 5179 4025
rect 5213 3991 5214 4025
rect 5034 3952 5214 3991
rect 5034 3918 5035 3952
rect 5069 3918 5107 3952
rect 5141 3918 5179 3952
rect 5213 3918 5214 3952
rect 5034 3879 5214 3918
rect 5034 3845 5035 3879
rect 5069 3845 5107 3879
rect 5141 3845 5179 3879
rect 5213 3845 5214 3879
rect 5034 3806 5214 3845
rect 5034 3772 5035 3806
rect 5069 3772 5107 3806
rect 5141 3772 5179 3806
rect 5213 3772 5214 3806
rect 5034 3733 5214 3772
rect 5034 3699 5035 3733
rect 5069 3699 5107 3733
rect 5141 3699 5179 3733
rect 5213 3699 5214 3733
rect 5034 3660 5214 3699
rect 5034 3626 5035 3660
rect 5069 3626 5107 3660
rect 5141 3626 5179 3660
rect 5213 3626 5214 3660
rect 5034 3587 5214 3626
rect 5034 3553 5035 3587
rect 5069 3553 5107 3587
rect 5141 3553 5179 3587
rect 5213 3553 5214 3587
rect 5034 3514 5214 3553
rect 5034 3480 5035 3514
rect 5069 3480 5107 3514
rect 5141 3480 5179 3514
rect 5213 3480 5214 3514
rect 5034 3441 5214 3480
rect 5034 3407 5035 3441
rect 5069 3407 5107 3441
rect 5141 3407 5179 3441
rect 5213 3407 5214 3441
rect 5034 3368 5214 3407
rect 5034 3334 5035 3368
rect 5069 3334 5107 3368
rect 5141 3334 5179 3368
rect 5213 3334 5214 3368
rect 5034 3295 5214 3334
rect 5034 3261 5035 3295
rect 5069 3261 5107 3295
rect 5141 3261 5179 3295
rect 5213 3261 5214 3295
rect 5034 3222 5214 3261
rect 5034 3188 5035 3222
rect 5069 3188 5107 3222
rect 5141 3188 5179 3222
rect 5213 3188 5214 3222
rect 5034 3149 5214 3188
rect 5034 3115 5035 3149
rect 5069 3115 5107 3149
rect 5141 3115 5179 3149
rect 5213 3115 5214 3149
rect 5034 3076 5214 3115
rect 5034 3042 5035 3076
rect 5069 3042 5107 3076
rect 5141 3042 5179 3076
rect 5213 3042 5214 3076
rect 5034 3003 5214 3042
rect 5034 2969 5035 3003
rect 5069 2969 5107 3003
rect 5141 2969 5179 3003
rect 5213 2969 5214 3003
rect 5034 2930 5214 2969
rect 5034 2896 5035 2930
rect 5069 2896 5107 2930
rect 5141 2896 5179 2930
rect 5213 2896 5214 2930
rect 5034 2857 5214 2896
rect 5034 2823 5035 2857
rect 5069 2823 5107 2857
rect 5141 2823 5179 2857
rect 5213 2823 5214 2857
rect 5034 2784 5214 2823
rect 5034 2750 5035 2784
rect 5069 2750 5107 2784
rect 5141 2750 5179 2784
rect 5213 2750 5214 2784
rect 5034 2711 5214 2750
rect 5034 2677 5035 2711
rect 5069 2677 5107 2711
rect 5141 2677 5179 2711
rect 5213 2677 5214 2711
rect 5034 2638 5214 2677
rect 5034 2604 5035 2638
rect 5069 2604 5107 2638
rect 5141 2604 5179 2638
rect 5213 2604 5214 2638
rect 5034 2565 5214 2604
rect 5034 2531 5035 2565
rect 5069 2531 5107 2565
rect 5141 2531 5179 2565
rect 5213 2531 5214 2565
rect 5034 2492 5214 2531
rect 5034 2458 5035 2492
rect 5069 2458 5107 2492
rect 5141 2458 5179 2492
rect 5213 2458 5214 2492
rect 5034 2419 5214 2458
rect 5034 2385 5035 2419
rect 5069 2385 5107 2419
rect 5141 2385 5179 2419
rect 5213 2385 5214 2419
rect 5034 2346 5214 2385
rect 5034 2312 5035 2346
rect 5069 2312 5107 2346
rect 5141 2312 5179 2346
rect 5213 2312 5214 2346
rect 5034 2273 5214 2312
rect 5034 2239 5035 2273
rect 5069 2239 5107 2273
rect 5141 2239 5179 2273
rect 5213 2239 5214 2273
rect 5034 2200 5214 2239
rect 5034 2166 5035 2200
rect 5069 2166 5107 2200
rect 5141 2166 5179 2200
rect 5213 2166 5214 2200
rect 5034 2126 5214 2166
rect 5034 2092 5035 2126
rect 5069 2092 5107 2126
rect 5141 2092 5179 2126
rect 5213 2092 5214 2126
rect 5034 2052 5214 2092
rect 5034 2018 5035 2052
rect 5069 2018 5107 2052
rect 5141 2018 5179 2052
rect 5213 2018 5214 2052
rect 5034 1978 5214 2018
rect 5034 1944 5035 1978
rect 5069 1944 5107 1978
rect 5141 1944 5179 1978
rect 5213 1944 5214 1978
rect 5034 1904 5214 1944
rect 5034 1870 5035 1904
rect 5069 1870 5107 1904
rect 5141 1870 5179 1904
rect 5213 1870 5214 1904
rect 5034 1830 5214 1870
rect 5034 1796 5035 1830
rect 5069 1796 5107 1830
rect 5141 1796 5179 1830
rect 5213 1796 5214 1830
rect 5034 1756 5214 1796
rect 5034 1722 5035 1756
rect 5069 1722 5107 1756
rect 5141 1722 5179 1756
rect 5213 1722 5214 1756
rect 5034 1682 5214 1722
rect 5034 1648 5035 1682
rect 5069 1648 5107 1682
rect 5141 1648 5179 1682
rect 5213 1648 5214 1682
rect 5034 1608 5214 1648
rect 5034 1574 5035 1608
rect 5069 1574 5107 1608
rect 5141 1574 5179 1608
rect 5213 1574 5214 1608
rect 5034 1548 5214 1574
rect 5279 3104 5399 4200
rect 5841 4308 5961 4324
rect 5841 4274 5884 4308
rect 5918 4274 5961 4308
rect 5841 4234 5961 4274
rect 5841 4200 5884 4234
rect 5918 4200 5961 4234
rect 5279 3070 5322 3104
rect 5356 3070 5399 3104
rect 5279 3026 5399 3070
rect 5279 2992 5322 3026
rect 5356 2992 5399 3026
rect 5279 2948 5399 2992
rect 5279 2914 5322 2948
rect 5356 2914 5399 2948
rect 5279 2870 5399 2914
rect 5279 2836 5322 2870
rect 5356 2836 5399 2870
rect 5279 2792 5399 2836
rect 5279 2758 5322 2792
rect 5356 2758 5399 2792
rect 5279 2713 5399 2758
rect 5279 2679 5322 2713
rect 5356 2679 5399 2713
rect 5279 2634 5399 2679
rect 5279 2600 5322 2634
rect 5356 2600 5399 2634
rect 4849 1470 4892 1504
rect 4926 1470 4969 1504
rect 4849 1430 4969 1470
rect 4849 1396 4892 1430
rect 4926 1396 4969 1430
rect 4849 1250 4969 1396
rect 4849 1144 4856 1250
rect 4962 1144 4969 1250
rect 5279 1504 5399 2600
rect 5501 4092 5739 4104
rect 5501 4058 5531 4092
rect 5565 4058 5675 4092
rect 5709 4058 5739 4092
rect 5501 4020 5739 4058
rect 5501 3986 5531 4020
rect 5565 3986 5675 4020
rect 5709 3986 5739 4020
rect 5501 3948 5739 3986
rect 5501 3914 5531 3948
rect 5565 3914 5675 3948
rect 5709 3914 5739 3948
rect 5501 3876 5739 3914
rect 5501 3842 5531 3876
rect 5565 3842 5675 3876
rect 5709 3842 5739 3876
rect 5501 3804 5739 3842
rect 5501 3770 5531 3804
rect 5565 3770 5675 3804
rect 5709 3770 5739 3804
rect 5501 3732 5739 3770
rect 5501 3698 5531 3732
rect 5565 3698 5675 3732
rect 5709 3698 5739 3732
rect 5501 3660 5739 3698
rect 5501 3626 5531 3660
rect 5565 3626 5675 3660
rect 5709 3626 5739 3660
rect 5501 3588 5739 3626
rect 5501 3554 5531 3588
rect 5565 3554 5675 3588
rect 5709 3554 5739 3588
rect 5501 3516 5739 3554
rect 5501 3482 5531 3516
rect 5565 3482 5675 3516
rect 5709 3482 5739 3516
rect 5501 3444 5739 3482
rect 5501 3410 5531 3444
rect 5565 3410 5675 3444
rect 5709 3410 5739 3444
rect 5501 3372 5739 3410
rect 5501 3338 5531 3372
rect 5565 3338 5675 3372
rect 5709 3338 5739 3372
rect 5501 3300 5739 3338
rect 5501 3266 5531 3300
rect 5565 3266 5675 3300
rect 5709 3266 5739 3300
rect 5501 3228 5739 3266
rect 5501 3194 5531 3228
rect 5565 3194 5675 3228
rect 5709 3194 5739 3228
rect 5501 3108 5739 3194
rect 5501 3074 5531 3108
rect 5565 3074 5603 3108
rect 5637 3074 5675 3108
rect 5709 3074 5739 3108
rect 5501 3044 5739 3074
rect 5501 3028 5569 3044
rect 5501 2994 5531 3028
rect 5565 3010 5569 3028
rect 5603 3028 5637 3044
rect 5565 2994 5603 3010
rect 5671 3028 5739 3044
rect 5671 3010 5675 3028
rect 5637 2994 5675 3010
rect 5709 2994 5739 3028
rect 5501 2974 5739 2994
rect 5501 2948 5569 2974
rect 5501 2914 5531 2948
rect 5565 2940 5569 2948
rect 5603 2948 5637 2974
rect 5565 2914 5603 2940
rect 5671 2948 5739 2974
rect 5671 2940 5675 2948
rect 5637 2914 5675 2940
rect 5709 2914 5739 2948
rect 5501 2904 5739 2914
rect 5501 2870 5569 2904
rect 5603 2870 5637 2904
rect 5671 2870 5739 2904
rect 5501 2868 5739 2870
rect 5501 2834 5531 2868
rect 5565 2834 5603 2868
rect 5637 2834 5675 2868
rect 5709 2834 5739 2868
rect 5501 2800 5569 2834
rect 5603 2800 5637 2834
rect 5671 2800 5739 2834
rect 5501 2788 5739 2800
rect 5501 2754 5531 2788
rect 5565 2764 5603 2788
rect 5565 2754 5569 2764
rect 5501 2730 5569 2754
rect 5637 2764 5675 2788
rect 5603 2730 5637 2754
rect 5671 2754 5675 2764
rect 5709 2754 5739 2788
rect 5671 2730 5739 2754
rect 5501 2708 5739 2730
rect 5501 2674 5531 2708
rect 5565 2694 5603 2708
rect 5565 2674 5569 2694
rect 5501 2660 5569 2674
rect 5637 2694 5675 2708
rect 5603 2660 5637 2674
rect 5671 2674 5675 2694
rect 5709 2674 5739 2708
rect 5671 2660 5739 2674
rect 5501 2628 5739 2660
rect 5501 2594 5531 2628
rect 5565 2594 5603 2628
rect 5637 2594 5675 2628
rect 5709 2594 5739 2628
rect 5501 2518 5739 2594
rect 5501 2484 5531 2518
rect 5565 2484 5675 2518
rect 5709 2484 5739 2518
rect 5501 2446 5739 2484
rect 5501 2412 5531 2446
rect 5565 2412 5675 2446
rect 5709 2412 5739 2446
rect 5501 2374 5739 2412
rect 5501 2340 5531 2374
rect 5565 2340 5675 2374
rect 5709 2340 5739 2374
rect 5501 2302 5739 2340
rect 5501 2268 5531 2302
rect 5565 2268 5675 2302
rect 5709 2268 5739 2302
rect 5501 2230 5739 2268
rect 5501 2196 5531 2230
rect 5565 2196 5675 2230
rect 5709 2196 5739 2230
rect 5501 2158 5739 2196
rect 5501 2124 5531 2158
rect 5565 2124 5675 2158
rect 5709 2124 5739 2158
rect 5501 2086 5739 2124
rect 5501 2052 5531 2086
rect 5565 2052 5675 2086
rect 5709 2052 5739 2086
rect 5501 2014 5739 2052
rect 5501 1980 5531 2014
rect 5565 1980 5675 2014
rect 5709 1980 5739 2014
rect 5501 1942 5739 1980
rect 5501 1908 5531 1942
rect 5565 1908 5675 1942
rect 5709 1908 5739 1942
rect 5501 1870 5739 1908
rect 5501 1836 5531 1870
rect 5565 1836 5675 1870
rect 5709 1836 5739 1870
rect 5501 1798 5739 1836
rect 5501 1764 5531 1798
rect 5565 1764 5675 1798
rect 5709 1764 5739 1798
rect 5501 1726 5739 1764
rect 5501 1692 5531 1726
rect 5565 1692 5675 1726
rect 5709 1692 5739 1726
rect 5501 1654 5739 1692
rect 5501 1620 5531 1654
rect 5565 1620 5675 1654
rect 5709 1620 5739 1654
rect 5501 1536 5739 1620
rect 5841 3104 5961 4200
rect 6271 4308 6391 4324
rect 6271 4274 6314 4308
rect 6348 4274 6391 4308
rect 6271 4234 6391 4274
rect 6271 4200 6314 4234
rect 6348 4200 6391 4234
rect 5841 3070 5884 3104
rect 5918 3070 5961 3104
rect 5841 3026 5961 3070
rect 5841 2992 5884 3026
rect 5918 2992 5961 3026
rect 5841 2948 5961 2992
rect 5841 2914 5884 2948
rect 5918 2914 5961 2948
rect 5841 2870 5961 2914
rect 5841 2836 5884 2870
rect 5918 2836 5961 2870
rect 5841 2792 5961 2836
rect 5841 2758 5884 2792
rect 5918 2758 5961 2792
rect 5841 2713 5961 2758
rect 5841 2679 5884 2713
rect 5918 2679 5961 2713
rect 5841 2634 5961 2679
rect 5841 2600 5884 2634
rect 5918 2600 5961 2634
rect 5279 1470 5322 1504
rect 5356 1470 5399 1504
rect 5279 1430 5399 1470
rect 5279 1396 5322 1430
rect 5356 1396 5399 1430
rect 5279 1250 5399 1396
rect 5279 1144 5286 1250
rect 5392 1144 5399 1250
rect 5841 1504 5961 2600
rect 6026 4064 6027 4098
rect 6061 4064 6099 4098
rect 6133 4064 6171 4098
rect 6205 4064 6206 4098
rect 6026 4025 6206 4064
rect 6026 3991 6027 4025
rect 6061 3991 6099 4025
rect 6133 3991 6171 4025
rect 6205 3991 6206 4025
rect 6026 3952 6206 3991
rect 6026 3918 6027 3952
rect 6061 3918 6099 3952
rect 6133 3918 6171 3952
rect 6205 3918 6206 3952
rect 6026 3879 6206 3918
rect 6026 3845 6027 3879
rect 6061 3845 6099 3879
rect 6133 3845 6171 3879
rect 6205 3845 6206 3879
rect 6026 3806 6206 3845
rect 6026 3772 6027 3806
rect 6061 3772 6099 3806
rect 6133 3772 6171 3806
rect 6205 3772 6206 3806
rect 6026 3733 6206 3772
rect 6026 3699 6027 3733
rect 6061 3699 6099 3733
rect 6133 3699 6171 3733
rect 6205 3699 6206 3733
rect 6026 3660 6206 3699
rect 6026 3626 6027 3660
rect 6061 3626 6099 3660
rect 6133 3626 6171 3660
rect 6205 3626 6206 3660
rect 6026 3587 6206 3626
rect 6026 3553 6027 3587
rect 6061 3553 6099 3587
rect 6133 3553 6171 3587
rect 6205 3553 6206 3587
rect 6026 3514 6206 3553
rect 6026 3480 6027 3514
rect 6061 3480 6099 3514
rect 6133 3480 6171 3514
rect 6205 3480 6206 3514
rect 6026 3441 6206 3480
rect 6026 3407 6027 3441
rect 6061 3407 6099 3441
rect 6133 3407 6171 3441
rect 6205 3407 6206 3441
rect 6026 3368 6206 3407
rect 6026 3334 6027 3368
rect 6061 3334 6099 3368
rect 6133 3334 6171 3368
rect 6205 3334 6206 3368
rect 6026 3295 6206 3334
rect 6026 3261 6027 3295
rect 6061 3261 6099 3295
rect 6133 3261 6171 3295
rect 6205 3261 6206 3295
rect 6026 3222 6206 3261
rect 6026 3188 6027 3222
rect 6061 3188 6099 3222
rect 6133 3188 6171 3222
rect 6205 3188 6206 3222
rect 6026 3149 6206 3188
rect 6026 3115 6027 3149
rect 6061 3115 6099 3149
rect 6133 3115 6171 3149
rect 6205 3115 6206 3149
rect 6026 3076 6206 3115
rect 6026 3042 6027 3076
rect 6061 3042 6099 3076
rect 6133 3042 6171 3076
rect 6205 3042 6206 3076
rect 6026 3003 6206 3042
rect 6026 2969 6027 3003
rect 6061 2969 6099 3003
rect 6133 2969 6171 3003
rect 6205 2969 6206 3003
rect 6026 2930 6206 2969
rect 6026 2896 6027 2930
rect 6061 2896 6099 2930
rect 6133 2896 6171 2930
rect 6205 2896 6206 2930
rect 6026 2857 6206 2896
rect 6026 2823 6027 2857
rect 6061 2823 6099 2857
rect 6133 2823 6171 2857
rect 6205 2823 6206 2857
rect 6026 2784 6206 2823
rect 6026 2750 6027 2784
rect 6061 2750 6099 2784
rect 6133 2750 6171 2784
rect 6205 2750 6206 2784
rect 6026 2711 6206 2750
rect 6026 2677 6027 2711
rect 6061 2677 6099 2711
rect 6133 2677 6171 2711
rect 6205 2677 6206 2711
rect 6026 2638 6206 2677
rect 6026 2604 6027 2638
rect 6061 2604 6099 2638
rect 6133 2604 6171 2638
rect 6205 2604 6206 2638
rect 6026 2565 6206 2604
rect 6026 2531 6027 2565
rect 6061 2531 6099 2565
rect 6133 2531 6171 2565
rect 6205 2531 6206 2565
rect 6026 2492 6206 2531
rect 6026 2458 6027 2492
rect 6061 2458 6099 2492
rect 6133 2458 6171 2492
rect 6205 2458 6206 2492
rect 6026 2419 6206 2458
rect 6026 2385 6027 2419
rect 6061 2385 6099 2419
rect 6133 2385 6171 2419
rect 6205 2385 6206 2419
rect 6026 2346 6206 2385
rect 6026 2312 6027 2346
rect 6061 2312 6099 2346
rect 6133 2312 6171 2346
rect 6205 2312 6206 2346
rect 6026 2273 6206 2312
rect 6026 2239 6027 2273
rect 6061 2239 6099 2273
rect 6133 2239 6171 2273
rect 6205 2239 6206 2273
rect 6026 2200 6206 2239
rect 6026 2166 6027 2200
rect 6061 2166 6099 2200
rect 6133 2166 6171 2200
rect 6205 2166 6206 2200
rect 6026 2126 6206 2166
rect 6026 2092 6027 2126
rect 6061 2092 6099 2126
rect 6133 2092 6171 2126
rect 6205 2092 6206 2126
rect 6026 2052 6206 2092
rect 6026 2018 6027 2052
rect 6061 2018 6099 2052
rect 6133 2018 6171 2052
rect 6205 2018 6206 2052
rect 6026 1978 6206 2018
rect 6026 1944 6027 1978
rect 6061 1944 6099 1978
rect 6133 1944 6171 1978
rect 6205 1944 6206 1978
rect 6026 1904 6206 1944
rect 6026 1870 6027 1904
rect 6061 1870 6099 1904
rect 6133 1870 6171 1904
rect 6205 1870 6206 1904
rect 6026 1830 6206 1870
rect 6026 1796 6027 1830
rect 6061 1796 6099 1830
rect 6133 1796 6171 1830
rect 6205 1796 6206 1830
rect 6026 1756 6206 1796
rect 6026 1722 6027 1756
rect 6061 1722 6099 1756
rect 6133 1722 6171 1756
rect 6205 1722 6206 1756
rect 6026 1682 6206 1722
rect 6026 1648 6027 1682
rect 6061 1648 6099 1682
rect 6133 1648 6171 1682
rect 6205 1648 6206 1682
rect 6026 1608 6206 1648
rect 6026 1574 6027 1608
rect 6061 1574 6099 1608
rect 6133 1574 6171 1608
rect 6205 1574 6206 1608
rect 6026 1548 6206 1574
rect 6271 3104 6391 4200
rect 6833 4308 6953 4324
rect 6833 4274 6876 4308
rect 6910 4274 6953 4308
rect 6833 4234 6953 4274
rect 6833 4200 6876 4234
rect 6910 4200 6953 4234
rect 6271 3070 6314 3104
rect 6348 3070 6391 3104
rect 6271 3026 6391 3070
rect 6271 2992 6314 3026
rect 6348 2992 6391 3026
rect 6271 2948 6391 2992
rect 6271 2914 6314 2948
rect 6348 2914 6391 2948
rect 6271 2870 6391 2914
rect 6271 2836 6314 2870
rect 6348 2836 6391 2870
rect 6271 2792 6391 2836
rect 6271 2758 6314 2792
rect 6348 2758 6391 2792
rect 6271 2713 6391 2758
rect 6271 2679 6314 2713
rect 6348 2679 6391 2713
rect 6271 2634 6391 2679
rect 6271 2600 6314 2634
rect 6348 2600 6391 2634
rect 5841 1470 5884 1504
rect 5918 1470 5961 1504
rect 5841 1430 5961 1470
rect 5841 1396 5884 1430
rect 5918 1396 5961 1430
rect 5841 1250 5961 1396
rect 5841 1144 5848 1250
rect 5954 1144 5961 1250
rect 6271 1504 6391 2600
rect 6493 4092 6731 4104
rect 6493 4058 6523 4092
rect 6557 4058 6667 4092
rect 6701 4058 6731 4092
rect 6493 4020 6731 4058
rect 6493 3986 6523 4020
rect 6557 3986 6667 4020
rect 6701 3986 6731 4020
rect 6493 3948 6731 3986
rect 6493 3914 6523 3948
rect 6557 3914 6667 3948
rect 6701 3914 6731 3948
rect 6493 3876 6731 3914
rect 6493 3842 6523 3876
rect 6557 3842 6667 3876
rect 6701 3842 6731 3876
rect 6493 3804 6731 3842
rect 6493 3770 6523 3804
rect 6557 3770 6667 3804
rect 6701 3770 6731 3804
rect 6493 3732 6731 3770
rect 6493 3698 6523 3732
rect 6557 3698 6667 3732
rect 6701 3698 6731 3732
rect 6493 3660 6731 3698
rect 6493 3626 6523 3660
rect 6557 3626 6667 3660
rect 6701 3626 6731 3660
rect 6493 3588 6731 3626
rect 6493 3554 6523 3588
rect 6557 3554 6667 3588
rect 6701 3554 6731 3588
rect 6493 3516 6731 3554
rect 6493 3482 6523 3516
rect 6557 3482 6667 3516
rect 6701 3482 6731 3516
rect 6493 3444 6731 3482
rect 6493 3410 6523 3444
rect 6557 3410 6667 3444
rect 6701 3410 6731 3444
rect 6493 3372 6731 3410
rect 6493 3338 6523 3372
rect 6557 3338 6667 3372
rect 6701 3338 6731 3372
rect 6493 3300 6731 3338
rect 6493 3266 6523 3300
rect 6557 3266 6667 3300
rect 6701 3266 6731 3300
rect 6493 3228 6731 3266
rect 6493 3194 6523 3228
rect 6557 3194 6667 3228
rect 6701 3194 6731 3228
rect 6493 3108 6731 3194
rect 6493 3074 6523 3108
rect 6557 3074 6595 3108
rect 6629 3074 6667 3108
rect 6701 3074 6731 3108
rect 6493 3044 6731 3074
rect 6493 3028 6561 3044
rect 6493 2994 6523 3028
rect 6557 3010 6561 3028
rect 6595 3028 6629 3044
rect 6557 2994 6595 3010
rect 6663 3028 6731 3044
rect 6663 3010 6667 3028
rect 6629 2994 6667 3010
rect 6701 2994 6731 3028
rect 6493 2974 6731 2994
rect 6493 2948 6561 2974
rect 6493 2914 6523 2948
rect 6557 2940 6561 2948
rect 6595 2948 6629 2974
rect 6557 2914 6595 2940
rect 6663 2948 6731 2974
rect 6663 2940 6667 2948
rect 6629 2914 6667 2940
rect 6701 2914 6731 2948
rect 6493 2904 6731 2914
rect 6493 2870 6561 2904
rect 6595 2870 6629 2904
rect 6663 2870 6731 2904
rect 6493 2868 6731 2870
rect 6493 2834 6523 2868
rect 6557 2834 6595 2868
rect 6629 2834 6667 2868
rect 6701 2834 6731 2868
rect 6493 2800 6561 2834
rect 6595 2800 6629 2834
rect 6663 2800 6731 2834
rect 6493 2788 6731 2800
rect 6493 2754 6523 2788
rect 6557 2764 6595 2788
rect 6557 2754 6561 2764
rect 6493 2730 6561 2754
rect 6629 2764 6667 2788
rect 6595 2730 6629 2754
rect 6663 2754 6667 2764
rect 6701 2754 6731 2788
rect 6663 2730 6731 2754
rect 6493 2708 6731 2730
rect 6493 2674 6523 2708
rect 6557 2694 6595 2708
rect 6557 2674 6561 2694
rect 6493 2660 6561 2674
rect 6629 2694 6667 2708
rect 6595 2660 6629 2674
rect 6663 2674 6667 2694
rect 6701 2674 6731 2708
rect 6663 2660 6731 2674
rect 6493 2628 6731 2660
rect 6493 2594 6523 2628
rect 6557 2594 6595 2628
rect 6629 2594 6667 2628
rect 6701 2594 6731 2628
rect 6493 2518 6731 2594
rect 6493 2484 6523 2518
rect 6557 2484 6667 2518
rect 6701 2484 6731 2518
rect 6493 2446 6731 2484
rect 6493 2412 6523 2446
rect 6557 2412 6667 2446
rect 6701 2412 6731 2446
rect 6493 2374 6731 2412
rect 6493 2340 6523 2374
rect 6557 2340 6667 2374
rect 6701 2340 6731 2374
rect 6493 2302 6731 2340
rect 6493 2268 6523 2302
rect 6557 2268 6667 2302
rect 6701 2268 6731 2302
rect 6493 2230 6731 2268
rect 6493 2196 6523 2230
rect 6557 2196 6667 2230
rect 6701 2196 6731 2230
rect 6493 2158 6731 2196
rect 6493 2124 6523 2158
rect 6557 2124 6667 2158
rect 6701 2124 6731 2158
rect 6493 2086 6731 2124
rect 6493 2052 6523 2086
rect 6557 2052 6667 2086
rect 6701 2052 6731 2086
rect 6493 2014 6731 2052
rect 6493 1980 6523 2014
rect 6557 1980 6667 2014
rect 6701 1980 6731 2014
rect 6493 1942 6731 1980
rect 6493 1908 6523 1942
rect 6557 1908 6667 1942
rect 6701 1908 6731 1942
rect 6493 1870 6731 1908
rect 6493 1836 6523 1870
rect 6557 1836 6667 1870
rect 6701 1836 6731 1870
rect 6493 1798 6731 1836
rect 6493 1764 6523 1798
rect 6557 1764 6667 1798
rect 6701 1764 6731 1798
rect 6493 1726 6731 1764
rect 6493 1692 6523 1726
rect 6557 1692 6667 1726
rect 6701 1692 6731 1726
rect 6493 1654 6731 1692
rect 6493 1620 6523 1654
rect 6557 1620 6667 1654
rect 6701 1620 6731 1654
rect 6493 1536 6731 1620
rect 6833 3104 6953 4200
rect 7263 4308 7383 4324
rect 7263 4274 7306 4308
rect 7340 4274 7383 4308
rect 7263 4234 7383 4274
rect 7263 4200 7306 4234
rect 7340 4200 7383 4234
rect 6833 3070 6876 3104
rect 6910 3070 6953 3104
rect 6833 3026 6953 3070
rect 6833 2992 6876 3026
rect 6910 2992 6953 3026
rect 6833 2948 6953 2992
rect 6833 2914 6876 2948
rect 6910 2914 6953 2948
rect 6833 2870 6953 2914
rect 6833 2836 6876 2870
rect 6910 2836 6953 2870
rect 6833 2792 6953 2836
rect 6833 2758 6876 2792
rect 6910 2758 6953 2792
rect 6833 2713 6953 2758
rect 6833 2679 6876 2713
rect 6910 2679 6953 2713
rect 6833 2634 6953 2679
rect 6833 2600 6876 2634
rect 6910 2600 6953 2634
rect 6271 1470 6314 1504
rect 6348 1470 6391 1504
rect 6271 1430 6391 1470
rect 6271 1396 6314 1430
rect 6348 1396 6391 1430
rect 6271 1250 6391 1396
rect 6271 1144 6278 1250
rect 6384 1144 6391 1250
rect 6833 1504 6953 2600
rect 7018 4064 7019 4098
rect 7053 4064 7091 4098
rect 7125 4064 7163 4098
rect 7197 4064 7198 4098
rect 7018 4025 7198 4064
rect 7018 3991 7019 4025
rect 7053 3991 7091 4025
rect 7125 3991 7163 4025
rect 7197 3991 7198 4025
rect 7018 3952 7198 3991
rect 7018 3918 7019 3952
rect 7053 3918 7091 3952
rect 7125 3918 7163 3952
rect 7197 3918 7198 3952
rect 7018 3879 7198 3918
rect 7018 3845 7019 3879
rect 7053 3845 7091 3879
rect 7125 3845 7163 3879
rect 7197 3845 7198 3879
rect 7018 3806 7198 3845
rect 7018 3772 7019 3806
rect 7053 3772 7091 3806
rect 7125 3772 7163 3806
rect 7197 3772 7198 3806
rect 7018 3733 7198 3772
rect 7018 3699 7019 3733
rect 7053 3699 7091 3733
rect 7125 3699 7163 3733
rect 7197 3699 7198 3733
rect 7018 3660 7198 3699
rect 7018 3626 7019 3660
rect 7053 3626 7091 3660
rect 7125 3626 7163 3660
rect 7197 3626 7198 3660
rect 7018 3587 7198 3626
rect 7018 3553 7019 3587
rect 7053 3553 7091 3587
rect 7125 3553 7163 3587
rect 7197 3553 7198 3587
rect 7018 3514 7198 3553
rect 7018 3480 7019 3514
rect 7053 3480 7091 3514
rect 7125 3480 7163 3514
rect 7197 3480 7198 3514
rect 7018 3441 7198 3480
rect 7018 3407 7019 3441
rect 7053 3407 7091 3441
rect 7125 3407 7163 3441
rect 7197 3407 7198 3441
rect 7018 3368 7198 3407
rect 7018 3334 7019 3368
rect 7053 3334 7091 3368
rect 7125 3334 7163 3368
rect 7197 3334 7198 3368
rect 7018 3295 7198 3334
rect 7018 3261 7019 3295
rect 7053 3261 7091 3295
rect 7125 3261 7163 3295
rect 7197 3261 7198 3295
rect 7018 3222 7198 3261
rect 7018 3188 7019 3222
rect 7053 3188 7091 3222
rect 7125 3188 7163 3222
rect 7197 3188 7198 3222
rect 7018 3149 7198 3188
rect 7018 3115 7019 3149
rect 7053 3115 7091 3149
rect 7125 3115 7163 3149
rect 7197 3115 7198 3149
rect 7018 3076 7198 3115
rect 7018 3042 7019 3076
rect 7053 3042 7091 3076
rect 7125 3042 7163 3076
rect 7197 3042 7198 3076
rect 7018 3003 7198 3042
rect 7018 2969 7019 3003
rect 7053 2969 7091 3003
rect 7125 2969 7163 3003
rect 7197 2969 7198 3003
rect 7018 2930 7198 2969
rect 7018 2896 7019 2930
rect 7053 2896 7091 2930
rect 7125 2896 7163 2930
rect 7197 2896 7198 2930
rect 7018 2857 7198 2896
rect 7018 2823 7019 2857
rect 7053 2823 7091 2857
rect 7125 2823 7163 2857
rect 7197 2823 7198 2857
rect 7018 2784 7198 2823
rect 7018 2750 7019 2784
rect 7053 2750 7091 2784
rect 7125 2750 7163 2784
rect 7197 2750 7198 2784
rect 7018 2711 7198 2750
rect 7018 2677 7019 2711
rect 7053 2677 7091 2711
rect 7125 2677 7163 2711
rect 7197 2677 7198 2711
rect 7018 2638 7198 2677
rect 7018 2604 7019 2638
rect 7053 2604 7091 2638
rect 7125 2604 7163 2638
rect 7197 2604 7198 2638
rect 7018 2565 7198 2604
rect 7018 2531 7019 2565
rect 7053 2531 7091 2565
rect 7125 2531 7163 2565
rect 7197 2531 7198 2565
rect 7018 2492 7198 2531
rect 7018 2458 7019 2492
rect 7053 2458 7091 2492
rect 7125 2458 7163 2492
rect 7197 2458 7198 2492
rect 7018 2419 7198 2458
rect 7018 2385 7019 2419
rect 7053 2385 7091 2419
rect 7125 2385 7163 2419
rect 7197 2385 7198 2419
rect 7018 2346 7198 2385
rect 7018 2312 7019 2346
rect 7053 2312 7091 2346
rect 7125 2312 7163 2346
rect 7197 2312 7198 2346
rect 7018 2273 7198 2312
rect 7018 2239 7019 2273
rect 7053 2239 7091 2273
rect 7125 2239 7163 2273
rect 7197 2239 7198 2273
rect 7018 2200 7198 2239
rect 7018 2166 7019 2200
rect 7053 2166 7091 2200
rect 7125 2166 7163 2200
rect 7197 2166 7198 2200
rect 7018 2126 7198 2166
rect 7018 2092 7019 2126
rect 7053 2092 7091 2126
rect 7125 2092 7163 2126
rect 7197 2092 7198 2126
rect 7018 2052 7198 2092
rect 7018 2018 7019 2052
rect 7053 2018 7091 2052
rect 7125 2018 7163 2052
rect 7197 2018 7198 2052
rect 7018 1978 7198 2018
rect 7018 1944 7019 1978
rect 7053 1944 7091 1978
rect 7125 1944 7163 1978
rect 7197 1944 7198 1978
rect 7018 1904 7198 1944
rect 7018 1870 7019 1904
rect 7053 1870 7091 1904
rect 7125 1870 7163 1904
rect 7197 1870 7198 1904
rect 7018 1830 7198 1870
rect 7018 1796 7019 1830
rect 7053 1796 7091 1830
rect 7125 1796 7163 1830
rect 7197 1796 7198 1830
rect 7018 1756 7198 1796
rect 7018 1722 7019 1756
rect 7053 1722 7091 1756
rect 7125 1722 7163 1756
rect 7197 1722 7198 1756
rect 7018 1682 7198 1722
rect 7018 1648 7019 1682
rect 7053 1648 7091 1682
rect 7125 1648 7163 1682
rect 7197 1648 7198 1682
rect 7018 1608 7198 1648
rect 7018 1574 7019 1608
rect 7053 1574 7091 1608
rect 7125 1574 7163 1608
rect 7197 1574 7198 1608
rect 7018 1548 7198 1574
rect 7263 3104 7383 4200
rect 7825 4308 7945 4324
rect 7825 4274 7868 4308
rect 7902 4274 7945 4308
rect 7825 4234 7945 4274
rect 7825 4200 7868 4234
rect 7902 4200 7945 4234
rect 7263 3070 7306 3104
rect 7340 3070 7383 3104
rect 7263 3026 7383 3070
rect 7263 2992 7306 3026
rect 7340 2992 7383 3026
rect 7263 2948 7383 2992
rect 7263 2914 7306 2948
rect 7340 2914 7383 2948
rect 7263 2870 7383 2914
rect 7263 2836 7306 2870
rect 7340 2836 7383 2870
rect 7263 2792 7383 2836
rect 7263 2758 7306 2792
rect 7340 2758 7383 2792
rect 7263 2713 7383 2758
rect 7263 2679 7306 2713
rect 7340 2679 7383 2713
rect 7263 2634 7383 2679
rect 7263 2600 7306 2634
rect 7340 2600 7383 2634
rect 6833 1470 6876 1504
rect 6910 1470 6953 1504
rect 6833 1430 6953 1470
rect 6833 1396 6876 1430
rect 6910 1396 6953 1430
rect 6833 1250 6953 1396
rect 6833 1144 6840 1250
rect 6946 1144 6953 1250
rect 7263 1504 7383 2600
rect 7485 4092 7723 4104
rect 7485 4058 7515 4092
rect 7549 4058 7659 4092
rect 7693 4058 7723 4092
rect 7485 4020 7723 4058
rect 7485 3986 7515 4020
rect 7549 3986 7659 4020
rect 7693 3986 7723 4020
rect 7485 3948 7723 3986
rect 7485 3914 7515 3948
rect 7549 3914 7659 3948
rect 7693 3914 7723 3948
rect 7485 3876 7723 3914
rect 7485 3842 7515 3876
rect 7549 3842 7659 3876
rect 7693 3842 7723 3876
rect 7485 3804 7723 3842
rect 7485 3770 7515 3804
rect 7549 3770 7659 3804
rect 7693 3770 7723 3804
rect 7485 3732 7723 3770
rect 7485 3698 7515 3732
rect 7549 3698 7659 3732
rect 7693 3698 7723 3732
rect 7485 3660 7723 3698
rect 7485 3626 7515 3660
rect 7549 3626 7659 3660
rect 7693 3626 7723 3660
rect 7485 3588 7723 3626
rect 7485 3554 7515 3588
rect 7549 3554 7659 3588
rect 7693 3554 7723 3588
rect 7485 3516 7723 3554
rect 7485 3482 7515 3516
rect 7549 3482 7659 3516
rect 7693 3482 7723 3516
rect 7485 3444 7723 3482
rect 7485 3410 7515 3444
rect 7549 3410 7659 3444
rect 7693 3410 7723 3444
rect 7485 3372 7723 3410
rect 7485 3338 7515 3372
rect 7549 3338 7659 3372
rect 7693 3338 7723 3372
rect 7485 3300 7723 3338
rect 7485 3266 7515 3300
rect 7549 3266 7659 3300
rect 7693 3266 7723 3300
rect 7485 3228 7723 3266
rect 7485 3194 7515 3228
rect 7549 3194 7659 3228
rect 7693 3194 7723 3228
rect 7485 3108 7723 3194
rect 7485 3074 7515 3108
rect 7549 3074 7587 3108
rect 7621 3074 7659 3108
rect 7693 3074 7723 3108
rect 7485 3044 7723 3074
rect 7485 3028 7553 3044
rect 7485 2994 7515 3028
rect 7549 3010 7553 3028
rect 7587 3028 7621 3044
rect 7549 2994 7587 3010
rect 7655 3028 7723 3044
rect 7655 3010 7659 3028
rect 7621 2994 7659 3010
rect 7693 2994 7723 3028
rect 7485 2974 7723 2994
rect 7485 2948 7553 2974
rect 7485 2914 7515 2948
rect 7549 2940 7553 2948
rect 7587 2948 7621 2974
rect 7549 2914 7587 2940
rect 7655 2948 7723 2974
rect 7655 2940 7659 2948
rect 7621 2914 7659 2940
rect 7693 2914 7723 2948
rect 7485 2904 7723 2914
rect 7485 2870 7553 2904
rect 7587 2870 7621 2904
rect 7655 2870 7723 2904
rect 7485 2868 7723 2870
rect 7485 2834 7515 2868
rect 7549 2834 7587 2868
rect 7621 2834 7659 2868
rect 7693 2834 7723 2868
rect 7485 2800 7553 2834
rect 7587 2800 7621 2834
rect 7655 2800 7723 2834
rect 7485 2788 7723 2800
rect 7485 2754 7515 2788
rect 7549 2764 7587 2788
rect 7549 2754 7553 2764
rect 7485 2730 7553 2754
rect 7621 2764 7659 2788
rect 7587 2730 7621 2754
rect 7655 2754 7659 2764
rect 7693 2754 7723 2788
rect 7655 2730 7723 2754
rect 7485 2708 7723 2730
rect 7485 2674 7515 2708
rect 7549 2694 7587 2708
rect 7549 2674 7553 2694
rect 7485 2660 7553 2674
rect 7621 2694 7659 2708
rect 7587 2660 7621 2674
rect 7655 2674 7659 2694
rect 7693 2674 7723 2708
rect 7655 2660 7723 2674
rect 7485 2628 7723 2660
rect 7485 2594 7515 2628
rect 7549 2594 7587 2628
rect 7621 2594 7659 2628
rect 7693 2594 7723 2628
rect 7485 2518 7723 2594
rect 7485 2484 7515 2518
rect 7549 2484 7659 2518
rect 7693 2484 7723 2518
rect 7485 2446 7723 2484
rect 7485 2412 7515 2446
rect 7549 2412 7659 2446
rect 7693 2412 7723 2446
rect 7485 2374 7723 2412
rect 7485 2340 7515 2374
rect 7549 2340 7659 2374
rect 7693 2340 7723 2374
rect 7485 2302 7723 2340
rect 7485 2268 7515 2302
rect 7549 2268 7659 2302
rect 7693 2268 7723 2302
rect 7485 2230 7723 2268
rect 7485 2196 7515 2230
rect 7549 2196 7659 2230
rect 7693 2196 7723 2230
rect 7485 2158 7723 2196
rect 7485 2124 7515 2158
rect 7549 2124 7659 2158
rect 7693 2124 7723 2158
rect 7485 2086 7723 2124
rect 7485 2052 7515 2086
rect 7549 2052 7659 2086
rect 7693 2052 7723 2086
rect 7485 2014 7723 2052
rect 7485 1980 7515 2014
rect 7549 1980 7659 2014
rect 7693 1980 7723 2014
rect 7485 1942 7723 1980
rect 7485 1908 7515 1942
rect 7549 1908 7659 1942
rect 7693 1908 7723 1942
rect 7485 1870 7723 1908
rect 7485 1836 7515 1870
rect 7549 1836 7659 1870
rect 7693 1836 7723 1870
rect 7485 1798 7723 1836
rect 7485 1764 7515 1798
rect 7549 1764 7659 1798
rect 7693 1764 7723 1798
rect 7485 1726 7723 1764
rect 7485 1692 7515 1726
rect 7549 1692 7659 1726
rect 7693 1692 7723 1726
rect 7485 1654 7723 1692
rect 7485 1620 7515 1654
rect 7549 1620 7659 1654
rect 7693 1620 7723 1654
rect 7485 1536 7723 1620
rect 7825 3104 7945 4200
rect 8255 4308 8375 4324
rect 8255 4274 8298 4308
rect 8332 4274 8375 4308
rect 8255 4234 8375 4274
rect 8255 4200 8298 4234
rect 8332 4200 8375 4234
rect 7825 3070 7868 3104
rect 7902 3070 7945 3104
rect 7825 3026 7945 3070
rect 7825 2992 7868 3026
rect 7902 2992 7945 3026
rect 7825 2948 7945 2992
rect 7825 2914 7868 2948
rect 7902 2914 7945 2948
rect 7825 2870 7945 2914
rect 7825 2836 7868 2870
rect 7902 2836 7945 2870
rect 7825 2792 7945 2836
rect 7825 2758 7868 2792
rect 7902 2758 7945 2792
rect 7825 2713 7945 2758
rect 7825 2679 7868 2713
rect 7902 2679 7945 2713
rect 7825 2634 7945 2679
rect 7825 2600 7868 2634
rect 7902 2600 7945 2634
rect 7263 1470 7306 1504
rect 7340 1470 7383 1504
rect 7263 1430 7383 1470
rect 7263 1396 7306 1430
rect 7340 1396 7383 1430
rect 7263 1250 7383 1396
rect 7263 1144 7270 1250
rect 7376 1144 7383 1250
rect 7825 1504 7945 2600
rect 8010 4064 8011 4098
rect 8045 4064 8083 4098
rect 8117 4064 8155 4098
rect 8189 4064 8190 4098
rect 8010 4025 8190 4064
rect 8010 3991 8011 4025
rect 8045 3991 8083 4025
rect 8117 3991 8155 4025
rect 8189 3991 8190 4025
rect 8010 3952 8190 3991
rect 8010 3918 8011 3952
rect 8045 3918 8083 3952
rect 8117 3918 8155 3952
rect 8189 3918 8190 3952
rect 8010 3879 8190 3918
rect 8010 3845 8011 3879
rect 8045 3845 8083 3879
rect 8117 3845 8155 3879
rect 8189 3845 8190 3879
rect 8010 3806 8190 3845
rect 8010 3772 8011 3806
rect 8045 3772 8083 3806
rect 8117 3772 8155 3806
rect 8189 3772 8190 3806
rect 8010 3733 8190 3772
rect 8010 3699 8011 3733
rect 8045 3699 8083 3733
rect 8117 3699 8155 3733
rect 8189 3699 8190 3733
rect 8010 3660 8190 3699
rect 8010 3626 8011 3660
rect 8045 3626 8083 3660
rect 8117 3626 8155 3660
rect 8189 3626 8190 3660
rect 8010 3587 8190 3626
rect 8010 3553 8011 3587
rect 8045 3553 8083 3587
rect 8117 3553 8155 3587
rect 8189 3553 8190 3587
rect 8010 3514 8190 3553
rect 8010 3480 8011 3514
rect 8045 3480 8083 3514
rect 8117 3480 8155 3514
rect 8189 3480 8190 3514
rect 8010 3441 8190 3480
rect 8010 3407 8011 3441
rect 8045 3407 8083 3441
rect 8117 3407 8155 3441
rect 8189 3407 8190 3441
rect 8010 3368 8190 3407
rect 8010 3334 8011 3368
rect 8045 3334 8083 3368
rect 8117 3334 8155 3368
rect 8189 3334 8190 3368
rect 8010 3295 8190 3334
rect 8010 3261 8011 3295
rect 8045 3261 8083 3295
rect 8117 3261 8155 3295
rect 8189 3261 8190 3295
rect 8010 3222 8190 3261
rect 8010 3188 8011 3222
rect 8045 3188 8083 3222
rect 8117 3188 8155 3222
rect 8189 3188 8190 3222
rect 8010 3149 8190 3188
rect 8010 3115 8011 3149
rect 8045 3115 8083 3149
rect 8117 3115 8155 3149
rect 8189 3115 8190 3149
rect 8010 3076 8190 3115
rect 8010 3042 8011 3076
rect 8045 3042 8083 3076
rect 8117 3042 8155 3076
rect 8189 3042 8190 3076
rect 8010 3003 8190 3042
rect 8010 2969 8011 3003
rect 8045 2969 8083 3003
rect 8117 2969 8155 3003
rect 8189 2969 8190 3003
rect 8010 2930 8190 2969
rect 8010 2896 8011 2930
rect 8045 2896 8083 2930
rect 8117 2896 8155 2930
rect 8189 2896 8190 2930
rect 8010 2857 8190 2896
rect 8010 2823 8011 2857
rect 8045 2823 8083 2857
rect 8117 2823 8155 2857
rect 8189 2823 8190 2857
rect 8010 2784 8190 2823
rect 8010 2750 8011 2784
rect 8045 2750 8083 2784
rect 8117 2750 8155 2784
rect 8189 2750 8190 2784
rect 8010 2711 8190 2750
rect 8010 2677 8011 2711
rect 8045 2677 8083 2711
rect 8117 2677 8155 2711
rect 8189 2677 8190 2711
rect 8010 2638 8190 2677
rect 8010 2604 8011 2638
rect 8045 2604 8083 2638
rect 8117 2604 8155 2638
rect 8189 2604 8190 2638
rect 8010 2565 8190 2604
rect 8010 2531 8011 2565
rect 8045 2531 8083 2565
rect 8117 2531 8155 2565
rect 8189 2531 8190 2565
rect 8010 2492 8190 2531
rect 8010 2458 8011 2492
rect 8045 2458 8083 2492
rect 8117 2458 8155 2492
rect 8189 2458 8190 2492
rect 8010 2419 8190 2458
rect 8010 2385 8011 2419
rect 8045 2385 8083 2419
rect 8117 2385 8155 2419
rect 8189 2385 8190 2419
rect 8010 2346 8190 2385
rect 8010 2312 8011 2346
rect 8045 2312 8083 2346
rect 8117 2312 8155 2346
rect 8189 2312 8190 2346
rect 8010 2273 8190 2312
rect 8010 2239 8011 2273
rect 8045 2239 8083 2273
rect 8117 2239 8155 2273
rect 8189 2239 8190 2273
rect 8010 2200 8190 2239
rect 8010 2166 8011 2200
rect 8045 2166 8083 2200
rect 8117 2166 8155 2200
rect 8189 2166 8190 2200
rect 8010 2126 8190 2166
rect 8010 2092 8011 2126
rect 8045 2092 8083 2126
rect 8117 2092 8155 2126
rect 8189 2092 8190 2126
rect 8010 2052 8190 2092
rect 8010 2018 8011 2052
rect 8045 2018 8083 2052
rect 8117 2018 8155 2052
rect 8189 2018 8190 2052
rect 8010 1978 8190 2018
rect 8010 1944 8011 1978
rect 8045 1944 8083 1978
rect 8117 1944 8155 1978
rect 8189 1944 8190 1978
rect 8010 1904 8190 1944
rect 8010 1870 8011 1904
rect 8045 1870 8083 1904
rect 8117 1870 8155 1904
rect 8189 1870 8190 1904
rect 8010 1830 8190 1870
rect 8010 1796 8011 1830
rect 8045 1796 8083 1830
rect 8117 1796 8155 1830
rect 8189 1796 8190 1830
rect 8010 1756 8190 1796
rect 8010 1722 8011 1756
rect 8045 1722 8083 1756
rect 8117 1722 8155 1756
rect 8189 1722 8190 1756
rect 8010 1682 8190 1722
rect 8010 1648 8011 1682
rect 8045 1648 8083 1682
rect 8117 1648 8155 1682
rect 8189 1648 8190 1682
rect 8010 1608 8190 1648
rect 8010 1574 8011 1608
rect 8045 1574 8083 1608
rect 8117 1574 8155 1608
rect 8189 1574 8190 1608
rect 8010 1548 8190 1574
rect 8255 3104 8375 4200
rect 8817 4308 8937 4324
rect 8817 4274 8860 4308
rect 8894 4274 8937 4308
rect 8817 4234 8937 4274
rect 8817 4200 8860 4234
rect 8894 4200 8937 4234
rect 8255 3070 8298 3104
rect 8332 3070 8375 3104
rect 8255 3026 8375 3070
rect 8255 2992 8298 3026
rect 8332 2992 8375 3026
rect 8255 2948 8375 2992
rect 8255 2914 8298 2948
rect 8332 2914 8375 2948
rect 8255 2870 8375 2914
rect 8255 2836 8298 2870
rect 8332 2836 8375 2870
rect 8255 2792 8375 2836
rect 8255 2758 8298 2792
rect 8332 2758 8375 2792
rect 8255 2713 8375 2758
rect 8255 2679 8298 2713
rect 8332 2679 8375 2713
rect 8255 2634 8375 2679
rect 8255 2600 8298 2634
rect 8332 2600 8375 2634
rect 7825 1470 7868 1504
rect 7902 1470 7945 1504
rect 7825 1430 7945 1470
rect 7825 1396 7868 1430
rect 7902 1396 7945 1430
rect 7825 1250 7945 1396
rect 7825 1144 7832 1250
rect 7938 1144 7945 1250
rect 8255 1504 8375 2600
rect 8477 4092 8715 4104
rect 8477 4058 8507 4092
rect 8541 4058 8651 4092
rect 8685 4058 8715 4092
rect 8477 4020 8715 4058
rect 8477 3986 8507 4020
rect 8541 3986 8651 4020
rect 8685 3986 8715 4020
rect 8477 3948 8715 3986
rect 8477 3914 8507 3948
rect 8541 3914 8651 3948
rect 8685 3914 8715 3948
rect 8477 3876 8715 3914
rect 8477 3842 8507 3876
rect 8541 3842 8651 3876
rect 8685 3842 8715 3876
rect 8477 3804 8715 3842
rect 8477 3770 8507 3804
rect 8541 3770 8651 3804
rect 8685 3770 8715 3804
rect 8477 3732 8715 3770
rect 8477 3698 8507 3732
rect 8541 3698 8651 3732
rect 8685 3698 8715 3732
rect 8477 3660 8715 3698
rect 8477 3626 8507 3660
rect 8541 3626 8651 3660
rect 8685 3626 8715 3660
rect 8477 3588 8715 3626
rect 8477 3554 8507 3588
rect 8541 3554 8651 3588
rect 8685 3554 8715 3588
rect 8477 3516 8715 3554
rect 8477 3482 8507 3516
rect 8541 3482 8651 3516
rect 8685 3482 8715 3516
rect 8477 3444 8715 3482
rect 8477 3410 8507 3444
rect 8541 3410 8651 3444
rect 8685 3410 8715 3444
rect 8477 3372 8715 3410
rect 8477 3338 8507 3372
rect 8541 3338 8651 3372
rect 8685 3338 8715 3372
rect 8477 3300 8715 3338
rect 8477 3266 8507 3300
rect 8541 3266 8651 3300
rect 8685 3266 8715 3300
rect 8477 3228 8715 3266
rect 8477 3194 8507 3228
rect 8541 3194 8651 3228
rect 8685 3194 8715 3228
rect 8477 3108 8715 3194
rect 8477 3074 8507 3108
rect 8541 3074 8579 3108
rect 8613 3074 8651 3108
rect 8685 3074 8715 3108
rect 8477 3044 8715 3074
rect 8477 3028 8545 3044
rect 8477 2994 8507 3028
rect 8541 3010 8545 3028
rect 8579 3028 8613 3044
rect 8541 2994 8579 3010
rect 8647 3028 8715 3044
rect 8647 3010 8651 3028
rect 8613 2994 8651 3010
rect 8685 2994 8715 3028
rect 8477 2974 8715 2994
rect 8477 2948 8545 2974
rect 8477 2914 8507 2948
rect 8541 2940 8545 2948
rect 8579 2948 8613 2974
rect 8541 2914 8579 2940
rect 8647 2948 8715 2974
rect 8647 2940 8651 2948
rect 8613 2914 8651 2940
rect 8685 2914 8715 2948
rect 8477 2904 8715 2914
rect 8477 2870 8545 2904
rect 8579 2870 8613 2904
rect 8647 2870 8715 2904
rect 8477 2868 8715 2870
rect 8477 2834 8507 2868
rect 8541 2834 8579 2868
rect 8613 2834 8651 2868
rect 8685 2834 8715 2868
rect 8477 2800 8545 2834
rect 8579 2800 8613 2834
rect 8647 2800 8715 2834
rect 8477 2788 8715 2800
rect 8477 2754 8507 2788
rect 8541 2764 8579 2788
rect 8541 2754 8545 2764
rect 8477 2730 8545 2754
rect 8613 2764 8651 2788
rect 8579 2730 8613 2754
rect 8647 2754 8651 2764
rect 8685 2754 8715 2788
rect 8647 2730 8715 2754
rect 8477 2708 8715 2730
rect 8477 2674 8507 2708
rect 8541 2694 8579 2708
rect 8541 2674 8545 2694
rect 8477 2660 8545 2674
rect 8613 2694 8651 2708
rect 8579 2660 8613 2674
rect 8647 2674 8651 2694
rect 8685 2674 8715 2708
rect 8647 2660 8715 2674
rect 8477 2628 8715 2660
rect 8477 2594 8507 2628
rect 8541 2594 8579 2628
rect 8613 2594 8651 2628
rect 8685 2594 8715 2628
rect 8477 2518 8715 2594
rect 8477 2484 8507 2518
rect 8541 2484 8651 2518
rect 8685 2484 8715 2518
rect 8477 2446 8715 2484
rect 8477 2412 8507 2446
rect 8541 2412 8651 2446
rect 8685 2412 8715 2446
rect 8477 2374 8715 2412
rect 8477 2340 8507 2374
rect 8541 2340 8651 2374
rect 8685 2340 8715 2374
rect 8477 2302 8715 2340
rect 8477 2268 8507 2302
rect 8541 2268 8651 2302
rect 8685 2268 8715 2302
rect 8477 2230 8715 2268
rect 8477 2196 8507 2230
rect 8541 2196 8651 2230
rect 8685 2196 8715 2230
rect 8477 2158 8715 2196
rect 8477 2124 8507 2158
rect 8541 2124 8651 2158
rect 8685 2124 8715 2158
rect 8477 2086 8715 2124
rect 8477 2052 8507 2086
rect 8541 2052 8651 2086
rect 8685 2052 8715 2086
rect 8477 2014 8715 2052
rect 8477 1980 8507 2014
rect 8541 1980 8651 2014
rect 8685 1980 8715 2014
rect 8477 1942 8715 1980
rect 8477 1908 8507 1942
rect 8541 1908 8651 1942
rect 8685 1908 8715 1942
rect 8477 1870 8715 1908
rect 8477 1836 8507 1870
rect 8541 1836 8651 1870
rect 8685 1836 8715 1870
rect 8477 1798 8715 1836
rect 8477 1764 8507 1798
rect 8541 1764 8651 1798
rect 8685 1764 8715 1798
rect 8477 1726 8715 1764
rect 8477 1692 8507 1726
rect 8541 1692 8651 1726
rect 8685 1692 8715 1726
rect 8477 1654 8715 1692
rect 8477 1620 8507 1654
rect 8541 1620 8651 1654
rect 8685 1620 8715 1654
rect 8477 1536 8715 1620
rect 8817 3104 8937 4200
rect 9247 4308 9367 4324
rect 9247 4274 9290 4308
rect 9324 4274 9367 4308
rect 9247 4234 9367 4274
rect 9247 4200 9290 4234
rect 9324 4200 9367 4234
rect 8817 3070 8860 3104
rect 8894 3070 8937 3104
rect 8817 3026 8937 3070
rect 8817 2992 8860 3026
rect 8894 2992 8937 3026
rect 8817 2948 8937 2992
rect 8817 2914 8860 2948
rect 8894 2914 8937 2948
rect 8817 2870 8937 2914
rect 8817 2836 8860 2870
rect 8894 2836 8937 2870
rect 8817 2792 8937 2836
rect 8817 2758 8860 2792
rect 8894 2758 8937 2792
rect 8817 2713 8937 2758
rect 8817 2679 8860 2713
rect 8894 2679 8937 2713
rect 8817 2634 8937 2679
rect 8817 2600 8860 2634
rect 8894 2600 8937 2634
rect 8255 1470 8298 1504
rect 8332 1470 8375 1504
rect 8255 1430 8375 1470
rect 8255 1396 8298 1430
rect 8332 1396 8375 1430
rect 8255 1250 8375 1396
rect 8255 1144 8262 1250
rect 8368 1144 8375 1250
rect 8817 1504 8937 2600
rect 9002 4098 9182 4099
rect 9002 4064 9003 4098
rect 9037 4064 9075 4098
rect 9109 4064 9147 4098
rect 9181 4064 9182 4098
rect 9002 4025 9182 4064
rect 9002 3991 9003 4025
rect 9037 3991 9075 4025
rect 9109 3991 9147 4025
rect 9181 3991 9182 4025
rect 9002 3952 9182 3991
rect 9002 3918 9003 3952
rect 9037 3918 9075 3952
rect 9109 3918 9147 3952
rect 9181 3918 9182 3952
rect 9002 3879 9182 3918
rect 9002 3845 9003 3879
rect 9037 3845 9075 3879
rect 9109 3845 9147 3879
rect 9181 3845 9182 3879
rect 9002 3806 9182 3845
rect 9002 3772 9003 3806
rect 9037 3772 9075 3806
rect 9109 3772 9147 3806
rect 9181 3772 9182 3806
rect 9002 3733 9182 3772
rect 9002 3699 9003 3733
rect 9037 3699 9075 3733
rect 9109 3699 9147 3733
rect 9181 3699 9182 3733
rect 9002 3660 9182 3699
rect 9002 3626 9003 3660
rect 9037 3626 9075 3660
rect 9109 3626 9147 3660
rect 9181 3626 9182 3660
rect 9002 3587 9182 3626
rect 9002 3553 9003 3587
rect 9037 3553 9075 3587
rect 9109 3553 9147 3587
rect 9181 3553 9182 3587
rect 9002 3514 9182 3553
rect 9002 3480 9003 3514
rect 9037 3480 9075 3514
rect 9109 3480 9147 3514
rect 9181 3480 9182 3514
rect 9002 3441 9182 3480
rect 9002 3407 9003 3441
rect 9037 3407 9075 3441
rect 9109 3407 9147 3441
rect 9181 3407 9182 3441
rect 9002 3368 9182 3407
rect 9002 3334 9003 3368
rect 9037 3334 9075 3368
rect 9109 3334 9147 3368
rect 9181 3334 9182 3368
rect 9002 3295 9182 3334
rect 9002 3261 9003 3295
rect 9037 3261 9075 3295
rect 9109 3261 9147 3295
rect 9181 3261 9182 3295
rect 9002 3222 9182 3261
rect 9002 3188 9003 3222
rect 9037 3188 9075 3222
rect 9109 3188 9147 3222
rect 9181 3188 9182 3222
rect 9002 3149 9182 3188
rect 9002 3115 9003 3149
rect 9037 3115 9075 3149
rect 9109 3115 9147 3149
rect 9181 3115 9182 3149
rect 9002 3076 9182 3115
rect 9002 3042 9003 3076
rect 9037 3042 9075 3076
rect 9109 3042 9147 3076
rect 9181 3042 9182 3076
rect 9002 3003 9182 3042
rect 9002 2969 9003 3003
rect 9037 2969 9075 3003
rect 9109 2969 9147 3003
rect 9181 2969 9182 3003
rect 9002 2930 9182 2969
rect 9002 2896 9003 2930
rect 9037 2896 9075 2930
rect 9109 2896 9147 2930
rect 9181 2896 9182 2930
rect 9002 2857 9182 2896
rect 9002 2823 9003 2857
rect 9037 2823 9075 2857
rect 9109 2823 9147 2857
rect 9181 2823 9182 2857
rect 9002 2784 9182 2823
rect 9002 2750 9003 2784
rect 9037 2750 9075 2784
rect 9109 2750 9147 2784
rect 9181 2750 9182 2784
rect 9002 2711 9182 2750
rect 9002 2677 9003 2711
rect 9037 2677 9075 2711
rect 9109 2677 9147 2711
rect 9181 2677 9182 2711
rect 9002 2638 9182 2677
rect 9002 2604 9003 2638
rect 9037 2604 9075 2638
rect 9109 2604 9147 2638
rect 9181 2604 9182 2638
rect 9002 2565 9182 2604
rect 9002 2531 9003 2565
rect 9037 2531 9075 2565
rect 9109 2531 9147 2565
rect 9181 2531 9182 2565
rect 9002 2492 9182 2531
rect 9002 2458 9003 2492
rect 9037 2458 9075 2492
rect 9109 2458 9147 2492
rect 9181 2458 9182 2492
rect 9002 2419 9182 2458
rect 9002 2385 9003 2419
rect 9037 2385 9075 2419
rect 9109 2385 9147 2419
rect 9181 2385 9182 2419
rect 9002 2346 9182 2385
rect 9002 2312 9003 2346
rect 9037 2312 9075 2346
rect 9109 2312 9147 2346
rect 9181 2312 9182 2346
rect 9002 2273 9182 2312
rect 9002 2239 9003 2273
rect 9037 2239 9075 2273
rect 9109 2239 9147 2273
rect 9181 2239 9182 2273
rect 9002 2200 9182 2239
rect 9002 2166 9003 2200
rect 9037 2166 9075 2200
rect 9109 2166 9147 2200
rect 9181 2166 9182 2200
rect 9002 2126 9182 2166
rect 9002 2092 9003 2126
rect 9037 2092 9075 2126
rect 9109 2092 9147 2126
rect 9181 2092 9182 2126
rect 9002 2052 9182 2092
rect 9002 2018 9003 2052
rect 9037 2018 9075 2052
rect 9109 2018 9147 2052
rect 9181 2018 9182 2052
rect 9002 1978 9182 2018
rect 9002 1944 9003 1978
rect 9037 1944 9075 1978
rect 9109 1944 9147 1978
rect 9181 1944 9182 1978
rect 9002 1904 9182 1944
rect 9002 1870 9003 1904
rect 9037 1870 9075 1904
rect 9109 1870 9147 1904
rect 9181 1870 9182 1904
rect 9002 1830 9182 1870
rect 9002 1796 9003 1830
rect 9037 1796 9075 1830
rect 9109 1796 9147 1830
rect 9181 1796 9182 1830
rect 9002 1756 9182 1796
rect 9002 1722 9003 1756
rect 9037 1722 9075 1756
rect 9109 1722 9147 1756
rect 9181 1722 9182 1756
rect 9002 1682 9182 1722
rect 9002 1648 9003 1682
rect 9037 1648 9075 1682
rect 9109 1648 9147 1682
rect 9181 1648 9182 1682
rect 9002 1608 9182 1648
rect 9002 1574 9003 1608
rect 9037 1574 9075 1608
rect 9109 1574 9147 1608
rect 9181 1574 9182 1608
rect 9002 1548 9182 1574
rect 9247 3104 9367 4200
rect 9809 4308 9929 4324
rect 9809 4274 9852 4308
rect 9886 4274 9929 4308
rect 9809 4234 9929 4274
rect 9809 4200 9852 4234
rect 9886 4200 9929 4234
rect 9247 3070 9290 3104
rect 9324 3070 9367 3104
rect 9247 3026 9367 3070
rect 9247 2992 9290 3026
rect 9324 2992 9367 3026
rect 9247 2948 9367 2992
rect 9247 2914 9290 2948
rect 9324 2914 9367 2948
rect 9247 2870 9367 2914
rect 9247 2836 9290 2870
rect 9324 2836 9367 2870
rect 9247 2792 9367 2836
rect 9247 2758 9290 2792
rect 9324 2758 9367 2792
rect 9247 2713 9367 2758
rect 9247 2679 9290 2713
rect 9324 2679 9367 2713
rect 9247 2634 9367 2679
rect 9247 2600 9290 2634
rect 9324 2600 9367 2634
rect 8817 1470 8860 1504
rect 8894 1470 8937 1504
rect 8817 1430 8937 1470
rect 8817 1396 8860 1430
rect 8894 1396 8937 1430
rect 8817 1250 8937 1396
rect 8817 1144 8824 1250
rect 8930 1144 8937 1250
rect 9247 1504 9367 2600
rect 9469 4092 9707 4104
rect 9469 4058 9499 4092
rect 9533 4058 9643 4092
rect 9677 4058 9707 4092
rect 9469 4020 9707 4058
rect 9469 3986 9499 4020
rect 9533 3986 9643 4020
rect 9677 3986 9707 4020
rect 9469 3948 9707 3986
rect 9469 3914 9499 3948
rect 9533 3914 9643 3948
rect 9677 3914 9707 3948
rect 9469 3876 9707 3914
rect 9469 3842 9499 3876
rect 9533 3842 9643 3876
rect 9677 3842 9707 3876
rect 9469 3804 9707 3842
rect 9469 3770 9499 3804
rect 9533 3770 9643 3804
rect 9677 3770 9707 3804
rect 9469 3732 9707 3770
rect 9469 3698 9499 3732
rect 9533 3698 9643 3732
rect 9677 3698 9707 3732
rect 9469 3660 9707 3698
rect 9469 3626 9499 3660
rect 9533 3626 9643 3660
rect 9677 3626 9707 3660
rect 9469 3588 9707 3626
rect 9469 3554 9499 3588
rect 9533 3554 9643 3588
rect 9677 3554 9707 3588
rect 9469 3516 9707 3554
rect 9469 3482 9499 3516
rect 9533 3482 9643 3516
rect 9677 3482 9707 3516
rect 9469 3444 9707 3482
rect 9469 3410 9499 3444
rect 9533 3410 9643 3444
rect 9677 3410 9707 3444
rect 9469 3372 9707 3410
rect 9469 3338 9499 3372
rect 9533 3338 9643 3372
rect 9677 3338 9707 3372
rect 9469 3300 9707 3338
rect 9469 3266 9499 3300
rect 9533 3266 9643 3300
rect 9677 3266 9707 3300
rect 9469 3228 9707 3266
rect 9469 3194 9499 3228
rect 9533 3194 9643 3228
rect 9677 3194 9707 3228
rect 9469 3108 9707 3194
rect 9469 3074 9499 3108
rect 9533 3074 9571 3108
rect 9605 3074 9643 3108
rect 9677 3074 9707 3108
rect 9469 3044 9707 3074
rect 9469 3028 9537 3044
rect 9469 2994 9499 3028
rect 9533 3010 9537 3028
rect 9571 3028 9605 3044
rect 9533 2994 9571 3010
rect 9639 3028 9707 3044
rect 9639 3010 9643 3028
rect 9605 2994 9643 3010
rect 9677 2994 9707 3028
rect 9469 2974 9707 2994
rect 9469 2948 9537 2974
rect 9469 2914 9499 2948
rect 9533 2940 9537 2948
rect 9571 2948 9605 2974
rect 9533 2914 9571 2940
rect 9639 2948 9707 2974
rect 9639 2940 9643 2948
rect 9605 2914 9643 2940
rect 9677 2914 9707 2948
rect 9469 2904 9707 2914
rect 9469 2870 9537 2904
rect 9571 2870 9605 2904
rect 9639 2870 9707 2904
rect 9469 2868 9707 2870
rect 9469 2834 9499 2868
rect 9533 2834 9571 2868
rect 9605 2834 9643 2868
rect 9677 2834 9707 2868
rect 9469 2800 9537 2834
rect 9571 2800 9605 2834
rect 9639 2800 9707 2834
rect 9469 2788 9707 2800
rect 9469 2754 9499 2788
rect 9533 2764 9571 2788
rect 9533 2754 9537 2764
rect 9469 2730 9537 2754
rect 9605 2764 9643 2788
rect 9571 2730 9605 2754
rect 9639 2754 9643 2764
rect 9677 2754 9707 2788
rect 9639 2730 9707 2754
rect 9469 2708 9707 2730
rect 9469 2674 9499 2708
rect 9533 2694 9571 2708
rect 9533 2674 9537 2694
rect 9469 2660 9537 2674
rect 9605 2694 9643 2708
rect 9571 2660 9605 2674
rect 9639 2674 9643 2694
rect 9677 2674 9707 2708
rect 9639 2660 9707 2674
rect 9469 2628 9707 2660
rect 9469 2594 9499 2628
rect 9533 2594 9571 2628
rect 9605 2594 9643 2628
rect 9677 2594 9707 2628
rect 9469 2518 9707 2594
rect 9469 2484 9499 2518
rect 9533 2484 9643 2518
rect 9677 2484 9707 2518
rect 9469 2446 9707 2484
rect 9469 2412 9499 2446
rect 9533 2412 9643 2446
rect 9677 2412 9707 2446
rect 9469 2374 9707 2412
rect 9469 2340 9499 2374
rect 9533 2340 9643 2374
rect 9677 2340 9707 2374
rect 9469 2302 9707 2340
rect 9469 2268 9499 2302
rect 9533 2268 9643 2302
rect 9677 2268 9707 2302
rect 9469 2230 9707 2268
rect 9469 2196 9499 2230
rect 9533 2196 9643 2230
rect 9677 2196 9707 2230
rect 9469 2158 9707 2196
rect 9469 2124 9499 2158
rect 9533 2124 9643 2158
rect 9677 2124 9707 2158
rect 9469 2086 9707 2124
rect 9469 2052 9499 2086
rect 9533 2052 9643 2086
rect 9677 2052 9707 2086
rect 9469 2014 9707 2052
rect 9469 1980 9499 2014
rect 9533 1980 9643 2014
rect 9677 1980 9707 2014
rect 9469 1942 9707 1980
rect 9469 1908 9499 1942
rect 9533 1908 9643 1942
rect 9677 1908 9707 1942
rect 9469 1870 9707 1908
rect 9469 1836 9499 1870
rect 9533 1836 9643 1870
rect 9677 1836 9707 1870
rect 9469 1798 9707 1836
rect 9469 1764 9499 1798
rect 9533 1764 9643 1798
rect 9677 1764 9707 1798
rect 9469 1726 9707 1764
rect 9469 1692 9499 1726
rect 9533 1692 9643 1726
rect 9677 1692 9707 1726
rect 9469 1654 9707 1692
rect 9469 1620 9499 1654
rect 9533 1620 9643 1654
rect 9677 1620 9707 1654
rect 9469 1536 9707 1620
rect 9809 3104 9929 4200
rect 10239 4308 10359 4324
rect 10239 4274 10282 4308
rect 10316 4274 10359 4308
rect 10239 4234 10359 4274
rect 10239 4200 10282 4234
rect 10316 4200 10359 4234
rect 9809 3070 9852 3104
rect 9886 3070 9929 3104
rect 9809 3026 9929 3070
rect 9809 2992 9852 3026
rect 9886 2992 9929 3026
rect 9809 2948 9929 2992
rect 9809 2914 9852 2948
rect 9886 2914 9929 2948
rect 9809 2870 9929 2914
rect 9809 2836 9852 2870
rect 9886 2836 9929 2870
rect 9809 2792 9929 2836
rect 9809 2758 9852 2792
rect 9886 2758 9929 2792
rect 9809 2713 9929 2758
rect 9809 2679 9852 2713
rect 9886 2679 9929 2713
rect 9809 2634 9929 2679
rect 9809 2600 9852 2634
rect 9886 2600 9929 2634
rect 9247 1470 9290 1504
rect 9324 1470 9367 1504
rect 9247 1430 9367 1470
rect 9247 1396 9290 1430
rect 9324 1396 9367 1430
rect 9247 1250 9367 1396
rect 9247 1144 9254 1250
rect 9360 1144 9367 1250
rect 9809 1504 9929 2600
rect 9994 4098 10174 4118
rect 9994 4064 9995 4098
rect 10029 4064 10067 4098
rect 10101 4064 10139 4098
rect 10173 4064 10174 4098
rect 9994 4025 10174 4064
rect 9994 3991 9995 4025
rect 10029 3991 10067 4025
rect 10101 3991 10139 4025
rect 10173 3991 10174 4025
rect 9994 3952 10174 3991
rect 9994 3918 9995 3952
rect 10029 3918 10067 3952
rect 10101 3918 10139 3952
rect 10173 3918 10174 3952
rect 9994 3879 10174 3918
rect 9994 3845 9995 3879
rect 10029 3845 10067 3879
rect 10101 3845 10139 3879
rect 10173 3845 10174 3879
rect 9994 3806 10174 3845
rect 9994 3772 9995 3806
rect 10029 3772 10067 3806
rect 10101 3772 10139 3806
rect 10173 3772 10174 3806
rect 9994 3733 10174 3772
rect 9994 3699 9995 3733
rect 10029 3699 10067 3733
rect 10101 3699 10139 3733
rect 10173 3699 10174 3733
rect 9994 3660 10174 3699
rect 9994 3626 9995 3660
rect 10029 3626 10067 3660
rect 10101 3626 10139 3660
rect 10173 3626 10174 3660
rect 9994 3587 10174 3626
rect 9994 3553 9995 3587
rect 10029 3553 10067 3587
rect 10101 3553 10139 3587
rect 10173 3553 10174 3587
rect 9994 3514 10174 3553
rect 9994 3480 9995 3514
rect 10029 3480 10067 3514
rect 10101 3480 10139 3514
rect 10173 3480 10174 3514
rect 9994 3441 10174 3480
rect 9994 3407 9995 3441
rect 10029 3407 10067 3441
rect 10101 3407 10139 3441
rect 10173 3407 10174 3441
rect 9994 3368 10174 3407
rect 9994 3334 9995 3368
rect 10029 3334 10067 3368
rect 10101 3334 10139 3368
rect 10173 3334 10174 3368
rect 9994 3295 10174 3334
rect 9994 3261 9995 3295
rect 10029 3261 10067 3295
rect 10101 3261 10139 3295
rect 10173 3261 10174 3295
rect 9994 3222 10174 3261
rect 9994 3188 9995 3222
rect 10029 3188 10067 3222
rect 10101 3188 10139 3222
rect 10173 3188 10174 3222
rect 9994 3149 10174 3188
rect 9994 3115 9995 3149
rect 10029 3115 10067 3149
rect 10101 3115 10139 3149
rect 10173 3115 10174 3149
rect 9994 3076 10174 3115
rect 9994 3042 9995 3076
rect 10029 3042 10067 3076
rect 10101 3042 10139 3076
rect 10173 3042 10174 3076
rect 9994 3003 10174 3042
rect 9994 2969 9995 3003
rect 10029 2969 10067 3003
rect 10101 2969 10139 3003
rect 10173 2969 10174 3003
rect 9994 2930 10174 2969
rect 9994 2896 9995 2930
rect 10029 2896 10067 2930
rect 10101 2896 10139 2930
rect 10173 2896 10174 2930
rect 9994 2857 10174 2896
rect 9994 2823 9995 2857
rect 10029 2823 10067 2857
rect 10101 2823 10139 2857
rect 10173 2823 10174 2857
rect 9994 2784 10174 2823
rect 9994 2750 9995 2784
rect 10029 2750 10067 2784
rect 10101 2750 10139 2784
rect 10173 2750 10174 2784
rect 9994 2711 10174 2750
rect 9994 2677 9995 2711
rect 10029 2677 10067 2711
rect 10101 2677 10139 2711
rect 10173 2677 10174 2711
rect 9994 2638 10174 2677
rect 9994 2604 9995 2638
rect 10029 2604 10067 2638
rect 10101 2604 10139 2638
rect 10173 2604 10174 2638
rect 9994 2565 10174 2604
rect 9994 2531 9995 2565
rect 10029 2531 10067 2565
rect 10101 2531 10139 2565
rect 10173 2531 10174 2565
rect 9994 2492 10174 2531
rect 9994 2458 9995 2492
rect 10029 2458 10067 2492
rect 10101 2458 10139 2492
rect 10173 2458 10174 2492
rect 9994 2419 10174 2458
rect 9994 2385 9995 2419
rect 10029 2385 10067 2419
rect 10101 2385 10139 2419
rect 10173 2385 10174 2419
rect 9994 2346 10174 2385
rect 9994 2312 9995 2346
rect 10029 2312 10067 2346
rect 10101 2312 10139 2346
rect 10173 2312 10174 2346
rect 9994 2273 10174 2312
rect 9994 2239 9995 2273
rect 10029 2239 10067 2273
rect 10101 2239 10139 2273
rect 10173 2239 10174 2273
rect 9994 2200 10174 2239
rect 9994 2166 9995 2200
rect 10029 2166 10067 2200
rect 10101 2166 10139 2200
rect 10173 2166 10174 2200
rect 9994 2126 10174 2166
rect 9994 2092 9995 2126
rect 10029 2092 10067 2126
rect 10101 2092 10139 2126
rect 10173 2092 10174 2126
rect 9994 2052 10174 2092
rect 9994 2018 9995 2052
rect 10029 2018 10067 2052
rect 10101 2018 10139 2052
rect 10173 2018 10174 2052
rect 9994 1978 10174 2018
rect 9994 1944 9995 1978
rect 10029 1944 10067 1978
rect 10101 1944 10139 1978
rect 10173 1944 10174 1978
rect 9994 1904 10174 1944
rect 9994 1870 9995 1904
rect 10029 1870 10067 1904
rect 10101 1870 10139 1904
rect 10173 1870 10174 1904
rect 9994 1830 10174 1870
rect 9994 1796 9995 1830
rect 10029 1796 10067 1830
rect 10101 1796 10139 1830
rect 10173 1796 10174 1830
rect 9994 1756 10174 1796
rect 9994 1722 9995 1756
rect 10029 1722 10067 1756
rect 10101 1722 10139 1756
rect 10173 1722 10174 1756
rect 9994 1682 10174 1722
rect 9994 1648 9995 1682
rect 10029 1648 10067 1682
rect 10101 1648 10139 1682
rect 10173 1648 10174 1682
rect 9994 1608 10174 1648
rect 9994 1574 9995 1608
rect 10029 1574 10067 1608
rect 10101 1574 10139 1608
rect 10173 1574 10174 1608
rect 9994 1548 10174 1574
rect 10239 3104 10359 4200
rect 10801 4308 10921 4324
rect 10801 4274 10844 4308
rect 10878 4274 10921 4308
rect 10801 4234 10921 4274
rect 10801 4200 10844 4234
rect 10878 4200 10921 4234
rect 10239 3070 10282 3104
rect 10316 3070 10359 3104
rect 10239 3026 10359 3070
rect 10239 2992 10282 3026
rect 10316 2992 10359 3026
rect 10239 2948 10359 2992
rect 10239 2914 10282 2948
rect 10316 2914 10359 2948
rect 10239 2870 10359 2914
rect 10239 2836 10282 2870
rect 10316 2836 10359 2870
rect 10239 2792 10359 2836
rect 10239 2758 10282 2792
rect 10316 2758 10359 2792
rect 10239 2713 10359 2758
rect 10239 2679 10282 2713
rect 10316 2679 10359 2713
rect 10239 2634 10359 2679
rect 10239 2600 10282 2634
rect 10316 2600 10359 2634
rect 9809 1470 9852 1504
rect 9886 1470 9929 1504
rect 9809 1430 9929 1470
rect 9809 1396 9852 1430
rect 9886 1396 9929 1430
rect 9809 1250 9929 1396
rect 9809 1144 9816 1250
rect 9922 1144 9929 1250
rect 10239 1504 10359 2600
rect 10461 4092 10699 4130
rect 10461 4058 10491 4092
rect 10525 4058 10635 4092
rect 10669 4058 10699 4092
rect 10461 4020 10699 4058
rect 10461 3986 10491 4020
rect 10525 3986 10635 4020
rect 10669 3986 10699 4020
rect 10461 3948 10699 3986
rect 10461 3914 10491 3948
rect 10525 3914 10635 3948
rect 10669 3914 10699 3948
rect 10461 3876 10699 3914
rect 10461 3842 10491 3876
rect 10525 3842 10635 3876
rect 10669 3842 10699 3876
rect 10461 3804 10699 3842
rect 10461 3770 10491 3804
rect 10525 3770 10635 3804
rect 10669 3770 10699 3804
rect 10461 3732 10699 3770
rect 10461 3698 10491 3732
rect 10525 3698 10635 3732
rect 10669 3698 10699 3732
rect 10461 3660 10699 3698
rect 10461 3626 10491 3660
rect 10525 3626 10635 3660
rect 10669 3626 10699 3660
rect 10461 3588 10699 3626
rect 10461 3554 10491 3588
rect 10525 3554 10635 3588
rect 10669 3554 10699 3588
rect 10461 3516 10699 3554
rect 10461 3482 10491 3516
rect 10525 3482 10635 3516
rect 10669 3482 10699 3516
rect 10461 3444 10699 3482
rect 10461 3410 10491 3444
rect 10525 3410 10635 3444
rect 10669 3410 10699 3444
rect 10461 3372 10699 3410
rect 10461 3338 10491 3372
rect 10525 3338 10635 3372
rect 10669 3338 10699 3372
rect 10461 3300 10699 3338
rect 10461 3266 10491 3300
rect 10525 3266 10635 3300
rect 10669 3266 10699 3300
rect 10461 3228 10699 3266
rect 10461 3194 10491 3228
rect 10525 3194 10635 3228
rect 10669 3194 10699 3228
rect 10461 3108 10699 3194
rect 10461 3074 10491 3108
rect 10525 3074 10563 3108
rect 10597 3074 10635 3108
rect 10669 3074 10699 3108
rect 10461 3044 10699 3074
rect 10461 3028 10529 3044
rect 10461 2994 10491 3028
rect 10525 3010 10529 3028
rect 10563 3028 10597 3044
rect 10525 2994 10563 3010
rect 10631 3028 10699 3044
rect 10631 3010 10635 3028
rect 10597 2994 10635 3010
rect 10669 2994 10699 3028
rect 10461 2974 10699 2994
rect 10461 2948 10529 2974
rect 10461 2914 10491 2948
rect 10525 2940 10529 2948
rect 10563 2948 10597 2974
rect 10525 2914 10563 2940
rect 10631 2948 10699 2974
rect 10631 2940 10635 2948
rect 10597 2914 10635 2940
rect 10669 2914 10699 2948
rect 10461 2904 10699 2914
rect 10461 2870 10529 2904
rect 10563 2870 10597 2904
rect 10631 2870 10699 2904
rect 10461 2868 10699 2870
rect 10461 2834 10491 2868
rect 10525 2834 10563 2868
rect 10597 2834 10635 2868
rect 10669 2834 10699 2868
rect 10461 2800 10529 2834
rect 10563 2800 10597 2834
rect 10631 2800 10699 2834
rect 10461 2788 10699 2800
rect 10461 2754 10491 2788
rect 10525 2764 10563 2788
rect 10525 2754 10529 2764
rect 10461 2730 10529 2754
rect 10597 2764 10635 2788
rect 10563 2730 10597 2754
rect 10631 2754 10635 2764
rect 10669 2754 10699 2788
rect 10631 2730 10699 2754
rect 10461 2708 10699 2730
rect 10461 2674 10491 2708
rect 10525 2694 10563 2708
rect 10525 2674 10529 2694
rect 10461 2660 10529 2674
rect 10597 2694 10635 2708
rect 10563 2660 10597 2674
rect 10631 2674 10635 2694
rect 10669 2674 10699 2708
rect 10631 2660 10699 2674
rect 10461 2628 10699 2660
rect 10461 2594 10491 2628
rect 10525 2594 10563 2628
rect 10597 2594 10635 2628
rect 10669 2594 10699 2628
rect 10461 2518 10699 2594
rect 10461 2484 10491 2518
rect 10525 2484 10635 2518
rect 10669 2484 10699 2518
rect 10461 2446 10699 2484
rect 10461 2412 10491 2446
rect 10525 2412 10635 2446
rect 10669 2412 10699 2446
rect 10461 2374 10699 2412
rect 10461 2340 10491 2374
rect 10525 2340 10635 2374
rect 10669 2340 10699 2374
rect 10461 2302 10699 2340
rect 10461 2268 10491 2302
rect 10525 2268 10635 2302
rect 10669 2268 10699 2302
rect 10461 2230 10699 2268
rect 10461 2196 10491 2230
rect 10525 2196 10635 2230
rect 10669 2196 10699 2230
rect 10461 2158 10699 2196
rect 10461 2124 10491 2158
rect 10525 2124 10635 2158
rect 10669 2124 10699 2158
rect 10461 2086 10699 2124
rect 10461 2052 10491 2086
rect 10525 2052 10635 2086
rect 10669 2052 10699 2086
rect 10461 2014 10699 2052
rect 10461 1980 10491 2014
rect 10525 1980 10635 2014
rect 10669 1980 10699 2014
rect 10461 1942 10699 1980
rect 10461 1908 10491 1942
rect 10525 1908 10635 1942
rect 10669 1908 10699 1942
rect 10461 1870 10699 1908
rect 10461 1836 10491 1870
rect 10525 1836 10635 1870
rect 10669 1836 10699 1870
rect 10461 1798 10699 1836
rect 10461 1764 10491 1798
rect 10525 1764 10635 1798
rect 10669 1764 10699 1798
rect 10461 1726 10699 1764
rect 10461 1692 10491 1726
rect 10525 1692 10635 1726
rect 10669 1692 10699 1726
rect 10461 1654 10699 1692
rect 10461 1620 10491 1654
rect 10525 1620 10635 1654
rect 10669 1620 10699 1654
rect 10461 1536 10699 1620
rect 10801 3104 10921 4200
rect 11231 4308 11351 4324
rect 11231 4274 11274 4308
rect 11308 4274 11351 4308
rect 11231 4234 11351 4274
rect 11231 4200 11274 4234
rect 11308 4200 11351 4234
rect 10801 3070 10844 3104
rect 10878 3070 10921 3104
rect 10801 3026 10921 3070
rect 10801 2992 10844 3026
rect 10878 2992 10921 3026
rect 10801 2948 10921 2992
rect 10801 2914 10844 2948
rect 10878 2914 10921 2948
rect 10801 2870 10921 2914
rect 10801 2836 10844 2870
rect 10878 2836 10921 2870
rect 10801 2792 10921 2836
rect 10801 2758 10844 2792
rect 10878 2758 10921 2792
rect 10801 2713 10921 2758
rect 10801 2679 10844 2713
rect 10878 2679 10921 2713
rect 10801 2634 10921 2679
rect 10801 2600 10844 2634
rect 10878 2600 10921 2634
rect 10239 1470 10282 1504
rect 10316 1470 10359 1504
rect 10239 1430 10359 1470
rect 10239 1396 10282 1430
rect 10316 1396 10359 1430
rect 10239 1250 10359 1396
rect 10239 1144 10246 1250
rect 10352 1144 10359 1250
rect 10801 1504 10921 2600
rect 10986 4064 10987 4098
rect 11021 4064 11059 4098
rect 11093 4064 11131 4098
rect 11165 4064 11166 4098
rect 10986 4025 11166 4064
rect 10986 3991 10987 4025
rect 11021 3991 11059 4025
rect 11093 3991 11131 4025
rect 11165 3991 11166 4025
rect 10986 3952 11166 3991
rect 10986 3918 10987 3952
rect 11021 3918 11059 3952
rect 11093 3918 11131 3952
rect 11165 3918 11166 3952
rect 10986 3879 11166 3918
rect 10986 3845 10987 3879
rect 11021 3845 11059 3879
rect 11093 3845 11131 3879
rect 11165 3845 11166 3879
rect 10986 3806 11166 3845
rect 10986 3772 10987 3806
rect 11021 3772 11059 3806
rect 11093 3772 11131 3806
rect 11165 3772 11166 3806
rect 10986 3733 11166 3772
rect 10986 3699 10987 3733
rect 11021 3699 11059 3733
rect 11093 3699 11131 3733
rect 11165 3699 11166 3733
rect 10986 3660 11166 3699
rect 10986 3626 10987 3660
rect 11021 3626 11059 3660
rect 11093 3626 11131 3660
rect 11165 3626 11166 3660
rect 10986 3587 11166 3626
rect 10986 3553 10987 3587
rect 11021 3553 11059 3587
rect 11093 3553 11131 3587
rect 11165 3553 11166 3587
rect 10986 3514 11166 3553
rect 10986 3480 10987 3514
rect 11021 3480 11059 3514
rect 11093 3480 11131 3514
rect 11165 3480 11166 3514
rect 10986 3441 11166 3480
rect 10986 3407 10987 3441
rect 11021 3407 11059 3441
rect 11093 3407 11131 3441
rect 11165 3407 11166 3441
rect 10986 3368 11166 3407
rect 10986 3334 10987 3368
rect 11021 3334 11059 3368
rect 11093 3334 11131 3368
rect 11165 3334 11166 3368
rect 10986 3295 11166 3334
rect 10986 3261 10987 3295
rect 11021 3261 11059 3295
rect 11093 3261 11131 3295
rect 11165 3261 11166 3295
rect 10986 3222 11166 3261
rect 10986 3188 10987 3222
rect 11021 3188 11059 3222
rect 11093 3188 11131 3222
rect 11165 3188 11166 3222
rect 10986 3149 11166 3188
rect 10986 3115 10987 3149
rect 11021 3115 11059 3149
rect 11093 3115 11131 3149
rect 11165 3115 11166 3149
rect 10986 3076 11166 3115
rect 10986 3042 10987 3076
rect 11021 3042 11059 3076
rect 11093 3042 11131 3076
rect 11165 3042 11166 3076
rect 10986 3003 11166 3042
rect 10986 2969 10987 3003
rect 11021 2969 11059 3003
rect 11093 2969 11131 3003
rect 11165 2969 11166 3003
rect 10986 2930 11166 2969
rect 10986 2896 10987 2930
rect 11021 2896 11059 2930
rect 11093 2896 11131 2930
rect 11165 2896 11166 2930
rect 10986 2857 11166 2896
rect 10986 2823 10987 2857
rect 11021 2823 11059 2857
rect 11093 2823 11131 2857
rect 11165 2823 11166 2857
rect 10986 2784 11166 2823
rect 10986 2750 10987 2784
rect 11021 2750 11059 2784
rect 11093 2750 11131 2784
rect 11165 2750 11166 2784
rect 10986 2711 11166 2750
rect 10986 2677 10987 2711
rect 11021 2677 11059 2711
rect 11093 2677 11131 2711
rect 11165 2677 11166 2711
rect 10986 2638 11166 2677
rect 10986 2604 10987 2638
rect 11021 2604 11059 2638
rect 11093 2604 11131 2638
rect 11165 2604 11166 2638
rect 10986 2565 11166 2604
rect 10986 2531 10987 2565
rect 11021 2531 11059 2565
rect 11093 2531 11131 2565
rect 11165 2531 11166 2565
rect 10986 2492 11166 2531
rect 10986 2458 10987 2492
rect 11021 2458 11059 2492
rect 11093 2458 11131 2492
rect 11165 2458 11166 2492
rect 10986 2419 11166 2458
rect 10986 2385 10987 2419
rect 11021 2385 11059 2419
rect 11093 2385 11131 2419
rect 11165 2385 11166 2419
rect 10986 2346 11166 2385
rect 10986 2312 10987 2346
rect 11021 2312 11059 2346
rect 11093 2312 11131 2346
rect 11165 2312 11166 2346
rect 10986 2273 11166 2312
rect 10986 2239 10987 2273
rect 11021 2239 11059 2273
rect 11093 2239 11131 2273
rect 11165 2239 11166 2273
rect 10986 2200 11166 2239
rect 10986 2166 10987 2200
rect 11021 2166 11059 2200
rect 11093 2166 11131 2200
rect 11165 2166 11166 2200
rect 10986 2126 11166 2166
rect 10986 2092 10987 2126
rect 11021 2092 11059 2126
rect 11093 2092 11131 2126
rect 11165 2092 11166 2126
rect 10986 2052 11166 2092
rect 10986 2018 10987 2052
rect 11021 2018 11059 2052
rect 11093 2018 11131 2052
rect 11165 2018 11166 2052
rect 10986 1978 11166 2018
rect 10986 1944 10987 1978
rect 11021 1944 11059 1978
rect 11093 1944 11131 1978
rect 11165 1944 11166 1978
rect 10986 1904 11166 1944
rect 10986 1870 10987 1904
rect 11021 1870 11059 1904
rect 11093 1870 11131 1904
rect 11165 1870 11166 1904
rect 10986 1830 11166 1870
rect 10986 1796 10987 1830
rect 11021 1796 11059 1830
rect 11093 1796 11131 1830
rect 11165 1796 11166 1830
rect 10986 1756 11166 1796
rect 10986 1722 10987 1756
rect 11021 1722 11059 1756
rect 11093 1722 11131 1756
rect 11165 1722 11166 1756
rect 10986 1682 11166 1722
rect 10986 1648 10987 1682
rect 11021 1648 11059 1682
rect 11093 1648 11131 1682
rect 11165 1648 11166 1682
rect 10986 1608 11166 1648
rect 10986 1574 10987 1608
rect 11021 1574 11059 1608
rect 11093 1574 11131 1608
rect 11165 1574 11166 1608
rect 10986 1548 11166 1574
rect 11231 3104 11351 4200
rect 11793 4308 11913 4324
rect 11793 4274 11836 4308
rect 11870 4274 11913 4308
rect 11793 4234 11913 4274
rect 11793 4200 11836 4234
rect 11870 4200 11913 4234
rect 11231 3070 11274 3104
rect 11308 3070 11351 3104
rect 11231 3026 11351 3070
rect 11231 2992 11274 3026
rect 11308 2992 11351 3026
rect 11231 2948 11351 2992
rect 11231 2914 11274 2948
rect 11308 2914 11351 2948
rect 11231 2870 11351 2914
rect 11231 2836 11274 2870
rect 11308 2836 11351 2870
rect 11231 2792 11351 2836
rect 11231 2758 11274 2792
rect 11308 2758 11351 2792
rect 11231 2713 11351 2758
rect 11231 2679 11274 2713
rect 11308 2679 11351 2713
rect 11231 2634 11351 2679
rect 11231 2600 11274 2634
rect 11308 2600 11351 2634
rect 10801 1470 10844 1504
rect 10878 1470 10921 1504
rect 10801 1430 10921 1470
rect 10801 1396 10844 1430
rect 10878 1396 10921 1430
rect 10801 1250 10921 1396
rect 10801 1144 10808 1250
rect 10914 1144 10921 1250
rect 11231 1504 11351 2600
rect 11453 4092 11691 4110
rect 11453 4058 11483 4092
rect 11517 4058 11627 4092
rect 11661 4058 11691 4092
rect 11453 4020 11691 4058
rect 11453 3986 11483 4020
rect 11517 3986 11627 4020
rect 11661 3986 11691 4020
rect 11453 3948 11691 3986
rect 11453 3914 11483 3948
rect 11517 3914 11627 3948
rect 11661 3914 11691 3948
rect 11453 3876 11691 3914
rect 11453 3842 11483 3876
rect 11517 3842 11627 3876
rect 11661 3842 11691 3876
rect 11453 3804 11691 3842
rect 11453 3770 11483 3804
rect 11517 3770 11627 3804
rect 11661 3770 11691 3804
rect 11453 3732 11691 3770
rect 11453 3698 11483 3732
rect 11517 3698 11627 3732
rect 11661 3698 11691 3732
rect 11453 3660 11691 3698
rect 11453 3626 11483 3660
rect 11517 3626 11627 3660
rect 11661 3626 11691 3660
rect 11453 3588 11691 3626
rect 11453 3554 11483 3588
rect 11517 3554 11627 3588
rect 11661 3554 11691 3588
rect 11453 3516 11691 3554
rect 11453 3482 11483 3516
rect 11517 3482 11627 3516
rect 11661 3482 11691 3516
rect 11453 3444 11691 3482
rect 11453 3410 11483 3444
rect 11517 3410 11627 3444
rect 11661 3410 11691 3444
rect 11453 3372 11691 3410
rect 11453 3338 11483 3372
rect 11517 3338 11627 3372
rect 11661 3338 11691 3372
rect 11453 3300 11691 3338
rect 11453 3266 11483 3300
rect 11517 3266 11627 3300
rect 11661 3266 11691 3300
rect 11453 3228 11691 3266
rect 11453 3194 11483 3228
rect 11517 3194 11627 3228
rect 11661 3194 11691 3228
rect 11453 3108 11691 3194
rect 11453 3074 11483 3108
rect 11517 3074 11555 3108
rect 11589 3074 11627 3108
rect 11661 3074 11691 3108
rect 11453 3044 11691 3074
rect 11453 3028 11521 3044
rect 11453 2994 11483 3028
rect 11517 3010 11521 3028
rect 11555 3028 11589 3044
rect 11517 2994 11555 3010
rect 11623 3028 11691 3044
rect 11623 3010 11627 3028
rect 11589 2994 11627 3010
rect 11661 2994 11691 3028
rect 11453 2974 11691 2994
rect 11453 2948 11521 2974
rect 11453 2914 11483 2948
rect 11517 2940 11521 2948
rect 11555 2948 11589 2974
rect 11517 2914 11555 2940
rect 11623 2948 11691 2974
rect 11623 2940 11627 2948
rect 11589 2914 11627 2940
rect 11661 2914 11691 2948
rect 11453 2904 11691 2914
rect 11453 2870 11521 2904
rect 11555 2870 11589 2904
rect 11623 2870 11691 2904
rect 11453 2868 11691 2870
rect 11453 2834 11483 2868
rect 11517 2834 11555 2868
rect 11589 2834 11627 2868
rect 11661 2834 11691 2868
rect 11453 2800 11521 2834
rect 11555 2800 11589 2834
rect 11623 2800 11691 2834
rect 11453 2788 11691 2800
rect 11453 2754 11483 2788
rect 11517 2764 11555 2788
rect 11517 2754 11521 2764
rect 11453 2730 11521 2754
rect 11589 2764 11627 2788
rect 11555 2730 11589 2754
rect 11623 2754 11627 2764
rect 11661 2754 11691 2788
rect 11623 2730 11691 2754
rect 11453 2708 11691 2730
rect 11453 2674 11483 2708
rect 11517 2694 11555 2708
rect 11517 2674 11521 2694
rect 11453 2660 11521 2674
rect 11589 2694 11627 2708
rect 11555 2660 11589 2674
rect 11623 2674 11627 2694
rect 11661 2674 11691 2708
rect 11623 2660 11691 2674
rect 11453 2628 11691 2660
rect 11453 2594 11483 2628
rect 11517 2594 11555 2628
rect 11589 2594 11627 2628
rect 11661 2594 11691 2628
rect 11453 2518 11691 2594
rect 11453 2484 11483 2518
rect 11517 2484 11627 2518
rect 11661 2484 11691 2518
rect 11453 2446 11691 2484
rect 11453 2412 11483 2446
rect 11517 2412 11627 2446
rect 11661 2412 11691 2446
rect 11453 2374 11691 2412
rect 11453 2340 11483 2374
rect 11517 2340 11627 2374
rect 11661 2340 11691 2374
rect 11453 2302 11691 2340
rect 11453 2268 11483 2302
rect 11517 2268 11627 2302
rect 11661 2268 11691 2302
rect 11453 2230 11691 2268
rect 11453 2196 11483 2230
rect 11517 2196 11627 2230
rect 11661 2196 11691 2230
rect 11453 2158 11691 2196
rect 11453 2124 11483 2158
rect 11517 2124 11627 2158
rect 11661 2124 11691 2158
rect 11453 2086 11691 2124
rect 11453 2052 11483 2086
rect 11517 2052 11627 2086
rect 11661 2052 11691 2086
rect 11453 2014 11691 2052
rect 11453 1980 11483 2014
rect 11517 1980 11627 2014
rect 11661 1980 11691 2014
rect 11453 1942 11691 1980
rect 11453 1908 11483 1942
rect 11517 1908 11627 1942
rect 11661 1908 11691 1942
rect 11453 1870 11691 1908
rect 11453 1836 11483 1870
rect 11517 1836 11627 1870
rect 11661 1836 11691 1870
rect 11453 1798 11691 1836
rect 11453 1764 11483 1798
rect 11517 1764 11627 1798
rect 11661 1764 11691 1798
rect 11453 1726 11691 1764
rect 11453 1692 11483 1726
rect 11517 1692 11627 1726
rect 11661 1692 11691 1726
rect 11453 1654 11691 1692
rect 11453 1620 11483 1654
rect 11517 1620 11627 1654
rect 11661 1620 11691 1654
rect 11453 1536 11691 1620
rect 11793 3104 11913 4200
rect 12223 4308 12343 4324
rect 12223 4274 12266 4308
rect 12300 4274 12343 4308
rect 12223 4234 12343 4274
rect 12223 4200 12266 4234
rect 12300 4200 12343 4234
rect 11793 3070 11836 3104
rect 11870 3070 11913 3104
rect 11793 3026 11913 3070
rect 11793 2992 11836 3026
rect 11870 2992 11913 3026
rect 11793 2948 11913 2992
rect 11793 2914 11836 2948
rect 11870 2914 11913 2948
rect 11793 2870 11913 2914
rect 11793 2836 11836 2870
rect 11870 2836 11913 2870
rect 11793 2792 11913 2836
rect 11793 2758 11836 2792
rect 11870 2758 11913 2792
rect 11793 2713 11913 2758
rect 11793 2679 11836 2713
rect 11870 2679 11913 2713
rect 11793 2634 11913 2679
rect 11793 2600 11836 2634
rect 11870 2600 11913 2634
rect 11231 1470 11274 1504
rect 11308 1470 11351 1504
rect 11231 1430 11351 1470
rect 11231 1396 11274 1430
rect 11308 1396 11351 1430
rect 11231 1250 11351 1396
rect 11231 1144 11238 1250
rect 11344 1144 11351 1250
rect 11793 1504 11913 2600
rect 11978 4064 11979 4098
rect 12013 4064 12051 4098
rect 12085 4064 12123 4098
rect 12157 4064 12158 4098
rect 11978 4025 12158 4064
rect 11978 3991 11979 4025
rect 12013 3991 12051 4025
rect 12085 3991 12123 4025
rect 12157 3991 12158 4025
rect 11978 3952 12158 3991
rect 11978 3918 11979 3952
rect 12013 3918 12051 3952
rect 12085 3918 12123 3952
rect 12157 3918 12158 3952
rect 11978 3879 12158 3918
rect 11978 3845 11979 3879
rect 12013 3845 12051 3879
rect 12085 3845 12123 3879
rect 12157 3845 12158 3879
rect 11978 3806 12158 3845
rect 11978 3772 11979 3806
rect 12013 3772 12051 3806
rect 12085 3772 12123 3806
rect 12157 3772 12158 3806
rect 11978 3733 12158 3772
rect 11978 3699 11979 3733
rect 12013 3699 12051 3733
rect 12085 3699 12123 3733
rect 12157 3699 12158 3733
rect 11978 3660 12158 3699
rect 11978 3626 11979 3660
rect 12013 3626 12051 3660
rect 12085 3626 12123 3660
rect 12157 3626 12158 3660
rect 11978 3587 12158 3626
rect 11978 3553 11979 3587
rect 12013 3553 12051 3587
rect 12085 3553 12123 3587
rect 12157 3553 12158 3587
rect 11978 3514 12158 3553
rect 11978 3480 11979 3514
rect 12013 3480 12051 3514
rect 12085 3480 12123 3514
rect 12157 3480 12158 3514
rect 11978 3441 12158 3480
rect 11978 3407 11979 3441
rect 12013 3407 12051 3441
rect 12085 3407 12123 3441
rect 12157 3407 12158 3441
rect 11978 3368 12158 3407
rect 11978 3334 11979 3368
rect 12013 3334 12051 3368
rect 12085 3334 12123 3368
rect 12157 3334 12158 3368
rect 11978 3295 12158 3334
rect 11978 3261 11979 3295
rect 12013 3261 12051 3295
rect 12085 3261 12123 3295
rect 12157 3261 12158 3295
rect 11978 3222 12158 3261
rect 11978 3188 11979 3222
rect 12013 3188 12051 3222
rect 12085 3188 12123 3222
rect 12157 3188 12158 3222
rect 11978 3149 12158 3188
rect 11978 3115 11979 3149
rect 12013 3115 12051 3149
rect 12085 3115 12123 3149
rect 12157 3115 12158 3149
rect 11978 3076 12158 3115
rect 11978 3042 11979 3076
rect 12013 3042 12051 3076
rect 12085 3042 12123 3076
rect 12157 3042 12158 3076
rect 11978 3003 12158 3042
rect 11978 2969 11979 3003
rect 12013 2969 12051 3003
rect 12085 2969 12123 3003
rect 12157 2969 12158 3003
rect 11978 2930 12158 2969
rect 11978 2896 11979 2930
rect 12013 2896 12051 2930
rect 12085 2896 12123 2930
rect 12157 2896 12158 2930
rect 11978 2857 12158 2896
rect 11978 2823 11979 2857
rect 12013 2823 12051 2857
rect 12085 2823 12123 2857
rect 12157 2823 12158 2857
rect 11978 2784 12158 2823
rect 11978 2750 11979 2784
rect 12013 2750 12051 2784
rect 12085 2750 12123 2784
rect 12157 2750 12158 2784
rect 11978 2711 12158 2750
rect 11978 2677 11979 2711
rect 12013 2677 12051 2711
rect 12085 2677 12123 2711
rect 12157 2677 12158 2711
rect 11978 2638 12158 2677
rect 11978 2604 11979 2638
rect 12013 2604 12051 2638
rect 12085 2604 12123 2638
rect 12157 2604 12158 2638
rect 11978 2565 12158 2604
rect 11978 2531 11979 2565
rect 12013 2531 12051 2565
rect 12085 2531 12123 2565
rect 12157 2531 12158 2565
rect 11978 2492 12158 2531
rect 11978 2458 11979 2492
rect 12013 2458 12051 2492
rect 12085 2458 12123 2492
rect 12157 2458 12158 2492
rect 11978 2419 12158 2458
rect 11978 2385 11979 2419
rect 12013 2385 12051 2419
rect 12085 2385 12123 2419
rect 12157 2385 12158 2419
rect 11978 2346 12158 2385
rect 11978 2312 11979 2346
rect 12013 2312 12051 2346
rect 12085 2312 12123 2346
rect 12157 2312 12158 2346
rect 11978 2273 12158 2312
rect 11978 2239 11979 2273
rect 12013 2239 12051 2273
rect 12085 2239 12123 2273
rect 12157 2239 12158 2273
rect 11978 2200 12158 2239
rect 11978 2166 11979 2200
rect 12013 2166 12051 2200
rect 12085 2166 12123 2200
rect 12157 2166 12158 2200
rect 11978 2126 12158 2166
rect 11978 2092 11979 2126
rect 12013 2092 12051 2126
rect 12085 2092 12123 2126
rect 12157 2092 12158 2126
rect 11978 2052 12158 2092
rect 11978 2018 11979 2052
rect 12013 2018 12051 2052
rect 12085 2018 12123 2052
rect 12157 2018 12158 2052
rect 11978 1978 12158 2018
rect 11978 1944 11979 1978
rect 12013 1944 12051 1978
rect 12085 1944 12123 1978
rect 12157 1944 12158 1978
rect 11978 1904 12158 1944
rect 11978 1870 11979 1904
rect 12013 1870 12051 1904
rect 12085 1870 12123 1904
rect 12157 1870 12158 1904
rect 11978 1830 12158 1870
rect 11978 1796 11979 1830
rect 12013 1796 12051 1830
rect 12085 1796 12123 1830
rect 12157 1796 12158 1830
rect 11978 1756 12158 1796
rect 11978 1722 11979 1756
rect 12013 1722 12051 1756
rect 12085 1722 12123 1756
rect 12157 1722 12158 1756
rect 11978 1682 12158 1722
rect 11978 1648 11979 1682
rect 12013 1648 12051 1682
rect 12085 1648 12123 1682
rect 12157 1648 12158 1682
rect 11978 1608 12158 1648
rect 11978 1574 11979 1608
rect 12013 1574 12051 1608
rect 12085 1574 12123 1608
rect 12157 1574 12158 1608
rect 11978 1548 12158 1574
rect 12223 3104 12343 4200
rect 12785 4308 12905 4324
rect 12785 4274 12828 4308
rect 12862 4274 12905 4308
rect 12785 4234 12905 4274
rect 12785 4200 12828 4234
rect 12862 4200 12905 4234
rect 12223 3070 12266 3104
rect 12300 3070 12343 3104
rect 12223 3026 12343 3070
rect 12223 2992 12266 3026
rect 12300 2992 12343 3026
rect 12223 2948 12343 2992
rect 12223 2914 12266 2948
rect 12300 2914 12343 2948
rect 12223 2870 12343 2914
rect 12223 2836 12266 2870
rect 12300 2836 12343 2870
rect 12223 2792 12343 2836
rect 12223 2758 12266 2792
rect 12300 2758 12343 2792
rect 12223 2713 12343 2758
rect 12223 2679 12266 2713
rect 12300 2679 12343 2713
rect 12223 2634 12343 2679
rect 12223 2600 12266 2634
rect 12300 2600 12343 2634
rect 11793 1470 11836 1504
rect 11870 1470 11913 1504
rect 11793 1430 11913 1470
rect 11793 1396 11836 1430
rect 11870 1396 11913 1430
rect 11793 1250 11913 1396
rect 11793 1144 11800 1250
rect 11906 1144 11913 1250
rect 12223 1504 12343 2600
rect 12445 4092 12683 4110
rect 12445 4058 12475 4092
rect 12509 4058 12619 4092
rect 12653 4058 12683 4092
rect 12445 4020 12683 4058
rect 12445 3986 12475 4020
rect 12509 3986 12619 4020
rect 12653 3986 12683 4020
rect 12445 3948 12683 3986
rect 12445 3914 12475 3948
rect 12509 3914 12619 3948
rect 12653 3914 12683 3948
rect 12445 3876 12683 3914
rect 12445 3842 12475 3876
rect 12509 3842 12619 3876
rect 12653 3842 12683 3876
rect 12445 3804 12683 3842
rect 12445 3770 12475 3804
rect 12509 3770 12619 3804
rect 12653 3770 12683 3804
rect 12445 3732 12683 3770
rect 12445 3698 12475 3732
rect 12509 3698 12619 3732
rect 12653 3698 12683 3732
rect 12445 3660 12683 3698
rect 12445 3626 12475 3660
rect 12509 3626 12619 3660
rect 12653 3626 12683 3660
rect 12445 3588 12683 3626
rect 12445 3554 12475 3588
rect 12509 3554 12619 3588
rect 12653 3554 12683 3588
rect 12445 3516 12683 3554
rect 12445 3482 12475 3516
rect 12509 3482 12619 3516
rect 12653 3482 12683 3516
rect 12445 3444 12683 3482
rect 12445 3410 12475 3444
rect 12509 3410 12619 3444
rect 12653 3410 12683 3444
rect 12445 3372 12683 3410
rect 12445 3338 12475 3372
rect 12509 3338 12619 3372
rect 12653 3338 12683 3372
rect 12445 3300 12683 3338
rect 12445 3266 12475 3300
rect 12509 3266 12619 3300
rect 12653 3266 12683 3300
rect 12445 3228 12683 3266
rect 12445 3194 12475 3228
rect 12509 3194 12619 3228
rect 12653 3194 12683 3228
rect 12445 3108 12683 3194
rect 12445 3074 12475 3108
rect 12509 3074 12547 3108
rect 12581 3074 12619 3108
rect 12653 3074 12683 3108
rect 12445 3044 12683 3074
rect 12445 3028 12513 3044
rect 12445 2994 12475 3028
rect 12509 3010 12513 3028
rect 12547 3028 12581 3044
rect 12509 2994 12547 3010
rect 12615 3028 12683 3044
rect 12615 3010 12619 3028
rect 12581 2994 12619 3010
rect 12653 2994 12683 3028
rect 12445 2974 12683 2994
rect 12445 2948 12513 2974
rect 12445 2914 12475 2948
rect 12509 2940 12513 2948
rect 12547 2948 12581 2974
rect 12509 2914 12547 2940
rect 12615 2948 12683 2974
rect 12615 2940 12619 2948
rect 12581 2914 12619 2940
rect 12653 2914 12683 2948
rect 12445 2904 12683 2914
rect 12445 2870 12513 2904
rect 12547 2870 12581 2904
rect 12615 2870 12683 2904
rect 12445 2868 12683 2870
rect 12445 2834 12475 2868
rect 12509 2834 12547 2868
rect 12581 2834 12619 2868
rect 12653 2834 12683 2868
rect 12445 2800 12513 2834
rect 12547 2800 12581 2834
rect 12615 2800 12683 2834
rect 12445 2788 12683 2800
rect 12445 2754 12475 2788
rect 12509 2764 12547 2788
rect 12509 2754 12513 2764
rect 12445 2730 12513 2754
rect 12581 2764 12619 2788
rect 12547 2730 12581 2754
rect 12615 2754 12619 2764
rect 12653 2754 12683 2788
rect 12615 2730 12683 2754
rect 12445 2708 12683 2730
rect 12445 2674 12475 2708
rect 12509 2694 12547 2708
rect 12509 2674 12513 2694
rect 12445 2660 12513 2674
rect 12581 2694 12619 2708
rect 12547 2660 12581 2674
rect 12615 2674 12619 2694
rect 12653 2674 12683 2708
rect 12615 2660 12683 2674
rect 12445 2628 12683 2660
rect 12445 2594 12475 2628
rect 12509 2594 12547 2628
rect 12581 2594 12619 2628
rect 12653 2594 12683 2628
rect 12445 2518 12683 2594
rect 12445 2484 12475 2518
rect 12509 2484 12619 2518
rect 12653 2484 12683 2518
rect 12445 2446 12683 2484
rect 12445 2412 12475 2446
rect 12509 2412 12619 2446
rect 12653 2412 12683 2446
rect 12445 2374 12683 2412
rect 12445 2340 12475 2374
rect 12509 2340 12619 2374
rect 12653 2340 12683 2374
rect 12445 2302 12683 2340
rect 12445 2268 12475 2302
rect 12509 2268 12619 2302
rect 12653 2268 12683 2302
rect 12445 2230 12683 2268
rect 12445 2196 12475 2230
rect 12509 2196 12619 2230
rect 12653 2196 12683 2230
rect 12445 2158 12683 2196
rect 12445 2124 12475 2158
rect 12509 2124 12619 2158
rect 12653 2124 12683 2158
rect 12445 2086 12683 2124
rect 12445 2052 12475 2086
rect 12509 2052 12619 2086
rect 12653 2052 12683 2086
rect 12445 2014 12683 2052
rect 12445 1980 12475 2014
rect 12509 1980 12619 2014
rect 12653 1980 12683 2014
rect 12445 1942 12683 1980
rect 12445 1908 12475 1942
rect 12509 1908 12619 1942
rect 12653 1908 12683 1942
rect 12445 1870 12683 1908
rect 12445 1836 12475 1870
rect 12509 1836 12619 1870
rect 12653 1836 12683 1870
rect 12445 1798 12683 1836
rect 12445 1764 12475 1798
rect 12509 1764 12619 1798
rect 12653 1764 12683 1798
rect 12445 1726 12683 1764
rect 12445 1692 12475 1726
rect 12509 1692 12619 1726
rect 12653 1692 12683 1726
rect 12445 1654 12683 1692
rect 12445 1620 12475 1654
rect 12509 1620 12619 1654
rect 12653 1620 12683 1654
rect 12445 1536 12683 1620
rect 12785 3104 12905 4200
rect 13215 4308 13335 4324
rect 13215 4274 13258 4308
rect 13292 4274 13335 4308
rect 13215 4234 13335 4274
rect 13215 4200 13258 4234
rect 13292 4200 13335 4234
rect 12785 3070 12828 3104
rect 12862 3070 12905 3104
rect 12785 3026 12905 3070
rect 12785 2992 12828 3026
rect 12862 2992 12905 3026
rect 12785 2948 12905 2992
rect 12785 2914 12828 2948
rect 12862 2914 12905 2948
rect 12785 2870 12905 2914
rect 12785 2836 12828 2870
rect 12862 2836 12905 2870
rect 12785 2792 12905 2836
rect 12785 2758 12828 2792
rect 12862 2758 12905 2792
rect 12785 2713 12905 2758
rect 12785 2679 12828 2713
rect 12862 2679 12905 2713
rect 12785 2634 12905 2679
rect 12785 2600 12828 2634
rect 12862 2600 12905 2634
rect 12223 1470 12266 1504
rect 12300 1470 12343 1504
rect 12223 1430 12343 1470
rect 12223 1396 12266 1430
rect 12300 1396 12343 1430
rect 12223 1250 12343 1396
rect 12223 1144 12230 1250
rect 12336 1144 12343 1250
rect 12785 1504 12905 2600
rect 12970 4064 12971 4098
rect 13005 4064 13043 4098
rect 13077 4064 13115 4098
rect 13149 4064 13150 4098
rect 12970 4025 13150 4064
rect 12970 3991 12971 4025
rect 13005 3991 13043 4025
rect 13077 3991 13115 4025
rect 13149 3991 13150 4025
rect 12970 3952 13150 3991
rect 12970 3918 12971 3952
rect 13005 3918 13043 3952
rect 13077 3918 13115 3952
rect 13149 3918 13150 3952
rect 12970 3879 13150 3918
rect 12970 3845 12971 3879
rect 13005 3845 13043 3879
rect 13077 3845 13115 3879
rect 13149 3845 13150 3879
rect 12970 3806 13150 3845
rect 12970 3772 12971 3806
rect 13005 3772 13043 3806
rect 13077 3772 13115 3806
rect 13149 3772 13150 3806
rect 12970 3733 13150 3772
rect 12970 3699 12971 3733
rect 13005 3699 13043 3733
rect 13077 3699 13115 3733
rect 13149 3699 13150 3733
rect 12970 3660 13150 3699
rect 12970 3626 12971 3660
rect 13005 3626 13043 3660
rect 13077 3626 13115 3660
rect 13149 3626 13150 3660
rect 12970 3587 13150 3626
rect 12970 3553 12971 3587
rect 13005 3553 13043 3587
rect 13077 3553 13115 3587
rect 13149 3553 13150 3587
rect 12970 3514 13150 3553
rect 12970 3480 12971 3514
rect 13005 3480 13043 3514
rect 13077 3480 13115 3514
rect 13149 3480 13150 3514
rect 12970 3441 13150 3480
rect 12970 3407 12971 3441
rect 13005 3407 13043 3441
rect 13077 3407 13115 3441
rect 13149 3407 13150 3441
rect 12970 3368 13150 3407
rect 12970 3334 12971 3368
rect 13005 3334 13043 3368
rect 13077 3334 13115 3368
rect 13149 3334 13150 3368
rect 12970 3295 13150 3334
rect 12970 3261 12971 3295
rect 13005 3261 13043 3295
rect 13077 3261 13115 3295
rect 13149 3261 13150 3295
rect 12970 3222 13150 3261
rect 12970 3188 12971 3222
rect 13005 3188 13043 3222
rect 13077 3188 13115 3222
rect 13149 3188 13150 3222
rect 12970 3149 13150 3188
rect 12970 3115 12971 3149
rect 13005 3115 13043 3149
rect 13077 3115 13115 3149
rect 13149 3115 13150 3149
rect 12970 3076 13150 3115
rect 12970 3042 12971 3076
rect 13005 3042 13043 3076
rect 13077 3042 13115 3076
rect 13149 3042 13150 3076
rect 12970 3003 13150 3042
rect 12970 2969 12971 3003
rect 13005 2969 13043 3003
rect 13077 2969 13115 3003
rect 13149 2969 13150 3003
rect 12970 2930 13150 2969
rect 12970 2896 12971 2930
rect 13005 2896 13043 2930
rect 13077 2896 13115 2930
rect 13149 2896 13150 2930
rect 12970 2857 13150 2896
rect 12970 2823 12971 2857
rect 13005 2823 13043 2857
rect 13077 2823 13115 2857
rect 13149 2823 13150 2857
rect 12970 2784 13150 2823
rect 12970 2750 12971 2784
rect 13005 2750 13043 2784
rect 13077 2750 13115 2784
rect 13149 2750 13150 2784
rect 12970 2711 13150 2750
rect 12970 2677 12971 2711
rect 13005 2677 13043 2711
rect 13077 2677 13115 2711
rect 13149 2677 13150 2711
rect 12970 2638 13150 2677
rect 12970 2604 12971 2638
rect 13005 2604 13043 2638
rect 13077 2604 13115 2638
rect 13149 2604 13150 2638
rect 12970 2565 13150 2604
rect 12970 2531 12971 2565
rect 13005 2531 13043 2565
rect 13077 2531 13115 2565
rect 13149 2531 13150 2565
rect 12970 2492 13150 2531
rect 12970 2458 12971 2492
rect 13005 2458 13043 2492
rect 13077 2458 13115 2492
rect 13149 2458 13150 2492
rect 12970 2419 13150 2458
rect 12970 2385 12971 2419
rect 13005 2385 13043 2419
rect 13077 2385 13115 2419
rect 13149 2385 13150 2419
rect 12970 2346 13150 2385
rect 12970 2312 12971 2346
rect 13005 2312 13043 2346
rect 13077 2312 13115 2346
rect 13149 2312 13150 2346
rect 12970 2273 13150 2312
rect 12970 2239 12971 2273
rect 13005 2239 13043 2273
rect 13077 2239 13115 2273
rect 13149 2239 13150 2273
rect 12970 2200 13150 2239
rect 12970 2166 12971 2200
rect 13005 2166 13043 2200
rect 13077 2166 13115 2200
rect 13149 2166 13150 2200
rect 12970 2126 13150 2166
rect 12970 2092 12971 2126
rect 13005 2092 13043 2126
rect 13077 2092 13115 2126
rect 13149 2092 13150 2126
rect 12970 2052 13150 2092
rect 12970 2018 12971 2052
rect 13005 2018 13043 2052
rect 13077 2018 13115 2052
rect 13149 2018 13150 2052
rect 12970 1978 13150 2018
rect 12970 1944 12971 1978
rect 13005 1944 13043 1978
rect 13077 1944 13115 1978
rect 13149 1944 13150 1978
rect 12970 1904 13150 1944
rect 12970 1870 12971 1904
rect 13005 1870 13043 1904
rect 13077 1870 13115 1904
rect 13149 1870 13150 1904
rect 12970 1830 13150 1870
rect 12970 1796 12971 1830
rect 13005 1796 13043 1830
rect 13077 1796 13115 1830
rect 13149 1796 13150 1830
rect 12970 1756 13150 1796
rect 12970 1722 12971 1756
rect 13005 1722 13043 1756
rect 13077 1722 13115 1756
rect 13149 1722 13150 1756
rect 12970 1682 13150 1722
rect 12970 1648 12971 1682
rect 13005 1648 13043 1682
rect 13077 1648 13115 1682
rect 13149 1648 13150 1682
rect 12970 1608 13150 1648
rect 12970 1574 12971 1608
rect 13005 1574 13043 1608
rect 13077 1574 13115 1608
rect 13149 1574 13150 1608
rect 12970 1548 13150 1574
rect 13215 3104 13335 4200
rect 13777 4308 13897 4324
rect 13777 4274 13820 4308
rect 13854 4274 13897 4308
rect 13777 4234 13897 4274
rect 13777 4200 13820 4234
rect 13854 4200 13897 4234
rect 13215 3070 13258 3104
rect 13292 3070 13335 3104
rect 13215 3026 13335 3070
rect 13215 2992 13258 3026
rect 13292 2992 13335 3026
rect 13215 2948 13335 2992
rect 13215 2914 13258 2948
rect 13292 2914 13335 2948
rect 13215 2870 13335 2914
rect 13215 2836 13258 2870
rect 13292 2836 13335 2870
rect 13215 2792 13335 2836
rect 13215 2758 13258 2792
rect 13292 2758 13335 2792
rect 13215 2713 13335 2758
rect 13215 2679 13258 2713
rect 13292 2679 13335 2713
rect 13215 2634 13335 2679
rect 13215 2600 13258 2634
rect 13292 2600 13335 2634
rect 12785 1470 12828 1504
rect 12862 1470 12905 1504
rect 12785 1430 12905 1470
rect 12785 1396 12828 1430
rect 12862 1396 12905 1430
rect 12785 1250 12905 1396
rect 12785 1144 12792 1250
rect 12898 1144 12905 1250
rect 13215 1504 13335 2600
rect 13437 4092 13675 4110
rect 13437 4058 13467 4092
rect 13501 4058 13611 4092
rect 13645 4058 13675 4092
rect 13437 4020 13675 4058
rect 13437 3986 13467 4020
rect 13501 3986 13611 4020
rect 13645 3986 13675 4020
rect 13437 3948 13675 3986
rect 13437 3914 13467 3948
rect 13501 3914 13611 3948
rect 13645 3914 13675 3948
rect 13437 3876 13675 3914
rect 13437 3842 13467 3876
rect 13501 3842 13611 3876
rect 13645 3842 13675 3876
rect 13437 3804 13675 3842
rect 13437 3770 13467 3804
rect 13501 3770 13611 3804
rect 13645 3770 13675 3804
rect 13437 3732 13675 3770
rect 13437 3698 13467 3732
rect 13501 3698 13611 3732
rect 13645 3698 13675 3732
rect 13437 3660 13675 3698
rect 13437 3626 13467 3660
rect 13501 3626 13611 3660
rect 13645 3626 13675 3660
rect 13437 3588 13675 3626
rect 13437 3554 13467 3588
rect 13501 3554 13611 3588
rect 13645 3554 13675 3588
rect 13437 3516 13675 3554
rect 13437 3482 13467 3516
rect 13501 3482 13611 3516
rect 13645 3482 13675 3516
rect 13437 3444 13675 3482
rect 13437 3410 13467 3444
rect 13501 3410 13611 3444
rect 13645 3410 13675 3444
rect 13437 3372 13675 3410
rect 13437 3338 13467 3372
rect 13501 3338 13611 3372
rect 13645 3338 13675 3372
rect 13437 3300 13675 3338
rect 13437 3266 13467 3300
rect 13501 3266 13611 3300
rect 13645 3266 13675 3300
rect 13437 3228 13675 3266
rect 13437 3194 13467 3228
rect 13501 3194 13611 3228
rect 13645 3194 13675 3228
rect 13437 3108 13675 3194
rect 13437 3074 13467 3108
rect 13501 3074 13539 3108
rect 13573 3074 13611 3108
rect 13645 3074 13675 3108
rect 13437 3044 13675 3074
rect 13437 3028 13505 3044
rect 13437 2994 13467 3028
rect 13501 3010 13505 3028
rect 13539 3028 13573 3044
rect 13501 2994 13539 3010
rect 13607 3028 13675 3044
rect 13607 3010 13611 3028
rect 13573 2994 13611 3010
rect 13645 2994 13675 3028
rect 13437 2974 13675 2994
rect 13437 2948 13505 2974
rect 13437 2914 13467 2948
rect 13501 2940 13505 2948
rect 13539 2948 13573 2974
rect 13501 2914 13539 2940
rect 13607 2948 13675 2974
rect 13607 2940 13611 2948
rect 13573 2914 13611 2940
rect 13645 2914 13675 2948
rect 13437 2904 13675 2914
rect 13437 2870 13505 2904
rect 13539 2870 13573 2904
rect 13607 2870 13675 2904
rect 13437 2868 13675 2870
rect 13437 2834 13467 2868
rect 13501 2834 13539 2868
rect 13573 2834 13611 2868
rect 13645 2834 13675 2868
rect 13437 2800 13505 2834
rect 13539 2800 13573 2834
rect 13607 2800 13675 2834
rect 13437 2788 13675 2800
rect 13437 2754 13467 2788
rect 13501 2764 13539 2788
rect 13501 2754 13505 2764
rect 13437 2730 13505 2754
rect 13573 2764 13611 2788
rect 13539 2730 13573 2754
rect 13607 2754 13611 2764
rect 13645 2754 13675 2788
rect 13607 2730 13675 2754
rect 13437 2708 13675 2730
rect 13437 2674 13467 2708
rect 13501 2694 13539 2708
rect 13501 2674 13505 2694
rect 13437 2660 13505 2674
rect 13573 2694 13611 2708
rect 13539 2660 13573 2674
rect 13607 2674 13611 2694
rect 13645 2674 13675 2708
rect 13607 2660 13675 2674
rect 13437 2628 13675 2660
rect 13437 2594 13467 2628
rect 13501 2594 13539 2628
rect 13573 2594 13611 2628
rect 13645 2594 13675 2628
rect 13437 2518 13675 2594
rect 13437 2484 13467 2518
rect 13501 2484 13611 2518
rect 13645 2484 13675 2518
rect 13437 2446 13675 2484
rect 13437 2412 13467 2446
rect 13501 2412 13611 2446
rect 13645 2412 13675 2446
rect 13437 2374 13675 2412
rect 13437 2340 13467 2374
rect 13501 2340 13611 2374
rect 13645 2340 13675 2374
rect 13437 2302 13675 2340
rect 13437 2268 13467 2302
rect 13501 2268 13611 2302
rect 13645 2268 13675 2302
rect 13437 2230 13675 2268
rect 13437 2196 13467 2230
rect 13501 2196 13611 2230
rect 13645 2196 13675 2230
rect 13437 2158 13675 2196
rect 13437 2124 13467 2158
rect 13501 2124 13611 2158
rect 13645 2124 13675 2158
rect 13437 2086 13675 2124
rect 13437 2052 13467 2086
rect 13501 2052 13611 2086
rect 13645 2052 13675 2086
rect 13437 2014 13675 2052
rect 13437 1980 13467 2014
rect 13501 1980 13611 2014
rect 13645 1980 13675 2014
rect 13437 1942 13675 1980
rect 13437 1908 13467 1942
rect 13501 1908 13611 1942
rect 13645 1908 13675 1942
rect 13437 1870 13675 1908
rect 13437 1836 13467 1870
rect 13501 1836 13611 1870
rect 13645 1836 13675 1870
rect 13437 1798 13675 1836
rect 13437 1764 13467 1798
rect 13501 1764 13611 1798
rect 13645 1764 13675 1798
rect 13437 1726 13675 1764
rect 13437 1692 13467 1726
rect 13501 1692 13611 1726
rect 13645 1692 13675 1726
rect 13437 1654 13675 1692
rect 13437 1620 13467 1654
rect 13501 1620 13611 1654
rect 13645 1620 13675 1654
rect 13437 1536 13675 1620
rect 13777 3104 13897 4200
rect 14135 4308 14255 4324
rect 14135 4274 14178 4308
rect 14212 4274 14255 4308
rect 14135 4234 14255 4274
rect 14135 4200 14178 4234
rect 14212 4200 14255 4234
rect 13777 3070 13820 3104
rect 13854 3070 13897 3104
rect 13777 3026 13897 3070
rect 13777 2992 13820 3026
rect 13854 2992 13897 3026
rect 13777 2948 13897 2992
rect 13777 2914 13820 2948
rect 13854 2914 13897 2948
rect 13777 2870 13897 2914
rect 13777 2836 13820 2870
rect 13854 2836 13897 2870
rect 13777 2792 13897 2836
rect 13777 2758 13820 2792
rect 13854 2758 13897 2792
rect 13777 2713 13897 2758
rect 13777 2679 13820 2713
rect 13854 2679 13897 2713
rect 13777 2634 13897 2679
rect 13777 2600 13820 2634
rect 13854 2600 13897 2634
rect 13215 1470 13258 1504
rect 13292 1470 13335 1504
rect 13215 1430 13335 1470
rect 13215 1396 13258 1430
rect 13292 1396 13335 1430
rect 13215 1250 13335 1396
rect 13215 1144 13222 1250
rect 13328 1144 13335 1250
rect 13777 1504 13897 2600
rect 13999 4025 14033 4064
rect 13999 3952 14033 3991
rect 13999 3879 14033 3918
rect 13999 3806 14033 3845
rect 13999 3733 14033 3772
rect 13999 3660 14033 3699
rect 13999 3587 14033 3626
rect 13999 3514 14033 3553
rect 13999 3441 14033 3480
rect 13999 3368 14033 3407
rect 13999 3295 14033 3334
rect 13999 3222 14033 3261
rect 13999 3149 14033 3188
rect 13999 3076 14033 3115
rect 13999 3003 14033 3042
rect 13999 2930 14033 2969
rect 13999 2857 14033 2896
rect 13999 2784 14033 2823
rect 13999 2711 14033 2750
rect 13999 2638 14033 2677
rect 13999 2565 14033 2604
rect 13999 2492 14033 2531
rect 13999 2419 14033 2458
rect 13999 2346 14033 2385
rect 13999 2273 14033 2312
rect 13999 2200 14033 2239
rect 13999 2126 14033 2166
rect 13999 2052 14033 2092
rect 13999 1978 14033 2018
rect 13999 1904 14033 1944
rect 13999 1830 14033 1870
rect 13999 1756 14033 1796
rect 13999 1682 14033 1722
rect 13999 1608 14033 1648
rect 14135 3104 14255 4200
rect 14135 3070 14178 3104
rect 14212 3070 14255 3104
rect 14135 3026 14255 3070
rect 14135 2992 14178 3026
rect 14212 2992 14255 3026
rect 14135 2948 14255 2992
rect 14135 2914 14178 2948
rect 14212 2914 14255 2948
rect 14135 2870 14255 2914
rect 14135 2836 14178 2870
rect 14212 2836 14255 2870
rect 14135 2792 14255 2836
rect 14135 2758 14178 2792
rect 14212 2758 14255 2792
rect 14135 2713 14255 2758
rect 14135 2679 14178 2713
rect 14212 2679 14255 2713
rect 14135 2634 14255 2679
rect 14135 2600 14178 2634
rect 14212 2600 14255 2634
rect 13777 1470 13820 1504
rect 13854 1470 13897 1504
rect 13777 1430 13897 1470
rect 13777 1396 13820 1430
rect 13854 1396 13897 1430
rect 13777 1250 13897 1396
rect 13777 1144 13784 1250
rect 13890 1144 13897 1250
rect 14135 1504 14255 2600
rect 14135 1470 14178 1504
rect 14212 1470 14255 1504
rect 14135 1430 14255 1470
rect 14135 1396 14178 1430
rect 14212 1396 14255 1430
rect 14135 1250 14255 1396
rect 14135 1144 14142 1250
rect 14248 1144 14255 1250
rect 14356 4286 14428 4325
rect 14390 4252 14428 4286
rect 14356 4213 14428 4252
rect 14390 4179 14428 4213
rect 14356 4140 14428 4179
rect 14390 4106 14428 4140
rect 14356 4067 14428 4106
rect 14390 4033 14428 4067
rect 14356 3994 14428 4033
rect 14390 3960 14428 3994
rect 14356 3957 14536 3960
rect 14356 3952 14468 3957
rect 14356 3921 14428 3952
rect 14390 3918 14428 3921
rect 14462 3923 14468 3952
rect 14502 3924 14536 3957
rect 14502 3923 14604 3924
rect 14462 3921 14604 3923
rect 14462 3918 14500 3921
rect 14390 3888 14500 3918
rect 14534 3889 14572 3921
rect 14638 3905 14653 4551
rect 14390 3887 14468 3888
rect 14534 3887 14536 3889
rect 14356 3880 14468 3887
rect 14356 3848 14428 3880
rect 14390 3846 14428 3848
rect 14462 3854 14468 3880
rect 14502 3855 14536 3887
rect 14570 3887 14572 3889
rect 14606 3887 14653 3905
rect 14570 3871 14653 3887
rect 14570 3855 14604 3871
rect 14502 3854 14604 3855
rect 14462 3848 14604 3854
rect 14462 3846 14500 3848
rect 14390 3819 14500 3846
rect 14534 3820 14572 3848
rect 14638 3837 14653 3871
rect 14390 3814 14468 3819
rect 14534 3814 14536 3820
rect 14356 3808 14468 3814
rect 14356 3775 14428 3808
rect 14390 3774 14428 3775
rect 14462 3785 14468 3808
rect 14502 3786 14536 3814
rect 14570 3814 14572 3820
rect 14606 3814 14653 3837
rect 14570 3803 14653 3814
rect 14570 3786 14604 3803
rect 14502 3785 14604 3786
rect 14462 3775 14604 3785
rect 14462 3774 14500 3775
rect 14390 3750 14500 3774
rect 14534 3751 14572 3775
rect 14638 3769 14653 3803
rect 14390 3741 14468 3750
rect 14534 3741 14536 3751
rect 14356 3736 14468 3741
rect 14356 3702 14428 3736
rect 14462 3716 14468 3736
rect 14502 3717 14536 3741
rect 14570 3741 14572 3751
rect 14606 3741 14653 3769
rect 14570 3735 14653 3741
rect 14570 3717 14604 3735
rect 14502 3716 14604 3717
rect 14462 3702 14604 3716
rect 14390 3681 14500 3702
rect 14534 3682 14572 3702
rect 14638 3701 14653 3735
rect 14390 3668 14468 3681
rect 14534 3668 14536 3682
rect 14356 3664 14468 3668
rect 14356 3630 14428 3664
rect 14462 3647 14468 3664
rect 14502 3648 14536 3668
rect 14570 3668 14572 3682
rect 14606 3668 14653 3701
rect 14570 3667 14653 3668
rect 14570 3648 14604 3667
rect 14502 3647 14604 3648
rect 14462 3633 14604 3647
rect 14638 3633 14653 3667
rect 14462 3630 14653 3633
rect 14356 3629 14653 3630
rect 14390 3612 14500 3629
rect 14534 3613 14572 3629
rect 14390 3595 14468 3612
rect 14534 3595 14536 3613
rect 14356 3592 14468 3595
rect 14356 3558 14428 3592
rect 14462 3578 14468 3592
rect 14502 3579 14536 3595
rect 14570 3595 14572 3613
rect 14606 3599 14653 3629
rect 14570 3579 14604 3595
rect 14502 3578 14604 3579
rect 14462 3565 14604 3578
rect 14638 3565 14653 3599
rect 14462 3558 14653 3565
rect 14356 3556 14653 3558
rect 14390 3543 14500 3556
rect 14534 3544 14572 3556
rect 14390 3522 14468 3543
rect 14534 3522 14536 3544
rect 14356 3520 14468 3522
rect 14356 3486 14428 3520
rect 14462 3509 14468 3520
rect 14502 3510 14536 3522
rect 14570 3522 14572 3544
rect 14606 3531 14653 3556
rect 14570 3510 14604 3522
rect 14502 3509 14604 3510
rect 14462 3497 14604 3509
rect 14638 3497 14653 3531
rect 14462 3486 14653 3497
rect 14356 3483 14653 3486
rect 14390 3474 14500 3483
rect 14534 3475 14572 3483
rect 14390 3449 14468 3474
rect 14534 3449 14536 3475
rect 14356 3448 14468 3449
rect 14356 3414 14428 3448
rect 14462 3440 14468 3448
rect 14502 3441 14536 3449
rect 14570 3449 14572 3475
rect 14606 3463 14653 3483
rect 14570 3441 14604 3449
rect 14502 3440 14604 3441
rect 14462 3429 14604 3440
rect 14638 3429 14653 3463
rect 14462 3414 14653 3429
rect 14356 3410 14653 3414
rect 14390 3405 14500 3410
rect 14534 3406 14572 3410
rect 14390 3376 14468 3405
rect 14534 3376 14536 3406
rect 14356 3342 14428 3376
rect 14462 3371 14468 3376
rect 14502 3372 14536 3376
rect 14570 3376 14572 3406
rect 14606 3395 14653 3410
rect 14570 3372 14604 3376
rect 14502 3371 14604 3372
rect 14462 3361 14604 3371
rect 14638 3361 14653 3395
rect 14462 3342 14653 3361
rect 14356 3337 14653 3342
rect 14390 3336 14500 3337
rect 14390 3304 14468 3336
rect 14390 3303 14428 3304
rect 14356 3270 14428 3303
rect 14462 3302 14468 3304
rect 14534 3303 14536 3337
rect 14570 3303 14572 3337
rect 14606 3327 14653 3337
rect 14502 3302 14604 3303
rect 14462 3293 14604 3302
rect 14638 3293 14653 3327
rect 14462 3270 14653 3293
rect 14356 3268 14653 3270
rect 14356 3267 14536 3268
rect 14356 3264 14468 3267
rect 14502 3264 14536 3267
rect 14390 3233 14468 3264
rect 14534 3234 14536 3264
rect 14570 3264 14653 3268
rect 14570 3234 14572 3264
rect 14606 3259 14653 3264
rect 14390 3232 14500 3233
rect 14390 3230 14428 3232
rect 14356 3198 14428 3230
rect 14462 3230 14500 3232
rect 14534 3230 14572 3234
rect 14462 3225 14604 3230
rect 14638 3225 14653 3259
rect 14462 3199 14653 3225
rect 14462 3198 14536 3199
rect 14356 3191 14468 3198
rect 14502 3191 14536 3198
rect 14390 3164 14468 3191
rect 14534 3165 14536 3191
rect 14570 3191 14653 3199
rect 14570 3165 14572 3191
rect 14390 3160 14500 3164
rect 14390 3157 14428 3160
rect 14356 3126 14428 3157
rect 14462 3157 14500 3160
rect 14534 3157 14572 3165
rect 14638 3157 14653 3191
rect 14462 3130 14653 3157
rect 14462 3129 14536 3130
rect 14462 3126 14468 3129
rect 14356 3118 14468 3126
rect 14502 3118 14536 3129
rect 14390 3095 14468 3118
rect 14534 3096 14536 3118
rect 14570 3123 14653 3130
rect 14570 3118 14604 3123
rect 14570 3096 14572 3118
rect 14390 3088 14500 3095
rect 14390 3084 14428 3088
rect 14356 3054 14428 3084
rect 14462 3084 14500 3088
rect 14534 3084 14572 3096
rect 14638 3089 14653 3123
rect 14606 3084 14653 3089
rect 14462 3061 14653 3084
rect 14462 3060 14536 3061
rect 14462 3054 14468 3060
rect 14356 3045 14468 3054
rect 14502 3045 14536 3060
rect 14390 3026 14468 3045
rect 14534 3027 14536 3045
rect 14570 3055 14653 3061
rect 14570 3045 14604 3055
rect 14570 3027 14572 3045
rect 14390 3016 14500 3026
rect 14390 3011 14428 3016
rect 14356 2982 14428 3011
rect 14462 3011 14500 3016
rect 14534 3011 14572 3027
rect 14638 3021 14653 3055
rect 14606 3011 14653 3021
rect 14462 2992 14653 3011
rect 14462 2991 14536 2992
rect 14462 2982 14468 2991
rect 14356 2972 14468 2982
rect 14502 2972 14536 2991
rect 14390 2957 14468 2972
rect 14534 2958 14536 2972
rect 14570 2987 14653 2992
rect 14570 2972 14604 2987
rect 14570 2958 14572 2972
rect 14390 2944 14500 2957
rect 14390 2938 14428 2944
rect 14356 2910 14428 2938
rect 14462 2938 14500 2944
rect 14534 2938 14572 2958
rect 14638 2953 14653 2987
rect 14606 2938 14653 2953
rect 14462 2923 14653 2938
rect 14462 2922 14536 2923
rect 14462 2910 14468 2922
rect 14356 2899 14468 2910
rect 14502 2899 14536 2922
rect 14390 2888 14468 2899
rect 14534 2889 14536 2899
rect 14570 2919 14653 2923
rect 14570 2899 14604 2919
rect 14570 2889 14572 2899
rect 14390 2872 14500 2888
rect 14390 2865 14428 2872
rect 14356 2838 14428 2865
rect 14462 2865 14500 2872
rect 14534 2865 14572 2889
rect 14638 2885 14653 2919
rect 14606 2865 14653 2885
rect 14462 2854 14653 2865
rect 14462 2853 14536 2854
rect 14462 2838 14468 2853
rect 14356 2826 14468 2838
rect 14502 2826 14536 2853
rect 14390 2819 14468 2826
rect 14534 2820 14536 2826
rect 14570 2851 14653 2854
rect 14570 2826 14604 2851
rect 14570 2820 14572 2826
rect 14390 2800 14500 2819
rect 14390 2792 14428 2800
rect 14356 2766 14428 2792
rect 14462 2792 14500 2800
rect 14534 2792 14572 2820
rect 14638 2817 14653 2851
rect 14606 2792 14653 2817
rect 14462 2785 14653 2792
rect 14462 2784 14536 2785
rect 14462 2766 14468 2784
rect 14356 2753 14468 2766
rect 14502 2753 14536 2784
rect 14390 2750 14468 2753
rect 14534 2751 14536 2753
rect 14570 2783 14653 2785
rect 14570 2753 14604 2783
rect 14570 2751 14572 2753
rect 14390 2728 14500 2750
rect 14390 2719 14428 2728
rect 14356 2694 14428 2719
rect 14462 2719 14500 2728
rect 14534 2719 14572 2751
rect 14638 2749 14653 2783
rect 14606 2719 14653 2749
rect 14462 2716 14653 2719
rect 14462 2715 14536 2716
rect 14462 2694 14468 2715
rect 14356 2681 14468 2694
rect 14502 2682 14536 2715
rect 14570 2715 14653 2716
rect 14570 2682 14604 2715
rect 14502 2681 14604 2682
rect 14638 2681 14653 2715
rect 14356 2680 14653 2681
rect 14390 2656 14500 2680
rect 14390 2646 14428 2656
rect 14356 2622 14428 2646
rect 14462 2646 14500 2656
rect 14534 2647 14572 2680
rect 14606 2647 14653 2680
rect 14534 2646 14536 2647
rect 14462 2622 14468 2646
rect 14356 2612 14468 2622
rect 14502 2613 14536 2646
rect 14570 2646 14572 2647
rect 14570 2613 14604 2646
rect 14638 2613 14653 2647
rect 14502 2612 14653 2613
rect 14356 2607 14653 2612
rect 14390 2584 14500 2607
rect 14390 2573 14428 2584
rect 14356 2550 14428 2573
rect 14462 2577 14500 2584
rect 14534 2578 14572 2607
rect 14606 2579 14653 2607
rect 14462 2550 14468 2577
rect 14534 2573 14536 2578
rect 14356 2543 14468 2550
rect 14502 2544 14536 2573
rect 14570 2573 14572 2578
rect 14570 2545 14604 2573
rect 14638 2545 14653 2579
rect 14570 2544 14653 2545
rect 14502 2543 14653 2544
rect 14356 2534 14653 2543
rect 14390 2512 14500 2534
rect 14390 2500 14428 2512
rect 14356 2478 14428 2500
rect 14462 2508 14500 2512
rect 14534 2509 14572 2534
rect 14606 2511 14653 2534
rect 14462 2478 14468 2508
rect 14534 2500 14536 2509
rect 14356 2474 14468 2478
rect 14502 2475 14536 2500
rect 14570 2500 14572 2509
rect 14570 2477 14604 2500
rect 14638 2477 14653 2511
rect 14570 2475 14653 2477
rect 14502 2474 14653 2475
rect 14356 2461 14653 2474
rect 14390 2440 14500 2461
rect 14390 2427 14428 2440
rect 14356 2406 14428 2427
rect 14462 2439 14500 2440
rect 14534 2440 14572 2461
rect 14606 2443 14653 2461
rect 14462 2406 14468 2439
rect 14534 2427 14536 2440
rect 14356 2405 14468 2406
rect 14502 2406 14536 2427
rect 14570 2427 14572 2440
rect 14570 2409 14604 2427
rect 14638 2409 14653 2443
rect 14570 2406 14653 2409
rect 14502 2405 14653 2406
rect 14356 2388 14653 2405
rect 14390 2370 14500 2388
rect 14534 2371 14572 2388
rect 14606 2375 14653 2388
rect 14390 2368 14468 2370
rect 14390 2354 14428 2368
rect 14356 2334 14428 2354
rect 14462 2336 14468 2368
rect 14534 2354 14536 2371
rect 14502 2337 14536 2354
rect 14570 2354 14572 2371
rect 14570 2341 14604 2354
rect 14638 2341 14653 2375
rect 14570 2337 14653 2341
rect 14502 2336 14653 2337
rect 14462 2334 14653 2336
rect 14356 2315 14653 2334
rect 14390 2301 14500 2315
rect 14534 2302 14572 2315
rect 14606 2307 14653 2315
rect 14390 2296 14468 2301
rect 14390 2281 14428 2296
rect 14356 2262 14428 2281
rect 14462 2267 14468 2296
rect 14534 2281 14536 2302
rect 14502 2268 14536 2281
rect 14570 2281 14572 2302
rect 14570 2273 14604 2281
rect 14638 2273 14653 2307
rect 14570 2268 14653 2273
rect 14502 2267 14653 2268
rect 14462 2262 14653 2267
rect 14356 2242 14653 2262
rect 14390 2232 14500 2242
rect 14534 2233 14572 2242
rect 14606 2239 14653 2242
rect 14390 2224 14468 2232
rect 14390 2208 14428 2224
rect 14356 2190 14428 2208
rect 14462 2198 14468 2224
rect 14534 2208 14536 2233
rect 14502 2199 14536 2208
rect 14570 2208 14572 2233
rect 14570 2205 14604 2208
rect 14638 2205 14653 2239
rect 14570 2199 14653 2205
rect 14502 2198 14653 2199
rect 14462 2190 14653 2198
rect 14356 2171 14653 2190
rect 14356 2169 14604 2171
rect 14390 2163 14500 2169
rect 14534 2164 14572 2169
rect 14390 2152 14468 2163
rect 14390 2135 14428 2152
rect 14356 2118 14428 2135
rect 14462 2129 14468 2152
rect 14534 2135 14536 2164
rect 14502 2130 14536 2135
rect 14570 2135 14572 2164
rect 14638 2137 14653 2171
rect 14606 2135 14653 2137
rect 14570 2130 14653 2135
rect 14502 2129 14653 2130
rect 14462 2118 14653 2129
rect 14356 2103 14653 2118
rect 14356 2096 14604 2103
rect 14390 2094 14500 2096
rect 14534 2095 14572 2096
rect 14390 2080 14468 2094
rect 14390 2062 14428 2080
rect 14356 2046 14428 2062
rect 14462 2060 14468 2080
rect 14534 2062 14536 2095
rect 14502 2061 14536 2062
rect 14570 2062 14572 2095
rect 14638 2069 14653 2103
rect 14606 2062 14653 2069
rect 14570 2061 14653 2062
rect 14502 2060 14653 2061
rect 14462 2046 14653 2060
rect 14356 2035 14653 2046
rect 14356 2026 14604 2035
rect 14356 2025 14536 2026
rect 14356 2023 14468 2025
rect 14502 2023 14536 2025
rect 14390 2008 14468 2023
rect 14390 1989 14428 2008
rect 14356 1974 14428 1989
rect 14462 1991 14468 2008
rect 14534 1992 14536 2023
rect 14570 2023 14604 2026
rect 14570 1992 14572 2023
rect 14638 2001 14653 2035
rect 14462 1989 14500 1991
rect 14534 1989 14572 1992
rect 14606 1989 14653 2001
rect 14462 1974 14653 1989
rect 14356 1967 14653 1974
rect 14356 1957 14604 1967
rect 14356 1956 14536 1957
rect 14356 1950 14468 1956
rect 14502 1950 14536 1956
rect 14390 1936 14468 1950
rect 14390 1916 14428 1936
rect 14356 1902 14428 1916
rect 14462 1922 14468 1936
rect 14534 1923 14536 1950
rect 14570 1950 14604 1957
rect 14570 1923 14572 1950
rect 14638 1933 14653 1967
rect 14462 1916 14500 1922
rect 14534 1916 14572 1923
rect 14606 1916 14653 1933
rect 14462 1902 14653 1916
rect 14356 1899 14653 1902
rect 14356 1888 14604 1899
rect 14356 1887 14536 1888
rect 14356 1877 14468 1887
rect 14502 1877 14536 1887
rect 14390 1864 14468 1877
rect 14390 1843 14428 1864
rect 14356 1830 14428 1843
rect 14462 1853 14468 1864
rect 14534 1854 14536 1877
rect 14570 1877 14604 1888
rect 14570 1854 14572 1877
rect 14638 1865 14653 1899
rect 14462 1843 14500 1853
rect 14534 1843 14572 1854
rect 14606 1843 14653 1865
rect 14462 1831 14653 1843
rect 14462 1830 14604 1831
rect 14356 1819 14604 1830
rect 14356 1818 14536 1819
rect 14356 1804 14468 1818
rect 14502 1804 14536 1818
rect 14390 1792 14468 1804
rect 14390 1770 14428 1792
rect 14356 1758 14428 1770
rect 14462 1784 14468 1792
rect 14534 1785 14536 1804
rect 14570 1804 14604 1819
rect 14570 1785 14572 1804
rect 14638 1797 14653 1831
rect 14462 1770 14500 1784
rect 14534 1770 14572 1785
rect 14606 1770 14653 1797
rect 14462 1763 14653 1770
rect 14462 1758 14604 1763
rect 14356 1750 14604 1758
rect 14356 1749 14536 1750
rect 14356 1731 14468 1749
rect 14502 1731 14536 1749
rect 14390 1720 14468 1731
rect 14390 1697 14428 1720
rect 14356 1686 14428 1697
rect 14462 1715 14468 1720
rect 14534 1716 14536 1731
rect 14570 1731 14604 1750
rect 14570 1716 14572 1731
rect 14638 1729 14653 1763
rect 14462 1697 14500 1715
rect 14534 1697 14572 1716
rect 14606 1697 14653 1729
rect 14462 1695 14653 1697
rect 14462 1686 14604 1695
rect 14356 1681 14604 1686
rect 14356 1680 14536 1681
rect 14356 1657 14468 1680
rect 14502 1658 14536 1680
rect 14390 1648 14468 1657
rect 14390 1623 14428 1648
rect 14356 1614 14428 1623
rect 14462 1646 14468 1648
rect 14534 1647 14536 1658
rect 14570 1661 14604 1681
rect 14638 1661 14653 1695
rect 14570 1658 14653 1661
rect 14570 1647 14572 1658
rect 14462 1624 14500 1646
rect 14534 1624 14572 1647
rect 14606 1627 14653 1658
rect 14462 1614 14604 1624
rect 14356 1612 14604 1614
rect 14356 1611 14536 1612
rect 14356 1583 14468 1611
rect 14502 1585 14536 1611
rect 14390 1577 14468 1583
rect 14534 1578 14536 1585
rect 14570 1593 14604 1612
rect 14638 1593 14653 1627
rect 14570 1585 14653 1593
rect 14570 1578 14572 1585
rect 14390 1576 14500 1577
rect 14390 1549 14428 1576
rect 14356 1542 14428 1549
rect 14462 1551 14500 1576
rect 14534 1551 14572 1578
rect 14606 1559 14653 1585
rect 14462 1543 14604 1551
rect 14462 1542 14536 1543
rect 14356 1509 14468 1542
rect 14502 1512 14536 1542
rect 14390 1508 14468 1509
rect 14534 1509 14536 1512
rect 14570 1525 14604 1543
rect 14638 1525 14653 1559
rect 14570 1512 14653 1525
rect 14570 1509 14572 1512
rect 14390 1504 14500 1508
rect 14390 1475 14428 1504
rect 14356 1470 14428 1475
rect 14462 1478 14500 1504
rect 14534 1478 14572 1509
rect 14606 1491 14653 1512
rect 14462 1474 14604 1478
rect 14462 1473 14536 1474
rect 14462 1470 14468 1473
rect 14356 1439 14468 1470
rect 14502 1440 14536 1473
rect 14570 1457 14604 1474
rect 14638 1457 14653 1491
rect 14570 1440 14653 1457
rect 14502 1439 14653 1440
rect 14356 1435 14500 1439
rect 14390 1432 14500 1435
rect 14390 1401 14428 1432
rect 14356 1398 14428 1401
rect 14462 1405 14500 1432
rect 14534 1405 14572 1439
rect 14606 1423 14653 1439
rect 14462 1404 14536 1405
rect 14462 1398 14468 1404
rect 14356 1370 14468 1398
rect 14502 1371 14536 1404
rect 14570 1389 14604 1405
rect 14638 1389 14653 1423
rect 14570 1371 14653 1389
rect 14502 1370 14653 1371
rect 14356 1366 14653 1370
rect 14356 1361 14500 1366
rect 14390 1360 14500 1361
rect 14390 1327 14428 1360
rect 14356 1326 14428 1327
rect 14462 1335 14500 1360
rect 14534 1336 14572 1366
rect 14606 1355 14653 1366
rect 14462 1326 14468 1335
rect 14534 1332 14536 1336
rect 14356 1301 14468 1326
rect 14502 1302 14536 1332
rect 14570 1332 14572 1336
rect 14570 1321 14604 1332
rect 14638 1321 14653 1355
rect 14570 1302 14653 1321
rect 14502 1301 14653 1302
rect 14356 1293 14653 1301
rect 14356 1288 14500 1293
rect 14356 1287 14428 1288
rect 14390 1254 14428 1287
rect 14462 1266 14500 1288
rect 14534 1267 14572 1293
rect 14606 1287 14653 1293
rect 14462 1254 14468 1266
rect 14534 1259 14536 1267
rect 14390 1253 14468 1254
rect 14356 1232 14468 1253
rect 14502 1233 14536 1259
rect 14570 1259 14572 1267
rect 14570 1253 14604 1259
rect 14638 1253 14653 1287
rect 14570 1233 14653 1253
rect 14502 1232 14653 1233
rect 14356 1220 14653 1232
rect 14356 1216 14500 1220
rect 14356 1213 14428 1216
rect 14390 1182 14428 1213
rect 14462 1197 14500 1216
rect 14534 1198 14572 1220
rect 14606 1218 14653 1220
rect 14462 1182 14468 1197
rect 14534 1186 14536 1198
rect 14390 1179 14468 1182
rect 14356 1163 14468 1179
rect 14502 1164 14536 1186
rect 14570 1186 14572 1198
rect 14570 1184 14604 1186
rect 14638 1184 14653 1218
rect 14570 1164 14653 1184
rect 14502 1163 14653 1164
rect 14356 1149 14653 1163
rect 14356 1147 14604 1149
rect 14356 1144 14500 1147
rect 667 883 746 894
rect 667 867 780 883
rect 14356 1139 14428 1144
rect 14390 1110 14428 1139
rect 14462 1128 14500 1144
rect 14534 1129 14572 1147
rect 14462 1110 14468 1128
rect 14534 1113 14536 1129
rect 14390 1105 14468 1110
rect 14356 1094 14468 1105
rect 14502 1095 14536 1113
rect 14570 1113 14572 1129
rect 14638 1115 14653 1149
rect 14606 1113 14653 1115
rect 14570 1095 14653 1113
rect 14502 1094 14653 1095
rect 14356 1080 14653 1094
rect 14356 1074 14604 1080
rect 14356 1072 14500 1074
rect 14356 1065 14428 1072
rect 14390 1038 14428 1065
rect 14462 1059 14500 1072
rect 14534 1060 14572 1074
rect 14462 1038 14468 1059
rect 14534 1040 14536 1060
rect 14390 1031 14468 1038
rect 14356 1025 14468 1031
rect 14502 1026 14536 1040
rect 14570 1040 14572 1060
rect 14638 1046 14653 1080
rect 14606 1040 14653 1046
rect 14570 1026 14653 1040
rect 14502 1025 14653 1026
rect 14356 1011 14653 1025
rect 14356 1001 14604 1011
rect 14356 1000 14500 1001
rect 14356 991 14428 1000
rect 14390 966 14428 991
rect 14462 990 14500 1000
rect 14534 991 14572 1001
rect 14462 966 14468 990
rect 14534 967 14536 991
rect 14390 957 14468 966
rect 14356 956 14468 957
rect 14502 957 14536 967
rect 14570 967 14572 991
rect 14638 977 14653 1011
rect 14606 967 14653 977
rect 14570 957 14653 967
rect 14502 956 14653 957
rect 14356 942 14653 956
rect 14356 928 14604 942
rect 14356 917 14428 928
rect 14390 894 14428 917
rect 14462 921 14500 928
rect 14534 922 14572 928
rect 14462 894 14468 921
rect 14534 894 14536 922
rect 14390 887 14468 894
rect 14502 888 14536 894
rect 14570 894 14572 922
rect 14638 908 14653 942
rect 14606 894 14653 908
rect 14570 888 14653 894
rect 14502 887 14653 888
rect 14390 883 14653 887
rect 14356 873 14653 883
rect 14356 867 14604 873
rect 667 853 14604 867
rect 667 852 14536 853
rect 667 818 702 852
rect 736 820 771 852
rect 805 820 840 852
rect 874 820 909 852
rect 943 820 978 852
rect 1012 820 1047 852
rect 1081 820 1116 852
rect 1150 820 1185 852
rect 1219 820 1254 852
rect 1288 820 1323 852
rect 1357 820 1392 852
rect 1426 820 1461 852
rect 1495 820 1530 852
rect 1564 820 1599 852
rect 1633 820 1668 852
rect 1702 820 1737 852
rect 1771 820 1806 852
rect 1840 820 1875 852
rect 1909 820 1944 852
rect 1978 820 2013 852
rect 2047 820 2082 852
rect 2116 820 2151 852
rect 2185 820 2220 852
rect 2254 820 2289 852
rect 2323 820 2358 852
rect 2392 820 2427 852
rect 2461 820 2496 852
rect 2530 820 2565 852
rect 2599 820 2634 852
rect 2668 820 2703 852
rect 2737 820 2772 852
rect 743 818 771 820
rect 816 818 840 820
rect 889 818 909 820
rect 599 786 709 818
rect 743 786 782 818
rect 816 786 855 818
rect 889 786 928 818
rect 599 784 928 786
rect 482 750 565 769
rect 599 750 634 784
rect 668 750 703 784
rect 737 750 772 784
rect 806 750 841 784
rect 875 750 910 784
rect 14502 819 14536 852
rect 14570 839 14604 853
rect 14638 839 14653 873
rect 14570 819 14653 839
rect 14502 804 14653 819
rect 14502 784 14604 804
rect 14570 770 14604 784
rect 14638 770 14653 804
rect 14570 750 14653 770
rect 482 748 928 750
rect 482 716 709 748
rect 743 716 782 748
rect 816 716 855 748
rect 889 716 928 748
rect 482 682 516 716
rect 550 682 585 716
rect 619 682 654 716
rect 688 714 709 716
rect 757 714 782 716
rect 826 714 855 716
rect 895 714 928 716
rect 14551 735 14653 750
rect 688 682 723 714
rect 757 682 792 714
rect 826 682 861 714
rect 895 682 930 714
rect 964 682 999 714
rect 1033 682 1068 714
rect 1102 682 1137 714
rect 1171 682 1206 714
rect 1240 682 1275 714
rect 1309 682 1344 714
rect 1378 682 1413 714
rect 1447 682 1482 714
rect 1516 682 1551 714
rect 1585 682 1620 714
rect 1654 682 1689 714
rect 1723 682 1758 714
rect 1792 682 1827 714
rect 1861 682 1896 714
rect 1930 682 1965 714
rect 1999 682 2034 714
rect 2068 682 2103 714
rect 2137 682 2172 714
rect 2206 682 2241 714
rect 2275 682 2310 714
rect 2344 682 2379 714
rect 2413 682 2448 714
rect 2482 682 2517 714
rect 2551 682 2586 714
rect 2620 682 2655 714
rect 2689 682 2724 714
rect 2758 682 2793 714
rect 2827 682 2862 714
rect 2896 682 2931 714
rect 2965 682 3000 714
rect 3034 682 3069 714
rect 3103 682 3138 714
rect 3172 682 3207 714
rect 3241 682 3276 714
rect 3310 682 3345 714
rect 3379 682 3414 714
rect 3448 682 3483 714
rect 3517 682 3552 714
rect 3586 682 3621 714
rect 3655 682 3690 714
rect 3724 682 3759 714
rect 3793 682 3828 714
rect 3862 682 3897 714
rect 3931 682 3966 714
rect 4000 682 4035 714
rect 4069 682 4104 714
rect 4138 682 4173 714
rect 4207 682 4242 714
rect 4276 682 4311 714
rect 4345 682 4380 714
rect 4414 682 4449 714
rect 4483 682 4518 714
rect 4552 682 4587 714
rect 4621 682 4656 714
rect 4690 682 4725 714
rect 14551 701 14604 735
rect 14638 701 14653 735
rect 14551 682 14653 701
rect 482 667 14653 682
rect 14807 4636 14832 4670
rect 14807 4598 14840 4636
rect 14807 4564 14832 4598
rect 14807 4526 14840 4564
rect 14807 4492 14832 4526
rect 14807 4454 14840 4492
rect 14807 4420 14832 4454
rect 14807 4382 14840 4420
rect 14807 4348 14832 4382
rect 14807 4310 14840 4348
rect 14807 4276 14832 4310
rect 14807 4238 14840 4276
rect 14807 4204 14832 4238
rect 14807 4166 14840 4204
rect 14807 4132 14832 4166
rect 14807 4094 14840 4132
rect 14807 4060 14832 4094
rect 14807 4022 14840 4060
rect 14807 3988 14832 4022
rect 14807 3950 14840 3988
rect 14807 3916 14832 3950
rect 14807 3878 14840 3916
rect 14807 3844 14832 3878
rect 14807 3806 14840 3844
rect 14807 3772 14832 3806
rect 14807 3734 14840 3772
rect 14807 3700 14832 3734
rect 14807 3662 14840 3700
rect 14807 3628 14832 3662
rect 14807 3590 14840 3628
rect 14807 3556 14832 3590
rect 14807 3518 14840 3556
rect 14807 3484 14832 3518
rect 14807 3446 14840 3484
rect 14807 3412 14832 3446
rect 14807 3374 14840 3412
rect 14807 3340 14832 3374
rect 14807 3302 14840 3340
rect 14807 3268 14832 3302
rect 14807 3230 14840 3268
rect 14807 3196 14832 3230
rect 14807 3158 14840 3196
rect 14807 3124 14832 3158
rect 14807 3086 14840 3124
rect 14807 3052 14832 3086
rect 14807 3014 14840 3052
rect 14807 2980 14832 3014
rect 14807 2942 14840 2980
rect 14807 2908 14832 2942
rect 14807 2870 14840 2908
rect 14807 2836 14832 2870
rect 14807 2798 14840 2836
rect 14807 2764 14832 2798
rect 14807 2726 14840 2764
rect 14807 2692 14832 2726
rect 14807 2654 14840 2692
rect 14807 2620 14832 2654
rect 14807 2582 14840 2620
rect 14807 2548 14832 2582
rect 14807 2510 14840 2548
rect 14807 2476 14832 2510
rect 14807 2438 14840 2476
rect 14807 2404 14832 2438
rect 14807 2366 14840 2404
rect 14807 2332 14832 2366
rect 14807 2294 14840 2332
rect 14807 2260 14832 2294
rect 14807 2222 14840 2260
rect 14807 2188 14832 2222
rect 14807 2150 14840 2188
rect 14807 2116 14832 2150
rect 14807 2078 14840 2116
rect 14807 2044 14832 2078
rect 14807 2006 14840 2044
rect 14807 1972 14832 2006
rect 14807 1934 14840 1972
rect 14807 1900 14832 1934
rect 14807 1862 14840 1900
rect 14807 1828 14832 1862
rect 14807 1790 14840 1828
rect 14807 1756 14832 1790
rect 14807 1718 14840 1756
rect 14807 1684 14832 1718
rect 14807 1646 14840 1684
rect 14807 1612 14832 1646
rect 14807 1574 14840 1612
rect 14807 1540 14832 1574
rect 14807 1502 14840 1540
rect 14807 1468 14832 1502
rect 14807 1429 14840 1468
rect 14807 1395 14832 1429
rect 14807 1356 14840 1395
rect 14807 1322 14832 1356
rect 14807 1283 14840 1322
rect 14807 1249 14832 1283
rect 14807 1210 14840 1249
rect 14807 1176 14832 1210
rect 14807 1137 14840 1176
rect 14807 1103 14832 1137
rect 14807 1064 14840 1103
rect 14807 1030 14832 1064
rect 14807 991 14840 1030
rect 14807 957 14832 991
rect 14807 918 14840 957
rect 14807 884 14832 918
rect 14807 845 14840 884
rect 14807 811 14832 845
rect 14807 772 14840 811
rect 14807 738 14832 772
rect 14807 699 14840 738
rect 229 609 262 643
rect 296 641 329 643
rect 229 607 269 609
rect 303 607 329 641
rect 229 575 329 607
rect 229 541 262 575
rect 296 567 329 575
rect 229 533 269 541
rect 303 533 329 567
rect 229 514 329 533
rect 14807 665 14832 699
rect 14807 626 14840 665
rect 14807 592 14832 626
rect 14807 553 14840 592
rect 14807 519 14832 553
rect 14807 514 14840 519
rect 267 499 305 514
rect 14832 499 14840 514
rect 121 329 223 363
rect 228 465 262 499
rect 296 465 331 499
rect 365 497 400 499
rect 434 497 469 499
rect 503 497 538 499
rect 572 497 607 499
rect 377 465 400 497
rect 453 465 469 497
rect 529 465 538 497
rect 605 465 607 497
rect 641 497 676 499
rect 641 465 648 497
rect 710 465 745 499
rect 779 465 814 499
rect 848 465 883 499
rect 917 465 952 499
rect 986 465 1021 499
rect 1055 465 1090 499
rect 1124 465 1159 499
rect 1193 465 1228 499
rect 1262 465 1297 499
rect 1331 465 1366 499
rect 1400 465 1435 499
rect 1469 465 1504 499
rect 1538 465 1573 499
rect 1607 465 1642 499
rect 1676 465 1711 499
rect 1745 465 1780 499
rect 1814 465 1849 499
rect 1883 465 1918 499
rect 1952 465 1987 499
rect 2021 465 2056 499
rect 228 463 343 465
rect 377 463 419 465
rect 453 463 495 465
rect 529 463 571 465
rect 605 463 648 465
rect 682 463 2056 465
rect 228 431 2056 463
rect 228 397 262 431
rect 296 397 331 431
rect 365 397 400 431
rect 434 397 469 431
rect 503 397 538 431
rect 572 397 607 431
rect 641 397 676 431
rect 710 397 745 431
rect 779 397 814 431
rect 848 397 883 431
rect 917 397 952 431
rect 986 397 1021 431
rect 1055 397 1090 431
rect 1124 397 1159 431
rect 1193 397 1228 431
rect 1262 397 1297 431
rect 1331 397 1366 431
rect 1400 397 1435 431
rect 1469 397 1504 431
rect 1538 397 1573 431
rect 1607 397 1642 431
rect 1676 397 1711 431
rect 1745 397 1780 431
rect 1814 397 1849 431
rect 1883 397 1918 431
rect 1952 397 1987 431
rect 2021 397 2056 431
rect 228 375 2056 397
rect 14942 375 15051 4965
rect 228 363 361 375
rect 395 363 434 375
rect 228 329 262 363
rect 296 329 331 363
rect 395 341 400 363
rect 365 329 400 341
rect 468 363 507 375
rect 541 363 580 375
rect 614 363 653 375
rect 687 363 726 375
rect 760 363 799 375
rect 833 363 872 375
rect 906 363 945 375
rect 979 363 1018 375
rect 1052 363 1091 375
rect 1125 363 1164 375
rect 1198 363 1237 375
rect 1271 363 1310 375
rect 1344 363 1383 375
rect 1417 363 1456 375
rect 1490 363 1529 375
rect 1563 363 1602 375
rect 1636 363 1675 375
rect 1709 363 1748 375
rect 1782 363 1821 375
rect 1855 363 1894 375
rect 1928 363 1967 375
rect 2001 363 2040 375
rect 468 341 469 363
rect 434 329 469 341
rect 503 341 507 363
rect 572 341 580 363
rect 641 341 653 363
rect 710 341 726 363
rect 779 341 799 363
rect 848 341 872 363
rect 917 341 945 363
rect 986 341 1018 363
rect 503 329 538 341
rect 572 329 607 341
rect 641 329 676 341
rect 710 329 745 341
rect 779 329 814 341
rect 848 329 883 341
rect 917 329 952 341
rect 986 329 1021 341
rect 1055 329 1090 363
rect 1125 341 1159 363
rect 1198 341 1228 363
rect 1271 341 1297 363
rect 1344 341 1366 363
rect 1417 341 1435 363
rect 1490 341 1504 363
rect 1563 341 1573 363
rect 1636 341 1642 363
rect 1709 341 1711 363
rect 1124 329 1159 341
rect 1193 329 1228 341
rect 1262 329 1297 341
rect 1331 329 1366 341
rect 1400 329 1435 341
rect 1469 329 1504 341
rect 1538 329 1573 341
rect 1607 329 1642 341
rect 1676 329 1711 341
rect 1745 341 1748 363
rect 1814 341 1821 363
rect 1883 341 1894 363
rect 1952 341 1967 363
rect 2021 341 2040 363
rect 14806 341 15051 375
rect 1745 329 1780 341
rect 1814 329 1849 341
rect 1883 329 1918 341
rect 1952 329 1987 341
rect 2021 329 2056 341
rect 14806 329 14840 341
rect 329 314 14807 329
rect 14927 -976 15051 341
<< viali >>
rect 361 5077 395 5111
rect 434 5077 468 5111
rect 507 5077 541 5111
rect 580 5077 614 5111
rect 653 5077 687 5111
rect 726 5077 760 5111
rect 799 5077 833 5111
rect 872 5077 906 5111
rect 945 5077 979 5111
rect 1018 5077 1052 5111
rect 1091 5077 1125 5111
rect 1164 5077 1198 5111
rect 1237 5077 1271 5111
rect 1310 5077 1344 5111
rect 1383 5077 1417 5111
rect 1456 5077 1490 5111
rect 1529 5077 1563 5111
rect 1602 5077 1636 5111
rect 1675 5077 1709 5111
rect 1748 5077 1782 5111
rect 1821 5077 1855 5111
rect 1894 5077 1928 5111
rect 1967 5077 2001 5111
rect 2040 5077 2074 5111
rect 2113 5077 2147 5111
rect 2186 5077 2220 5111
rect 2259 5077 2293 5111
rect 2332 5077 2366 5111
rect 2405 5077 2439 5111
rect 2478 5077 2512 5111
rect 2551 5077 2585 5111
rect 2624 5077 2658 5111
rect 2697 5077 2731 5111
rect 2770 5077 2804 5111
rect 2843 5077 2877 5111
rect 2916 5077 2950 5111
rect 2989 5077 3023 5111
rect 3062 5077 3096 5111
rect 3135 5077 3169 5111
rect 3208 5077 3242 5111
rect 3281 5077 3315 5111
rect 3354 5077 3388 5111
rect 3427 5077 3461 5111
rect 3500 5077 3534 5111
rect 3573 5077 3607 5111
rect 3646 5077 3680 5111
rect 3719 5077 3753 5111
rect 3792 5077 3826 5111
rect 3865 5077 3899 5111
rect 3938 5077 3972 5111
rect 4011 5077 4045 5111
rect 4084 5077 4118 5111
rect 4157 5077 4191 5111
rect 4229 5077 4263 5111
rect 4301 5077 4335 5111
rect 4373 5077 4407 5111
rect 4445 5077 4479 5111
rect 4517 5077 4551 5111
rect 4589 5077 4623 5111
rect 4661 5077 4695 5111
rect 4733 5077 4767 5111
rect 4805 5077 4839 5111
rect 4877 5077 4911 5111
rect 4949 5077 4983 5111
rect 5021 5077 5055 5111
rect 5093 5077 5127 5111
rect 5165 5077 5199 5111
rect 5237 5077 5271 5111
rect 5309 5077 5343 5111
rect 5381 5077 5415 5111
rect 5453 5077 5487 5111
rect 5525 5077 5559 5111
rect 5597 5077 5631 5111
rect 5669 5077 5703 5111
rect 5741 5077 5775 5111
rect 5813 5077 5847 5111
rect 5885 5077 5919 5111
rect 5957 5077 5991 5111
rect 6029 5077 6063 5111
rect 6101 5077 6135 5111
rect 6173 5077 6207 5111
rect 6245 5077 6279 5111
rect 6317 5077 6351 5111
rect 6389 5077 6423 5111
rect 6461 5077 6495 5111
rect 6533 5077 6567 5111
rect 6605 5077 6639 5111
rect 6677 5077 6711 5111
rect 6749 5077 6783 5111
rect 6821 5077 6855 5111
rect 6893 5077 6927 5111
rect 6965 5077 6999 5111
rect 7037 5077 7071 5111
rect 7109 5077 7143 5111
rect 7181 5077 7215 5111
rect 7253 5077 7287 5111
rect 7325 5077 7359 5111
rect 7397 5077 7431 5111
rect 7469 5077 7503 5111
rect 7541 5077 7575 5111
rect 7613 5077 7647 5111
rect 7685 5077 7719 5111
rect 7757 5077 7791 5111
rect 7829 5077 7863 5111
rect 7901 5077 7935 5111
rect 7973 5077 8007 5111
rect 8045 5077 8079 5111
rect 8117 5077 8151 5111
rect 8189 5077 8223 5111
rect 8261 5077 8295 5111
rect 8333 5077 8367 5111
rect 8405 5077 8439 5111
rect 8477 5077 8511 5111
rect 8549 5077 8583 5111
rect 8621 5077 8655 5111
rect 8693 5077 8727 5111
rect 8765 5077 8799 5111
rect 8837 5077 8871 5111
rect 8909 5077 8943 5111
rect 8981 5077 9015 5111
rect 9053 5077 9087 5111
rect 9125 5077 9159 5111
rect 9197 5077 9231 5111
rect 9269 5077 9303 5111
rect 9341 5077 9375 5111
rect 9413 5077 9447 5111
rect 9485 5077 9519 5111
rect 9557 5077 9591 5111
rect 9629 5077 9663 5111
rect 9701 5077 9735 5111
rect 9773 5077 9807 5111
rect 9845 5077 9879 5111
rect 9917 5077 9951 5111
rect 9989 5077 10023 5111
rect 10061 5077 10095 5111
rect 10133 5077 10167 5111
rect 10205 5077 10239 5111
rect 10277 5077 10311 5111
rect 10349 5077 10383 5111
rect 10421 5077 10455 5111
rect 10493 5077 10527 5111
rect 10565 5077 10599 5111
rect 10637 5077 10671 5111
rect 10709 5077 10743 5111
rect 10781 5077 10815 5111
rect 10853 5077 10887 5111
rect 10925 5077 10959 5111
rect 10997 5077 11031 5111
rect 11069 5077 11103 5111
rect 11141 5077 11175 5111
rect 11213 5077 11247 5111
rect 11285 5077 11319 5111
rect 11357 5077 11391 5111
rect 11429 5077 11463 5111
rect 11501 5077 11535 5111
rect 11573 5077 11607 5111
rect 11645 5077 11679 5111
rect 11717 5077 11751 5111
rect 11789 5077 11823 5111
rect 11861 5077 11895 5111
rect 11933 5077 11967 5111
rect 12005 5077 12039 5111
rect 12077 5077 12111 5111
rect 12149 5077 12183 5111
rect 12221 5077 12255 5111
rect 12293 5077 12327 5111
rect 12365 5077 12399 5111
rect 12437 5077 12471 5111
rect 12509 5077 12543 5111
rect 12581 5077 12615 5111
rect 12653 5077 12687 5111
rect 12725 5077 12759 5111
rect 12797 5077 12831 5111
rect 12869 5077 12903 5111
rect 12941 5077 12975 5111
rect 13013 5077 13047 5111
rect 13085 5077 13119 5111
rect 13157 5077 13191 5111
rect 13229 5077 13263 5111
rect 13301 5077 13335 5111
rect 13373 5077 13407 5111
rect 13445 5077 13479 5111
rect 13517 5077 13551 5111
rect 13589 5077 13623 5111
rect 13661 5077 13695 5111
rect 13733 5077 13767 5111
rect 13805 5077 13839 5111
rect 13877 5077 13911 5111
rect 13949 5077 13983 5111
rect 14021 5077 14055 5111
rect 14093 5077 14127 5111
rect 14165 5077 14199 5111
rect 14237 5077 14271 5111
rect 14309 5077 14343 5111
rect 14381 5077 14415 5111
rect 14453 5077 14487 5111
rect 14525 5077 14559 5111
rect 14597 5077 14631 5111
rect 14669 5077 14703 5111
rect 14741 5077 14775 5111
rect 269 4995 303 5029
rect 361 5001 395 5035
rect 434 5001 468 5035
rect 507 5001 541 5035
rect 580 5001 614 5035
rect 653 5001 687 5035
rect 726 5001 760 5035
rect 799 5001 833 5035
rect 872 5001 906 5035
rect 945 5001 979 5035
rect 1018 5001 1052 5035
rect 1091 5001 1125 5035
rect 1164 5001 1198 5035
rect 1237 5001 1271 5035
rect 1310 5001 1344 5035
rect 1383 5001 1417 5035
rect 1456 5001 1490 5035
rect 1529 5001 1563 5035
rect 1602 5001 1636 5035
rect 1675 5001 1709 5035
rect 1748 5001 1782 5035
rect 1821 5001 1855 5035
rect 1894 5001 1928 5035
rect 1967 5001 2001 5035
rect 2040 5001 2074 5035
rect 2113 5001 2147 5035
rect 2186 5001 2220 5035
rect 2259 5001 2293 5035
rect 2332 5001 2366 5035
rect 2405 5001 2439 5035
rect 2478 5001 2512 5035
rect 2551 5001 2585 5035
rect 2624 5001 2658 5035
rect 2697 5001 2731 5035
rect 2770 5001 2804 5035
rect 2843 5001 2877 5035
rect 2916 5001 2950 5035
rect 2989 5001 3023 5035
rect 3062 5001 3096 5035
rect 3135 5001 3169 5035
rect 3208 5001 3242 5035
rect 3281 5001 3315 5035
rect 3354 5001 3388 5035
rect 3427 5001 3461 5035
rect 3500 5001 3534 5035
rect 3573 5001 3607 5035
rect 3646 5001 3680 5035
rect 3719 5001 3753 5035
rect 3792 5001 3826 5035
rect 3865 5001 3899 5035
rect 3938 5001 3972 5035
rect 4011 5001 4045 5035
rect 4084 5001 4118 5035
rect 4157 5001 4191 5035
rect 4229 5001 4263 5035
rect 4301 5001 4335 5035
rect 4373 5001 4407 5035
rect 4445 5001 4479 5035
rect 4517 5001 4551 5035
rect 4589 5001 4623 5035
rect 4661 5001 4695 5035
rect 4733 5001 4767 5035
rect 4805 5001 4839 5035
rect 4877 5001 4911 5035
rect 4949 5001 4983 5035
rect 5021 5001 5055 5035
rect 5093 5001 5127 5035
rect 5165 5001 5199 5035
rect 5237 5001 5271 5035
rect 5309 5001 5343 5035
rect 5381 5001 5415 5035
rect 5453 5001 5487 5035
rect 5525 5001 5559 5035
rect 5597 5001 5631 5035
rect 5669 5001 5703 5035
rect 5741 5001 5775 5035
rect 5813 5001 5847 5035
rect 5885 5001 5919 5035
rect 5957 5001 5991 5035
rect 6029 5001 6063 5035
rect 6101 5001 6135 5035
rect 6173 5001 6207 5035
rect 6245 5001 6279 5035
rect 6317 5001 6351 5035
rect 6389 5001 6423 5035
rect 6461 5001 6495 5035
rect 6533 5001 6567 5035
rect 6605 5001 6639 5035
rect 6677 5001 6711 5035
rect 6749 5001 6783 5035
rect 6821 5001 6855 5035
rect 6893 5001 6927 5035
rect 6965 5001 6999 5035
rect 7037 5001 7071 5035
rect 7109 5001 7143 5035
rect 7181 5001 7215 5035
rect 7253 5001 7287 5035
rect 7325 5001 7359 5035
rect 7397 5001 7431 5035
rect 7469 5001 7503 5035
rect 7541 5001 7575 5035
rect 7613 5001 7647 5035
rect 7685 5001 7719 5035
rect 7757 5001 7791 5035
rect 7829 5001 7863 5035
rect 7901 5001 7935 5035
rect 7973 5001 8007 5035
rect 8045 5001 8079 5035
rect 8117 5001 8151 5035
rect 8189 5001 8223 5035
rect 8261 5001 8295 5035
rect 8333 5001 8367 5035
rect 8405 5001 8439 5035
rect 8477 5001 8511 5035
rect 8549 5001 8583 5035
rect 8621 5001 8655 5035
rect 8693 5001 8727 5035
rect 8765 5001 8799 5035
rect 8837 5001 8871 5035
rect 8909 5001 8943 5035
rect 8981 5001 9015 5035
rect 9053 5001 9087 5035
rect 9125 5001 9159 5035
rect 9197 5001 9231 5035
rect 9269 5001 9303 5035
rect 9341 5001 9375 5035
rect 9413 5001 9447 5035
rect 9485 5001 9519 5035
rect 9557 5001 9591 5035
rect 9629 5001 9663 5035
rect 9701 5001 9735 5035
rect 9773 5001 9807 5035
rect 9845 5001 9879 5035
rect 9917 5001 9951 5035
rect 9989 5001 10023 5035
rect 10061 5001 10095 5035
rect 10133 5001 10167 5035
rect 10205 5001 10239 5035
rect 10277 5001 10311 5035
rect 10349 5001 10383 5035
rect 10421 5001 10455 5035
rect 10493 5001 10527 5035
rect 10565 5001 10599 5035
rect 10637 5001 10671 5035
rect 10709 5001 10743 5035
rect 10781 5001 10815 5035
rect 10853 5001 10887 5035
rect 10925 5001 10959 5035
rect 10997 5001 11031 5035
rect 11069 5001 11103 5035
rect 11141 5001 11175 5035
rect 11213 5001 11247 5035
rect 11285 5001 11319 5035
rect 11357 5001 11391 5035
rect 11429 5001 11463 5035
rect 11501 5001 11535 5035
rect 11573 5001 11607 5035
rect 11645 5001 11679 5035
rect 11717 5001 11751 5035
rect 11789 5001 11823 5035
rect 11861 5001 11895 5035
rect 11933 5001 11967 5035
rect 12005 5001 12039 5035
rect 12077 5001 12111 5035
rect 12149 5001 12183 5035
rect 12221 5001 12255 5035
rect 12293 5001 12327 5035
rect 12365 5001 12399 5035
rect 12437 5001 12471 5035
rect 12509 5001 12543 5035
rect 12581 5001 12615 5035
rect 12653 5001 12687 5035
rect 12725 5001 12759 5035
rect 12797 5001 12831 5035
rect 12869 5001 12903 5035
rect 12941 5001 12975 5035
rect 13013 5001 13047 5035
rect 13085 5001 13119 5035
rect 13157 5001 13191 5035
rect 13229 5001 13263 5035
rect 13301 5001 13335 5035
rect 13373 5001 13407 5035
rect 13445 5001 13479 5035
rect 13517 5001 13551 5035
rect 13589 5001 13600 5035
rect 13600 5001 13623 5035
rect 13661 5034 13669 5035
rect 13669 5034 13695 5035
rect 13733 5034 13738 5035
rect 13738 5034 13767 5035
rect 13805 5034 13807 5035
rect 13807 5034 13839 5035
rect 13661 5001 13695 5034
rect 13733 5001 13767 5034
rect 13805 5001 13839 5034
rect 13877 5001 13911 5035
rect 13949 5034 13980 5035
rect 13980 5034 13983 5035
rect 14021 5034 14049 5035
rect 14049 5034 14055 5035
rect 14093 5034 14118 5035
rect 14118 5034 14127 5035
rect 14165 5034 14187 5035
rect 14187 5034 14199 5035
rect 14237 5034 14256 5035
rect 14256 5034 14271 5035
rect 14309 5034 14325 5035
rect 14325 5034 14343 5035
rect 14381 5034 14394 5035
rect 14394 5034 14415 5035
rect 14453 5034 14463 5035
rect 14463 5034 14487 5035
rect 14525 5034 14532 5035
rect 14532 5034 14559 5035
rect 14597 5034 14601 5035
rect 14601 5034 14631 5035
rect 14669 5034 14670 5035
rect 14670 5034 14703 5035
rect 14741 5034 14773 5035
rect 14773 5034 14775 5035
rect 13949 5001 13983 5034
rect 14021 5001 14055 5034
rect 14093 5001 14127 5034
rect 14165 5001 14199 5034
rect 14237 5001 14271 5034
rect 14309 5001 14343 5034
rect 14381 5001 14415 5034
rect 14453 5001 14487 5034
rect 14525 5001 14559 5034
rect 14597 5001 14631 5034
rect 14669 5001 14703 5034
rect 14741 5001 14775 5034
rect 14832 4999 14840 5030
rect 14840 4999 14866 5030
rect 14832 4996 14866 4999
rect 269 4922 303 4956
rect 361 4925 395 4959
rect 434 4925 468 4959
rect 507 4925 541 4959
rect 580 4925 614 4959
rect 653 4925 687 4959
rect 726 4925 760 4959
rect 799 4925 833 4959
rect 872 4925 906 4959
rect 945 4925 979 4959
rect 1018 4925 1052 4959
rect 1091 4925 1125 4959
rect 1164 4925 1198 4959
rect 1237 4925 1271 4959
rect 1310 4925 1344 4959
rect 1383 4925 1417 4959
rect 1456 4925 1490 4959
rect 1529 4925 1563 4959
rect 1602 4925 1636 4959
rect 1675 4925 1709 4959
rect 1748 4925 1782 4959
rect 1821 4925 1855 4959
rect 1894 4925 1928 4959
rect 1967 4925 2001 4959
rect 2040 4925 2074 4959
rect 2113 4925 2147 4959
rect 2186 4925 2220 4959
rect 2259 4925 2293 4959
rect 2332 4925 2366 4959
rect 2405 4925 2439 4959
rect 2478 4925 2512 4959
rect 2551 4925 2585 4959
rect 2624 4925 2658 4959
rect 2697 4925 2731 4959
rect 2770 4925 2804 4959
rect 2843 4925 2877 4959
rect 2916 4925 2950 4959
rect 2989 4925 3023 4959
rect 3062 4925 3096 4959
rect 3135 4925 3169 4959
rect 3208 4925 3242 4959
rect 3281 4925 3315 4959
rect 3354 4925 3388 4959
rect 3427 4925 3461 4959
rect 3500 4925 3534 4959
rect 3573 4925 3607 4959
rect 3646 4925 3680 4959
rect 3719 4925 3753 4959
rect 3792 4925 3826 4959
rect 3865 4925 3899 4959
rect 3938 4925 3972 4959
rect 4011 4925 4045 4959
rect 4084 4925 4118 4959
rect 4157 4925 4191 4959
rect 4229 4925 4263 4959
rect 4301 4925 4335 4959
rect 4373 4925 4407 4959
rect 4445 4925 4479 4959
rect 4517 4925 4551 4959
rect 4589 4925 4623 4959
rect 4661 4925 4695 4959
rect 4733 4925 4767 4959
rect 4805 4925 4839 4959
rect 4877 4925 4911 4959
rect 4949 4925 4983 4959
rect 5021 4925 5055 4959
rect 5093 4925 5127 4959
rect 5165 4925 5199 4959
rect 5237 4925 5271 4959
rect 5309 4925 5343 4959
rect 5381 4925 5415 4959
rect 5453 4925 5487 4959
rect 5525 4925 5559 4959
rect 5597 4925 5631 4959
rect 5669 4925 5703 4959
rect 5741 4925 5775 4959
rect 5813 4925 5847 4959
rect 5885 4925 5919 4959
rect 5957 4925 5991 4959
rect 6029 4925 6063 4959
rect 6101 4925 6135 4959
rect 6173 4925 6207 4959
rect 6245 4925 6279 4959
rect 6317 4925 6351 4959
rect 6389 4925 6423 4959
rect 6461 4925 6495 4959
rect 6533 4925 6567 4959
rect 6605 4925 6639 4959
rect 6677 4925 6711 4959
rect 6749 4925 6783 4959
rect 6821 4925 6855 4959
rect 6893 4925 6927 4959
rect 6965 4925 6999 4959
rect 7037 4925 7071 4959
rect 7109 4925 7143 4959
rect 7181 4925 7215 4959
rect 7253 4925 7287 4959
rect 7325 4925 7359 4959
rect 7397 4925 7431 4959
rect 7469 4925 7503 4959
rect 7541 4925 7575 4959
rect 7613 4925 7647 4959
rect 7685 4925 7719 4959
rect 7757 4925 7791 4959
rect 7829 4925 7863 4959
rect 7901 4925 7935 4959
rect 7973 4925 8007 4959
rect 8045 4925 8079 4959
rect 8117 4925 8151 4959
rect 8189 4925 8223 4959
rect 8261 4925 8295 4959
rect 8333 4925 8367 4959
rect 8405 4925 8439 4959
rect 8477 4925 8511 4959
rect 8549 4925 8583 4959
rect 8621 4925 8655 4959
rect 8693 4925 8727 4959
rect 8765 4925 8799 4959
rect 8837 4925 8871 4959
rect 8909 4925 8943 4959
rect 8981 4925 9015 4959
rect 9053 4925 9087 4959
rect 9125 4925 9159 4959
rect 9197 4925 9231 4959
rect 9269 4925 9303 4959
rect 9341 4925 9375 4959
rect 9413 4925 9447 4959
rect 9485 4925 9519 4959
rect 9557 4925 9591 4959
rect 9629 4925 9663 4959
rect 9701 4925 9735 4959
rect 9773 4925 9807 4959
rect 9845 4925 9879 4959
rect 9917 4925 9951 4959
rect 9989 4925 10023 4959
rect 10061 4925 10095 4959
rect 10133 4925 10167 4959
rect 10205 4925 10239 4959
rect 10277 4925 10311 4959
rect 10349 4925 10383 4959
rect 10421 4925 10455 4959
rect 10493 4925 10527 4959
rect 10565 4925 10599 4959
rect 10637 4925 10671 4959
rect 10709 4925 10743 4959
rect 10781 4925 10815 4959
rect 10853 4925 10887 4959
rect 10925 4925 10959 4959
rect 10997 4925 11031 4959
rect 11069 4925 11103 4959
rect 11141 4925 11175 4959
rect 11213 4925 11247 4959
rect 11285 4925 11319 4959
rect 11357 4925 11391 4959
rect 11429 4925 11463 4959
rect 11501 4925 11535 4959
rect 11573 4925 11607 4959
rect 11645 4925 11679 4959
rect 11717 4925 11751 4959
rect 11789 4925 11823 4959
rect 11861 4925 11895 4959
rect 11933 4925 11967 4959
rect 12005 4925 12039 4959
rect 12077 4925 12111 4959
rect 12149 4925 12183 4959
rect 12221 4925 12255 4959
rect 12293 4925 12327 4959
rect 12365 4925 12399 4959
rect 12437 4925 12471 4959
rect 12509 4925 12543 4959
rect 12581 4925 12615 4959
rect 12653 4925 12687 4959
rect 12725 4925 12759 4959
rect 12797 4925 12831 4959
rect 12869 4925 12903 4959
rect 12941 4925 12975 4959
rect 13013 4925 13047 4959
rect 13085 4925 13119 4959
rect 13157 4925 13191 4959
rect 13229 4925 13263 4959
rect 13301 4925 13335 4959
rect 13373 4925 13407 4959
rect 13445 4925 13479 4959
rect 13517 4925 13551 4959
rect 13589 4925 13600 4959
rect 13600 4925 13623 4959
rect 13661 4932 13695 4959
rect 13733 4932 13767 4959
rect 13805 4932 13839 4959
rect 13661 4925 13669 4932
rect 13669 4925 13695 4932
rect 13733 4925 13738 4932
rect 13738 4925 13767 4932
rect 13805 4925 13807 4932
rect 13807 4925 13839 4932
rect 13877 4925 13911 4959
rect 13949 4932 13983 4959
rect 14021 4932 14055 4959
rect 14093 4932 14127 4959
rect 14165 4932 14199 4959
rect 14237 4932 14271 4959
rect 14309 4932 14343 4959
rect 14381 4932 14415 4959
rect 14453 4932 14487 4959
rect 14525 4932 14559 4959
rect 14597 4932 14631 4959
rect 14669 4932 14703 4959
rect 14741 4932 14775 4959
rect 13949 4925 13980 4932
rect 13980 4925 13983 4932
rect 14021 4925 14049 4932
rect 14049 4925 14055 4932
rect 14093 4925 14118 4932
rect 14118 4925 14127 4932
rect 14165 4925 14187 4932
rect 14187 4925 14199 4932
rect 14237 4925 14256 4932
rect 14256 4925 14271 4932
rect 14309 4925 14325 4932
rect 14325 4925 14343 4932
rect 14381 4925 14394 4932
rect 14394 4925 14415 4932
rect 14453 4925 14463 4932
rect 14463 4925 14487 4932
rect 14525 4925 14532 4932
rect 14532 4925 14559 4932
rect 14597 4925 14601 4932
rect 14601 4925 14631 4932
rect 14669 4925 14670 4932
rect 14670 4925 14703 4932
rect 14741 4925 14773 4932
rect 14773 4925 14775 4932
rect 14832 4924 14840 4958
rect 14840 4924 14866 4958
rect 269 4859 303 4883
rect 269 4849 296 4859
rect 296 4849 303 4859
rect 269 4791 303 4810
rect 269 4776 296 4791
rect 296 4776 303 4791
rect 269 4723 303 4737
rect 269 4703 296 4723
rect 296 4703 303 4723
rect 269 4655 303 4664
rect 269 4630 296 4655
rect 296 4630 303 4655
rect 14832 4852 14840 4886
rect 14840 4852 14866 4886
rect 14832 4780 14840 4814
rect 14840 4780 14866 4814
rect 14832 4708 14840 4742
rect 14840 4708 14866 4742
rect 269 4587 303 4591
rect 269 4557 296 4587
rect 296 4557 303 4587
rect 269 4485 296 4518
rect 296 4485 303 4518
rect 269 4484 303 4485
rect 269 4417 296 4445
rect 296 4417 303 4445
rect 269 4411 303 4417
rect 269 4349 296 4372
rect 296 4349 303 4372
rect 269 4338 303 4349
rect 269 4281 296 4299
rect 296 4281 303 4299
rect 269 4265 303 4281
rect 269 4213 296 4226
rect 296 4213 303 4226
rect 269 4192 303 4213
rect 269 4145 296 4153
rect 296 4145 303 4153
rect 269 4119 303 4145
rect 269 4077 296 4080
rect 296 4077 303 4080
rect 269 4046 303 4077
rect 269 3975 303 4007
rect 269 3973 296 3975
rect 296 3973 303 3975
rect 269 3907 303 3934
rect 269 3900 296 3907
rect 296 3900 303 3907
rect 269 3839 303 3861
rect 269 3827 296 3839
rect 296 3827 303 3839
rect 269 3771 303 3788
rect 269 3754 296 3771
rect 296 3754 303 3771
rect 269 3703 303 3715
rect 269 3681 296 3703
rect 296 3681 303 3703
rect 269 3635 303 3642
rect 269 3608 296 3635
rect 296 3608 303 3635
rect 269 3567 303 3569
rect 269 3535 296 3567
rect 296 3535 303 3567
rect 269 3465 296 3496
rect 296 3465 303 3496
rect 269 3462 303 3465
rect 269 3397 296 3423
rect 296 3397 303 3423
rect 269 3389 303 3397
rect 269 3329 296 3350
rect 296 3329 303 3350
rect 269 3316 303 3329
rect 269 3261 296 3277
rect 296 3261 303 3277
rect 269 3243 303 3261
rect 269 3193 296 3204
rect 296 3193 303 3204
rect 269 3170 303 3193
rect 269 3125 296 3131
rect 296 3125 303 3131
rect 269 3097 303 3125
rect 269 3057 296 3058
rect 296 3057 303 3058
rect 269 3024 303 3057
rect 269 2955 303 2985
rect 269 2951 296 2955
rect 296 2951 303 2955
rect 269 2887 303 2912
rect 269 2878 296 2887
rect 296 2878 303 2887
rect 269 2819 303 2839
rect 269 2805 296 2819
rect 296 2805 303 2819
rect 269 2751 303 2766
rect 269 2732 296 2751
rect 296 2732 303 2751
rect 269 2683 303 2693
rect 269 2659 296 2683
rect 296 2659 303 2683
rect 269 2615 303 2620
rect 269 2586 296 2615
rect 296 2586 303 2615
rect 269 2513 296 2547
rect 296 2513 303 2547
rect 269 2445 296 2474
rect 296 2445 303 2474
rect 269 2440 303 2445
rect 269 2377 296 2401
rect 296 2377 303 2401
rect 269 2367 303 2377
rect 269 2309 296 2328
rect 296 2309 303 2328
rect 269 2294 303 2309
rect 269 2241 296 2255
rect 296 2241 303 2255
rect 269 2221 303 2241
rect 269 2173 296 2182
rect 296 2173 303 2182
rect 269 2148 303 2173
rect 269 2105 296 2109
rect 296 2105 303 2109
rect 269 2075 303 2105
rect 269 2003 303 2036
rect 269 2002 296 2003
rect 296 2002 303 2003
rect 269 1935 303 1963
rect 269 1929 296 1935
rect 296 1929 303 1935
rect 269 1867 303 1890
rect 269 1856 296 1867
rect 296 1856 303 1867
rect 269 1799 303 1817
rect 269 1783 296 1799
rect 296 1783 303 1799
rect 269 1731 303 1744
rect 269 1710 296 1731
rect 296 1710 303 1731
rect 269 1663 303 1671
rect 269 1637 296 1663
rect 296 1637 303 1663
rect 269 1595 303 1598
rect 269 1564 296 1595
rect 296 1564 303 1595
rect 269 1493 296 1525
rect 296 1493 303 1525
rect 269 1491 303 1493
rect 269 1425 296 1452
rect 296 1425 303 1452
rect 269 1418 303 1425
rect 269 1357 296 1379
rect 296 1357 303 1379
rect 269 1345 303 1357
rect 269 1289 296 1306
rect 296 1289 303 1306
rect 269 1272 303 1289
rect 269 1221 296 1233
rect 296 1221 303 1233
rect 269 1199 303 1221
rect 269 1153 296 1159
rect 296 1153 303 1159
rect 269 1125 303 1153
rect 269 1051 303 1085
rect 269 983 303 1011
rect 269 977 296 983
rect 296 977 303 983
rect 269 915 303 937
rect 269 903 296 915
rect 296 903 303 915
rect 269 847 303 863
rect 269 829 296 847
rect 296 829 303 847
rect 269 779 303 789
rect 269 755 296 779
rect 296 755 303 779
rect 269 711 303 715
rect 269 681 296 711
rect 296 681 303 711
rect 709 4570 10410 4606
rect 10410 4604 10445 4606
rect 10445 4604 10479 4606
rect 10479 4604 10514 4606
rect 10514 4604 10548 4606
rect 10548 4604 10583 4606
rect 10583 4604 10617 4606
rect 10617 4604 10652 4606
rect 10652 4604 10686 4606
rect 10686 4604 10721 4606
rect 10721 4604 10755 4606
rect 10755 4604 10790 4606
rect 10790 4604 10824 4606
rect 10824 4604 10859 4606
rect 10859 4604 10893 4606
rect 10893 4604 10928 4606
rect 10928 4604 10962 4606
rect 10962 4604 10997 4606
rect 10997 4604 11031 4606
rect 11031 4604 11066 4606
rect 11066 4604 11100 4606
rect 11100 4604 11135 4606
rect 11135 4604 11169 4606
rect 11169 4604 11204 4606
rect 11204 4604 11238 4606
rect 11238 4604 11273 4606
rect 11273 4604 11307 4606
rect 11307 4604 11342 4606
rect 11342 4604 11376 4606
rect 11376 4604 11411 4606
rect 11411 4604 11445 4606
rect 11445 4604 11480 4606
rect 11480 4604 11514 4606
rect 11514 4604 11549 4606
rect 11549 4604 11583 4606
rect 11583 4604 11618 4606
rect 11618 4604 11652 4606
rect 11652 4604 11687 4606
rect 11687 4604 11721 4606
rect 11721 4604 11756 4606
rect 11756 4604 11790 4606
rect 11790 4604 11825 4606
rect 11825 4604 11859 4606
rect 11859 4604 11894 4606
rect 11894 4604 11928 4606
rect 11928 4604 11963 4606
rect 11963 4604 11997 4606
rect 11997 4604 12032 4606
rect 12032 4604 12066 4606
rect 12066 4604 12101 4606
rect 12101 4604 12135 4606
rect 12135 4604 12170 4606
rect 12170 4604 12204 4606
rect 12204 4604 12239 4606
rect 12239 4604 12273 4606
rect 12273 4604 12308 4606
rect 12308 4604 12342 4606
rect 12342 4604 12377 4606
rect 12377 4604 12411 4606
rect 12411 4604 12446 4606
rect 12446 4604 12480 4606
rect 12480 4604 12515 4606
rect 12515 4604 12549 4606
rect 12549 4604 12584 4606
rect 12584 4604 12618 4606
rect 12618 4604 12653 4606
rect 12653 4604 12687 4606
rect 12687 4604 12722 4606
rect 12722 4604 12756 4606
rect 12756 4604 12791 4606
rect 12791 4604 12825 4606
rect 12825 4604 12860 4606
rect 12860 4604 12894 4606
rect 12894 4604 12929 4606
rect 12929 4604 12963 4606
rect 12963 4604 12998 4606
rect 12998 4604 13032 4606
rect 13032 4604 13067 4606
rect 13067 4604 13101 4606
rect 13101 4604 13136 4606
rect 13136 4604 13170 4606
rect 13170 4604 13205 4606
rect 13205 4604 13239 4606
rect 13239 4604 13274 4606
rect 13274 4604 13308 4606
rect 13308 4604 13343 4606
rect 13343 4604 13377 4606
rect 13377 4604 13412 4606
rect 13412 4604 13446 4606
rect 13446 4604 13481 4606
rect 13481 4604 13515 4606
rect 13515 4604 13550 4606
rect 13550 4604 13584 4606
rect 13584 4604 13619 4606
rect 13619 4604 13653 4606
rect 13653 4604 13688 4606
rect 13688 4604 13722 4606
rect 13722 4604 13757 4606
rect 13757 4604 13791 4606
rect 13791 4604 13826 4606
rect 13826 4604 13860 4606
rect 13860 4604 13895 4606
rect 13895 4604 13929 4606
rect 13929 4604 13964 4606
rect 13964 4604 13998 4606
rect 13998 4604 14033 4606
rect 14033 4604 14067 4606
rect 14067 4604 14102 4606
rect 14102 4604 14136 4606
rect 14136 4604 14171 4606
rect 14171 4604 14205 4606
rect 14205 4604 14207 4606
rect 14246 4604 14274 4606
rect 14274 4604 14280 4606
rect 14319 4604 14343 4606
rect 14343 4604 14353 4606
rect 14392 4604 14412 4606
rect 14412 4604 14426 4606
rect 10410 4570 14207 4604
rect 14246 4572 14280 4604
rect 14319 4572 14353 4604
rect 14392 4572 14426 4604
rect 709 4500 12363 4570
rect 12363 4536 12397 4570
rect 12397 4536 12431 4570
rect 12431 4536 12466 4570
rect 12466 4536 12500 4570
rect 12500 4536 12535 4570
rect 12535 4536 12569 4570
rect 12569 4536 12604 4570
rect 12604 4536 12638 4570
rect 12638 4536 12673 4570
rect 12673 4536 12707 4570
rect 12707 4536 12742 4570
rect 12742 4536 12776 4570
rect 12776 4536 12811 4570
rect 12811 4536 12845 4570
rect 12845 4536 12880 4570
rect 12880 4536 12914 4570
rect 12914 4536 12949 4570
rect 12949 4536 12983 4570
rect 12983 4536 13018 4570
rect 13018 4536 13052 4570
rect 13052 4536 13087 4570
rect 13087 4536 13121 4570
rect 13121 4536 13156 4570
rect 13156 4536 13190 4570
rect 13190 4536 13225 4570
rect 13225 4536 13259 4570
rect 13259 4536 13294 4570
rect 13294 4536 13328 4570
rect 13328 4536 13363 4570
rect 13363 4536 13397 4570
rect 13397 4536 13432 4570
rect 13432 4536 13466 4570
rect 13466 4536 13501 4570
rect 13501 4536 13535 4570
rect 13535 4536 13570 4570
rect 13570 4536 13604 4570
rect 13604 4536 13639 4570
rect 13639 4536 13673 4570
rect 13673 4536 13708 4570
rect 13708 4536 13742 4570
rect 13742 4536 13777 4570
rect 13777 4536 13811 4570
rect 13811 4536 13846 4570
rect 13846 4536 13880 4570
rect 13880 4536 13915 4570
rect 13915 4536 13949 4570
rect 13949 4536 13984 4570
rect 13984 4536 14018 4570
rect 14018 4536 14053 4570
rect 14053 4536 14087 4570
rect 14087 4536 14122 4570
rect 14122 4536 14156 4570
rect 14156 4536 14191 4570
rect 14191 4536 14207 4570
rect 12363 4502 14207 4536
rect 14246 4502 14280 4534
rect 14319 4502 14353 4534
rect 14392 4502 14426 4534
rect 12363 4500 12398 4502
rect 12398 4500 12432 4502
rect 12432 4500 12467 4502
rect 12467 4500 12501 4502
rect 12501 4500 12536 4502
rect 12536 4500 12570 4502
rect 12570 4500 12605 4502
rect 12605 4500 12639 4502
rect 12639 4500 12674 4502
rect 12674 4500 12708 4502
rect 12708 4500 12743 4502
rect 12743 4500 12777 4502
rect 12777 4500 12812 4502
rect 12812 4500 12846 4502
rect 12846 4500 12881 4502
rect 12881 4500 12915 4502
rect 12915 4500 12950 4502
rect 12950 4500 12984 4502
rect 12984 4500 13019 4502
rect 13019 4500 13053 4502
rect 13053 4500 13088 4502
rect 13088 4500 13122 4502
rect 13122 4500 13157 4502
rect 13157 4500 13191 4502
rect 13191 4500 13226 4502
rect 13226 4500 13260 4502
rect 13260 4500 13295 4502
rect 13295 4500 13329 4502
rect 13329 4500 13364 4502
rect 13364 4500 13398 4502
rect 13398 4500 13433 4502
rect 13433 4500 13467 4502
rect 13467 4500 13502 4502
rect 13502 4500 13536 4502
rect 13536 4500 13571 4502
rect 13571 4500 13605 4502
rect 13605 4500 13640 4502
rect 13640 4500 13674 4502
rect 13674 4500 13709 4502
rect 13709 4500 13743 4502
rect 13743 4500 13778 4502
rect 13778 4500 13812 4502
rect 13812 4500 13847 4502
rect 13847 4500 13881 4502
rect 13881 4500 13916 4502
rect 13916 4500 13950 4502
rect 13950 4500 13985 4502
rect 13985 4500 14019 4502
rect 14019 4500 14054 4502
rect 14054 4500 14088 4502
rect 14088 4500 14123 4502
rect 14123 4500 14157 4502
rect 14157 4500 14192 4502
rect 14192 4500 14207 4502
rect 14246 4500 14261 4502
rect 14261 4500 14280 4502
rect 14319 4500 14330 4502
rect 14330 4500 14353 4502
rect 14392 4500 14399 4502
rect 14399 4500 14426 4502
rect 674 4445 708 4456
rect 529 4409 563 4426
rect 529 4392 531 4409
rect 531 4392 563 4409
rect 601 4395 633 4426
rect 633 4395 635 4426
rect 601 4392 635 4395
rect 529 4339 563 4351
rect 529 4317 531 4339
rect 531 4317 563 4339
rect 601 4322 633 4351
rect 633 4322 635 4351
rect 601 4317 635 4322
rect 529 4269 563 4276
rect 529 4242 531 4269
rect 531 4242 563 4269
rect 601 4249 633 4276
rect 633 4249 635 4276
rect 601 4242 635 4249
rect 529 4199 563 4201
rect 529 4167 531 4199
rect 531 4167 563 4199
rect 601 4177 633 4201
rect 633 4177 635 4201
rect 601 4167 635 4177
rect 529 4095 531 4126
rect 531 4095 563 4126
rect 601 4105 633 4126
rect 633 4105 635 4126
rect 529 4092 563 4095
rect 601 4092 635 4105
rect 529 4025 531 4052
rect 531 4025 563 4052
rect 601 4033 633 4052
rect 633 4033 635 4052
rect 529 4018 563 4025
rect 601 4018 635 4033
rect 529 3955 531 3978
rect 531 3955 563 3978
rect 601 3961 633 3978
rect 633 3961 635 3978
rect 529 3944 563 3955
rect 601 3944 635 3961
rect 529 3886 531 3904
rect 531 3886 563 3904
rect 601 3889 633 3904
rect 633 3889 635 3904
rect 529 3870 563 3886
rect 601 3870 635 3889
rect 529 3760 563 3794
rect 601 3760 635 3794
rect 529 3715 531 3720
rect 531 3715 563 3720
rect 601 3715 633 3720
rect 633 3715 635 3720
rect 529 3686 563 3715
rect 601 3686 635 3715
rect 529 3612 563 3646
rect 601 3612 635 3646
rect 529 3542 563 3572
rect 601 3542 635 3572
rect 529 3538 531 3542
rect 531 3538 563 3542
rect 601 3538 633 3542
rect 633 3538 635 3542
rect 529 3473 563 3498
rect 601 3473 635 3498
rect 529 3464 531 3473
rect 531 3464 563 3473
rect 601 3464 633 3473
rect 633 3464 635 3473
rect 529 3404 563 3424
rect 601 3404 635 3424
rect 529 3390 531 3404
rect 531 3390 563 3404
rect 601 3390 633 3404
rect 633 3390 635 3404
rect 529 3335 563 3350
rect 601 3335 635 3350
rect 529 3316 531 3335
rect 531 3316 563 3335
rect 601 3316 633 3335
rect 633 3316 635 3335
rect 529 3266 563 3276
rect 601 3266 635 3276
rect 529 3242 531 3266
rect 531 3242 563 3266
rect 601 3242 633 3266
rect 633 3242 635 3266
rect 529 3197 563 3202
rect 601 3197 635 3202
rect 529 3168 531 3197
rect 531 3168 563 3197
rect 601 3168 633 3197
rect 633 3168 635 3197
rect 529 3094 531 3128
rect 531 3094 563 3128
rect 601 3094 633 3128
rect 633 3094 635 3128
rect 529 3025 531 3054
rect 531 3025 563 3054
rect 601 3025 633 3054
rect 633 3025 635 3054
rect 529 3020 563 3025
rect 601 3020 635 3025
rect 529 2956 531 2980
rect 531 2956 563 2980
rect 601 2956 633 2980
rect 633 2956 635 2980
rect 529 2946 563 2956
rect 601 2946 635 2956
rect 529 2887 531 2906
rect 531 2887 563 2906
rect 601 2887 633 2906
rect 633 2887 635 2906
rect 529 2872 563 2887
rect 601 2872 635 2887
rect 529 2818 531 2832
rect 531 2818 563 2832
rect 601 2818 633 2832
rect 633 2818 635 2832
rect 529 2798 563 2818
rect 601 2798 635 2818
rect 529 2749 531 2758
rect 531 2749 563 2758
rect 601 2749 633 2758
rect 633 2749 635 2758
rect 529 2724 563 2749
rect 601 2724 635 2749
rect 529 2680 531 2684
rect 531 2680 563 2684
rect 601 2680 633 2684
rect 633 2680 635 2684
rect 529 2650 563 2680
rect 601 2650 635 2680
rect 529 2576 563 2610
rect 601 2576 635 2610
rect 529 2507 563 2536
rect 601 2507 635 2536
rect 529 2502 531 2507
rect 531 2502 563 2507
rect 601 2502 633 2507
rect 633 2502 635 2507
rect 529 2438 563 2462
rect 601 2438 635 2462
rect 529 2428 531 2438
rect 531 2428 563 2438
rect 601 2428 633 2438
rect 633 2428 635 2438
rect 529 2369 563 2389
rect 601 2369 635 2389
rect 529 2355 531 2369
rect 531 2355 563 2369
rect 601 2355 633 2369
rect 633 2355 635 2369
rect 529 2300 563 2316
rect 601 2300 635 2316
rect 529 2282 531 2300
rect 531 2282 563 2300
rect 601 2282 633 2300
rect 633 2282 635 2300
rect 529 2231 563 2243
rect 601 2231 635 2243
rect 529 2209 531 2231
rect 531 2209 563 2231
rect 601 2209 633 2231
rect 633 2209 635 2231
rect 529 2163 563 2170
rect 529 2136 531 2163
rect 531 2136 563 2163
rect 601 2162 635 2170
rect 601 2136 633 2162
rect 633 2136 635 2162
rect 529 2095 563 2097
rect 529 2063 531 2095
rect 531 2063 563 2095
rect 601 2093 635 2097
rect 601 2063 633 2093
rect 633 2063 635 2093
rect 529 1993 531 2024
rect 531 1993 563 2024
rect 529 1990 563 1993
rect 601 1990 633 2024
rect 633 1990 635 2024
rect 529 1925 531 1951
rect 531 1925 563 1951
rect 529 1917 563 1925
rect 601 1921 633 1951
rect 633 1921 635 1951
rect 601 1917 635 1921
rect 529 1857 531 1878
rect 531 1857 563 1878
rect 529 1844 563 1857
rect 601 1852 633 1878
rect 633 1852 635 1878
rect 601 1844 635 1852
rect 529 1789 531 1805
rect 531 1789 563 1805
rect 529 1771 563 1789
rect 601 1783 633 1805
rect 633 1783 635 1805
rect 601 1771 635 1783
rect 529 1721 531 1732
rect 531 1721 563 1732
rect 529 1698 563 1721
rect 601 1714 633 1732
rect 633 1714 635 1732
rect 601 1698 635 1714
rect 529 1653 531 1659
rect 531 1653 563 1659
rect 529 1625 563 1653
rect 601 1645 633 1659
rect 633 1645 635 1659
rect 601 1625 635 1645
rect 529 1585 531 1586
rect 531 1585 563 1586
rect 529 1552 563 1585
rect 601 1576 633 1586
rect 633 1576 635 1586
rect 601 1552 635 1576
rect 529 1483 563 1513
rect 601 1507 633 1513
rect 633 1507 635 1513
rect 529 1479 531 1483
rect 531 1479 563 1483
rect 601 1479 635 1507
rect 529 1415 563 1440
rect 601 1438 633 1440
rect 633 1438 635 1440
rect 529 1406 531 1415
rect 531 1406 563 1415
rect 601 1406 635 1438
rect 529 1347 563 1367
rect 529 1333 531 1347
rect 531 1333 563 1347
rect 601 1334 635 1367
rect 601 1333 633 1334
rect 633 1333 635 1334
rect 529 1279 563 1294
rect 529 1260 531 1279
rect 531 1260 563 1279
rect 601 1265 635 1294
rect 601 1260 633 1265
rect 633 1260 635 1265
rect 529 1211 563 1221
rect 529 1187 531 1211
rect 531 1187 563 1211
rect 601 1196 635 1221
rect 601 1187 633 1196
rect 633 1187 635 1196
rect 529 1143 563 1148
rect 529 1114 531 1143
rect 531 1114 563 1143
rect 601 1127 635 1148
rect 601 1114 633 1127
rect 633 1114 635 1127
rect 529 1041 531 1075
rect 531 1041 563 1075
rect 601 1058 635 1075
rect 601 1041 633 1058
rect 633 1041 635 1058
rect 529 973 531 1002
rect 531 973 563 1002
rect 601 989 635 1002
rect 529 968 563 973
rect 601 968 633 989
rect 633 968 635 989
rect 529 920 531 929
rect 531 920 563 929
rect 601 920 635 929
rect 529 895 563 920
rect 601 895 635 920
rect 674 894 780 4445
rect 14356 4398 14390 4432
rect 14428 4426 14462 4456
rect 14356 4325 14390 4359
rect 1067 4064 1101 4098
rect 1139 4064 1173 4098
rect 1211 4064 1245 4098
rect 1067 3991 1101 4025
rect 1139 3991 1173 4025
rect 1211 3991 1245 4025
rect 1067 3918 1101 3952
rect 1139 3918 1173 3952
rect 1211 3918 1245 3952
rect 1067 3845 1101 3879
rect 1139 3845 1173 3879
rect 1211 3845 1245 3879
rect 1067 3772 1101 3806
rect 1139 3772 1173 3806
rect 1211 3772 1245 3806
rect 1067 3699 1101 3733
rect 1139 3699 1173 3733
rect 1211 3699 1245 3733
rect 1067 3626 1101 3660
rect 1139 3626 1173 3660
rect 1211 3626 1245 3660
rect 1067 3553 1101 3587
rect 1139 3553 1173 3587
rect 1211 3553 1245 3587
rect 1067 3480 1101 3514
rect 1139 3480 1173 3514
rect 1211 3480 1245 3514
rect 1067 3407 1101 3441
rect 1139 3407 1173 3441
rect 1211 3407 1245 3441
rect 1067 3334 1101 3368
rect 1139 3334 1173 3368
rect 1211 3334 1245 3368
rect 1067 3261 1101 3295
rect 1139 3261 1173 3295
rect 1211 3261 1245 3295
rect 1067 3188 1101 3222
rect 1139 3188 1173 3222
rect 1211 3188 1245 3222
rect 1067 3115 1101 3149
rect 1139 3115 1173 3149
rect 1211 3115 1245 3149
rect 1067 3042 1101 3076
rect 1139 3042 1173 3076
rect 1211 3042 1245 3076
rect 1067 2969 1101 3003
rect 1139 2969 1173 3003
rect 1211 2969 1245 3003
rect 1067 2896 1101 2930
rect 1139 2896 1173 2930
rect 1211 2896 1245 2930
rect 1067 2823 1101 2857
rect 1139 2823 1173 2857
rect 1211 2823 1245 2857
rect 1067 2750 1101 2784
rect 1139 2750 1173 2784
rect 1211 2750 1245 2784
rect 1067 2677 1101 2711
rect 1139 2677 1173 2711
rect 1211 2677 1245 2711
rect 1067 2604 1101 2638
rect 1139 2604 1173 2638
rect 1211 2604 1245 2638
rect 1067 2531 1101 2565
rect 1139 2531 1173 2565
rect 1211 2531 1245 2565
rect 1067 2458 1101 2492
rect 1139 2458 1173 2492
rect 1211 2458 1245 2492
rect 1067 2385 1101 2419
rect 1139 2385 1173 2419
rect 1211 2385 1245 2419
rect 1067 2312 1101 2346
rect 1139 2312 1173 2346
rect 1211 2312 1245 2346
rect 1067 2239 1101 2273
rect 1139 2239 1173 2273
rect 1211 2239 1245 2273
rect 1067 2166 1101 2200
rect 1139 2166 1173 2200
rect 1211 2166 1245 2200
rect 1067 2092 1101 2126
rect 1139 2092 1173 2126
rect 1211 2092 1245 2126
rect 1067 2018 1101 2052
rect 1139 2018 1173 2052
rect 1211 2018 1245 2052
rect 1067 1944 1101 1978
rect 1139 1944 1173 1978
rect 1211 1944 1245 1978
rect 1067 1870 1101 1904
rect 1139 1870 1173 1904
rect 1211 1870 1245 1904
rect 1067 1796 1101 1830
rect 1139 1796 1173 1830
rect 1211 1796 1245 1830
rect 1067 1722 1101 1756
rect 1139 1722 1173 1756
rect 1211 1722 1245 1756
rect 1067 1648 1101 1682
rect 1139 1648 1173 1682
rect 1211 1648 1245 1682
rect 1067 1574 1101 1608
rect 1139 1574 1173 1608
rect 1211 1574 1245 1608
rect 924 1216 958 1250
rect 924 1144 958 1178
rect 1563 4058 1597 4092
rect 1707 4058 1741 4092
rect 1563 3986 1597 4020
rect 1707 3986 1741 4020
rect 1563 3914 1597 3948
rect 1707 3914 1741 3948
rect 1563 3842 1597 3876
rect 1707 3842 1741 3876
rect 1563 3770 1597 3804
rect 1707 3770 1741 3804
rect 1563 3698 1597 3732
rect 1707 3698 1741 3732
rect 1563 3626 1597 3660
rect 1707 3626 1741 3660
rect 1563 3554 1597 3588
rect 1707 3554 1741 3588
rect 1563 3482 1597 3516
rect 1707 3482 1741 3516
rect 1563 3410 1597 3444
rect 1707 3410 1741 3444
rect 1563 3338 1597 3372
rect 1707 3338 1741 3372
rect 1563 3266 1597 3300
rect 1707 3266 1741 3300
rect 1563 3194 1597 3228
rect 1707 3194 1741 3228
rect 1563 3074 1597 3108
rect 1635 3074 1669 3108
rect 1707 3074 1741 3108
rect 1563 2994 1597 3028
rect 1635 2994 1669 3028
rect 1707 2994 1741 3028
rect 1563 2914 1597 2948
rect 1635 2914 1669 2948
rect 1707 2914 1741 2948
rect 1563 2834 1597 2868
rect 1635 2834 1669 2868
rect 1707 2834 1741 2868
rect 1563 2754 1597 2788
rect 1635 2754 1669 2788
rect 1707 2754 1741 2788
rect 1563 2674 1597 2708
rect 1635 2674 1669 2708
rect 1707 2674 1741 2708
rect 1563 2594 1597 2628
rect 1635 2594 1669 2628
rect 1707 2594 1741 2628
rect 1563 2484 1597 2518
rect 1707 2484 1741 2518
rect 1563 2412 1597 2446
rect 1707 2412 1741 2446
rect 1563 2340 1597 2374
rect 1707 2340 1741 2374
rect 1563 2268 1597 2302
rect 1707 2268 1741 2302
rect 1563 2196 1597 2230
rect 1707 2196 1741 2230
rect 1563 2124 1597 2158
rect 1707 2124 1741 2158
rect 1563 2052 1597 2086
rect 1707 2052 1741 2086
rect 1563 1980 1597 2014
rect 1707 1980 1741 2014
rect 1563 1908 1597 1942
rect 1707 1908 1741 1942
rect 1563 1836 1597 1870
rect 1707 1836 1741 1870
rect 1563 1764 1597 1798
rect 1707 1764 1741 1798
rect 1563 1692 1597 1726
rect 1707 1692 1741 1726
rect 1563 1620 1597 1654
rect 1707 1620 1741 1654
rect 1318 1144 1424 1250
rect 2059 4064 2093 4098
rect 2131 4064 2165 4098
rect 2203 4064 2237 4098
rect 2059 3991 2093 4025
rect 2131 3991 2165 4025
rect 2203 3991 2237 4025
rect 2059 3918 2093 3952
rect 2131 3918 2165 3952
rect 2203 3918 2237 3952
rect 2059 3845 2093 3879
rect 2131 3845 2165 3879
rect 2203 3845 2237 3879
rect 2059 3772 2093 3806
rect 2131 3772 2165 3806
rect 2203 3772 2237 3806
rect 2059 3699 2093 3733
rect 2131 3699 2165 3733
rect 2203 3699 2237 3733
rect 2059 3626 2093 3660
rect 2131 3626 2165 3660
rect 2203 3626 2237 3660
rect 2059 3553 2093 3587
rect 2131 3553 2165 3587
rect 2203 3553 2237 3587
rect 2059 3480 2093 3514
rect 2131 3480 2165 3514
rect 2203 3480 2237 3514
rect 2059 3407 2093 3441
rect 2131 3407 2165 3441
rect 2203 3407 2237 3441
rect 2059 3334 2093 3368
rect 2131 3334 2165 3368
rect 2203 3334 2237 3368
rect 2059 3261 2093 3295
rect 2131 3261 2165 3295
rect 2203 3261 2237 3295
rect 2059 3188 2093 3222
rect 2131 3188 2165 3222
rect 2203 3188 2237 3222
rect 2059 3115 2093 3149
rect 2131 3115 2165 3149
rect 2203 3115 2237 3149
rect 2059 3042 2093 3076
rect 2131 3042 2165 3076
rect 2203 3042 2237 3076
rect 2059 2969 2093 3003
rect 2131 2969 2165 3003
rect 2203 2969 2237 3003
rect 2059 2896 2093 2930
rect 2131 2896 2165 2930
rect 2203 2896 2237 2930
rect 2059 2823 2093 2857
rect 2131 2823 2165 2857
rect 2203 2823 2237 2857
rect 2059 2750 2093 2784
rect 2131 2750 2165 2784
rect 2203 2750 2237 2784
rect 2059 2677 2093 2711
rect 2131 2677 2165 2711
rect 2203 2677 2237 2711
rect 2059 2604 2093 2638
rect 2131 2604 2165 2638
rect 2203 2604 2237 2638
rect 2059 2531 2093 2565
rect 2131 2531 2165 2565
rect 2203 2531 2237 2565
rect 2059 2458 2093 2492
rect 2131 2458 2165 2492
rect 2203 2458 2237 2492
rect 2059 2385 2093 2419
rect 2131 2385 2165 2419
rect 2203 2385 2237 2419
rect 2059 2312 2093 2346
rect 2131 2312 2165 2346
rect 2203 2312 2237 2346
rect 2059 2239 2093 2273
rect 2131 2239 2165 2273
rect 2203 2239 2237 2273
rect 2059 2166 2093 2200
rect 2131 2166 2165 2200
rect 2203 2166 2237 2200
rect 2059 2092 2093 2126
rect 2131 2092 2165 2126
rect 2203 2092 2237 2126
rect 2059 2018 2093 2052
rect 2131 2018 2165 2052
rect 2203 2018 2237 2052
rect 2059 1944 2093 1978
rect 2131 1944 2165 1978
rect 2203 1944 2237 1978
rect 2059 1870 2093 1904
rect 2131 1870 2165 1904
rect 2203 1870 2237 1904
rect 2059 1796 2093 1830
rect 2131 1796 2165 1830
rect 2203 1796 2237 1830
rect 2059 1722 2093 1756
rect 2131 1722 2165 1756
rect 2203 1722 2237 1756
rect 2059 1648 2093 1682
rect 2131 1648 2165 1682
rect 2203 1648 2237 1682
rect 2059 1574 2093 1608
rect 2131 1574 2165 1608
rect 2203 1574 2237 1608
rect 1880 1144 1986 1250
rect 2555 4058 2589 4092
rect 2699 4058 2733 4092
rect 2555 3986 2589 4020
rect 2699 3986 2733 4020
rect 2555 3914 2589 3948
rect 2699 3914 2733 3948
rect 2555 3842 2589 3876
rect 2699 3842 2733 3876
rect 2555 3770 2589 3804
rect 2699 3770 2733 3804
rect 2555 3698 2589 3732
rect 2699 3698 2733 3732
rect 2555 3626 2589 3660
rect 2699 3626 2733 3660
rect 2555 3554 2589 3588
rect 2699 3554 2733 3588
rect 2555 3482 2589 3516
rect 2699 3482 2733 3516
rect 2555 3410 2589 3444
rect 2699 3410 2733 3444
rect 2555 3338 2589 3372
rect 2699 3338 2733 3372
rect 2555 3266 2589 3300
rect 2699 3266 2733 3300
rect 2555 3194 2589 3228
rect 2699 3194 2733 3228
rect 2555 3074 2589 3108
rect 2627 3074 2661 3108
rect 2699 3074 2733 3108
rect 2555 2994 2589 3028
rect 2627 2994 2661 3028
rect 2699 2994 2733 3028
rect 2555 2914 2589 2948
rect 2627 2914 2661 2948
rect 2699 2914 2733 2948
rect 2555 2834 2589 2868
rect 2627 2834 2661 2868
rect 2699 2834 2733 2868
rect 2555 2754 2589 2788
rect 2627 2754 2661 2788
rect 2699 2754 2733 2788
rect 2555 2674 2589 2708
rect 2627 2674 2661 2708
rect 2699 2674 2733 2708
rect 2555 2594 2589 2628
rect 2627 2594 2661 2628
rect 2699 2594 2733 2628
rect 2555 2484 2589 2518
rect 2699 2484 2733 2518
rect 2555 2412 2589 2446
rect 2699 2412 2733 2446
rect 2555 2340 2589 2374
rect 2699 2340 2733 2374
rect 2555 2268 2589 2302
rect 2699 2268 2733 2302
rect 2555 2196 2589 2230
rect 2699 2196 2733 2230
rect 2555 2124 2589 2158
rect 2699 2124 2733 2158
rect 2555 2052 2589 2086
rect 2699 2052 2733 2086
rect 2555 1980 2589 2014
rect 2699 1980 2733 2014
rect 2555 1908 2589 1942
rect 2699 1908 2733 1942
rect 2555 1836 2589 1870
rect 2699 1836 2733 1870
rect 2555 1764 2589 1798
rect 2699 1764 2733 1798
rect 2555 1692 2589 1726
rect 2699 1692 2733 1726
rect 2555 1620 2589 1654
rect 2699 1620 2733 1654
rect 2310 1144 2416 1250
rect 3051 4064 3085 4098
rect 3123 4064 3157 4098
rect 3195 4064 3229 4098
rect 3051 3991 3085 4025
rect 3123 3991 3157 4025
rect 3195 3991 3229 4025
rect 3051 3918 3085 3952
rect 3123 3918 3157 3952
rect 3195 3918 3229 3952
rect 3051 3845 3085 3879
rect 3123 3845 3157 3879
rect 3195 3845 3229 3879
rect 3051 3772 3085 3806
rect 3123 3772 3157 3806
rect 3195 3772 3229 3806
rect 3051 3699 3085 3733
rect 3123 3699 3157 3733
rect 3195 3699 3229 3733
rect 3051 3626 3085 3660
rect 3123 3626 3157 3660
rect 3195 3626 3229 3660
rect 3051 3553 3085 3587
rect 3123 3553 3157 3587
rect 3195 3553 3229 3587
rect 3051 3480 3085 3514
rect 3123 3480 3157 3514
rect 3195 3480 3229 3514
rect 3051 3407 3085 3441
rect 3123 3407 3157 3441
rect 3195 3407 3229 3441
rect 3051 3334 3085 3368
rect 3123 3334 3157 3368
rect 3195 3334 3229 3368
rect 3051 3261 3085 3295
rect 3123 3261 3157 3295
rect 3195 3261 3229 3295
rect 3051 3188 3085 3222
rect 3123 3188 3157 3222
rect 3195 3188 3229 3222
rect 3051 3115 3085 3149
rect 3123 3115 3157 3149
rect 3195 3115 3229 3149
rect 3051 3042 3085 3076
rect 3123 3042 3157 3076
rect 3195 3042 3229 3076
rect 3051 2969 3085 3003
rect 3123 2969 3157 3003
rect 3195 2969 3229 3003
rect 3051 2896 3085 2930
rect 3123 2896 3157 2930
rect 3195 2896 3229 2930
rect 3051 2823 3085 2857
rect 3123 2823 3157 2857
rect 3195 2823 3229 2857
rect 3051 2750 3085 2784
rect 3123 2750 3157 2784
rect 3195 2750 3229 2784
rect 3051 2677 3085 2711
rect 3123 2677 3157 2711
rect 3195 2677 3229 2711
rect 3051 2604 3085 2638
rect 3123 2604 3157 2638
rect 3195 2604 3229 2638
rect 3051 2531 3085 2565
rect 3123 2531 3157 2565
rect 3195 2531 3229 2565
rect 3051 2458 3085 2492
rect 3123 2458 3157 2492
rect 3195 2458 3229 2492
rect 3051 2385 3085 2419
rect 3123 2385 3157 2419
rect 3195 2385 3229 2419
rect 3051 2312 3085 2346
rect 3123 2312 3157 2346
rect 3195 2312 3229 2346
rect 3051 2239 3085 2273
rect 3123 2239 3157 2273
rect 3195 2239 3229 2273
rect 3051 2166 3085 2200
rect 3123 2166 3157 2200
rect 3195 2166 3229 2200
rect 3051 2092 3085 2126
rect 3123 2092 3157 2126
rect 3195 2092 3229 2126
rect 3051 2018 3085 2052
rect 3123 2018 3157 2052
rect 3195 2018 3229 2052
rect 3051 1944 3085 1978
rect 3123 1944 3157 1978
rect 3195 1944 3229 1978
rect 3051 1870 3085 1904
rect 3123 1870 3157 1904
rect 3195 1870 3229 1904
rect 3051 1796 3085 1830
rect 3123 1796 3157 1830
rect 3195 1796 3229 1830
rect 3051 1722 3085 1756
rect 3123 1722 3157 1756
rect 3195 1722 3229 1756
rect 3051 1648 3085 1682
rect 3123 1648 3157 1682
rect 3195 1648 3229 1682
rect 3051 1574 3085 1608
rect 3123 1574 3157 1608
rect 3195 1574 3229 1608
rect 2872 1144 2978 1250
rect 3547 4058 3581 4092
rect 3691 4058 3725 4092
rect 3547 3986 3581 4020
rect 3691 3986 3725 4020
rect 3547 3914 3581 3948
rect 3691 3914 3725 3948
rect 3547 3842 3581 3876
rect 3691 3842 3725 3876
rect 3547 3770 3581 3804
rect 3691 3770 3725 3804
rect 3547 3698 3581 3732
rect 3691 3698 3725 3732
rect 3547 3626 3581 3660
rect 3691 3626 3725 3660
rect 3547 3554 3581 3588
rect 3691 3554 3725 3588
rect 3547 3482 3581 3516
rect 3691 3482 3725 3516
rect 3547 3410 3581 3444
rect 3691 3410 3725 3444
rect 3547 3338 3581 3372
rect 3691 3338 3725 3372
rect 3547 3266 3581 3300
rect 3691 3266 3725 3300
rect 3547 3194 3581 3228
rect 3691 3194 3725 3228
rect 3547 3074 3581 3108
rect 3619 3074 3653 3108
rect 3691 3074 3725 3108
rect 3547 2994 3581 3028
rect 3619 2994 3653 3028
rect 3691 2994 3725 3028
rect 3547 2914 3581 2948
rect 3619 2914 3653 2948
rect 3691 2914 3725 2948
rect 3547 2834 3581 2868
rect 3619 2834 3653 2868
rect 3691 2834 3725 2868
rect 3547 2754 3581 2788
rect 3619 2754 3653 2788
rect 3691 2754 3725 2788
rect 3547 2674 3581 2708
rect 3619 2674 3653 2708
rect 3691 2674 3725 2708
rect 3547 2594 3581 2628
rect 3619 2594 3653 2628
rect 3691 2594 3725 2628
rect 3547 2484 3581 2518
rect 3691 2484 3725 2518
rect 3547 2412 3581 2446
rect 3691 2412 3725 2446
rect 3547 2340 3581 2374
rect 3691 2340 3725 2374
rect 3547 2268 3581 2302
rect 3691 2268 3725 2302
rect 3547 2196 3581 2230
rect 3691 2196 3725 2230
rect 3547 2124 3581 2158
rect 3691 2124 3725 2158
rect 3547 2052 3581 2086
rect 3691 2052 3725 2086
rect 3547 1980 3581 2014
rect 3691 1980 3725 2014
rect 3547 1908 3581 1942
rect 3691 1908 3725 1942
rect 3547 1836 3581 1870
rect 3691 1836 3725 1870
rect 3547 1764 3581 1798
rect 3691 1764 3725 1798
rect 3547 1692 3581 1726
rect 3691 1692 3725 1726
rect 3547 1620 3581 1654
rect 3691 1620 3725 1654
rect 3302 1144 3408 1250
rect 4043 4064 4077 4098
rect 4115 4064 4149 4098
rect 4187 4064 4221 4098
rect 4043 3991 4077 4025
rect 4115 3991 4149 4025
rect 4187 3991 4221 4025
rect 4043 3918 4077 3952
rect 4115 3918 4149 3952
rect 4187 3918 4221 3952
rect 4043 3845 4077 3879
rect 4115 3845 4149 3879
rect 4187 3845 4221 3879
rect 4043 3772 4077 3806
rect 4115 3772 4149 3806
rect 4187 3772 4221 3806
rect 4043 3699 4077 3733
rect 4115 3699 4149 3733
rect 4187 3699 4221 3733
rect 4043 3626 4077 3660
rect 4115 3626 4149 3660
rect 4187 3626 4221 3660
rect 4043 3553 4077 3587
rect 4115 3553 4149 3587
rect 4187 3553 4221 3587
rect 4043 3480 4077 3514
rect 4115 3480 4149 3514
rect 4187 3480 4221 3514
rect 4043 3407 4077 3441
rect 4115 3407 4149 3441
rect 4187 3407 4221 3441
rect 4043 3334 4077 3368
rect 4115 3334 4149 3368
rect 4187 3334 4221 3368
rect 4043 3261 4077 3295
rect 4115 3261 4149 3295
rect 4187 3261 4221 3295
rect 4043 3188 4077 3222
rect 4115 3188 4149 3222
rect 4187 3188 4221 3222
rect 4043 3115 4077 3149
rect 4115 3115 4149 3149
rect 4187 3115 4221 3149
rect 4043 3042 4077 3076
rect 4115 3042 4149 3076
rect 4187 3042 4221 3076
rect 4043 2969 4077 3003
rect 4115 2969 4149 3003
rect 4187 2969 4221 3003
rect 4043 2896 4077 2930
rect 4115 2896 4149 2930
rect 4187 2896 4221 2930
rect 4043 2823 4077 2857
rect 4115 2823 4149 2857
rect 4187 2823 4221 2857
rect 4043 2750 4077 2784
rect 4115 2750 4149 2784
rect 4187 2750 4221 2784
rect 4043 2677 4077 2711
rect 4115 2677 4149 2711
rect 4187 2677 4221 2711
rect 4043 2604 4077 2638
rect 4115 2604 4149 2638
rect 4187 2604 4221 2638
rect 4043 2531 4077 2565
rect 4115 2531 4149 2565
rect 4187 2531 4221 2565
rect 4043 2458 4077 2492
rect 4115 2458 4149 2492
rect 4187 2458 4221 2492
rect 4043 2385 4077 2419
rect 4115 2385 4149 2419
rect 4187 2385 4221 2419
rect 4043 2312 4077 2346
rect 4115 2312 4149 2346
rect 4187 2312 4221 2346
rect 4043 2239 4077 2273
rect 4115 2239 4149 2273
rect 4187 2239 4221 2273
rect 4043 2166 4077 2200
rect 4115 2166 4149 2200
rect 4187 2166 4221 2200
rect 4043 2092 4077 2126
rect 4115 2092 4149 2126
rect 4187 2092 4221 2126
rect 4043 2018 4077 2052
rect 4115 2018 4149 2052
rect 4187 2018 4221 2052
rect 4043 1944 4077 1978
rect 4115 1944 4149 1978
rect 4187 1944 4221 1978
rect 4043 1870 4077 1904
rect 4115 1870 4149 1904
rect 4187 1870 4221 1904
rect 4043 1796 4077 1830
rect 4115 1796 4149 1830
rect 4187 1796 4221 1830
rect 4043 1722 4077 1756
rect 4115 1722 4149 1756
rect 4187 1722 4221 1756
rect 4043 1648 4077 1682
rect 4115 1648 4149 1682
rect 4187 1648 4221 1682
rect 4043 1574 4077 1608
rect 4115 1574 4149 1608
rect 4187 1574 4221 1608
rect 3864 1144 3970 1250
rect 4539 4058 4573 4092
rect 4683 4058 4717 4092
rect 4539 3986 4573 4020
rect 4683 3986 4717 4020
rect 4539 3914 4573 3948
rect 4683 3914 4717 3948
rect 4539 3842 4573 3876
rect 4683 3842 4717 3876
rect 4539 3770 4573 3804
rect 4683 3770 4717 3804
rect 4539 3698 4573 3732
rect 4683 3698 4717 3732
rect 4539 3626 4573 3660
rect 4683 3626 4717 3660
rect 4539 3554 4573 3588
rect 4683 3554 4717 3588
rect 4539 3482 4573 3516
rect 4683 3482 4717 3516
rect 4539 3410 4573 3444
rect 4683 3410 4717 3444
rect 4539 3338 4573 3372
rect 4683 3338 4717 3372
rect 4539 3266 4573 3300
rect 4683 3266 4717 3300
rect 4539 3194 4573 3228
rect 4683 3194 4717 3228
rect 4539 3074 4573 3108
rect 4611 3074 4645 3108
rect 4683 3074 4717 3108
rect 4539 2994 4573 3028
rect 4611 2994 4645 3028
rect 4683 2994 4717 3028
rect 4539 2914 4573 2948
rect 4611 2914 4645 2948
rect 4683 2914 4717 2948
rect 4539 2834 4573 2868
rect 4611 2834 4645 2868
rect 4683 2834 4717 2868
rect 4539 2754 4573 2788
rect 4611 2754 4645 2788
rect 4683 2754 4717 2788
rect 4539 2674 4573 2708
rect 4611 2674 4645 2708
rect 4683 2674 4717 2708
rect 4539 2594 4573 2628
rect 4611 2594 4645 2628
rect 4683 2594 4717 2628
rect 4539 2484 4573 2518
rect 4683 2484 4717 2518
rect 4539 2412 4573 2446
rect 4683 2412 4717 2446
rect 4539 2340 4573 2374
rect 4683 2340 4717 2374
rect 4539 2268 4573 2302
rect 4683 2268 4717 2302
rect 4539 2196 4573 2230
rect 4683 2196 4717 2230
rect 4539 2124 4573 2158
rect 4683 2124 4717 2158
rect 4539 2052 4573 2086
rect 4683 2052 4717 2086
rect 4539 1980 4573 2014
rect 4683 1980 4717 2014
rect 4539 1908 4573 1942
rect 4683 1908 4717 1942
rect 4539 1836 4573 1870
rect 4683 1836 4717 1870
rect 4539 1764 4573 1798
rect 4683 1764 4717 1798
rect 4539 1692 4573 1726
rect 4683 1692 4717 1726
rect 4539 1620 4573 1654
rect 4683 1620 4717 1654
rect 4294 1144 4400 1250
rect 5035 4064 5069 4098
rect 5107 4064 5141 4098
rect 5179 4064 5213 4098
rect 5035 3991 5069 4025
rect 5107 3991 5141 4025
rect 5179 3991 5213 4025
rect 5035 3918 5069 3952
rect 5107 3918 5141 3952
rect 5179 3918 5213 3952
rect 5035 3845 5069 3879
rect 5107 3845 5141 3879
rect 5179 3845 5213 3879
rect 5035 3772 5069 3806
rect 5107 3772 5141 3806
rect 5179 3772 5213 3806
rect 5035 3699 5069 3733
rect 5107 3699 5141 3733
rect 5179 3699 5213 3733
rect 5035 3626 5069 3660
rect 5107 3626 5141 3660
rect 5179 3626 5213 3660
rect 5035 3553 5069 3587
rect 5107 3553 5141 3587
rect 5179 3553 5213 3587
rect 5035 3480 5069 3514
rect 5107 3480 5141 3514
rect 5179 3480 5213 3514
rect 5035 3407 5069 3441
rect 5107 3407 5141 3441
rect 5179 3407 5213 3441
rect 5035 3334 5069 3368
rect 5107 3334 5141 3368
rect 5179 3334 5213 3368
rect 5035 3261 5069 3295
rect 5107 3261 5141 3295
rect 5179 3261 5213 3295
rect 5035 3188 5069 3222
rect 5107 3188 5141 3222
rect 5179 3188 5213 3222
rect 5035 3115 5069 3149
rect 5107 3115 5141 3149
rect 5179 3115 5213 3149
rect 5035 3042 5069 3076
rect 5107 3042 5141 3076
rect 5179 3042 5213 3076
rect 5035 2969 5069 3003
rect 5107 2969 5141 3003
rect 5179 2969 5213 3003
rect 5035 2896 5069 2930
rect 5107 2896 5141 2930
rect 5179 2896 5213 2930
rect 5035 2823 5069 2857
rect 5107 2823 5141 2857
rect 5179 2823 5213 2857
rect 5035 2750 5069 2784
rect 5107 2750 5141 2784
rect 5179 2750 5213 2784
rect 5035 2677 5069 2711
rect 5107 2677 5141 2711
rect 5179 2677 5213 2711
rect 5035 2604 5069 2638
rect 5107 2604 5141 2638
rect 5179 2604 5213 2638
rect 5035 2531 5069 2565
rect 5107 2531 5141 2565
rect 5179 2531 5213 2565
rect 5035 2458 5069 2492
rect 5107 2458 5141 2492
rect 5179 2458 5213 2492
rect 5035 2385 5069 2419
rect 5107 2385 5141 2419
rect 5179 2385 5213 2419
rect 5035 2312 5069 2346
rect 5107 2312 5141 2346
rect 5179 2312 5213 2346
rect 5035 2239 5069 2273
rect 5107 2239 5141 2273
rect 5179 2239 5213 2273
rect 5035 2166 5069 2200
rect 5107 2166 5141 2200
rect 5179 2166 5213 2200
rect 5035 2092 5069 2126
rect 5107 2092 5141 2126
rect 5179 2092 5213 2126
rect 5035 2018 5069 2052
rect 5107 2018 5141 2052
rect 5179 2018 5213 2052
rect 5035 1944 5069 1978
rect 5107 1944 5141 1978
rect 5179 1944 5213 1978
rect 5035 1870 5069 1904
rect 5107 1870 5141 1904
rect 5179 1870 5213 1904
rect 5035 1796 5069 1830
rect 5107 1796 5141 1830
rect 5179 1796 5213 1830
rect 5035 1722 5069 1756
rect 5107 1722 5141 1756
rect 5179 1722 5213 1756
rect 5035 1648 5069 1682
rect 5107 1648 5141 1682
rect 5179 1648 5213 1682
rect 5035 1574 5069 1608
rect 5107 1574 5141 1608
rect 5179 1574 5213 1608
rect 4856 1144 4962 1250
rect 5531 4058 5565 4092
rect 5675 4058 5709 4092
rect 5531 3986 5565 4020
rect 5675 3986 5709 4020
rect 5531 3914 5565 3948
rect 5675 3914 5709 3948
rect 5531 3842 5565 3876
rect 5675 3842 5709 3876
rect 5531 3770 5565 3804
rect 5675 3770 5709 3804
rect 5531 3698 5565 3732
rect 5675 3698 5709 3732
rect 5531 3626 5565 3660
rect 5675 3626 5709 3660
rect 5531 3554 5565 3588
rect 5675 3554 5709 3588
rect 5531 3482 5565 3516
rect 5675 3482 5709 3516
rect 5531 3410 5565 3444
rect 5675 3410 5709 3444
rect 5531 3338 5565 3372
rect 5675 3338 5709 3372
rect 5531 3266 5565 3300
rect 5675 3266 5709 3300
rect 5531 3194 5565 3228
rect 5675 3194 5709 3228
rect 5531 3074 5565 3108
rect 5603 3074 5637 3108
rect 5675 3074 5709 3108
rect 5531 2994 5565 3028
rect 5603 2994 5637 3028
rect 5675 2994 5709 3028
rect 5531 2914 5565 2948
rect 5603 2914 5637 2948
rect 5675 2914 5709 2948
rect 5531 2834 5565 2868
rect 5603 2834 5637 2868
rect 5675 2834 5709 2868
rect 5531 2754 5565 2788
rect 5603 2754 5637 2788
rect 5675 2754 5709 2788
rect 5531 2674 5565 2708
rect 5603 2674 5637 2708
rect 5675 2674 5709 2708
rect 5531 2594 5565 2628
rect 5603 2594 5637 2628
rect 5675 2594 5709 2628
rect 5531 2484 5565 2518
rect 5675 2484 5709 2518
rect 5531 2412 5565 2446
rect 5675 2412 5709 2446
rect 5531 2340 5565 2374
rect 5675 2340 5709 2374
rect 5531 2268 5565 2302
rect 5675 2268 5709 2302
rect 5531 2196 5565 2230
rect 5675 2196 5709 2230
rect 5531 2124 5565 2158
rect 5675 2124 5709 2158
rect 5531 2052 5565 2086
rect 5675 2052 5709 2086
rect 5531 1980 5565 2014
rect 5675 1980 5709 2014
rect 5531 1908 5565 1942
rect 5675 1908 5709 1942
rect 5531 1836 5565 1870
rect 5675 1836 5709 1870
rect 5531 1764 5565 1798
rect 5675 1764 5709 1798
rect 5531 1692 5565 1726
rect 5675 1692 5709 1726
rect 5531 1620 5565 1654
rect 5675 1620 5709 1654
rect 5286 1144 5392 1250
rect 6027 4064 6061 4098
rect 6099 4064 6133 4098
rect 6171 4064 6205 4098
rect 6027 3991 6061 4025
rect 6099 3991 6133 4025
rect 6171 3991 6205 4025
rect 6027 3918 6061 3952
rect 6099 3918 6133 3952
rect 6171 3918 6205 3952
rect 6027 3845 6061 3879
rect 6099 3845 6133 3879
rect 6171 3845 6205 3879
rect 6027 3772 6061 3806
rect 6099 3772 6133 3806
rect 6171 3772 6205 3806
rect 6027 3699 6061 3733
rect 6099 3699 6133 3733
rect 6171 3699 6205 3733
rect 6027 3626 6061 3660
rect 6099 3626 6133 3660
rect 6171 3626 6205 3660
rect 6027 3553 6061 3587
rect 6099 3553 6133 3587
rect 6171 3553 6205 3587
rect 6027 3480 6061 3514
rect 6099 3480 6133 3514
rect 6171 3480 6205 3514
rect 6027 3407 6061 3441
rect 6099 3407 6133 3441
rect 6171 3407 6205 3441
rect 6027 3334 6061 3368
rect 6099 3334 6133 3368
rect 6171 3334 6205 3368
rect 6027 3261 6061 3295
rect 6099 3261 6133 3295
rect 6171 3261 6205 3295
rect 6027 3188 6061 3222
rect 6099 3188 6133 3222
rect 6171 3188 6205 3222
rect 6027 3115 6061 3149
rect 6099 3115 6133 3149
rect 6171 3115 6205 3149
rect 6027 3042 6061 3076
rect 6099 3042 6133 3076
rect 6171 3042 6205 3076
rect 6027 2969 6061 3003
rect 6099 2969 6133 3003
rect 6171 2969 6205 3003
rect 6027 2896 6061 2930
rect 6099 2896 6133 2930
rect 6171 2896 6205 2930
rect 6027 2823 6061 2857
rect 6099 2823 6133 2857
rect 6171 2823 6205 2857
rect 6027 2750 6061 2784
rect 6099 2750 6133 2784
rect 6171 2750 6205 2784
rect 6027 2677 6061 2711
rect 6099 2677 6133 2711
rect 6171 2677 6205 2711
rect 6027 2604 6061 2638
rect 6099 2604 6133 2638
rect 6171 2604 6205 2638
rect 6027 2531 6061 2565
rect 6099 2531 6133 2565
rect 6171 2531 6205 2565
rect 6027 2458 6061 2492
rect 6099 2458 6133 2492
rect 6171 2458 6205 2492
rect 6027 2385 6061 2419
rect 6099 2385 6133 2419
rect 6171 2385 6205 2419
rect 6027 2312 6061 2346
rect 6099 2312 6133 2346
rect 6171 2312 6205 2346
rect 6027 2239 6061 2273
rect 6099 2239 6133 2273
rect 6171 2239 6205 2273
rect 6027 2166 6061 2200
rect 6099 2166 6133 2200
rect 6171 2166 6205 2200
rect 6027 2092 6061 2126
rect 6099 2092 6133 2126
rect 6171 2092 6205 2126
rect 6027 2018 6061 2052
rect 6099 2018 6133 2052
rect 6171 2018 6205 2052
rect 6027 1944 6061 1978
rect 6099 1944 6133 1978
rect 6171 1944 6205 1978
rect 6027 1870 6061 1904
rect 6099 1870 6133 1904
rect 6171 1870 6205 1904
rect 6027 1796 6061 1830
rect 6099 1796 6133 1830
rect 6171 1796 6205 1830
rect 6027 1722 6061 1756
rect 6099 1722 6133 1756
rect 6171 1722 6205 1756
rect 6027 1648 6061 1682
rect 6099 1648 6133 1682
rect 6171 1648 6205 1682
rect 6027 1574 6061 1608
rect 6099 1574 6133 1608
rect 6171 1574 6205 1608
rect 5848 1144 5954 1250
rect 6523 4058 6557 4092
rect 6667 4058 6701 4092
rect 6523 3986 6557 4020
rect 6667 3986 6701 4020
rect 6523 3914 6557 3948
rect 6667 3914 6701 3948
rect 6523 3842 6557 3876
rect 6667 3842 6701 3876
rect 6523 3770 6557 3804
rect 6667 3770 6701 3804
rect 6523 3698 6557 3732
rect 6667 3698 6701 3732
rect 6523 3626 6557 3660
rect 6667 3626 6701 3660
rect 6523 3554 6557 3588
rect 6667 3554 6701 3588
rect 6523 3482 6557 3516
rect 6667 3482 6701 3516
rect 6523 3410 6557 3444
rect 6667 3410 6701 3444
rect 6523 3338 6557 3372
rect 6667 3338 6701 3372
rect 6523 3266 6557 3300
rect 6667 3266 6701 3300
rect 6523 3194 6557 3228
rect 6667 3194 6701 3228
rect 6523 3074 6557 3108
rect 6595 3074 6629 3108
rect 6667 3074 6701 3108
rect 6523 2994 6557 3028
rect 6595 2994 6629 3028
rect 6667 2994 6701 3028
rect 6523 2914 6557 2948
rect 6595 2914 6629 2948
rect 6667 2914 6701 2948
rect 6523 2834 6557 2868
rect 6595 2834 6629 2868
rect 6667 2834 6701 2868
rect 6523 2754 6557 2788
rect 6595 2754 6629 2788
rect 6667 2754 6701 2788
rect 6523 2674 6557 2708
rect 6595 2674 6629 2708
rect 6667 2674 6701 2708
rect 6523 2594 6557 2628
rect 6595 2594 6629 2628
rect 6667 2594 6701 2628
rect 6523 2484 6557 2518
rect 6667 2484 6701 2518
rect 6523 2412 6557 2446
rect 6667 2412 6701 2446
rect 6523 2340 6557 2374
rect 6667 2340 6701 2374
rect 6523 2268 6557 2302
rect 6667 2268 6701 2302
rect 6523 2196 6557 2230
rect 6667 2196 6701 2230
rect 6523 2124 6557 2158
rect 6667 2124 6701 2158
rect 6523 2052 6557 2086
rect 6667 2052 6701 2086
rect 6523 1980 6557 2014
rect 6667 1980 6701 2014
rect 6523 1908 6557 1942
rect 6667 1908 6701 1942
rect 6523 1836 6557 1870
rect 6667 1836 6701 1870
rect 6523 1764 6557 1798
rect 6667 1764 6701 1798
rect 6523 1692 6557 1726
rect 6667 1692 6701 1726
rect 6523 1620 6557 1654
rect 6667 1620 6701 1654
rect 6278 1144 6384 1250
rect 7019 4064 7053 4098
rect 7091 4064 7125 4098
rect 7163 4064 7197 4098
rect 7019 3991 7053 4025
rect 7091 3991 7125 4025
rect 7163 3991 7197 4025
rect 7019 3918 7053 3952
rect 7091 3918 7125 3952
rect 7163 3918 7197 3952
rect 7019 3845 7053 3879
rect 7091 3845 7125 3879
rect 7163 3845 7197 3879
rect 7019 3772 7053 3806
rect 7091 3772 7125 3806
rect 7163 3772 7197 3806
rect 7019 3699 7053 3733
rect 7091 3699 7125 3733
rect 7163 3699 7197 3733
rect 7019 3626 7053 3660
rect 7091 3626 7125 3660
rect 7163 3626 7197 3660
rect 7019 3553 7053 3587
rect 7091 3553 7125 3587
rect 7163 3553 7197 3587
rect 7019 3480 7053 3514
rect 7091 3480 7125 3514
rect 7163 3480 7197 3514
rect 7019 3407 7053 3441
rect 7091 3407 7125 3441
rect 7163 3407 7197 3441
rect 7019 3334 7053 3368
rect 7091 3334 7125 3368
rect 7163 3334 7197 3368
rect 7019 3261 7053 3295
rect 7091 3261 7125 3295
rect 7163 3261 7197 3295
rect 7019 3188 7053 3222
rect 7091 3188 7125 3222
rect 7163 3188 7197 3222
rect 7019 3115 7053 3149
rect 7091 3115 7125 3149
rect 7163 3115 7197 3149
rect 7019 3042 7053 3076
rect 7091 3042 7125 3076
rect 7163 3042 7197 3076
rect 7019 2969 7053 3003
rect 7091 2969 7125 3003
rect 7163 2969 7197 3003
rect 7019 2896 7053 2930
rect 7091 2896 7125 2930
rect 7163 2896 7197 2930
rect 7019 2823 7053 2857
rect 7091 2823 7125 2857
rect 7163 2823 7197 2857
rect 7019 2750 7053 2784
rect 7091 2750 7125 2784
rect 7163 2750 7197 2784
rect 7019 2677 7053 2711
rect 7091 2677 7125 2711
rect 7163 2677 7197 2711
rect 7019 2604 7053 2638
rect 7091 2604 7125 2638
rect 7163 2604 7197 2638
rect 7019 2531 7053 2565
rect 7091 2531 7125 2565
rect 7163 2531 7197 2565
rect 7019 2458 7053 2492
rect 7091 2458 7125 2492
rect 7163 2458 7197 2492
rect 7019 2385 7053 2419
rect 7091 2385 7125 2419
rect 7163 2385 7197 2419
rect 7019 2312 7053 2346
rect 7091 2312 7125 2346
rect 7163 2312 7197 2346
rect 7019 2239 7053 2273
rect 7091 2239 7125 2273
rect 7163 2239 7197 2273
rect 7019 2166 7053 2200
rect 7091 2166 7125 2200
rect 7163 2166 7197 2200
rect 7019 2092 7053 2126
rect 7091 2092 7125 2126
rect 7163 2092 7197 2126
rect 7019 2018 7053 2052
rect 7091 2018 7125 2052
rect 7163 2018 7197 2052
rect 7019 1944 7053 1978
rect 7091 1944 7125 1978
rect 7163 1944 7197 1978
rect 7019 1870 7053 1904
rect 7091 1870 7125 1904
rect 7163 1870 7197 1904
rect 7019 1796 7053 1830
rect 7091 1796 7125 1830
rect 7163 1796 7197 1830
rect 7019 1722 7053 1756
rect 7091 1722 7125 1756
rect 7163 1722 7197 1756
rect 7019 1648 7053 1682
rect 7091 1648 7125 1682
rect 7163 1648 7197 1682
rect 7019 1574 7053 1608
rect 7091 1574 7125 1608
rect 7163 1574 7197 1608
rect 6840 1144 6946 1250
rect 7515 4058 7549 4092
rect 7659 4058 7693 4092
rect 7515 3986 7549 4020
rect 7659 3986 7693 4020
rect 7515 3914 7549 3948
rect 7659 3914 7693 3948
rect 7515 3842 7549 3876
rect 7659 3842 7693 3876
rect 7515 3770 7549 3804
rect 7659 3770 7693 3804
rect 7515 3698 7549 3732
rect 7659 3698 7693 3732
rect 7515 3626 7549 3660
rect 7659 3626 7693 3660
rect 7515 3554 7549 3588
rect 7659 3554 7693 3588
rect 7515 3482 7549 3516
rect 7659 3482 7693 3516
rect 7515 3410 7549 3444
rect 7659 3410 7693 3444
rect 7515 3338 7549 3372
rect 7659 3338 7693 3372
rect 7515 3266 7549 3300
rect 7659 3266 7693 3300
rect 7515 3194 7549 3228
rect 7659 3194 7693 3228
rect 7515 3074 7549 3108
rect 7587 3074 7621 3108
rect 7659 3074 7693 3108
rect 7515 2994 7549 3028
rect 7587 2994 7621 3028
rect 7659 2994 7693 3028
rect 7515 2914 7549 2948
rect 7587 2914 7621 2948
rect 7659 2914 7693 2948
rect 7515 2834 7549 2868
rect 7587 2834 7621 2868
rect 7659 2834 7693 2868
rect 7515 2754 7549 2788
rect 7587 2754 7621 2788
rect 7659 2754 7693 2788
rect 7515 2674 7549 2708
rect 7587 2674 7621 2708
rect 7659 2674 7693 2708
rect 7515 2594 7549 2628
rect 7587 2594 7621 2628
rect 7659 2594 7693 2628
rect 7515 2484 7549 2518
rect 7659 2484 7693 2518
rect 7515 2412 7549 2446
rect 7659 2412 7693 2446
rect 7515 2340 7549 2374
rect 7659 2340 7693 2374
rect 7515 2268 7549 2302
rect 7659 2268 7693 2302
rect 7515 2196 7549 2230
rect 7659 2196 7693 2230
rect 7515 2124 7549 2158
rect 7659 2124 7693 2158
rect 7515 2052 7549 2086
rect 7659 2052 7693 2086
rect 7515 1980 7549 2014
rect 7659 1980 7693 2014
rect 7515 1908 7549 1942
rect 7659 1908 7693 1942
rect 7515 1836 7549 1870
rect 7659 1836 7693 1870
rect 7515 1764 7549 1798
rect 7659 1764 7693 1798
rect 7515 1692 7549 1726
rect 7659 1692 7693 1726
rect 7515 1620 7549 1654
rect 7659 1620 7693 1654
rect 7270 1144 7376 1250
rect 8011 4064 8045 4098
rect 8083 4064 8117 4098
rect 8155 4064 8189 4098
rect 8011 3991 8045 4025
rect 8083 3991 8117 4025
rect 8155 3991 8189 4025
rect 8011 3918 8045 3952
rect 8083 3918 8117 3952
rect 8155 3918 8189 3952
rect 8011 3845 8045 3879
rect 8083 3845 8117 3879
rect 8155 3845 8189 3879
rect 8011 3772 8045 3806
rect 8083 3772 8117 3806
rect 8155 3772 8189 3806
rect 8011 3699 8045 3733
rect 8083 3699 8117 3733
rect 8155 3699 8189 3733
rect 8011 3626 8045 3660
rect 8083 3626 8117 3660
rect 8155 3626 8189 3660
rect 8011 3553 8045 3587
rect 8083 3553 8117 3587
rect 8155 3553 8189 3587
rect 8011 3480 8045 3514
rect 8083 3480 8117 3514
rect 8155 3480 8189 3514
rect 8011 3407 8045 3441
rect 8083 3407 8117 3441
rect 8155 3407 8189 3441
rect 8011 3334 8045 3368
rect 8083 3334 8117 3368
rect 8155 3334 8189 3368
rect 8011 3261 8045 3295
rect 8083 3261 8117 3295
rect 8155 3261 8189 3295
rect 8011 3188 8045 3222
rect 8083 3188 8117 3222
rect 8155 3188 8189 3222
rect 8011 3115 8045 3149
rect 8083 3115 8117 3149
rect 8155 3115 8189 3149
rect 8011 3042 8045 3076
rect 8083 3042 8117 3076
rect 8155 3042 8189 3076
rect 8011 2969 8045 3003
rect 8083 2969 8117 3003
rect 8155 2969 8189 3003
rect 8011 2896 8045 2930
rect 8083 2896 8117 2930
rect 8155 2896 8189 2930
rect 8011 2823 8045 2857
rect 8083 2823 8117 2857
rect 8155 2823 8189 2857
rect 8011 2750 8045 2784
rect 8083 2750 8117 2784
rect 8155 2750 8189 2784
rect 8011 2677 8045 2711
rect 8083 2677 8117 2711
rect 8155 2677 8189 2711
rect 8011 2604 8045 2638
rect 8083 2604 8117 2638
rect 8155 2604 8189 2638
rect 8011 2531 8045 2565
rect 8083 2531 8117 2565
rect 8155 2531 8189 2565
rect 8011 2458 8045 2492
rect 8083 2458 8117 2492
rect 8155 2458 8189 2492
rect 8011 2385 8045 2419
rect 8083 2385 8117 2419
rect 8155 2385 8189 2419
rect 8011 2312 8045 2346
rect 8083 2312 8117 2346
rect 8155 2312 8189 2346
rect 8011 2239 8045 2273
rect 8083 2239 8117 2273
rect 8155 2239 8189 2273
rect 8011 2166 8045 2200
rect 8083 2166 8117 2200
rect 8155 2166 8189 2200
rect 8011 2092 8045 2126
rect 8083 2092 8117 2126
rect 8155 2092 8189 2126
rect 8011 2018 8045 2052
rect 8083 2018 8117 2052
rect 8155 2018 8189 2052
rect 8011 1944 8045 1978
rect 8083 1944 8117 1978
rect 8155 1944 8189 1978
rect 8011 1870 8045 1904
rect 8083 1870 8117 1904
rect 8155 1870 8189 1904
rect 8011 1796 8045 1830
rect 8083 1796 8117 1830
rect 8155 1796 8189 1830
rect 8011 1722 8045 1756
rect 8083 1722 8117 1756
rect 8155 1722 8189 1756
rect 8011 1648 8045 1682
rect 8083 1648 8117 1682
rect 8155 1648 8189 1682
rect 8011 1574 8045 1608
rect 8083 1574 8117 1608
rect 8155 1574 8189 1608
rect 7832 1144 7938 1250
rect 8507 4058 8541 4092
rect 8651 4058 8685 4092
rect 8507 3986 8541 4020
rect 8651 3986 8685 4020
rect 8507 3914 8541 3948
rect 8651 3914 8685 3948
rect 8507 3842 8541 3876
rect 8651 3842 8685 3876
rect 8507 3770 8541 3804
rect 8651 3770 8685 3804
rect 8507 3698 8541 3732
rect 8651 3698 8685 3732
rect 8507 3626 8541 3660
rect 8651 3626 8685 3660
rect 8507 3554 8541 3588
rect 8651 3554 8685 3588
rect 8507 3482 8541 3516
rect 8651 3482 8685 3516
rect 8507 3410 8541 3444
rect 8651 3410 8685 3444
rect 8507 3338 8541 3372
rect 8651 3338 8685 3372
rect 8507 3266 8541 3300
rect 8651 3266 8685 3300
rect 8507 3194 8541 3228
rect 8651 3194 8685 3228
rect 8507 3074 8541 3108
rect 8579 3074 8613 3108
rect 8651 3074 8685 3108
rect 8507 2994 8541 3028
rect 8579 2994 8613 3028
rect 8651 2994 8685 3028
rect 8507 2914 8541 2948
rect 8579 2914 8613 2948
rect 8651 2914 8685 2948
rect 8507 2834 8541 2868
rect 8579 2834 8613 2868
rect 8651 2834 8685 2868
rect 8507 2754 8541 2788
rect 8579 2754 8613 2788
rect 8651 2754 8685 2788
rect 8507 2674 8541 2708
rect 8579 2674 8613 2708
rect 8651 2674 8685 2708
rect 8507 2594 8541 2628
rect 8579 2594 8613 2628
rect 8651 2594 8685 2628
rect 8507 2484 8541 2518
rect 8651 2484 8685 2518
rect 8507 2412 8541 2446
rect 8651 2412 8685 2446
rect 8507 2340 8541 2374
rect 8651 2340 8685 2374
rect 8507 2268 8541 2302
rect 8651 2268 8685 2302
rect 8507 2196 8541 2230
rect 8651 2196 8685 2230
rect 8507 2124 8541 2158
rect 8651 2124 8685 2158
rect 8507 2052 8541 2086
rect 8651 2052 8685 2086
rect 8507 1980 8541 2014
rect 8651 1980 8685 2014
rect 8507 1908 8541 1942
rect 8651 1908 8685 1942
rect 8507 1836 8541 1870
rect 8651 1836 8685 1870
rect 8507 1764 8541 1798
rect 8651 1764 8685 1798
rect 8507 1692 8541 1726
rect 8651 1692 8685 1726
rect 8507 1620 8541 1654
rect 8651 1620 8685 1654
rect 8262 1144 8368 1250
rect 9003 4064 9037 4098
rect 9075 4064 9109 4098
rect 9147 4064 9181 4098
rect 9003 3991 9037 4025
rect 9075 3991 9109 4025
rect 9147 3991 9181 4025
rect 9003 3918 9037 3952
rect 9075 3918 9109 3952
rect 9147 3918 9181 3952
rect 9003 3845 9037 3879
rect 9075 3845 9109 3879
rect 9147 3845 9181 3879
rect 9003 3772 9037 3806
rect 9075 3772 9109 3806
rect 9147 3772 9181 3806
rect 9003 3699 9037 3733
rect 9075 3699 9109 3733
rect 9147 3699 9181 3733
rect 9003 3626 9037 3660
rect 9075 3626 9109 3660
rect 9147 3626 9181 3660
rect 9003 3553 9037 3587
rect 9075 3553 9109 3587
rect 9147 3553 9181 3587
rect 9003 3480 9037 3514
rect 9075 3480 9109 3514
rect 9147 3480 9181 3514
rect 9003 3407 9037 3441
rect 9075 3407 9109 3441
rect 9147 3407 9181 3441
rect 9003 3334 9037 3368
rect 9075 3334 9109 3368
rect 9147 3334 9181 3368
rect 9003 3261 9037 3295
rect 9075 3261 9109 3295
rect 9147 3261 9181 3295
rect 9003 3188 9037 3222
rect 9075 3188 9109 3222
rect 9147 3188 9181 3222
rect 9003 3115 9037 3149
rect 9075 3115 9109 3149
rect 9147 3115 9181 3149
rect 9003 3042 9037 3076
rect 9075 3042 9109 3076
rect 9147 3042 9181 3076
rect 9003 2969 9037 3003
rect 9075 2969 9109 3003
rect 9147 2969 9181 3003
rect 9003 2896 9037 2930
rect 9075 2896 9109 2930
rect 9147 2896 9181 2930
rect 9003 2823 9037 2857
rect 9075 2823 9109 2857
rect 9147 2823 9181 2857
rect 9003 2750 9037 2784
rect 9075 2750 9109 2784
rect 9147 2750 9181 2784
rect 9003 2677 9037 2711
rect 9075 2677 9109 2711
rect 9147 2677 9181 2711
rect 9003 2604 9037 2638
rect 9075 2604 9109 2638
rect 9147 2604 9181 2638
rect 9003 2531 9037 2565
rect 9075 2531 9109 2565
rect 9147 2531 9181 2565
rect 9003 2458 9037 2492
rect 9075 2458 9109 2492
rect 9147 2458 9181 2492
rect 9003 2385 9037 2419
rect 9075 2385 9109 2419
rect 9147 2385 9181 2419
rect 9003 2312 9037 2346
rect 9075 2312 9109 2346
rect 9147 2312 9181 2346
rect 9003 2239 9037 2273
rect 9075 2239 9109 2273
rect 9147 2239 9181 2273
rect 9003 2166 9037 2200
rect 9075 2166 9109 2200
rect 9147 2166 9181 2200
rect 9003 2092 9037 2126
rect 9075 2092 9109 2126
rect 9147 2092 9181 2126
rect 9003 2018 9037 2052
rect 9075 2018 9109 2052
rect 9147 2018 9181 2052
rect 9003 1944 9037 1978
rect 9075 1944 9109 1978
rect 9147 1944 9181 1978
rect 9003 1870 9037 1904
rect 9075 1870 9109 1904
rect 9147 1870 9181 1904
rect 9003 1796 9037 1830
rect 9075 1796 9109 1830
rect 9147 1796 9181 1830
rect 9003 1722 9037 1756
rect 9075 1722 9109 1756
rect 9147 1722 9181 1756
rect 9003 1648 9037 1682
rect 9075 1648 9109 1682
rect 9147 1648 9181 1682
rect 9003 1574 9037 1608
rect 9075 1574 9109 1608
rect 9147 1574 9181 1608
rect 8824 1144 8930 1250
rect 9499 4058 9533 4092
rect 9643 4058 9677 4092
rect 9499 3986 9533 4020
rect 9643 3986 9677 4020
rect 9499 3914 9533 3948
rect 9643 3914 9677 3948
rect 9499 3842 9533 3876
rect 9643 3842 9677 3876
rect 9499 3770 9533 3804
rect 9643 3770 9677 3804
rect 9499 3698 9533 3732
rect 9643 3698 9677 3732
rect 9499 3626 9533 3660
rect 9643 3626 9677 3660
rect 9499 3554 9533 3588
rect 9643 3554 9677 3588
rect 9499 3482 9533 3516
rect 9643 3482 9677 3516
rect 9499 3410 9533 3444
rect 9643 3410 9677 3444
rect 9499 3338 9533 3372
rect 9643 3338 9677 3372
rect 9499 3266 9533 3300
rect 9643 3266 9677 3300
rect 9499 3194 9533 3228
rect 9643 3194 9677 3228
rect 9499 3074 9533 3108
rect 9571 3074 9605 3108
rect 9643 3074 9677 3108
rect 9499 2994 9533 3028
rect 9571 2994 9605 3028
rect 9643 2994 9677 3028
rect 9499 2914 9533 2948
rect 9571 2914 9605 2948
rect 9643 2914 9677 2948
rect 9499 2834 9533 2868
rect 9571 2834 9605 2868
rect 9643 2834 9677 2868
rect 9499 2754 9533 2788
rect 9571 2754 9605 2788
rect 9643 2754 9677 2788
rect 9499 2674 9533 2708
rect 9571 2674 9605 2708
rect 9643 2674 9677 2708
rect 9499 2594 9533 2628
rect 9571 2594 9605 2628
rect 9643 2594 9677 2628
rect 9499 2484 9533 2518
rect 9643 2484 9677 2518
rect 9499 2412 9533 2446
rect 9643 2412 9677 2446
rect 9499 2340 9533 2374
rect 9643 2340 9677 2374
rect 9499 2268 9533 2302
rect 9643 2268 9677 2302
rect 9499 2196 9533 2230
rect 9643 2196 9677 2230
rect 9499 2124 9533 2158
rect 9643 2124 9677 2158
rect 9499 2052 9533 2086
rect 9643 2052 9677 2086
rect 9499 1980 9533 2014
rect 9643 1980 9677 2014
rect 9499 1908 9533 1942
rect 9643 1908 9677 1942
rect 9499 1836 9533 1870
rect 9643 1836 9677 1870
rect 9499 1764 9533 1798
rect 9643 1764 9677 1798
rect 9499 1692 9533 1726
rect 9643 1692 9677 1726
rect 9499 1620 9533 1654
rect 9643 1620 9677 1654
rect 9254 1144 9360 1250
rect 9995 4064 10029 4098
rect 10067 4064 10101 4098
rect 10139 4064 10173 4098
rect 9995 3991 10029 4025
rect 10067 3991 10101 4025
rect 10139 3991 10173 4025
rect 9995 3918 10029 3952
rect 10067 3918 10101 3952
rect 10139 3918 10173 3952
rect 9995 3845 10029 3879
rect 10067 3845 10101 3879
rect 10139 3845 10173 3879
rect 9995 3772 10029 3806
rect 10067 3772 10101 3806
rect 10139 3772 10173 3806
rect 9995 3699 10029 3733
rect 10067 3699 10101 3733
rect 10139 3699 10173 3733
rect 9995 3626 10029 3660
rect 10067 3626 10101 3660
rect 10139 3626 10173 3660
rect 9995 3553 10029 3587
rect 10067 3553 10101 3587
rect 10139 3553 10173 3587
rect 9995 3480 10029 3514
rect 10067 3480 10101 3514
rect 10139 3480 10173 3514
rect 9995 3407 10029 3441
rect 10067 3407 10101 3441
rect 10139 3407 10173 3441
rect 9995 3334 10029 3368
rect 10067 3334 10101 3368
rect 10139 3334 10173 3368
rect 9995 3261 10029 3295
rect 10067 3261 10101 3295
rect 10139 3261 10173 3295
rect 9995 3188 10029 3222
rect 10067 3188 10101 3222
rect 10139 3188 10173 3222
rect 9995 3115 10029 3149
rect 10067 3115 10101 3149
rect 10139 3115 10173 3149
rect 9995 3042 10029 3076
rect 10067 3042 10101 3076
rect 10139 3042 10173 3076
rect 9995 2969 10029 3003
rect 10067 2969 10101 3003
rect 10139 2969 10173 3003
rect 9995 2896 10029 2930
rect 10067 2896 10101 2930
rect 10139 2896 10173 2930
rect 9995 2823 10029 2857
rect 10067 2823 10101 2857
rect 10139 2823 10173 2857
rect 9995 2750 10029 2784
rect 10067 2750 10101 2784
rect 10139 2750 10173 2784
rect 9995 2677 10029 2711
rect 10067 2677 10101 2711
rect 10139 2677 10173 2711
rect 9995 2604 10029 2638
rect 10067 2604 10101 2638
rect 10139 2604 10173 2638
rect 9995 2531 10029 2565
rect 10067 2531 10101 2565
rect 10139 2531 10173 2565
rect 9995 2458 10029 2492
rect 10067 2458 10101 2492
rect 10139 2458 10173 2492
rect 9995 2385 10029 2419
rect 10067 2385 10101 2419
rect 10139 2385 10173 2419
rect 9995 2312 10029 2346
rect 10067 2312 10101 2346
rect 10139 2312 10173 2346
rect 9995 2239 10029 2273
rect 10067 2239 10101 2273
rect 10139 2239 10173 2273
rect 9995 2166 10029 2200
rect 10067 2166 10101 2200
rect 10139 2166 10173 2200
rect 9995 2092 10029 2126
rect 10067 2092 10101 2126
rect 10139 2092 10173 2126
rect 9995 2018 10029 2052
rect 10067 2018 10101 2052
rect 10139 2018 10173 2052
rect 9995 1944 10029 1978
rect 10067 1944 10101 1978
rect 10139 1944 10173 1978
rect 9995 1870 10029 1904
rect 10067 1870 10101 1904
rect 10139 1870 10173 1904
rect 9995 1796 10029 1830
rect 10067 1796 10101 1830
rect 10139 1796 10173 1830
rect 9995 1722 10029 1756
rect 10067 1722 10101 1756
rect 10139 1722 10173 1756
rect 9995 1648 10029 1682
rect 10067 1648 10101 1682
rect 10139 1648 10173 1682
rect 9995 1574 10029 1608
rect 10067 1574 10101 1608
rect 10139 1574 10173 1608
rect 9816 1144 9922 1250
rect 10491 4058 10525 4092
rect 10635 4058 10669 4092
rect 10491 3986 10525 4020
rect 10635 3986 10669 4020
rect 10491 3914 10525 3948
rect 10635 3914 10669 3948
rect 10491 3842 10525 3876
rect 10635 3842 10669 3876
rect 10491 3770 10525 3804
rect 10635 3770 10669 3804
rect 10491 3698 10525 3732
rect 10635 3698 10669 3732
rect 10491 3626 10525 3660
rect 10635 3626 10669 3660
rect 10491 3554 10525 3588
rect 10635 3554 10669 3588
rect 10491 3482 10525 3516
rect 10635 3482 10669 3516
rect 10491 3410 10525 3444
rect 10635 3410 10669 3444
rect 10491 3338 10525 3372
rect 10635 3338 10669 3372
rect 10491 3266 10525 3300
rect 10635 3266 10669 3300
rect 10491 3194 10525 3228
rect 10635 3194 10669 3228
rect 10491 3074 10525 3108
rect 10563 3074 10597 3108
rect 10635 3074 10669 3108
rect 10491 2994 10525 3028
rect 10563 2994 10597 3028
rect 10635 2994 10669 3028
rect 10491 2914 10525 2948
rect 10563 2914 10597 2948
rect 10635 2914 10669 2948
rect 10491 2834 10525 2868
rect 10563 2834 10597 2868
rect 10635 2834 10669 2868
rect 10491 2754 10525 2788
rect 10563 2754 10597 2788
rect 10635 2754 10669 2788
rect 10491 2674 10525 2708
rect 10563 2674 10597 2708
rect 10635 2674 10669 2708
rect 10491 2594 10525 2628
rect 10563 2594 10597 2628
rect 10635 2594 10669 2628
rect 10491 2484 10525 2518
rect 10635 2484 10669 2518
rect 10491 2412 10525 2446
rect 10635 2412 10669 2446
rect 10491 2340 10525 2374
rect 10635 2340 10669 2374
rect 10491 2268 10525 2302
rect 10635 2268 10669 2302
rect 10491 2196 10525 2230
rect 10635 2196 10669 2230
rect 10491 2124 10525 2158
rect 10635 2124 10669 2158
rect 10491 2052 10525 2086
rect 10635 2052 10669 2086
rect 10491 1980 10525 2014
rect 10635 1980 10669 2014
rect 10491 1908 10525 1942
rect 10635 1908 10669 1942
rect 10491 1836 10525 1870
rect 10635 1836 10669 1870
rect 10491 1764 10525 1798
rect 10635 1764 10669 1798
rect 10491 1692 10525 1726
rect 10635 1692 10669 1726
rect 10491 1620 10525 1654
rect 10635 1620 10669 1654
rect 10246 1144 10352 1250
rect 10987 4064 11021 4098
rect 11059 4064 11093 4098
rect 11131 4064 11165 4098
rect 10987 3991 11021 4025
rect 11059 3991 11093 4025
rect 11131 3991 11165 4025
rect 10987 3918 11021 3952
rect 11059 3918 11093 3952
rect 11131 3918 11165 3952
rect 10987 3845 11021 3879
rect 11059 3845 11093 3879
rect 11131 3845 11165 3879
rect 10987 3772 11021 3806
rect 11059 3772 11093 3806
rect 11131 3772 11165 3806
rect 10987 3699 11021 3733
rect 11059 3699 11093 3733
rect 11131 3699 11165 3733
rect 10987 3626 11021 3660
rect 11059 3626 11093 3660
rect 11131 3626 11165 3660
rect 10987 3553 11021 3587
rect 11059 3553 11093 3587
rect 11131 3553 11165 3587
rect 10987 3480 11021 3514
rect 11059 3480 11093 3514
rect 11131 3480 11165 3514
rect 10987 3407 11021 3441
rect 11059 3407 11093 3441
rect 11131 3407 11165 3441
rect 10987 3334 11021 3368
rect 11059 3334 11093 3368
rect 11131 3334 11165 3368
rect 10987 3261 11021 3295
rect 11059 3261 11093 3295
rect 11131 3261 11165 3295
rect 10987 3188 11021 3222
rect 11059 3188 11093 3222
rect 11131 3188 11165 3222
rect 10987 3115 11021 3149
rect 11059 3115 11093 3149
rect 11131 3115 11165 3149
rect 10987 3042 11021 3076
rect 11059 3042 11093 3076
rect 11131 3042 11165 3076
rect 10987 2969 11021 3003
rect 11059 2969 11093 3003
rect 11131 2969 11165 3003
rect 10987 2896 11021 2930
rect 11059 2896 11093 2930
rect 11131 2896 11165 2930
rect 10987 2823 11021 2857
rect 11059 2823 11093 2857
rect 11131 2823 11165 2857
rect 10987 2750 11021 2784
rect 11059 2750 11093 2784
rect 11131 2750 11165 2784
rect 10987 2677 11021 2711
rect 11059 2677 11093 2711
rect 11131 2677 11165 2711
rect 10987 2604 11021 2638
rect 11059 2604 11093 2638
rect 11131 2604 11165 2638
rect 10987 2531 11021 2565
rect 11059 2531 11093 2565
rect 11131 2531 11165 2565
rect 10987 2458 11021 2492
rect 11059 2458 11093 2492
rect 11131 2458 11165 2492
rect 10987 2385 11021 2419
rect 11059 2385 11093 2419
rect 11131 2385 11165 2419
rect 10987 2312 11021 2346
rect 11059 2312 11093 2346
rect 11131 2312 11165 2346
rect 10987 2239 11021 2273
rect 11059 2239 11093 2273
rect 11131 2239 11165 2273
rect 10987 2166 11021 2200
rect 11059 2166 11093 2200
rect 11131 2166 11165 2200
rect 10987 2092 11021 2126
rect 11059 2092 11093 2126
rect 11131 2092 11165 2126
rect 10987 2018 11021 2052
rect 11059 2018 11093 2052
rect 11131 2018 11165 2052
rect 10987 1944 11021 1978
rect 11059 1944 11093 1978
rect 11131 1944 11165 1978
rect 10987 1870 11021 1904
rect 11059 1870 11093 1904
rect 11131 1870 11165 1904
rect 10987 1796 11021 1830
rect 11059 1796 11093 1830
rect 11131 1796 11165 1830
rect 10987 1722 11021 1756
rect 11059 1722 11093 1756
rect 11131 1722 11165 1756
rect 10987 1648 11021 1682
rect 11059 1648 11093 1682
rect 11131 1648 11165 1682
rect 10987 1574 11021 1608
rect 11059 1574 11093 1608
rect 11131 1574 11165 1608
rect 10808 1144 10914 1250
rect 11483 4058 11517 4092
rect 11627 4058 11661 4092
rect 11483 3986 11517 4020
rect 11627 3986 11661 4020
rect 11483 3914 11517 3948
rect 11627 3914 11661 3948
rect 11483 3842 11517 3876
rect 11627 3842 11661 3876
rect 11483 3770 11517 3804
rect 11627 3770 11661 3804
rect 11483 3698 11517 3732
rect 11627 3698 11661 3732
rect 11483 3626 11517 3660
rect 11627 3626 11661 3660
rect 11483 3554 11517 3588
rect 11627 3554 11661 3588
rect 11483 3482 11517 3516
rect 11627 3482 11661 3516
rect 11483 3410 11517 3444
rect 11627 3410 11661 3444
rect 11483 3338 11517 3372
rect 11627 3338 11661 3372
rect 11483 3266 11517 3300
rect 11627 3266 11661 3300
rect 11483 3194 11517 3228
rect 11627 3194 11661 3228
rect 11483 3074 11517 3108
rect 11555 3074 11589 3108
rect 11627 3074 11661 3108
rect 11483 2994 11517 3028
rect 11555 2994 11589 3028
rect 11627 2994 11661 3028
rect 11483 2914 11517 2948
rect 11555 2914 11589 2948
rect 11627 2914 11661 2948
rect 11483 2834 11517 2868
rect 11555 2834 11589 2868
rect 11627 2834 11661 2868
rect 11483 2754 11517 2788
rect 11555 2754 11589 2788
rect 11627 2754 11661 2788
rect 11483 2674 11517 2708
rect 11555 2674 11589 2708
rect 11627 2674 11661 2708
rect 11483 2594 11517 2628
rect 11555 2594 11589 2628
rect 11627 2594 11661 2628
rect 11483 2484 11517 2518
rect 11627 2484 11661 2518
rect 11483 2412 11517 2446
rect 11627 2412 11661 2446
rect 11483 2340 11517 2374
rect 11627 2340 11661 2374
rect 11483 2268 11517 2302
rect 11627 2268 11661 2302
rect 11483 2196 11517 2230
rect 11627 2196 11661 2230
rect 11483 2124 11517 2158
rect 11627 2124 11661 2158
rect 11483 2052 11517 2086
rect 11627 2052 11661 2086
rect 11483 1980 11517 2014
rect 11627 1980 11661 2014
rect 11483 1908 11517 1942
rect 11627 1908 11661 1942
rect 11483 1836 11517 1870
rect 11627 1836 11661 1870
rect 11483 1764 11517 1798
rect 11627 1764 11661 1798
rect 11483 1692 11517 1726
rect 11627 1692 11661 1726
rect 11483 1620 11517 1654
rect 11627 1620 11661 1654
rect 11238 1144 11344 1250
rect 11979 4064 12013 4098
rect 12051 4064 12085 4098
rect 12123 4064 12157 4098
rect 11979 3991 12013 4025
rect 12051 3991 12085 4025
rect 12123 3991 12157 4025
rect 11979 3918 12013 3952
rect 12051 3918 12085 3952
rect 12123 3918 12157 3952
rect 11979 3845 12013 3879
rect 12051 3845 12085 3879
rect 12123 3845 12157 3879
rect 11979 3772 12013 3806
rect 12051 3772 12085 3806
rect 12123 3772 12157 3806
rect 11979 3699 12013 3733
rect 12051 3699 12085 3733
rect 12123 3699 12157 3733
rect 11979 3626 12013 3660
rect 12051 3626 12085 3660
rect 12123 3626 12157 3660
rect 11979 3553 12013 3587
rect 12051 3553 12085 3587
rect 12123 3553 12157 3587
rect 11979 3480 12013 3514
rect 12051 3480 12085 3514
rect 12123 3480 12157 3514
rect 11979 3407 12013 3441
rect 12051 3407 12085 3441
rect 12123 3407 12157 3441
rect 11979 3334 12013 3368
rect 12051 3334 12085 3368
rect 12123 3334 12157 3368
rect 11979 3261 12013 3295
rect 12051 3261 12085 3295
rect 12123 3261 12157 3295
rect 11979 3188 12013 3222
rect 12051 3188 12085 3222
rect 12123 3188 12157 3222
rect 11979 3115 12013 3149
rect 12051 3115 12085 3149
rect 12123 3115 12157 3149
rect 11979 3042 12013 3076
rect 12051 3042 12085 3076
rect 12123 3042 12157 3076
rect 11979 2969 12013 3003
rect 12051 2969 12085 3003
rect 12123 2969 12157 3003
rect 11979 2896 12013 2930
rect 12051 2896 12085 2930
rect 12123 2896 12157 2930
rect 11979 2823 12013 2857
rect 12051 2823 12085 2857
rect 12123 2823 12157 2857
rect 11979 2750 12013 2784
rect 12051 2750 12085 2784
rect 12123 2750 12157 2784
rect 11979 2677 12013 2711
rect 12051 2677 12085 2711
rect 12123 2677 12157 2711
rect 11979 2604 12013 2638
rect 12051 2604 12085 2638
rect 12123 2604 12157 2638
rect 11979 2531 12013 2565
rect 12051 2531 12085 2565
rect 12123 2531 12157 2565
rect 11979 2458 12013 2492
rect 12051 2458 12085 2492
rect 12123 2458 12157 2492
rect 11979 2385 12013 2419
rect 12051 2385 12085 2419
rect 12123 2385 12157 2419
rect 11979 2312 12013 2346
rect 12051 2312 12085 2346
rect 12123 2312 12157 2346
rect 11979 2239 12013 2273
rect 12051 2239 12085 2273
rect 12123 2239 12157 2273
rect 11979 2166 12013 2200
rect 12051 2166 12085 2200
rect 12123 2166 12157 2200
rect 11979 2092 12013 2126
rect 12051 2092 12085 2126
rect 12123 2092 12157 2126
rect 11979 2018 12013 2052
rect 12051 2018 12085 2052
rect 12123 2018 12157 2052
rect 11979 1944 12013 1978
rect 12051 1944 12085 1978
rect 12123 1944 12157 1978
rect 11979 1870 12013 1904
rect 12051 1870 12085 1904
rect 12123 1870 12157 1904
rect 11979 1796 12013 1830
rect 12051 1796 12085 1830
rect 12123 1796 12157 1830
rect 11979 1722 12013 1756
rect 12051 1722 12085 1756
rect 12123 1722 12157 1756
rect 11979 1648 12013 1682
rect 12051 1648 12085 1682
rect 12123 1648 12157 1682
rect 11979 1574 12013 1608
rect 12051 1574 12085 1608
rect 12123 1574 12157 1608
rect 11800 1144 11906 1250
rect 12475 4058 12509 4092
rect 12619 4058 12653 4092
rect 12475 3986 12509 4020
rect 12619 3986 12653 4020
rect 12475 3914 12509 3948
rect 12619 3914 12653 3948
rect 12475 3842 12509 3876
rect 12619 3842 12653 3876
rect 12475 3770 12509 3804
rect 12619 3770 12653 3804
rect 12475 3698 12509 3732
rect 12619 3698 12653 3732
rect 12475 3626 12509 3660
rect 12619 3626 12653 3660
rect 12475 3554 12509 3588
rect 12619 3554 12653 3588
rect 12475 3482 12509 3516
rect 12619 3482 12653 3516
rect 12475 3410 12509 3444
rect 12619 3410 12653 3444
rect 12475 3338 12509 3372
rect 12619 3338 12653 3372
rect 12475 3266 12509 3300
rect 12619 3266 12653 3300
rect 12475 3194 12509 3228
rect 12619 3194 12653 3228
rect 12475 3074 12509 3108
rect 12547 3074 12581 3108
rect 12619 3074 12653 3108
rect 12475 2994 12509 3028
rect 12547 2994 12581 3028
rect 12619 2994 12653 3028
rect 12475 2914 12509 2948
rect 12547 2914 12581 2948
rect 12619 2914 12653 2948
rect 12475 2834 12509 2868
rect 12547 2834 12581 2868
rect 12619 2834 12653 2868
rect 12475 2754 12509 2788
rect 12547 2754 12581 2788
rect 12619 2754 12653 2788
rect 12475 2674 12509 2708
rect 12547 2674 12581 2708
rect 12619 2674 12653 2708
rect 12475 2594 12509 2628
rect 12547 2594 12581 2628
rect 12619 2594 12653 2628
rect 12475 2484 12509 2518
rect 12619 2484 12653 2518
rect 12475 2412 12509 2446
rect 12619 2412 12653 2446
rect 12475 2340 12509 2374
rect 12619 2340 12653 2374
rect 12475 2268 12509 2302
rect 12619 2268 12653 2302
rect 12475 2196 12509 2230
rect 12619 2196 12653 2230
rect 12475 2124 12509 2158
rect 12619 2124 12653 2158
rect 12475 2052 12509 2086
rect 12619 2052 12653 2086
rect 12475 1980 12509 2014
rect 12619 1980 12653 2014
rect 12475 1908 12509 1942
rect 12619 1908 12653 1942
rect 12475 1836 12509 1870
rect 12619 1836 12653 1870
rect 12475 1764 12509 1798
rect 12619 1764 12653 1798
rect 12475 1692 12509 1726
rect 12619 1692 12653 1726
rect 12475 1620 12509 1654
rect 12619 1620 12653 1654
rect 12230 1144 12336 1250
rect 12971 4064 13005 4098
rect 13043 4064 13077 4098
rect 13115 4064 13149 4098
rect 12971 3991 13005 4025
rect 13043 3991 13077 4025
rect 13115 3991 13149 4025
rect 12971 3918 13005 3952
rect 13043 3918 13077 3952
rect 13115 3918 13149 3952
rect 12971 3845 13005 3879
rect 13043 3845 13077 3879
rect 13115 3845 13149 3879
rect 12971 3772 13005 3806
rect 13043 3772 13077 3806
rect 13115 3772 13149 3806
rect 12971 3699 13005 3733
rect 13043 3699 13077 3733
rect 13115 3699 13149 3733
rect 12971 3626 13005 3660
rect 13043 3626 13077 3660
rect 13115 3626 13149 3660
rect 12971 3553 13005 3587
rect 13043 3553 13077 3587
rect 13115 3553 13149 3587
rect 12971 3480 13005 3514
rect 13043 3480 13077 3514
rect 13115 3480 13149 3514
rect 12971 3407 13005 3441
rect 13043 3407 13077 3441
rect 13115 3407 13149 3441
rect 12971 3334 13005 3368
rect 13043 3334 13077 3368
rect 13115 3334 13149 3368
rect 12971 3261 13005 3295
rect 13043 3261 13077 3295
rect 13115 3261 13149 3295
rect 12971 3188 13005 3222
rect 13043 3188 13077 3222
rect 13115 3188 13149 3222
rect 12971 3115 13005 3149
rect 13043 3115 13077 3149
rect 13115 3115 13149 3149
rect 12971 3042 13005 3076
rect 13043 3042 13077 3076
rect 13115 3042 13149 3076
rect 12971 2969 13005 3003
rect 13043 2969 13077 3003
rect 13115 2969 13149 3003
rect 12971 2896 13005 2930
rect 13043 2896 13077 2930
rect 13115 2896 13149 2930
rect 12971 2823 13005 2857
rect 13043 2823 13077 2857
rect 13115 2823 13149 2857
rect 12971 2750 13005 2784
rect 13043 2750 13077 2784
rect 13115 2750 13149 2784
rect 12971 2677 13005 2711
rect 13043 2677 13077 2711
rect 13115 2677 13149 2711
rect 12971 2604 13005 2638
rect 13043 2604 13077 2638
rect 13115 2604 13149 2638
rect 12971 2531 13005 2565
rect 13043 2531 13077 2565
rect 13115 2531 13149 2565
rect 12971 2458 13005 2492
rect 13043 2458 13077 2492
rect 13115 2458 13149 2492
rect 12971 2385 13005 2419
rect 13043 2385 13077 2419
rect 13115 2385 13149 2419
rect 12971 2312 13005 2346
rect 13043 2312 13077 2346
rect 13115 2312 13149 2346
rect 12971 2239 13005 2273
rect 13043 2239 13077 2273
rect 13115 2239 13149 2273
rect 12971 2166 13005 2200
rect 13043 2166 13077 2200
rect 13115 2166 13149 2200
rect 12971 2092 13005 2126
rect 13043 2092 13077 2126
rect 13115 2092 13149 2126
rect 12971 2018 13005 2052
rect 13043 2018 13077 2052
rect 13115 2018 13149 2052
rect 12971 1944 13005 1978
rect 13043 1944 13077 1978
rect 13115 1944 13149 1978
rect 12971 1870 13005 1904
rect 13043 1870 13077 1904
rect 13115 1870 13149 1904
rect 12971 1796 13005 1830
rect 13043 1796 13077 1830
rect 13115 1796 13149 1830
rect 12971 1722 13005 1756
rect 13043 1722 13077 1756
rect 13115 1722 13149 1756
rect 12971 1648 13005 1682
rect 13043 1648 13077 1682
rect 13115 1648 13149 1682
rect 12971 1574 13005 1608
rect 13043 1574 13077 1608
rect 13115 1574 13149 1608
rect 12792 1144 12898 1250
rect 13467 4058 13501 4092
rect 13611 4058 13645 4092
rect 13467 3986 13501 4020
rect 13611 3986 13645 4020
rect 13467 3914 13501 3948
rect 13611 3914 13645 3948
rect 13467 3842 13501 3876
rect 13611 3842 13645 3876
rect 13467 3770 13501 3804
rect 13611 3770 13645 3804
rect 13467 3698 13501 3732
rect 13611 3698 13645 3732
rect 13467 3626 13501 3660
rect 13611 3626 13645 3660
rect 13467 3554 13501 3588
rect 13611 3554 13645 3588
rect 13467 3482 13501 3516
rect 13611 3482 13645 3516
rect 13467 3410 13501 3444
rect 13611 3410 13645 3444
rect 13467 3338 13501 3372
rect 13611 3338 13645 3372
rect 13467 3266 13501 3300
rect 13611 3266 13645 3300
rect 13467 3194 13501 3228
rect 13611 3194 13645 3228
rect 13467 3074 13501 3108
rect 13539 3074 13573 3108
rect 13611 3074 13645 3108
rect 13467 2994 13501 3028
rect 13539 2994 13573 3028
rect 13611 2994 13645 3028
rect 13467 2914 13501 2948
rect 13539 2914 13573 2948
rect 13611 2914 13645 2948
rect 13467 2834 13501 2868
rect 13539 2834 13573 2868
rect 13611 2834 13645 2868
rect 13467 2754 13501 2788
rect 13539 2754 13573 2788
rect 13611 2754 13645 2788
rect 13467 2674 13501 2708
rect 13539 2674 13573 2708
rect 13611 2674 13645 2708
rect 13467 2594 13501 2628
rect 13539 2594 13573 2628
rect 13611 2594 13645 2628
rect 13467 2484 13501 2518
rect 13611 2484 13645 2518
rect 13467 2412 13501 2446
rect 13611 2412 13645 2446
rect 13467 2340 13501 2374
rect 13611 2340 13645 2374
rect 13467 2268 13501 2302
rect 13611 2268 13645 2302
rect 13467 2196 13501 2230
rect 13611 2196 13645 2230
rect 13467 2124 13501 2158
rect 13611 2124 13645 2158
rect 13467 2052 13501 2086
rect 13611 2052 13645 2086
rect 13467 1980 13501 2014
rect 13611 1980 13645 2014
rect 13467 1908 13501 1942
rect 13611 1908 13645 1942
rect 13467 1836 13501 1870
rect 13611 1836 13645 1870
rect 13467 1764 13501 1798
rect 13611 1764 13645 1798
rect 13467 1692 13501 1726
rect 13611 1692 13645 1726
rect 13467 1620 13501 1654
rect 13611 1620 13645 1654
rect 13222 1144 13328 1250
rect 13999 4064 14033 4098
rect 13999 3991 14033 4025
rect 13999 3918 14033 3952
rect 13999 3845 14033 3879
rect 13999 3772 14033 3806
rect 13999 3699 14033 3733
rect 13999 3626 14033 3660
rect 13999 3553 14033 3587
rect 13999 3480 14033 3514
rect 13999 3407 14033 3441
rect 13999 3334 14033 3368
rect 13999 3261 14033 3295
rect 13999 3188 14033 3222
rect 13999 3115 14033 3149
rect 13999 3042 14033 3076
rect 13999 2969 14033 3003
rect 13999 2896 14033 2930
rect 13999 2823 14033 2857
rect 13999 2750 14033 2784
rect 13999 2677 14033 2711
rect 13999 2604 14033 2638
rect 13999 2531 14033 2565
rect 13999 2458 14033 2492
rect 13999 2385 14033 2419
rect 13999 2312 14033 2346
rect 13999 2239 14033 2273
rect 13999 2166 14033 2200
rect 13999 2092 14033 2126
rect 13999 2018 14033 2052
rect 13999 1944 14033 1978
rect 13999 1870 14033 1904
rect 13999 1796 14033 1830
rect 13999 1722 14033 1756
rect 13999 1648 14033 1682
rect 13999 1574 14033 1608
rect 13784 1144 13890 1250
rect 14142 1144 14248 1250
rect 14356 4252 14390 4286
rect 14356 4179 14390 4213
rect 14356 4106 14390 4140
rect 14356 4033 14390 4067
rect 14356 3960 14390 3994
rect 14428 3992 14468 4426
rect 14468 3992 14606 4426
rect 14428 3960 14536 3992
rect 14536 3960 14606 3992
rect 14356 3887 14390 3921
rect 14428 3918 14462 3952
rect 14500 3888 14534 3921
rect 14572 3905 14604 3921
rect 14604 3905 14606 3921
rect 14500 3887 14502 3888
rect 14502 3887 14534 3888
rect 14356 3814 14390 3848
rect 14428 3846 14462 3880
rect 14572 3887 14606 3905
rect 14500 3819 14534 3848
rect 14572 3837 14604 3848
rect 14604 3837 14606 3848
rect 14500 3814 14502 3819
rect 14502 3814 14534 3819
rect 14356 3741 14390 3775
rect 14428 3774 14462 3808
rect 14572 3814 14606 3837
rect 14500 3750 14534 3775
rect 14572 3769 14604 3775
rect 14604 3769 14606 3775
rect 14500 3741 14502 3750
rect 14502 3741 14534 3750
rect 14428 3702 14462 3736
rect 14572 3741 14606 3769
rect 14356 3668 14390 3702
rect 14500 3681 14534 3702
rect 14572 3701 14604 3702
rect 14604 3701 14606 3702
rect 14500 3668 14502 3681
rect 14502 3668 14534 3681
rect 14428 3630 14462 3664
rect 14572 3668 14606 3701
rect 14356 3595 14390 3629
rect 14500 3612 14534 3629
rect 14500 3595 14502 3612
rect 14502 3595 14534 3612
rect 14428 3558 14462 3592
rect 14572 3599 14606 3629
rect 14572 3595 14604 3599
rect 14604 3595 14606 3599
rect 14356 3522 14390 3556
rect 14500 3543 14534 3556
rect 14500 3522 14502 3543
rect 14502 3522 14534 3543
rect 14428 3486 14462 3520
rect 14572 3531 14606 3556
rect 14572 3522 14604 3531
rect 14604 3522 14606 3531
rect 14356 3449 14390 3483
rect 14500 3474 14534 3483
rect 14500 3449 14502 3474
rect 14502 3449 14534 3474
rect 14428 3414 14462 3448
rect 14572 3463 14606 3483
rect 14572 3449 14604 3463
rect 14604 3449 14606 3463
rect 14356 3376 14390 3410
rect 14500 3405 14534 3410
rect 14500 3376 14502 3405
rect 14502 3376 14534 3405
rect 14428 3342 14462 3376
rect 14572 3395 14606 3410
rect 14572 3376 14604 3395
rect 14604 3376 14606 3395
rect 14356 3303 14390 3337
rect 14500 3336 14534 3337
rect 14428 3270 14462 3304
rect 14500 3303 14502 3336
rect 14502 3303 14534 3336
rect 14572 3327 14606 3337
rect 14572 3303 14604 3327
rect 14604 3303 14606 3327
rect 14356 3230 14390 3264
rect 14500 3233 14502 3264
rect 14502 3233 14534 3264
rect 14572 3259 14606 3264
rect 14428 3198 14462 3232
rect 14500 3230 14534 3233
rect 14572 3230 14604 3259
rect 14604 3230 14606 3259
rect 14356 3157 14390 3191
rect 14500 3164 14502 3191
rect 14502 3164 14534 3191
rect 14428 3126 14462 3160
rect 14500 3157 14534 3164
rect 14572 3157 14604 3191
rect 14604 3157 14606 3191
rect 14356 3084 14390 3118
rect 14500 3095 14502 3118
rect 14502 3095 14534 3118
rect 14428 3054 14462 3088
rect 14500 3084 14534 3095
rect 14572 3089 14604 3118
rect 14604 3089 14606 3118
rect 14572 3084 14606 3089
rect 14356 3011 14390 3045
rect 14500 3026 14502 3045
rect 14502 3026 14534 3045
rect 14428 2982 14462 3016
rect 14500 3011 14534 3026
rect 14572 3021 14604 3045
rect 14604 3021 14606 3045
rect 14572 3011 14606 3021
rect 14356 2938 14390 2972
rect 14500 2957 14502 2972
rect 14502 2957 14534 2972
rect 14428 2910 14462 2944
rect 14500 2938 14534 2957
rect 14572 2953 14604 2972
rect 14604 2953 14606 2972
rect 14572 2938 14606 2953
rect 14356 2865 14390 2899
rect 14500 2888 14502 2899
rect 14502 2888 14534 2899
rect 14428 2838 14462 2872
rect 14500 2865 14534 2888
rect 14572 2885 14604 2899
rect 14604 2885 14606 2899
rect 14572 2865 14606 2885
rect 14356 2792 14390 2826
rect 14500 2819 14502 2826
rect 14502 2819 14534 2826
rect 14428 2766 14462 2800
rect 14500 2792 14534 2819
rect 14572 2817 14604 2826
rect 14604 2817 14606 2826
rect 14572 2792 14606 2817
rect 14356 2719 14390 2753
rect 14500 2750 14502 2753
rect 14502 2750 14534 2753
rect 14428 2694 14462 2728
rect 14500 2719 14534 2750
rect 14572 2749 14604 2753
rect 14604 2749 14606 2753
rect 14572 2719 14606 2749
rect 14356 2646 14390 2680
rect 14428 2622 14462 2656
rect 14500 2646 14534 2680
rect 14572 2647 14606 2680
rect 14572 2646 14604 2647
rect 14604 2646 14606 2647
rect 14356 2573 14390 2607
rect 14428 2550 14462 2584
rect 14500 2577 14534 2607
rect 14572 2579 14606 2607
rect 14500 2573 14502 2577
rect 14502 2573 14534 2577
rect 14572 2573 14604 2579
rect 14604 2573 14606 2579
rect 14356 2500 14390 2534
rect 14428 2478 14462 2512
rect 14500 2508 14534 2534
rect 14572 2511 14606 2534
rect 14500 2500 14502 2508
rect 14502 2500 14534 2508
rect 14572 2500 14604 2511
rect 14604 2500 14606 2511
rect 14356 2427 14390 2461
rect 14428 2406 14462 2440
rect 14500 2439 14534 2461
rect 14572 2443 14606 2461
rect 14500 2427 14502 2439
rect 14502 2427 14534 2439
rect 14572 2427 14604 2443
rect 14604 2427 14606 2443
rect 14356 2354 14390 2388
rect 14500 2370 14534 2388
rect 14572 2375 14606 2388
rect 14428 2334 14462 2368
rect 14500 2354 14502 2370
rect 14502 2354 14534 2370
rect 14572 2354 14604 2375
rect 14604 2354 14606 2375
rect 14356 2281 14390 2315
rect 14500 2301 14534 2315
rect 14572 2307 14606 2315
rect 14428 2262 14462 2296
rect 14500 2281 14502 2301
rect 14502 2281 14534 2301
rect 14572 2281 14604 2307
rect 14604 2281 14606 2307
rect 14356 2208 14390 2242
rect 14500 2232 14534 2242
rect 14572 2239 14606 2242
rect 14428 2190 14462 2224
rect 14500 2208 14502 2232
rect 14502 2208 14534 2232
rect 14572 2208 14604 2239
rect 14604 2208 14606 2239
rect 14356 2135 14390 2169
rect 14500 2163 14534 2169
rect 14428 2118 14462 2152
rect 14500 2135 14502 2163
rect 14502 2135 14534 2163
rect 14572 2137 14604 2169
rect 14604 2137 14606 2169
rect 14572 2135 14606 2137
rect 14356 2062 14390 2096
rect 14500 2094 14534 2096
rect 14428 2046 14462 2080
rect 14500 2062 14502 2094
rect 14502 2062 14534 2094
rect 14572 2069 14604 2096
rect 14604 2069 14606 2096
rect 14572 2062 14606 2069
rect 14356 1989 14390 2023
rect 14428 1974 14462 2008
rect 14500 1991 14502 2023
rect 14502 1991 14534 2023
rect 14572 2001 14604 2023
rect 14604 2001 14606 2023
rect 14500 1989 14534 1991
rect 14572 1989 14606 2001
rect 14356 1916 14390 1950
rect 14428 1902 14462 1936
rect 14500 1922 14502 1950
rect 14502 1922 14534 1950
rect 14572 1933 14604 1950
rect 14604 1933 14606 1950
rect 14500 1916 14534 1922
rect 14572 1916 14606 1933
rect 14356 1843 14390 1877
rect 14428 1830 14462 1864
rect 14500 1853 14502 1877
rect 14502 1853 14534 1877
rect 14572 1865 14604 1877
rect 14604 1865 14606 1877
rect 14500 1843 14534 1853
rect 14572 1843 14606 1865
rect 14356 1770 14390 1804
rect 14428 1758 14462 1792
rect 14500 1784 14502 1804
rect 14502 1784 14534 1804
rect 14572 1797 14604 1804
rect 14604 1797 14606 1804
rect 14500 1770 14534 1784
rect 14572 1770 14606 1797
rect 14356 1697 14390 1731
rect 14428 1686 14462 1720
rect 14500 1715 14502 1731
rect 14502 1715 14534 1731
rect 14572 1729 14604 1731
rect 14604 1729 14606 1731
rect 14500 1697 14534 1715
rect 14572 1697 14606 1729
rect 14356 1623 14390 1657
rect 14428 1614 14462 1648
rect 14500 1646 14502 1658
rect 14502 1646 14534 1658
rect 14500 1624 14534 1646
rect 14572 1627 14606 1658
rect 14572 1624 14604 1627
rect 14604 1624 14606 1627
rect 14356 1549 14390 1583
rect 14500 1577 14502 1585
rect 14502 1577 14534 1585
rect 14428 1542 14462 1576
rect 14500 1551 14534 1577
rect 14572 1559 14606 1585
rect 14572 1551 14604 1559
rect 14604 1551 14606 1559
rect 14356 1475 14390 1509
rect 14500 1508 14502 1512
rect 14502 1508 14534 1512
rect 14428 1470 14462 1504
rect 14500 1478 14534 1508
rect 14572 1491 14606 1512
rect 14572 1478 14604 1491
rect 14604 1478 14606 1491
rect 14356 1401 14390 1435
rect 14428 1398 14462 1432
rect 14500 1405 14534 1439
rect 14572 1423 14606 1439
rect 14572 1405 14604 1423
rect 14604 1405 14606 1423
rect 14356 1327 14390 1361
rect 14428 1326 14462 1360
rect 14500 1335 14534 1366
rect 14572 1355 14606 1366
rect 14500 1332 14502 1335
rect 14502 1332 14534 1335
rect 14572 1332 14604 1355
rect 14604 1332 14606 1355
rect 14356 1253 14390 1287
rect 14428 1254 14462 1288
rect 14500 1266 14534 1293
rect 14572 1287 14606 1293
rect 14500 1259 14502 1266
rect 14502 1259 14534 1266
rect 14572 1259 14604 1287
rect 14604 1259 14606 1287
rect 14356 1179 14390 1213
rect 14428 1182 14462 1216
rect 14500 1197 14534 1220
rect 14572 1218 14606 1220
rect 14500 1186 14502 1197
rect 14502 1186 14534 1197
rect 14572 1186 14604 1218
rect 14604 1186 14606 1218
rect 746 883 780 894
rect 14356 1105 14390 1139
rect 14428 1110 14462 1144
rect 14500 1128 14534 1147
rect 14500 1113 14502 1128
rect 14502 1113 14534 1128
rect 14572 1115 14604 1147
rect 14604 1115 14606 1147
rect 14572 1113 14606 1115
rect 14356 1031 14390 1065
rect 14428 1038 14462 1072
rect 14500 1059 14534 1074
rect 14500 1040 14502 1059
rect 14502 1040 14534 1059
rect 14572 1046 14604 1074
rect 14604 1046 14606 1074
rect 14572 1040 14606 1046
rect 14356 957 14390 991
rect 14428 966 14462 1000
rect 14500 990 14534 1001
rect 14500 967 14502 990
rect 14502 967 14534 990
rect 14572 977 14604 1001
rect 14604 977 14606 1001
rect 14572 967 14606 977
rect 14356 883 14390 917
rect 14428 894 14462 928
rect 14500 921 14534 928
rect 14500 894 14502 921
rect 14502 894 14534 921
rect 14572 908 14604 928
rect 14604 908 14606 928
rect 14572 894 14606 908
rect 709 818 736 820
rect 736 818 743 820
rect 782 818 805 820
rect 805 818 816 820
rect 855 818 874 820
rect 874 818 889 820
rect 928 818 943 820
rect 943 818 978 820
rect 978 818 1012 820
rect 1012 818 1047 820
rect 1047 818 1081 820
rect 1081 818 1116 820
rect 1116 818 1150 820
rect 1150 818 1185 820
rect 1185 818 1219 820
rect 1219 818 1254 820
rect 1254 818 1288 820
rect 1288 818 1323 820
rect 1323 818 1357 820
rect 1357 818 1392 820
rect 1392 818 1426 820
rect 1426 818 1461 820
rect 1461 818 1495 820
rect 1495 818 1530 820
rect 1530 818 1564 820
rect 1564 818 1599 820
rect 1599 818 1633 820
rect 1633 818 1668 820
rect 1668 818 1702 820
rect 1702 818 1737 820
rect 1737 818 1771 820
rect 1771 818 1806 820
rect 1806 818 1840 820
rect 1840 818 1875 820
rect 1875 818 1909 820
rect 1909 818 1944 820
rect 1944 818 1978 820
rect 1978 818 2013 820
rect 2013 818 2047 820
rect 2047 818 2082 820
rect 2082 818 2116 820
rect 2116 818 2151 820
rect 2151 818 2185 820
rect 2185 818 2220 820
rect 2220 818 2254 820
rect 2254 818 2289 820
rect 2289 818 2323 820
rect 2323 818 2358 820
rect 2358 818 2392 820
rect 2392 818 2427 820
rect 2427 818 2461 820
rect 2461 818 2496 820
rect 2496 818 2530 820
rect 2530 818 2565 820
rect 2565 818 2599 820
rect 2599 818 2634 820
rect 2634 818 2668 820
rect 2668 818 2703 820
rect 2703 818 2737 820
rect 2737 818 2772 820
rect 709 786 743 818
rect 782 786 816 818
rect 855 786 889 818
rect 928 784 2772 818
rect 928 750 944 784
rect 944 750 979 784
rect 979 750 1013 784
rect 1013 750 1048 784
rect 1048 750 1082 784
rect 1082 750 1117 784
rect 1117 750 1151 784
rect 1151 750 1186 784
rect 1186 750 1220 784
rect 1220 750 1255 784
rect 1255 750 1289 784
rect 1289 750 1324 784
rect 1324 750 1358 784
rect 1358 750 1393 784
rect 1393 750 1427 784
rect 1427 750 1462 784
rect 1462 750 1496 784
rect 1496 750 1531 784
rect 1531 750 1565 784
rect 1565 750 1600 784
rect 1600 750 1634 784
rect 1634 750 1669 784
rect 1669 750 1703 784
rect 1703 750 1738 784
rect 1738 750 1772 784
rect 1772 750 1807 784
rect 1807 750 1841 784
rect 1841 750 1876 784
rect 1876 750 1910 784
rect 1910 750 1945 784
rect 1945 750 1979 784
rect 1979 750 2014 784
rect 2014 750 2048 784
rect 2048 750 2083 784
rect 2083 750 2117 784
rect 2117 750 2152 784
rect 2152 750 2186 784
rect 2186 750 2221 784
rect 2221 750 2255 784
rect 2255 750 2290 784
rect 2290 750 2324 784
rect 2324 750 2359 784
rect 2359 750 2393 784
rect 2393 750 2428 784
rect 2428 750 2462 784
rect 2462 750 2497 784
rect 2497 750 2531 784
rect 2531 750 2566 784
rect 2566 750 2600 784
rect 2600 750 2635 784
rect 2635 750 2669 784
rect 2669 750 2704 784
rect 2704 750 2738 784
rect 2738 750 2772 784
rect 2772 750 14426 820
rect 709 716 743 748
rect 782 716 816 748
rect 855 716 889 748
rect 928 716 4725 750
rect 709 714 723 716
rect 723 714 743 716
rect 782 714 792 716
rect 792 714 816 716
rect 855 714 861 716
rect 861 714 889 716
rect 928 714 930 716
rect 930 714 964 716
rect 964 714 999 716
rect 999 714 1033 716
rect 1033 714 1068 716
rect 1068 714 1102 716
rect 1102 714 1137 716
rect 1137 714 1171 716
rect 1171 714 1206 716
rect 1206 714 1240 716
rect 1240 714 1275 716
rect 1275 714 1309 716
rect 1309 714 1344 716
rect 1344 714 1378 716
rect 1378 714 1413 716
rect 1413 714 1447 716
rect 1447 714 1482 716
rect 1482 714 1516 716
rect 1516 714 1551 716
rect 1551 714 1585 716
rect 1585 714 1620 716
rect 1620 714 1654 716
rect 1654 714 1689 716
rect 1689 714 1723 716
rect 1723 714 1758 716
rect 1758 714 1792 716
rect 1792 714 1827 716
rect 1827 714 1861 716
rect 1861 714 1896 716
rect 1896 714 1930 716
rect 1930 714 1965 716
rect 1965 714 1999 716
rect 1999 714 2034 716
rect 2034 714 2068 716
rect 2068 714 2103 716
rect 2103 714 2137 716
rect 2137 714 2172 716
rect 2172 714 2206 716
rect 2206 714 2241 716
rect 2241 714 2275 716
rect 2275 714 2310 716
rect 2310 714 2344 716
rect 2344 714 2379 716
rect 2379 714 2413 716
rect 2413 714 2448 716
rect 2448 714 2482 716
rect 2482 714 2517 716
rect 2517 714 2551 716
rect 2551 714 2586 716
rect 2586 714 2620 716
rect 2620 714 2655 716
rect 2655 714 2689 716
rect 2689 714 2724 716
rect 2724 714 2758 716
rect 2758 714 2793 716
rect 2793 714 2827 716
rect 2827 714 2862 716
rect 2862 714 2896 716
rect 2896 714 2931 716
rect 2931 714 2965 716
rect 2965 714 3000 716
rect 3000 714 3034 716
rect 3034 714 3069 716
rect 3069 714 3103 716
rect 3103 714 3138 716
rect 3138 714 3172 716
rect 3172 714 3207 716
rect 3207 714 3241 716
rect 3241 714 3276 716
rect 3276 714 3310 716
rect 3310 714 3345 716
rect 3345 714 3379 716
rect 3379 714 3414 716
rect 3414 714 3448 716
rect 3448 714 3483 716
rect 3483 714 3517 716
rect 3517 714 3552 716
rect 3552 714 3586 716
rect 3586 714 3621 716
rect 3621 714 3655 716
rect 3655 714 3690 716
rect 3690 714 3724 716
rect 3724 714 3759 716
rect 3759 714 3793 716
rect 3793 714 3828 716
rect 3828 714 3862 716
rect 3862 714 3897 716
rect 3897 714 3931 716
rect 3931 714 3966 716
rect 3966 714 4000 716
rect 4000 714 4035 716
rect 4035 714 4069 716
rect 4069 714 4104 716
rect 4104 714 4138 716
rect 4138 714 4173 716
rect 4173 714 4207 716
rect 4207 714 4242 716
rect 4242 714 4276 716
rect 4276 714 4311 716
rect 4311 714 4345 716
rect 4345 714 4380 716
rect 4380 714 4414 716
rect 4414 714 4449 716
rect 4449 714 4483 716
rect 4483 714 4518 716
rect 4518 714 4552 716
rect 4552 714 4587 716
rect 4587 714 4621 716
rect 4621 714 4656 716
rect 4656 714 4690 716
rect 4690 714 4725 716
rect 4725 714 14426 750
rect 14832 4636 14840 4670
rect 14840 4636 14866 4670
rect 14832 4564 14840 4598
rect 14840 4564 14866 4598
rect 14832 4492 14840 4526
rect 14840 4492 14866 4526
rect 14832 4420 14840 4454
rect 14840 4420 14866 4454
rect 14832 4348 14840 4382
rect 14840 4348 14866 4382
rect 14832 4276 14840 4310
rect 14840 4276 14866 4310
rect 14832 4204 14840 4238
rect 14840 4204 14866 4238
rect 14832 4132 14840 4166
rect 14840 4132 14866 4166
rect 14832 4060 14840 4094
rect 14840 4060 14866 4094
rect 14832 3988 14840 4022
rect 14840 3988 14866 4022
rect 14832 3916 14840 3950
rect 14840 3916 14866 3950
rect 14832 3844 14840 3878
rect 14840 3844 14866 3878
rect 14832 3772 14840 3806
rect 14840 3772 14866 3806
rect 14832 3700 14840 3734
rect 14840 3700 14866 3734
rect 14832 3628 14840 3662
rect 14840 3628 14866 3662
rect 14832 3556 14840 3590
rect 14840 3556 14866 3590
rect 14832 3484 14840 3518
rect 14840 3484 14866 3518
rect 14832 3412 14840 3446
rect 14840 3412 14866 3446
rect 14832 3340 14840 3374
rect 14840 3340 14866 3374
rect 14832 3268 14840 3302
rect 14840 3268 14866 3302
rect 14832 3196 14840 3230
rect 14840 3196 14866 3230
rect 14832 3124 14840 3158
rect 14840 3124 14866 3158
rect 14832 3052 14840 3086
rect 14840 3052 14866 3086
rect 14832 2980 14840 3014
rect 14840 2980 14866 3014
rect 14832 2908 14840 2942
rect 14840 2908 14866 2942
rect 14832 2836 14840 2870
rect 14840 2836 14866 2870
rect 14832 2764 14840 2798
rect 14840 2764 14866 2798
rect 14832 2692 14840 2726
rect 14840 2692 14866 2726
rect 14832 2620 14840 2654
rect 14840 2620 14866 2654
rect 14832 2548 14840 2582
rect 14840 2548 14866 2582
rect 14832 2476 14840 2510
rect 14840 2476 14866 2510
rect 14832 2404 14840 2438
rect 14840 2404 14866 2438
rect 14832 2332 14840 2366
rect 14840 2332 14866 2366
rect 14832 2260 14840 2294
rect 14840 2260 14866 2294
rect 14832 2188 14840 2222
rect 14840 2188 14866 2222
rect 14832 2116 14840 2150
rect 14840 2116 14866 2150
rect 14832 2044 14840 2078
rect 14840 2044 14866 2078
rect 14832 1972 14840 2006
rect 14840 1972 14866 2006
rect 14832 1900 14840 1934
rect 14840 1900 14866 1934
rect 14832 1828 14840 1862
rect 14840 1828 14866 1862
rect 14832 1756 14840 1790
rect 14840 1756 14866 1790
rect 14832 1684 14840 1718
rect 14840 1684 14866 1718
rect 14832 1612 14840 1646
rect 14840 1612 14866 1646
rect 14832 1540 14840 1574
rect 14840 1540 14866 1574
rect 14832 1468 14840 1502
rect 14840 1468 14866 1502
rect 14832 1395 14840 1429
rect 14840 1395 14866 1429
rect 14832 1322 14840 1356
rect 14840 1322 14866 1356
rect 14832 1249 14840 1283
rect 14840 1249 14866 1283
rect 14832 1176 14840 1210
rect 14840 1176 14866 1210
rect 14832 1103 14840 1137
rect 14840 1103 14866 1137
rect 14832 1030 14840 1064
rect 14840 1030 14866 1064
rect 14832 957 14840 991
rect 14840 957 14866 991
rect 14832 884 14840 918
rect 14840 884 14866 918
rect 14832 811 14840 845
rect 14840 811 14866 845
rect 14832 738 14840 772
rect 14840 738 14866 772
rect 269 609 296 641
rect 296 609 303 641
rect 269 607 303 609
rect 269 541 296 567
rect 296 541 303 567
rect 269 533 303 541
rect 14832 665 14840 699
rect 14840 665 14866 699
rect 14832 592 14840 626
rect 14840 592 14866 626
rect 14832 519 14840 553
rect 14840 519 14866 553
rect 343 465 365 497
rect 365 465 377 497
rect 419 465 434 497
rect 434 465 453 497
rect 495 465 503 497
rect 503 465 529 497
rect 571 465 572 497
rect 572 465 605 497
rect 648 465 676 497
rect 676 465 682 497
rect 343 463 377 465
rect 419 463 453 465
rect 495 463 529 465
rect 571 463 605 465
rect 648 463 682 465
rect 14465 447 14499 481
rect 14539 447 14573 481
rect 14613 447 14647 481
rect 14686 447 14720 481
rect 14759 447 14793 481
rect 361 363 395 375
rect 361 341 365 363
rect 365 341 395 363
rect 434 341 468 375
rect 507 363 541 375
rect 580 363 614 375
rect 653 363 687 375
rect 726 363 760 375
rect 799 363 833 375
rect 872 363 906 375
rect 945 363 979 375
rect 1018 363 1052 375
rect 1091 363 1125 375
rect 1164 363 1198 375
rect 1237 363 1271 375
rect 1310 363 1344 375
rect 1383 363 1417 375
rect 1456 363 1490 375
rect 1529 363 1563 375
rect 1602 363 1636 375
rect 1675 363 1709 375
rect 1748 363 1782 375
rect 1821 363 1855 375
rect 1894 363 1928 375
rect 1967 363 2001 375
rect 507 341 538 363
rect 538 341 541 363
rect 580 341 607 363
rect 607 341 614 363
rect 653 341 676 363
rect 676 341 687 363
rect 726 341 745 363
rect 745 341 760 363
rect 799 341 814 363
rect 814 341 833 363
rect 872 341 883 363
rect 883 341 906 363
rect 945 341 952 363
rect 952 341 979 363
rect 1018 341 1021 363
rect 1021 341 1052 363
rect 1091 341 1124 363
rect 1124 341 1125 363
rect 1164 341 1193 363
rect 1193 341 1198 363
rect 1237 341 1262 363
rect 1262 341 1271 363
rect 1310 341 1331 363
rect 1331 341 1344 363
rect 1383 341 1400 363
rect 1400 341 1417 363
rect 1456 341 1469 363
rect 1469 341 1490 363
rect 1529 341 1538 363
rect 1538 341 1563 363
rect 1602 341 1607 363
rect 1607 341 1636 363
rect 1675 341 1676 363
rect 1676 341 1709 363
rect 1748 341 1780 363
rect 1780 341 1782 363
rect 1821 341 1849 363
rect 1849 341 1855 363
rect 1894 341 1918 363
rect 1918 341 1928 363
rect 1967 341 1987 363
rect 1987 341 2001 363
rect 2040 341 2056 375
rect 2056 341 2074 375
rect 2113 341 2147 375
rect 2186 341 2220 375
rect 2259 341 2293 375
rect 2332 341 2366 375
rect 2405 341 2439 375
rect 2478 341 2512 375
rect 2551 341 2585 375
rect 2624 341 2658 375
rect 2697 341 2731 375
rect 2770 341 2804 375
rect 2843 341 2877 375
rect 2916 341 2950 375
rect 2989 341 3023 375
rect 3062 341 3096 375
rect 3135 341 3169 375
rect 3208 341 3242 375
rect 3281 341 3315 375
rect 3354 341 3388 375
rect 3427 341 3461 375
rect 3500 341 3534 375
rect 3573 341 3607 375
rect 3646 341 3680 375
rect 3719 341 3753 375
rect 3792 341 3826 375
rect 3865 341 3899 375
rect 3938 341 3972 375
rect 4011 341 4045 375
rect 4084 341 4118 375
rect 4157 341 4191 375
rect 4229 341 4263 375
rect 4301 341 4335 375
rect 4373 341 4407 375
rect 4445 341 4479 375
rect 4517 341 4551 375
rect 4589 341 4623 375
rect 4661 341 4695 375
rect 4733 341 4767 375
rect 4805 341 4839 375
rect 4877 341 4911 375
rect 4949 341 4983 375
rect 5021 341 5055 375
rect 5093 341 5127 375
rect 5165 341 5199 375
rect 5237 341 5271 375
rect 5309 341 5343 375
rect 5381 341 5415 375
rect 5453 341 5487 375
rect 5525 341 5559 375
rect 5597 341 5631 375
rect 5669 341 5703 375
rect 5741 341 5775 375
rect 5813 341 5847 375
rect 5885 341 5919 375
rect 5957 341 5991 375
rect 6029 341 6063 375
rect 6101 341 6135 375
rect 6173 341 6207 375
rect 6245 341 6279 375
rect 6317 341 6351 375
rect 6389 341 6423 375
rect 6461 341 6495 375
rect 6533 341 6567 375
rect 6605 341 6639 375
rect 6677 341 6711 375
rect 6749 341 6783 375
rect 6821 341 6855 375
rect 6893 341 6927 375
rect 6965 341 6999 375
rect 7037 341 7071 375
rect 7109 341 7143 375
rect 7181 341 7215 375
rect 7253 341 7287 375
rect 7325 341 7359 375
rect 7397 341 7431 375
rect 7469 341 7503 375
rect 7541 341 7575 375
rect 7613 341 7647 375
rect 7685 341 7719 375
rect 7757 341 7791 375
rect 7829 341 7863 375
rect 7901 341 7935 375
rect 7973 341 8007 375
rect 8045 341 8079 375
rect 8117 341 8151 375
rect 8189 341 8223 375
rect 8261 341 8295 375
rect 8333 341 8367 375
rect 8405 341 8439 375
rect 8477 341 8511 375
rect 8549 341 8583 375
rect 8621 341 8655 375
rect 8693 341 8727 375
rect 8765 341 8799 375
rect 8837 341 8871 375
rect 8909 341 8943 375
rect 8981 341 9015 375
rect 9053 341 9087 375
rect 9125 341 9159 375
rect 9197 341 9231 375
rect 9269 341 9303 375
rect 9341 341 9375 375
rect 9413 341 9447 375
rect 9485 341 9519 375
rect 9557 341 9591 375
rect 9629 341 9663 375
rect 9701 341 9735 375
rect 9773 341 9807 375
rect 9845 341 9879 375
rect 9917 341 9951 375
rect 9989 341 10023 375
rect 10061 341 10095 375
rect 10133 341 10167 375
rect 10205 341 10239 375
rect 10277 341 10311 375
rect 10349 341 10383 375
rect 10421 341 10455 375
rect 10493 341 10527 375
rect 10565 341 10599 375
rect 10637 341 10671 375
rect 10709 341 10743 375
rect 10781 341 10815 375
rect 10853 341 10887 375
rect 10925 341 10959 375
rect 10997 341 11031 375
rect 11069 341 11103 375
rect 11141 341 11175 375
rect 11213 341 11247 375
rect 11285 341 11319 375
rect 11357 341 11391 375
rect 11429 341 11463 375
rect 11501 341 11535 375
rect 11573 341 11607 375
rect 11645 341 11679 375
rect 11717 341 11751 375
rect 11789 341 11823 375
rect 11861 341 11895 375
rect 11933 341 11967 375
rect 12005 341 12039 375
rect 12077 341 12111 375
rect 12149 341 12183 375
rect 12221 341 12255 375
rect 12293 341 12327 375
rect 12365 341 12399 375
rect 12437 341 12471 375
rect 12509 341 12543 375
rect 12581 341 12615 375
rect 12653 341 12687 375
rect 12725 341 12759 375
rect 12797 341 12831 375
rect 12869 341 12903 375
rect 12941 341 12975 375
rect 13013 341 13047 375
rect 13085 341 13119 375
rect 13157 341 13191 375
rect 13229 341 13263 375
rect 13301 341 13335 375
rect 13373 341 13407 375
rect 13445 341 13479 375
rect 13517 341 13551 375
rect 13589 341 13623 375
rect 13661 341 13695 375
rect 13733 341 13767 375
rect 13805 341 13839 375
rect 13877 341 13911 375
rect 13949 341 13983 375
rect 14021 341 14055 375
rect 14093 341 14127 375
rect 14165 341 14199 375
rect 14237 341 14271 375
rect 14309 341 14343 375
rect 14381 341 14415 375
rect 14453 341 14487 375
rect 14525 341 14559 375
rect 14597 341 14631 375
rect 14669 341 14703 375
rect 14741 341 14775 375
<< metal1 >>
rect 39 5111 15097 5118
rect 39 5077 361 5111
rect 395 5077 434 5111
rect 468 5077 507 5111
rect 541 5077 580 5111
rect 614 5077 653 5111
rect 687 5077 726 5111
rect 760 5077 799 5111
rect 833 5077 872 5111
rect 906 5077 945 5111
rect 979 5077 1018 5111
rect 1052 5077 1091 5111
rect 1125 5077 1164 5111
rect 1198 5077 1237 5111
rect 1271 5077 1310 5111
rect 1344 5077 1383 5111
rect 1417 5077 1456 5111
rect 1490 5077 1529 5111
rect 1563 5077 1602 5111
rect 1636 5077 1675 5111
rect 1709 5077 1748 5111
rect 1782 5077 1821 5111
rect 1855 5077 1894 5111
rect 1928 5077 1967 5111
rect 2001 5077 2040 5111
rect 2074 5077 2113 5111
rect 2147 5077 2186 5111
rect 2220 5077 2259 5111
rect 2293 5077 2332 5111
rect 2366 5077 2405 5111
rect 2439 5077 2478 5111
rect 2512 5077 2551 5111
rect 2585 5077 2624 5111
rect 2658 5077 2697 5111
rect 2731 5077 2770 5111
rect 2804 5077 2843 5111
rect 2877 5077 2916 5111
rect 2950 5077 2989 5111
rect 3023 5077 3062 5111
rect 3096 5077 3135 5111
rect 3169 5077 3208 5111
rect 3242 5077 3281 5111
rect 3315 5077 3354 5111
rect 3388 5077 3427 5111
rect 3461 5077 3500 5111
rect 3534 5077 3573 5111
rect 3607 5077 3646 5111
rect 3680 5077 3719 5111
rect 3753 5077 3792 5111
rect 3826 5077 3865 5111
rect 3899 5077 3938 5111
rect 3972 5077 4011 5111
rect 4045 5077 4084 5111
rect 4118 5077 4157 5111
rect 4191 5077 4229 5111
rect 4263 5077 4301 5111
rect 4335 5077 4373 5111
rect 4407 5077 4445 5111
rect 4479 5077 4517 5111
rect 4551 5077 4589 5111
rect 4623 5077 4661 5111
rect 4695 5077 4733 5111
rect 4767 5077 4805 5111
rect 4839 5077 4877 5111
rect 4911 5077 4949 5111
rect 4983 5077 5021 5111
rect 5055 5077 5093 5111
rect 5127 5077 5165 5111
rect 5199 5077 5237 5111
rect 5271 5077 5309 5111
rect 5343 5077 5381 5111
rect 5415 5077 5453 5111
rect 5487 5077 5525 5111
rect 5559 5077 5597 5111
rect 5631 5077 5669 5111
rect 5703 5077 5741 5111
rect 5775 5077 5813 5111
rect 5847 5077 5885 5111
rect 5919 5077 5957 5111
rect 5991 5077 6029 5111
rect 6063 5077 6101 5111
rect 6135 5077 6173 5111
rect 6207 5077 6245 5111
rect 6279 5077 6317 5111
rect 6351 5077 6389 5111
rect 6423 5077 6461 5111
rect 6495 5077 6533 5111
rect 6567 5077 6605 5111
rect 6639 5077 6677 5111
rect 6711 5077 6749 5111
rect 6783 5077 6821 5111
rect 6855 5077 6893 5111
rect 6927 5077 6965 5111
rect 6999 5077 7037 5111
rect 7071 5077 7109 5111
rect 7143 5077 7181 5111
rect 7215 5077 7253 5111
rect 7287 5077 7325 5111
rect 7359 5077 7397 5111
rect 7431 5077 7469 5111
rect 7503 5077 7541 5111
rect 7575 5077 7613 5111
rect 7647 5077 7685 5111
rect 7719 5077 7757 5111
rect 7791 5077 7829 5111
rect 7863 5077 7901 5111
rect 7935 5077 7973 5111
rect 8007 5077 8045 5111
rect 8079 5077 8117 5111
rect 8151 5077 8189 5111
rect 8223 5077 8261 5111
rect 8295 5077 8333 5111
rect 8367 5077 8405 5111
rect 8439 5077 8477 5111
rect 8511 5077 8549 5111
rect 8583 5077 8621 5111
rect 8655 5077 8693 5111
rect 8727 5077 8765 5111
rect 8799 5077 8837 5111
rect 8871 5077 8909 5111
rect 8943 5077 8981 5111
rect 9015 5077 9053 5111
rect 9087 5077 9125 5111
rect 9159 5077 9197 5111
rect 9231 5077 9269 5111
rect 9303 5077 9341 5111
rect 9375 5077 9413 5111
rect 9447 5077 9485 5111
rect 9519 5077 9557 5111
rect 9591 5077 9629 5111
rect 9663 5077 9701 5111
rect 9735 5077 9773 5111
rect 9807 5077 9845 5111
rect 9879 5077 9917 5111
rect 9951 5077 9989 5111
rect 10023 5077 10061 5111
rect 10095 5077 10133 5111
rect 10167 5077 10205 5111
rect 10239 5077 10277 5111
rect 10311 5077 10349 5111
rect 10383 5077 10421 5111
rect 10455 5077 10493 5111
rect 10527 5077 10565 5111
rect 10599 5077 10637 5111
rect 10671 5077 10709 5111
rect 10743 5077 10781 5111
rect 10815 5077 10853 5111
rect 10887 5077 10925 5111
rect 10959 5077 10997 5111
rect 11031 5077 11069 5111
rect 11103 5077 11141 5111
rect 11175 5077 11213 5111
rect 11247 5077 11285 5111
rect 11319 5077 11357 5111
rect 11391 5077 11429 5111
rect 11463 5077 11501 5111
rect 11535 5077 11573 5111
rect 11607 5077 11645 5111
rect 11679 5077 11717 5111
rect 11751 5077 11789 5111
rect 11823 5077 11861 5111
rect 11895 5077 11933 5111
rect 11967 5077 12005 5111
rect 12039 5077 12077 5111
rect 12111 5077 12149 5111
rect 12183 5077 12221 5111
rect 12255 5077 12293 5111
rect 12327 5077 12365 5111
rect 12399 5077 12437 5111
rect 12471 5077 12509 5111
rect 12543 5077 12581 5111
rect 12615 5077 12653 5111
rect 12687 5077 12725 5111
rect 12759 5077 12797 5111
rect 12831 5077 12869 5111
rect 12903 5077 12941 5111
rect 12975 5077 13013 5111
rect 13047 5077 13085 5111
rect 13119 5077 13157 5111
rect 13191 5077 13229 5111
rect 13263 5077 13301 5111
rect 13335 5077 13373 5111
rect 13407 5077 13445 5111
rect 13479 5077 13517 5111
rect 13551 5077 13589 5111
rect 13623 5077 13661 5111
rect 13695 5077 13733 5111
rect 13767 5077 13805 5111
rect 13839 5077 13877 5111
rect 13911 5077 13949 5111
rect 13983 5077 14021 5111
rect 14055 5077 14093 5111
rect 14127 5077 14165 5111
rect 14199 5077 14237 5111
rect 14271 5077 14309 5111
rect 14343 5077 14381 5111
rect 14415 5077 14453 5111
rect 14487 5077 14525 5111
rect 14559 5077 14597 5111
rect 14631 5077 14669 5111
rect 14703 5077 14741 5111
rect 14775 5077 15097 5111
rect 39 5035 15097 5077
rect 39 5029 361 5035
rect 39 4995 269 5029
rect 303 5001 361 5029
rect 395 5001 434 5035
rect 468 5001 507 5035
rect 541 5001 580 5035
rect 614 5001 653 5035
rect 687 5001 726 5035
rect 760 5001 799 5035
rect 833 5001 872 5035
rect 906 5001 945 5035
rect 979 5001 1018 5035
rect 1052 5001 1091 5035
rect 1125 5001 1164 5035
rect 1198 5001 1237 5035
rect 1271 5001 1310 5035
rect 1344 5001 1383 5035
rect 1417 5001 1456 5035
rect 1490 5001 1529 5035
rect 1563 5001 1602 5035
rect 1636 5001 1675 5035
rect 1709 5001 1748 5035
rect 1782 5001 1821 5035
rect 1855 5001 1894 5035
rect 1928 5001 1967 5035
rect 2001 5001 2040 5035
rect 2074 5001 2113 5035
rect 2147 5001 2186 5035
rect 2220 5001 2259 5035
rect 2293 5001 2332 5035
rect 2366 5001 2405 5035
rect 2439 5001 2478 5035
rect 2512 5001 2551 5035
rect 2585 5001 2624 5035
rect 2658 5001 2697 5035
rect 2731 5001 2770 5035
rect 2804 5001 2843 5035
rect 2877 5001 2916 5035
rect 2950 5001 2989 5035
rect 3023 5001 3062 5035
rect 3096 5001 3135 5035
rect 3169 5001 3208 5035
rect 3242 5001 3281 5035
rect 3315 5001 3354 5035
rect 3388 5001 3427 5035
rect 3461 5001 3500 5035
rect 3534 5001 3573 5035
rect 3607 5001 3646 5035
rect 3680 5001 3719 5035
rect 3753 5001 3792 5035
rect 3826 5001 3865 5035
rect 3899 5001 3938 5035
rect 3972 5001 4011 5035
rect 4045 5001 4084 5035
rect 4118 5001 4157 5035
rect 4191 5001 4229 5035
rect 4263 5001 4301 5035
rect 4335 5001 4373 5035
rect 4407 5001 4445 5035
rect 4479 5001 4517 5035
rect 4551 5001 4589 5035
rect 4623 5001 4661 5035
rect 4695 5001 4733 5035
rect 4767 5001 4805 5035
rect 4839 5001 4877 5035
rect 4911 5001 4949 5035
rect 4983 5001 5021 5035
rect 5055 5001 5093 5035
rect 5127 5001 5165 5035
rect 5199 5001 5237 5035
rect 5271 5001 5309 5035
rect 5343 5001 5381 5035
rect 5415 5001 5453 5035
rect 5487 5001 5525 5035
rect 5559 5001 5597 5035
rect 5631 5001 5669 5035
rect 5703 5001 5741 5035
rect 5775 5001 5813 5035
rect 5847 5001 5885 5035
rect 5919 5001 5957 5035
rect 5991 5001 6029 5035
rect 6063 5001 6101 5035
rect 6135 5001 6173 5035
rect 6207 5001 6245 5035
rect 6279 5001 6317 5035
rect 6351 5001 6389 5035
rect 6423 5001 6461 5035
rect 6495 5001 6533 5035
rect 6567 5001 6605 5035
rect 6639 5001 6677 5035
rect 6711 5001 6749 5035
rect 6783 5001 6821 5035
rect 6855 5001 6893 5035
rect 6927 5001 6965 5035
rect 6999 5001 7037 5035
rect 7071 5001 7109 5035
rect 7143 5001 7181 5035
rect 7215 5001 7253 5035
rect 7287 5001 7325 5035
rect 7359 5001 7397 5035
rect 7431 5001 7469 5035
rect 7503 5001 7541 5035
rect 7575 5001 7613 5035
rect 7647 5001 7685 5035
rect 7719 5001 7757 5035
rect 7791 5001 7829 5035
rect 7863 5001 7901 5035
rect 7935 5001 7973 5035
rect 8007 5001 8045 5035
rect 8079 5001 8117 5035
rect 8151 5001 8189 5035
rect 8223 5001 8261 5035
rect 8295 5001 8333 5035
rect 8367 5001 8405 5035
rect 8439 5001 8477 5035
rect 8511 5001 8549 5035
rect 8583 5001 8621 5035
rect 8655 5001 8693 5035
rect 8727 5001 8765 5035
rect 8799 5001 8837 5035
rect 8871 5001 8909 5035
rect 8943 5001 8981 5035
rect 9015 5001 9053 5035
rect 9087 5001 9125 5035
rect 9159 5001 9197 5035
rect 9231 5001 9269 5035
rect 9303 5001 9341 5035
rect 9375 5001 9413 5035
rect 9447 5001 9485 5035
rect 9519 5001 9557 5035
rect 9591 5001 9629 5035
rect 9663 5001 9701 5035
rect 9735 5001 9773 5035
rect 9807 5001 9845 5035
rect 9879 5001 9917 5035
rect 9951 5001 9989 5035
rect 10023 5001 10061 5035
rect 10095 5001 10133 5035
rect 10167 5001 10205 5035
rect 10239 5001 10277 5035
rect 10311 5001 10349 5035
rect 10383 5001 10421 5035
rect 10455 5001 10493 5035
rect 10527 5001 10565 5035
rect 10599 5001 10637 5035
rect 10671 5001 10709 5035
rect 10743 5001 10781 5035
rect 10815 5001 10853 5035
rect 10887 5001 10925 5035
rect 10959 5001 10997 5035
rect 11031 5001 11069 5035
rect 11103 5001 11141 5035
rect 11175 5001 11213 5035
rect 11247 5001 11285 5035
rect 11319 5001 11357 5035
rect 11391 5001 11429 5035
rect 11463 5001 11501 5035
rect 11535 5001 11573 5035
rect 11607 5001 11645 5035
rect 11679 5001 11717 5035
rect 11751 5001 11789 5035
rect 11823 5001 11861 5035
rect 11895 5001 11933 5035
rect 11967 5001 12005 5035
rect 12039 5001 12077 5035
rect 12111 5001 12149 5035
rect 12183 5001 12221 5035
rect 12255 5001 12293 5035
rect 12327 5001 12365 5035
rect 12399 5001 12437 5035
rect 12471 5001 12509 5035
rect 12543 5001 12581 5035
rect 12615 5001 12653 5035
rect 12687 5001 12725 5035
rect 12759 5001 12797 5035
rect 12831 5001 12869 5035
rect 12903 5001 12941 5035
rect 12975 5001 13013 5035
rect 13047 5001 13085 5035
rect 13119 5001 13157 5035
rect 13191 5001 13229 5035
rect 13263 5001 13301 5035
rect 13335 5001 13373 5035
rect 13407 5001 13445 5035
rect 13479 5001 13517 5035
rect 13551 5001 13589 5035
rect 13623 5001 13661 5035
rect 13695 5001 13733 5035
rect 13767 5001 13805 5035
rect 13839 5001 13877 5035
rect 13911 5001 13949 5035
rect 13983 5001 14021 5035
rect 14055 5001 14093 5035
rect 14127 5001 14165 5035
rect 14199 5001 14237 5035
rect 14271 5001 14309 5035
rect 14343 5001 14381 5035
rect 14415 5001 14453 5035
rect 14487 5001 14525 5035
rect 14559 5001 14597 5035
rect 14631 5001 14669 5035
rect 14703 5001 14741 5035
rect 14775 5030 15097 5035
rect 14775 5001 14832 5030
rect 303 4996 14832 5001
rect 14866 4996 15097 5030
rect 303 4995 15097 4996
rect 39 4959 15097 4995
rect 39 4956 361 4959
rect 39 4922 269 4956
rect 303 4925 361 4956
rect 395 4925 434 4959
rect 468 4925 507 4959
rect 541 4925 580 4959
rect 614 4925 653 4959
rect 687 4925 726 4959
rect 760 4925 799 4959
rect 833 4925 872 4959
rect 906 4925 945 4959
rect 979 4925 1018 4959
rect 1052 4925 1091 4959
rect 1125 4925 1164 4959
rect 1198 4925 1237 4959
rect 1271 4925 1310 4959
rect 1344 4925 1383 4959
rect 1417 4925 1456 4959
rect 1490 4925 1529 4959
rect 1563 4925 1602 4959
rect 1636 4925 1675 4959
rect 1709 4925 1748 4959
rect 1782 4925 1821 4959
rect 1855 4925 1894 4959
rect 1928 4925 1967 4959
rect 2001 4925 2040 4959
rect 2074 4925 2113 4959
rect 2147 4925 2186 4959
rect 2220 4925 2259 4959
rect 2293 4925 2332 4959
rect 2366 4925 2405 4959
rect 2439 4925 2478 4959
rect 2512 4925 2551 4959
rect 2585 4925 2624 4959
rect 2658 4925 2697 4959
rect 2731 4925 2770 4959
rect 2804 4925 2843 4959
rect 2877 4925 2916 4959
rect 2950 4925 2989 4959
rect 3023 4925 3062 4959
rect 3096 4925 3135 4959
rect 3169 4925 3208 4959
rect 3242 4925 3281 4959
rect 3315 4925 3354 4959
rect 3388 4925 3427 4959
rect 3461 4925 3500 4959
rect 3534 4925 3573 4959
rect 3607 4925 3646 4959
rect 3680 4925 3719 4959
rect 3753 4925 3792 4959
rect 3826 4925 3865 4959
rect 3899 4925 3938 4959
rect 3972 4925 4011 4959
rect 4045 4925 4084 4959
rect 4118 4925 4157 4959
rect 4191 4925 4229 4959
rect 4263 4925 4301 4959
rect 4335 4925 4373 4959
rect 4407 4925 4445 4959
rect 4479 4925 4517 4959
rect 4551 4925 4589 4959
rect 4623 4925 4661 4959
rect 4695 4925 4733 4959
rect 4767 4925 4805 4959
rect 4839 4925 4877 4959
rect 4911 4925 4949 4959
rect 4983 4925 5021 4959
rect 5055 4925 5093 4959
rect 5127 4925 5165 4959
rect 5199 4925 5237 4959
rect 5271 4925 5309 4959
rect 5343 4925 5381 4959
rect 5415 4925 5453 4959
rect 5487 4925 5525 4959
rect 5559 4925 5597 4959
rect 5631 4925 5669 4959
rect 5703 4925 5741 4959
rect 5775 4925 5813 4959
rect 5847 4925 5885 4959
rect 5919 4925 5957 4959
rect 5991 4925 6029 4959
rect 6063 4925 6101 4959
rect 6135 4925 6173 4959
rect 6207 4925 6245 4959
rect 6279 4925 6317 4959
rect 6351 4925 6389 4959
rect 6423 4925 6461 4959
rect 6495 4925 6533 4959
rect 6567 4925 6605 4959
rect 6639 4925 6677 4959
rect 6711 4925 6749 4959
rect 6783 4925 6821 4959
rect 6855 4925 6893 4959
rect 6927 4925 6965 4959
rect 6999 4925 7037 4959
rect 7071 4925 7109 4959
rect 7143 4925 7181 4959
rect 7215 4925 7253 4959
rect 7287 4925 7325 4959
rect 7359 4925 7397 4959
rect 7431 4925 7469 4959
rect 7503 4925 7541 4959
rect 7575 4925 7613 4959
rect 7647 4925 7685 4959
rect 7719 4925 7757 4959
rect 7791 4925 7829 4959
rect 7863 4925 7901 4959
rect 7935 4925 7973 4959
rect 8007 4925 8045 4959
rect 8079 4925 8117 4959
rect 8151 4925 8189 4959
rect 8223 4925 8261 4959
rect 8295 4925 8333 4959
rect 8367 4925 8405 4959
rect 8439 4925 8477 4959
rect 8511 4925 8549 4959
rect 8583 4925 8621 4959
rect 8655 4925 8693 4959
rect 8727 4925 8765 4959
rect 8799 4925 8837 4959
rect 8871 4925 8909 4959
rect 8943 4925 8981 4959
rect 9015 4925 9053 4959
rect 9087 4925 9125 4959
rect 9159 4925 9197 4959
rect 9231 4925 9269 4959
rect 9303 4925 9341 4959
rect 9375 4925 9413 4959
rect 9447 4925 9485 4959
rect 9519 4925 9557 4959
rect 9591 4925 9629 4959
rect 9663 4925 9701 4959
rect 9735 4925 9773 4959
rect 9807 4925 9845 4959
rect 9879 4925 9917 4959
rect 9951 4925 9989 4959
rect 10023 4925 10061 4959
rect 10095 4925 10133 4959
rect 10167 4925 10205 4959
rect 10239 4925 10277 4959
rect 10311 4925 10349 4959
rect 10383 4925 10421 4959
rect 10455 4925 10493 4959
rect 10527 4925 10565 4959
rect 10599 4925 10637 4959
rect 10671 4925 10709 4959
rect 10743 4925 10781 4959
rect 10815 4925 10853 4959
rect 10887 4925 10925 4959
rect 10959 4925 10997 4959
rect 11031 4925 11069 4959
rect 11103 4925 11141 4959
rect 11175 4925 11213 4959
rect 11247 4925 11285 4959
rect 11319 4925 11357 4959
rect 11391 4925 11429 4959
rect 11463 4925 11501 4959
rect 11535 4925 11573 4959
rect 11607 4925 11645 4959
rect 11679 4925 11717 4959
rect 11751 4925 11789 4959
rect 11823 4925 11861 4959
rect 11895 4925 11933 4959
rect 11967 4925 12005 4959
rect 12039 4925 12077 4959
rect 12111 4925 12149 4959
rect 12183 4925 12221 4959
rect 12255 4925 12293 4959
rect 12327 4925 12365 4959
rect 12399 4925 12437 4959
rect 12471 4925 12509 4959
rect 12543 4925 12581 4959
rect 12615 4925 12653 4959
rect 12687 4925 12725 4959
rect 12759 4925 12797 4959
rect 12831 4925 12869 4959
rect 12903 4925 12941 4959
rect 12975 4925 13013 4959
rect 13047 4925 13085 4959
rect 13119 4925 13157 4959
rect 13191 4925 13229 4959
rect 13263 4925 13301 4959
rect 13335 4925 13373 4959
rect 13407 4925 13445 4959
rect 13479 4925 13517 4959
rect 13551 4925 13589 4959
rect 13623 4925 13661 4959
rect 13695 4925 13733 4959
rect 13767 4925 13805 4959
rect 13839 4925 13877 4959
rect 13911 4925 13949 4959
rect 13983 4925 14021 4959
rect 14055 4925 14093 4959
rect 14127 4925 14165 4959
rect 14199 4925 14237 4959
rect 14271 4925 14309 4959
rect 14343 4925 14381 4959
rect 14415 4925 14453 4959
rect 14487 4925 14525 4959
rect 14559 4925 14597 4959
rect 14631 4925 14669 4959
rect 14703 4925 14741 4959
rect 14775 4958 15097 4959
rect 14775 4925 14832 4958
rect 303 4924 14832 4925
rect 14866 4924 15097 4958
rect 303 4922 15097 4924
rect 39 4918 15097 4922
rect 39 4886 759 4918
tri 759 4886 791 4918 nw
tri 14335 4886 14367 4918 ne
rect 14367 4886 15097 4918
rect 39 4883 725 4886
rect 39 4849 269 4883
rect 303 4852 725 4883
tri 725 4852 759 4886 nw
tri 14367 4852 14401 4886 ne
rect 14401 4852 14832 4886
rect 14866 4852 15097 4886
rect 303 4849 687 4852
rect 39 4814 687 4849
tri 687 4814 725 4852 nw
tri 14401 4814 14439 4852 ne
rect 14439 4814 15097 4852
rect 39 4810 653 4814
rect 39 4776 269 4810
rect 303 4780 653 4810
tri 653 4780 687 4814 nw
tri 14439 4780 14473 4814 ne
rect 14473 4780 14832 4814
rect 14866 4780 15097 4814
rect 303 4776 615 4780
rect 39 4742 615 4776
tri 615 4742 653 4780 nw
tri 14473 4742 14511 4780 ne
rect 14511 4742 15097 4780
rect 39 4737 581 4742
rect 39 4703 269 4737
rect 303 4708 581 4737
tri 581 4708 615 4742 nw
tri 14511 4708 14545 4742 ne
rect 14545 4708 14832 4742
rect 14866 4708 15097 4742
rect 303 4703 543 4708
rect 39 4670 543 4703
tri 543 4670 581 4708 nw
tri 14545 4670 14583 4708 ne
rect 14583 4670 15097 4708
rect 39 4664 509 4670
rect 39 4630 269 4664
rect 303 4636 509 4664
tri 509 4636 543 4670 nw
tri 14583 4636 14617 4670 ne
rect 14617 4636 14832 4670
rect 14866 4636 15097 4670
rect 303 4630 491 4636
rect 39 4618 491 4630
tri 491 4618 509 4636 nw
tri 14617 4618 14635 4636 ne
rect 14635 4618 15097 4636
rect 39 4606 479 4618
tri 479 4606 491 4618 nw
tri 621 4606 633 4618 se
rect 633 4606 14502 4618
rect 39 4591 373 4606
rect 39 4557 269 4591
rect 303 4557 373 4591
rect 39 4518 373 4557
rect 39 4484 269 4518
rect 303 4500 373 4518
tri 373 4500 479 4606 nw
tri 517 4502 621 4606 se
rect 621 4502 709 4606
rect 517 4500 709 4502
rect 14207 4572 14246 4606
rect 14280 4572 14319 4606
rect 14353 4572 14392 4606
rect 14426 4598 14502 4606
tri 14502 4598 14522 4618 sw
tri 14635 4598 14655 4618 ne
rect 14655 4598 15097 4618
rect 14426 4572 14522 4598
rect 14207 4564 14522 4572
tri 14522 4564 14556 4598 sw
tri 14655 4564 14689 4598 ne
rect 14689 4564 14832 4598
rect 14866 4564 15097 4598
rect 14207 4534 14556 4564
rect 14207 4500 14246 4534
rect 14280 4500 14319 4534
rect 14353 4500 14392 4534
rect 14426 4526 14556 4534
tri 14556 4526 14594 4564 sw
tri 14689 4526 14727 4564 ne
rect 14727 4526 15097 4564
rect 14426 4502 14594 4526
tri 14594 4502 14618 4526 sw
rect 14426 4500 14618 4502
rect 303 4492 365 4500
tri 365 4492 373 4500 nw
rect 303 4484 329 4492
rect 39 4445 329 4484
tri 329 4456 365 4492 nw
rect 517 4488 14618 4500
tri 14727 4492 14761 4526 ne
rect 14761 4492 14832 4526
rect 14866 4492 15097 4526
rect 517 4456 946 4488
tri 946 4456 978 4488 nw
tri 14157 4456 14189 4488 ne
rect 14189 4456 14618 4488
rect 39 4411 269 4445
rect 303 4411 329 4445
rect 39 4372 329 4411
rect 39 4338 269 4372
rect 303 4338 329 4372
rect 39 4299 329 4338
rect 39 4265 269 4299
rect 303 4265 329 4299
rect 39 4226 329 4265
rect 39 4192 269 4226
rect 303 4192 329 4226
rect 39 4153 329 4192
rect 39 4119 269 4153
rect 303 4119 329 4153
rect 39 4080 329 4119
rect 39 4046 269 4080
rect 303 4046 329 4080
rect 39 4007 329 4046
rect 39 3973 269 4007
rect 303 3973 329 4007
rect 39 3934 329 3973
rect 39 3900 269 3934
rect 303 3900 329 3934
rect 39 3861 329 3900
rect 39 3827 269 3861
rect 303 3827 329 3861
rect 39 3788 329 3827
rect 39 3754 269 3788
rect 303 3754 329 3788
rect 39 3715 329 3754
rect 39 3681 269 3715
rect 303 3681 329 3715
rect 39 3642 329 3681
rect 39 3608 269 3642
rect 303 3608 329 3642
rect 39 3569 329 3608
rect 39 3535 269 3569
rect 303 3535 329 3569
rect 39 3496 329 3535
rect 39 3462 269 3496
rect 303 3462 329 3496
rect 39 3423 329 3462
rect 39 3389 269 3423
rect 303 3389 329 3423
rect 39 3350 329 3389
rect 39 3316 269 3350
rect 303 3316 329 3350
rect 39 3277 329 3316
rect 39 3243 269 3277
rect 303 3243 329 3277
rect 39 3204 329 3243
rect 39 3170 269 3204
rect 303 3170 329 3204
rect 39 3131 329 3170
rect 39 3097 269 3131
rect 303 3097 329 3131
rect 39 3058 329 3097
rect 39 3024 269 3058
rect 303 3024 329 3058
rect 39 2985 329 3024
rect 39 2951 269 2985
rect 303 2951 329 2985
rect 39 2912 329 2951
rect 39 2878 269 2912
rect 303 2878 329 2912
rect 39 2839 329 2878
rect 39 2805 269 2839
rect 303 2805 329 2839
rect 39 2766 329 2805
rect 39 2732 269 2766
rect 303 2732 329 2766
rect 39 2693 329 2732
rect 39 2659 269 2693
rect 303 2659 329 2693
rect 39 2620 329 2659
rect 39 2586 269 2620
rect 303 2586 329 2620
rect 39 2547 329 2586
rect 39 2513 269 2547
rect 303 2513 329 2547
rect 39 2474 329 2513
rect 39 2440 269 2474
rect 303 2440 329 2474
rect 39 2401 329 2440
rect 39 2367 269 2401
rect 303 2367 329 2401
rect 39 2328 329 2367
rect 39 2294 269 2328
rect 303 2294 329 2328
rect 39 2255 329 2294
rect 39 2221 269 2255
rect 303 2221 329 2255
rect 39 2182 329 2221
rect 39 2148 269 2182
rect 303 2148 329 2182
rect 39 2109 329 2148
rect 39 2075 269 2109
rect 303 2075 329 2109
rect 39 2036 329 2075
rect 39 2002 269 2036
rect 303 2002 329 2036
rect 39 1963 329 2002
rect 39 1929 269 1963
rect 303 1929 329 1963
rect 39 1890 329 1929
rect 39 1856 269 1890
rect 303 1856 329 1890
rect 39 1817 329 1856
rect 39 1783 269 1817
rect 303 1783 329 1817
rect 39 1744 329 1783
rect 39 1710 269 1744
rect 303 1710 329 1744
rect 39 1671 329 1710
rect 39 1637 269 1671
rect 303 1637 329 1671
rect 39 1598 329 1637
rect 39 1564 269 1598
rect 303 1564 329 1598
rect 39 1525 329 1564
rect 39 1491 269 1525
rect 303 1491 329 1525
rect 39 1452 329 1491
rect 39 1418 269 1452
rect 303 1418 329 1452
rect 39 1379 329 1418
rect 39 1345 269 1379
rect 303 1345 329 1379
rect 39 1306 329 1345
rect 39 1272 269 1306
rect 303 1272 329 1306
rect 39 1233 329 1272
rect 39 1199 269 1233
rect 303 1199 329 1233
rect 39 1159 329 1199
rect 39 1125 269 1159
rect 303 1125 329 1159
rect 39 1085 329 1125
rect 39 1051 269 1085
rect 303 1051 329 1085
rect 39 1011 329 1051
rect 39 977 269 1011
rect 303 977 329 1011
rect 39 937 329 977
rect 39 903 269 937
rect 303 903 329 937
rect 39 863 329 903
rect 517 4404 518 4456
rect 570 4404 590 4456
rect 642 4404 662 4456
rect 714 4445 734 4456
rect 786 4432 922 4456
tri 922 4432 946 4456 nw
tri 14189 4446 14199 4456 ne
rect 14199 4446 14428 4456
tri 14199 4432 14213 4446 ne
rect 14213 4432 14428 4446
rect 786 4404 888 4432
rect 517 4392 529 4404
rect 563 4392 601 4404
rect 635 4392 674 4404
rect 517 4390 674 4392
rect 780 4398 888 4404
tri 888 4398 922 4432 nw
tri 14213 4398 14247 4432 ne
rect 14247 4398 14356 4432
rect 14390 4398 14428 4432
rect 14462 4426 14618 4456
tri 14761 4454 14799 4492 ne
rect 14799 4454 15097 4492
tri 14799 4446 14807 4454 ne
rect 780 4390 849 4398
rect 517 4338 518 4390
rect 570 4338 590 4390
rect 642 4338 662 4390
rect 786 4359 849 4390
tri 849 4359 888 4398 nw
tri 14247 4359 14286 4398 ne
rect 14286 4359 14428 4398
rect 786 4338 815 4359
rect 517 4325 529 4338
rect 563 4325 601 4338
rect 635 4325 674 4338
rect 780 4325 815 4338
tri 815 4325 849 4359 nw
tri 14286 4325 14320 4359 ne
rect 14320 4325 14356 4359
rect 14390 4325 14428 4359
rect 517 4273 518 4325
rect 570 4273 590 4325
rect 642 4273 662 4325
tri 786 4296 815 4325 nw
tri 14320 4296 14349 4325 ne
rect 14349 4296 14428 4325
tri 14349 4295 14350 4296 ne
rect 517 4260 529 4273
rect 563 4260 601 4273
rect 635 4260 674 4273
rect 780 4260 786 4273
rect 517 4208 518 4260
rect 570 4208 590 4260
rect 642 4208 662 4260
rect 517 4201 674 4208
rect 517 4195 529 4201
rect 563 4195 601 4201
rect 635 4195 674 4201
rect 780 4195 786 4208
rect 517 4143 518 4195
rect 570 4143 590 4195
rect 642 4143 662 4195
rect 517 4130 674 4143
rect 780 4130 786 4143
rect 14350 4286 14428 4296
rect 14350 4252 14356 4286
rect 14390 4252 14428 4286
rect 14350 4213 14428 4252
rect 14350 4179 14356 4213
rect 14390 4179 14428 4213
rect 14350 4140 14428 4179
rect 517 4078 518 4130
rect 570 4078 590 4130
rect 642 4078 662 4130
rect 517 4065 674 4078
rect 780 4065 786 4078
rect 517 4013 518 4065
rect 570 4013 590 4065
rect 642 4013 662 4065
rect 517 4000 674 4013
rect 780 4000 786 4013
rect 517 3948 518 4000
rect 570 3948 590 4000
rect 642 3948 662 4000
rect 517 3944 529 3948
rect 563 3944 601 3948
rect 635 3944 674 3948
rect 517 3935 674 3944
rect 780 3935 786 3948
rect 517 3883 518 3935
rect 570 3883 590 3935
rect 642 3883 662 3935
rect 517 3870 529 3883
rect 563 3870 601 3883
rect 635 3870 674 3883
rect 780 3870 786 3883
rect 517 3818 518 3870
rect 570 3818 590 3870
rect 642 3818 662 3870
rect 517 3805 674 3818
rect 780 3805 786 3818
rect 517 3753 518 3805
rect 570 3753 590 3805
rect 642 3753 662 3805
rect 517 3740 674 3753
rect 780 3740 786 3753
rect 517 3688 518 3740
rect 570 3688 590 3740
rect 642 3688 662 3740
rect 517 3686 529 3688
rect 563 3686 601 3688
rect 635 3686 674 3688
rect 517 3675 674 3686
rect 780 3675 786 3688
rect 517 3623 518 3675
rect 570 3623 590 3675
rect 642 3623 662 3675
rect 517 3612 529 3623
rect 563 3612 601 3623
rect 635 3612 674 3623
rect 517 3610 674 3612
rect 780 3610 786 3623
rect 517 3558 518 3610
rect 570 3558 590 3610
rect 642 3558 662 3610
rect 517 3545 529 3558
rect 563 3545 601 3558
rect 635 3545 674 3558
rect 780 3545 786 3558
rect 517 3493 518 3545
rect 570 3493 590 3545
rect 642 3493 662 3545
rect 517 3480 529 3493
rect 563 3480 601 3493
rect 635 3480 674 3493
rect 780 3480 786 3493
rect 517 3428 518 3480
rect 570 3428 590 3480
rect 642 3428 662 3480
rect 517 3424 674 3428
rect 517 3415 529 3424
rect 563 3415 601 3424
rect 635 3415 674 3424
rect 780 3415 786 3428
rect 517 3363 518 3415
rect 570 3363 590 3415
rect 642 3363 662 3415
rect 517 3350 674 3363
rect 780 3350 786 3363
rect 517 3298 518 3350
rect 570 3298 590 3350
rect 642 3298 662 3350
rect 517 3285 674 3298
rect 780 3285 786 3298
rect 517 3233 518 3285
rect 570 3233 590 3285
rect 642 3233 662 3285
rect 517 3220 674 3233
rect 780 3220 786 3233
rect 517 3168 518 3220
rect 570 3168 590 3220
rect 642 3168 662 3220
rect 517 3155 674 3168
rect 780 3155 786 3168
rect 517 3103 518 3155
rect 570 3103 590 3155
rect 642 3103 662 3155
rect 517 3094 529 3103
rect 563 3094 601 3103
rect 635 3094 674 3103
rect 517 3090 674 3094
rect 780 3090 786 3103
rect 517 3038 518 3090
rect 570 3038 590 3090
rect 642 3038 662 3090
rect 517 3025 529 3038
rect 563 3025 601 3038
rect 635 3025 674 3038
rect 780 3025 786 3038
rect 517 2973 518 3025
rect 570 2973 590 3025
rect 642 2973 662 3025
rect 517 2960 529 2973
rect 563 2960 601 2973
rect 635 2960 674 2973
rect 780 2960 786 2973
rect 517 2908 518 2960
rect 570 2908 590 2960
rect 642 2908 662 2960
rect 517 2906 674 2908
rect 517 2895 529 2906
rect 563 2895 601 2906
rect 635 2895 674 2906
rect 780 2895 786 2908
rect 517 2843 518 2895
rect 570 2843 590 2895
rect 642 2843 662 2895
rect 517 2832 674 2843
rect 517 2830 529 2832
rect 563 2830 601 2832
rect 635 2830 674 2832
rect 780 2830 786 2843
rect 517 2778 518 2830
rect 570 2778 590 2830
rect 642 2778 662 2830
rect 517 2765 674 2778
rect 780 2765 786 2778
rect 517 2713 518 2765
rect 570 2713 590 2765
rect 642 2713 662 2765
rect 517 2700 674 2713
rect 780 2700 786 2713
rect 517 2648 518 2700
rect 570 2648 590 2700
rect 642 2648 662 2700
rect 517 2635 674 2648
rect 780 2635 786 2648
rect 517 2583 518 2635
rect 570 2583 590 2635
rect 642 2583 662 2635
rect 517 2576 529 2583
rect 563 2576 601 2583
rect 635 2576 674 2583
rect 517 2570 674 2576
rect 780 2570 786 2583
rect 517 2518 518 2570
rect 570 2518 590 2570
rect 642 2518 662 2570
rect 517 2505 529 2518
rect 563 2505 601 2518
rect 635 2505 674 2518
rect 780 2505 786 2518
rect 517 2453 518 2505
rect 570 2453 590 2505
rect 642 2453 662 2505
rect 517 2440 529 2453
rect 563 2440 601 2453
rect 635 2440 674 2453
rect 780 2440 786 2453
rect 517 2388 518 2440
rect 570 2388 590 2440
rect 642 2388 662 2440
rect 517 2375 529 2388
rect 563 2375 601 2388
rect 635 2375 674 2388
rect 780 2375 786 2388
rect 517 2323 518 2375
rect 570 2323 590 2375
rect 642 2323 662 2375
rect 517 2316 674 2323
rect 517 2310 529 2316
rect 563 2310 601 2316
rect 635 2310 674 2316
rect 780 2310 786 2323
rect 517 2258 518 2310
rect 570 2258 590 2310
rect 642 2258 662 2310
rect 517 2245 674 2258
rect 780 2245 786 2258
rect 517 2193 518 2245
rect 570 2193 590 2245
rect 642 2193 662 2245
rect 517 2180 674 2193
rect 780 2180 786 2193
rect 517 2128 518 2180
rect 570 2128 590 2180
rect 642 2128 662 2180
rect 517 2115 674 2128
rect 780 2115 786 2128
rect 517 2063 518 2115
rect 570 2063 590 2115
rect 642 2063 662 2115
rect 517 2050 674 2063
rect 780 2050 786 2063
rect 517 1998 518 2050
rect 570 1998 590 2050
rect 642 1998 662 2050
rect 517 1990 529 1998
rect 563 1990 601 1998
rect 635 1990 674 1998
rect 517 1985 674 1990
rect 780 1985 786 1998
rect 517 1933 518 1985
rect 570 1933 590 1985
rect 642 1933 662 1985
rect 517 1920 529 1933
rect 563 1920 601 1933
rect 635 1920 674 1933
rect 780 1920 786 1933
rect 517 1868 518 1920
rect 570 1868 590 1920
rect 642 1868 662 1920
rect 517 1855 529 1868
rect 563 1855 601 1868
rect 635 1855 674 1868
rect 780 1855 786 1868
rect 517 1803 518 1855
rect 570 1803 590 1855
rect 642 1803 662 1855
rect 517 1790 529 1803
rect 563 1790 601 1803
rect 635 1790 674 1803
rect 780 1790 786 1803
rect 517 1738 518 1790
rect 570 1738 590 1790
rect 642 1738 662 1790
rect 517 1732 674 1738
rect 517 1725 529 1732
rect 563 1725 601 1732
rect 635 1725 674 1732
rect 780 1725 786 1738
rect 517 1673 518 1725
rect 570 1673 590 1725
rect 642 1673 662 1725
rect 517 1660 674 1673
rect 780 1660 786 1673
rect 517 1608 518 1660
rect 570 1608 590 1660
rect 642 1608 662 1660
rect 517 1595 674 1608
rect 780 1595 786 1608
rect 517 1543 518 1595
rect 570 1543 590 1595
rect 642 1543 662 1595
rect 1060 4119 1252 4125
rect 1060 4067 1066 4119
rect 1118 4067 1130 4119
rect 1182 4067 1194 4119
rect 1246 4067 1252 4119
rect 1060 4064 1067 4067
rect 1101 4064 1139 4067
rect 1173 4064 1211 4067
rect 1245 4064 1252 4067
rect 1060 4054 1252 4064
rect 1060 4002 1066 4054
rect 1118 4002 1130 4054
rect 1182 4002 1194 4054
rect 1246 4002 1252 4054
rect 1060 3991 1067 4002
rect 1101 3991 1139 4002
rect 1173 3991 1211 4002
rect 1245 3991 1252 4002
rect 1060 3989 1252 3991
rect 1060 3937 1066 3989
rect 1118 3937 1130 3989
rect 1182 3937 1194 3989
rect 1246 3937 1252 3989
rect 1060 3924 1067 3937
rect 1101 3924 1139 3937
rect 1173 3924 1211 3937
rect 1245 3924 1252 3937
rect 1060 1568 1066 3924
rect 1246 1568 1252 3924
rect 1060 1562 1252 1568
rect 1556 4124 1748 4130
rect 1556 4072 1562 4124
rect 1614 4072 1626 4124
rect 1678 4072 1690 4124
rect 1742 4072 1748 4124
rect 1556 4059 1563 4072
rect 1597 4059 1707 4072
rect 1741 4059 1748 4072
rect 1556 4007 1562 4059
rect 1614 4007 1626 4059
rect 1678 4007 1690 4059
rect 1742 4007 1748 4059
rect 1556 3994 1563 4007
rect 1597 3994 1707 4007
rect 1741 3994 1748 4007
rect 1556 3942 1562 3994
rect 1614 3942 1626 3994
rect 1678 3942 1690 3994
rect 1742 3942 1748 3994
rect 1556 3929 1563 3942
rect 1597 3929 1707 3942
rect 1741 3929 1748 3942
rect 1556 3877 1562 3929
rect 1614 3877 1626 3929
rect 1678 3877 1690 3929
rect 1742 3877 1748 3929
rect 1556 3876 1748 3877
rect 1556 3864 1563 3876
rect 1597 3864 1707 3876
rect 1741 3864 1748 3876
rect 1556 3812 1562 3864
rect 1614 3812 1626 3864
rect 1678 3812 1690 3864
rect 1742 3812 1748 3864
rect 1556 3804 1748 3812
rect 1556 3799 1563 3804
rect 1597 3799 1707 3804
rect 1741 3799 1748 3804
rect 1556 3747 1562 3799
rect 1614 3747 1626 3799
rect 1678 3747 1690 3799
rect 1742 3747 1748 3799
rect 1556 3734 1748 3747
rect 1556 3682 1562 3734
rect 1614 3682 1626 3734
rect 1678 3682 1690 3734
rect 1742 3682 1748 3734
rect 1556 3669 1748 3682
rect 1556 3617 1562 3669
rect 1614 3617 1626 3669
rect 1678 3617 1690 3669
rect 1742 3617 1748 3669
rect 1556 3604 1748 3617
rect 1556 1568 1562 3604
rect 1742 1568 1748 3604
rect 1556 1562 1748 1568
rect 2052 4119 2244 4125
rect 2052 4067 2058 4119
rect 2110 4067 2122 4119
rect 2174 4067 2186 4119
rect 2238 4067 2244 4119
rect 2052 4064 2059 4067
rect 2093 4064 2131 4067
rect 2165 4064 2203 4067
rect 2237 4064 2244 4067
rect 2052 4054 2244 4064
rect 2052 4002 2058 4054
rect 2110 4002 2122 4054
rect 2174 4002 2186 4054
rect 2238 4002 2244 4054
rect 2052 3991 2059 4002
rect 2093 3991 2131 4002
rect 2165 3991 2203 4002
rect 2237 3991 2244 4002
rect 2052 3989 2244 3991
rect 2052 3937 2058 3989
rect 2110 3937 2122 3989
rect 2174 3937 2186 3989
rect 2238 3937 2244 3989
rect 2052 3924 2059 3937
rect 2093 3924 2131 3937
rect 2165 3924 2203 3937
rect 2237 3924 2244 3937
rect 2052 1568 2058 3924
rect 2238 1568 2244 3924
rect 2052 1562 2244 1568
rect 2548 4124 2740 4130
rect 2548 4072 2554 4124
rect 2606 4072 2618 4124
rect 2670 4072 2682 4124
rect 2734 4072 2740 4124
rect 2548 4059 2555 4072
rect 2589 4059 2699 4072
rect 2733 4059 2740 4072
rect 2548 4007 2554 4059
rect 2606 4007 2618 4059
rect 2670 4007 2682 4059
rect 2734 4007 2740 4059
rect 2548 3994 2555 4007
rect 2589 3994 2699 4007
rect 2733 3994 2740 4007
rect 2548 3942 2554 3994
rect 2606 3942 2618 3994
rect 2670 3942 2682 3994
rect 2734 3942 2740 3994
rect 2548 3929 2555 3942
rect 2589 3929 2699 3942
rect 2733 3929 2740 3942
rect 2548 3877 2554 3929
rect 2606 3877 2618 3929
rect 2670 3877 2682 3929
rect 2734 3877 2740 3929
rect 2548 3876 2740 3877
rect 2548 3864 2555 3876
rect 2589 3864 2699 3876
rect 2733 3864 2740 3876
rect 2548 3812 2554 3864
rect 2606 3812 2618 3864
rect 2670 3812 2682 3864
rect 2734 3812 2740 3864
rect 2548 3804 2740 3812
rect 2548 3799 2555 3804
rect 2589 3799 2699 3804
rect 2733 3799 2740 3804
rect 2548 3747 2554 3799
rect 2606 3747 2618 3799
rect 2670 3747 2682 3799
rect 2734 3747 2740 3799
rect 2548 3734 2740 3747
rect 2548 3682 2554 3734
rect 2606 3682 2618 3734
rect 2670 3682 2682 3734
rect 2734 3682 2740 3734
rect 2548 3669 2740 3682
rect 2548 3617 2554 3669
rect 2606 3617 2618 3669
rect 2670 3617 2682 3669
rect 2734 3617 2740 3669
rect 2548 3604 2740 3617
rect 2548 1568 2554 3604
rect 2734 1568 2740 3604
rect 2548 1562 2740 1568
rect 3044 4119 3236 4125
rect 3044 4067 3050 4119
rect 3102 4067 3114 4119
rect 3166 4067 3178 4119
rect 3230 4067 3236 4119
rect 3044 4064 3051 4067
rect 3085 4064 3123 4067
rect 3157 4064 3195 4067
rect 3229 4064 3236 4067
rect 3044 4054 3236 4064
rect 3044 4002 3050 4054
rect 3102 4002 3114 4054
rect 3166 4002 3178 4054
rect 3230 4002 3236 4054
rect 3044 3991 3051 4002
rect 3085 3991 3123 4002
rect 3157 3991 3195 4002
rect 3229 3991 3236 4002
rect 3044 3989 3236 3991
rect 3044 3937 3050 3989
rect 3102 3937 3114 3989
rect 3166 3937 3178 3989
rect 3230 3937 3236 3989
rect 3044 3924 3051 3937
rect 3085 3924 3123 3937
rect 3157 3924 3195 3937
rect 3229 3924 3236 3937
rect 3044 1568 3050 3924
rect 3230 1568 3236 3924
rect 3044 1562 3236 1568
rect 3540 4124 3732 4130
rect 3540 4072 3546 4124
rect 3598 4072 3610 4124
rect 3662 4072 3674 4124
rect 3726 4072 3732 4124
rect 3540 4059 3547 4072
rect 3581 4059 3691 4072
rect 3725 4059 3732 4072
rect 3540 4007 3546 4059
rect 3598 4007 3610 4059
rect 3662 4007 3674 4059
rect 3726 4007 3732 4059
rect 3540 3994 3547 4007
rect 3581 3994 3691 4007
rect 3725 3994 3732 4007
rect 3540 3942 3546 3994
rect 3598 3942 3610 3994
rect 3662 3942 3674 3994
rect 3726 3942 3732 3994
rect 3540 3929 3547 3942
rect 3581 3929 3691 3942
rect 3725 3929 3732 3942
rect 3540 3877 3546 3929
rect 3598 3877 3610 3929
rect 3662 3877 3674 3929
rect 3726 3877 3732 3929
rect 3540 3876 3732 3877
rect 3540 3864 3547 3876
rect 3581 3864 3691 3876
rect 3725 3864 3732 3876
rect 3540 3812 3546 3864
rect 3598 3812 3610 3864
rect 3662 3812 3674 3864
rect 3726 3812 3732 3864
rect 3540 3804 3732 3812
rect 3540 3799 3547 3804
rect 3581 3799 3691 3804
rect 3725 3799 3732 3804
rect 3540 3747 3546 3799
rect 3598 3747 3610 3799
rect 3662 3747 3674 3799
rect 3726 3747 3732 3799
rect 3540 3734 3732 3747
rect 3540 3682 3546 3734
rect 3598 3682 3610 3734
rect 3662 3682 3674 3734
rect 3726 3682 3732 3734
rect 3540 3669 3732 3682
rect 3540 3617 3546 3669
rect 3598 3617 3610 3669
rect 3662 3617 3674 3669
rect 3726 3617 3732 3669
rect 3540 3604 3732 3617
rect 3540 1568 3546 3604
rect 3726 1568 3732 3604
rect 3540 1562 3732 1568
rect 4036 4119 4228 4125
rect 4036 4067 4042 4119
rect 4094 4067 4106 4119
rect 4158 4067 4170 4119
rect 4222 4067 4228 4119
rect 4036 4064 4043 4067
rect 4077 4064 4115 4067
rect 4149 4064 4187 4067
rect 4221 4064 4228 4067
rect 4036 4054 4228 4064
rect 4036 4002 4042 4054
rect 4094 4002 4106 4054
rect 4158 4002 4170 4054
rect 4222 4002 4228 4054
rect 4036 3991 4043 4002
rect 4077 3991 4115 4002
rect 4149 3991 4187 4002
rect 4221 3991 4228 4002
rect 4036 3989 4228 3991
rect 4036 3937 4042 3989
rect 4094 3937 4106 3989
rect 4158 3937 4170 3989
rect 4222 3937 4228 3989
rect 4036 3924 4043 3937
rect 4077 3924 4115 3937
rect 4149 3924 4187 3937
rect 4221 3924 4228 3937
rect 4036 1568 4042 3924
rect 4222 1568 4228 3924
rect 4036 1562 4228 1568
rect 4532 4124 4724 4130
rect 4532 4072 4538 4124
rect 4590 4072 4602 4124
rect 4654 4072 4666 4124
rect 4718 4072 4724 4124
rect 4532 4059 4539 4072
rect 4573 4059 4683 4072
rect 4717 4059 4724 4072
rect 4532 4007 4538 4059
rect 4590 4007 4602 4059
rect 4654 4007 4666 4059
rect 4718 4007 4724 4059
rect 4532 3994 4539 4007
rect 4573 3994 4683 4007
rect 4717 3994 4724 4007
rect 4532 3942 4538 3994
rect 4590 3942 4602 3994
rect 4654 3942 4666 3994
rect 4718 3942 4724 3994
rect 4532 3929 4539 3942
rect 4573 3929 4683 3942
rect 4717 3929 4724 3942
rect 4532 3877 4538 3929
rect 4590 3877 4602 3929
rect 4654 3877 4666 3929
rect 4718 3877 4724 3929
rect 4532 3876 4724 3877
rect 4532 3864 4539 3876
rect 4573 3864 4683 3876
rect 4717 3864 4724 3876
rect 4532 3812 4538 3864
rect 4590 3812 4602 3864
rect 4654 3812 4666 3864
rect 4718 3812 4724 3864
rect 4532 3804 4724 3812
rect 4532 3799 4539 3804
rect 4573 3799 4683 3804
rect 4717 3799 4724 3804
rect 4532 3747 4538 3799
rect 4590 3747 4602 3799
rect 4654 3747 4666 3799
rect 4718 3747 4724 3799
rect 4532 3734 4724 3747
rect 4532 3682 4538 3734
rect 4590 3682 4602 3734
rect 4654 3682 4666 3734
rect 4718 3682 4724 3734
rect 4532 3669 4724 3682
rect 4532 3617 4538 3669
rect 4590 3617 4602 3669
rect 4654 3617 4666 3669
rect 4718 3617 4724 3669
rect 4532 3604 4724 3617
rect 4532 1568 4538 3604
rect 4718 1568 4724 3604
rect 4532 1562 4724 1568
rect 5028 4119 5220 4125
rect 5028 4067 5034 4119
rect 5086 4067 5098 4119
rect 5150 4067 5162 4119
rect 5214 4067 5220 4119
rect 5028 4064 5035 4067
rect 5069 4064 5107 4067
rect 5141 4064 5179 4067
rect 5213 4064 5220 4067
rect 5028 4054 5220 4064
rect 5028 4002 5034 4054
rect 5086 4002 5098 4054
rect 5150 4002 5162 4054
rect 5214 4002 5220 4054
rect 5028 3991 5035 4002
rect 5069 3991 5107 4002
rect 5141 3991 5179 4002
rect 5213 3991 5220 4002
rect 5028 3989 5220 3991
rect 5028 3937 5034 3989
rect 5086 3937 5098 3989
rect 5150 3937 5162 3989
rect 5214 3937 5220 3989
rect 5028 3924 5035 3937
rect 5069 3924 5107 3937
rect 5141 3924 5179 3937
rect 5213 3924 5220 3937
rect 5028 1568 5034 3924
rect 5214 1568 5220 3924
rect 5028 1562 5220 1568
rect 5524 4124 5716 4130
rect 5524 4072 5530 4124
rect 5582 4072 5594 4124
rect 5646 4072 5658 4124
rect 5710 4072 5716 4124
rect 5524 4059 5531 4072
rect 5565 4059 5675 4072
rect 5709 4059 5716 4072
rect 5524 4007 5530 4059
rect 5582 4007 5594 4059
rect 5646 4007 5658 4059
rect 5710 4007 5716 4059
rect 5524 3994 5531 4007
rect 5565 3994 5675 4007
rect 5709 3994 5716 4007
rect 5524 3942 5530 3994
rect 5582 3942 5594 3994
rect 5646 3942 5658 3994
rect 5710 3942 5716 3994
rect 5524 3929 5531 3942
rect 5565 3929 5675 3942
rect 5709 3929 5716 3942
rect 5524 3877 5530 3929
rect 5582 3877 5594 3929
rect 5646 3877 5658 3929
rect 5710 3877 5716 3929
rect 5524 3876 5716 3877
rect 5524 3864 5531 3876
rect 5565 3864 5675 3876
rect 5709 3864 5716 3876
rect 5524 3812 5530 3864
rect 5582 3812 5594 3864
rect 5646 3812 5658 3864
rect 5710 3812 5716 3864
rect 5524 3804 5716 3812
rect 5524 3799 5531 3804
rect 5565 3799 5675 3804
rect 5709 3799 5716 3804
rect 5524 3747 5530 3799
rect 5582 3747 5594 3799
rect 5646 3747 5658 3799
rect 5710 3747 5716 3799
rect 5524 3734 5716 3747
rect 5524 3682 5530 3734
rect 5582 3682 5594 3734
rect 5646 3682 5658 3734
rect 5710 3682 5716 3734
rect 5524 3669 5716 3682
rect 5524 3617 5530 3669
rect 5582 3617 5594 3669
rect 5646 3617 5658 3669
rect 5710 3617 5716 3669
rect 5524 3604 5716 3617
rect 5524 1568 5530 3604
rect 5710 1568 5716 3604
rect 5524 1562 5716 1568
rect 6020 4119 6212 4125
rect 6020 4067 6026 4119
rect 6078 4067 6090 4119
rect 6142 4067 6154 4119
rect 6206 4067 6212 4119
rect 6020 4064 6027 4067
rect 6061 4064 6099 4067
rect 6133 4064 6171 4067
rect 6205 4064 6212 4067
rect 6020 4054 6212 4064
rect 6020 4002 6026 4054
rect 6078 4002 6090 4054
rect 6142 4002 6154 4054
rect 6206 4002 6212 4054
rect 6020 3991 6027 4002
rect 6061 3991 6099 4002
rect 6133 3991 6171 4002
rect 6205 3991 6212 4002
rect 6020 3989 6212 3991
rect 6020 3937 6026 3989
rect 6078 3937 6090 3989
rect 6142 3937 6154 3989
rect 6206 3937 6212 3989
rect 6020 3924 6027 3937
rect 6061 3924 6099 3937
rect 6133 3924 6171 3937
rect 6205 3924 6212 3937
rect 6020 1568 6026 3924
rect 6206 1568 6212 3924
rect 6020 1562 6212 1568
rect 6516 4124 6708 4130
rect 6516 4072 6522 4124
rect 6574 4072 6586 4124
rect 6638 4072 6650 4124
rect 6702 4072 6708 4124
rect 6516 4059 6523 4072
rect 6557 4059 6667 4072
rect 6701 4059 6708 4072
rect 6516 4007 6522 4059
rect 6574 4007 6586 4059
rect 6638 4007 6650 4059
rect 6702 4007 6708 4059
rect 6516 3994 6523 4007
rect 6557 3994 6667 4007
rect 6701 3994 6708 4007
rect 6516 3942 6522 3994
rect 6574 3942 6586 3994
rect 6638 3942 6650 3994
rect 6702 3942 6708 3994
rect 6516 3929 6523 3942
rect 6557 3929 6667 3942
rect 6701 3929 6708 3942
rect 6516 3877 6522 3929
rect 6574 3877 6586 3929
rect 6638 3877 6650 3929
rect 6702 3877 6708 3929
rect 6516 3876 6708 3877
rect 6516 3864 6523 3876
rect 6557 3864 6667 3876
rect 6701 3864 6708 3876
rect 6516 3812 6522 3864
rect 6574 3812 6586 3864
rect 6638 3812 6650 3864
rect 6702 3812 6708 3864
rect 6516 3804 6708 3812
rect 6516 3799 6523 3804
rect 6557 3799 6667 3804
rect 6701 3799 6708 3804
rect 6516 3747 6522 3799
rect 6574 3747 6586 3799
rect 6638 3747 6650 3799
rect 6702 3747 6708 3799
rect 6516 3734 6708 3747
rect 6516 3682 6522 3734
rect 6574 3682 6586 3734
rect 6638 3682 6650 3734
rect 6702 3682 6708 3734
rect 6516 3669 6708 3682
rect 6516 3617 6522 3669
rect 6574 3617 6586 3669
rect 6638 3617 6650 3669
rect 6702 3617 6708 3669
rect 6516 3604 6708 3617
rect 6516 1568 6522 3604
rect 6702 1568 6708 3604
rect 6516 1562 6708 1568
rect 7012 4119 7204 4125
rect 7012 4067 7018 4119
rect 7070 4067 7082 4119
rect 7134 4067 7146 4119
rect 7198 4067 7204 4119
rect 7012 4064 7019 4067
rect 7053 4064 7091 4067
rect 7125 4064 7163 4067
rect 7197 4064 7204 4067
rect 7012 4054 7204 4064
rect 7012 4002 7018 4054
rect 7070 4002 7082 4054
rect 7134 4002 7146 4054
rect 7198 4002 7204 4054
rect 7012 3991 7019 4002
rect 7053 3991 7091 4002
rect 7125 3991 7163 4002
rect 7197 3991 7204 4002
rect 7012 3989 7204 3991
rect 7012 3937 7018 3989
rect 7070 3937 7082 3989
rect 7134 3937 7146 3989
rect 7198 3937 7204 3989
rect 7012 3924 7019 3937
rect 7053 3924 7091 3937
rect 7125 3924 7163 3937
rect 7197 3924 7204 3937
rect 7012 1568 7018 3924
rect 7198 1568 7204 3924
rect 7012 1562 7204 1568
rect 7508 4124 7700 4130
rect 7508 4072 7514 4124
rect 7566 4072 7578 4124
rect 7630 4072 7642 4124
rect 7694 4072 7700 4124
rect 7508 4059 7515 4072
rect 7549 4059 7659 4072
rect 7693 4059 7700 4072
rect 7508 4007 7514 4059
rect 7566 4007 7578 4059
rect 7630 4007 7642 4059
rect 7694 4007 7700 4059
rect 7508 3994 7515 4007
rect 7549 3994 7659 4007
rect 7693 3994 7700 4007
rect 7508 3942 7514 3994
rect 7566 3942 7578 3994
rect 7630 3942 7642 3994
rect 7694 3942 7700 3994
rect 7508 3929 7515 3942
rect 7549 3929 7659 3942
rect 7693 3929 7700 3942
rect 7508 3877 7514 3929
rect 7566 3877 7578 3929
rect 7630 3877 7642 3929
rect 7694 3877 7700 3929
rect 7508 3876 7700 3877
rect 7508 3864 7515 3876
rect 7549 3864 7659 3876
rect 7693 3864 7700 3876
rect 7508 3812 7514 3864
rect 7566 3812 7578 3864
rect 7630 3812 7642 3864
rect 7694 3812 7700 3864
rect 7508 3804 7700 3812
rect 7508 3799 7515 3804
rect 7549 3799 7659 3804
rect 7693 3799 7700 3804
rect 7508 3747 7514 3799
rect 7566 3747 7578 3799
rect 7630 3747 7642 3799
rect 7694 3747 7700 3799
rect 7508 3734 7700 3747
rect 7508 3682 7514 3734
rect 7566 3682 7578 3734
rect 7630 3682 7642 3734
rect 7694 3682 7700 3734
rect 7508 3669 7700 3682
rect 7508 3617 7514 3669
rect 7566 3617 7578 3669
rect 7630 3617 7642 3669
rect 7694 3617 7700 3669
rect 7508 3604 7700 3617
rect 7508 1568 7514 3604
rect 7694 1568 7700 3604
rect 7508 1562 7700 1568
rect 8004 4119 8196 4125
rect 8004 4067 8010 4119
rect 8062 4067 8074 4119
rect 8126 4067 8138 4119
rect 8190 4067 8196 4119
rect 8004 4064 8011 4067
rect 8045 4064 8083 4067
rect 8117 4064 8155 4067
rect 8189 4064 8196 4067
rect 8004 4054 8196 4064
rect 8004 4002 8010 4054
rect 8062 4002 8074 4054
rect 8126 4002 8138 4054
rect 8190 4002 8196 4054
rect 8004 3991 8011 4002
rect 8045 3991 8083 4002
rect 8117 3991 8155 4002
rect 8189 3991 8196 4002
rect 8004 3989 8196 3991
rect 8004 3937 8010 3989
rect 8062 3937 8074 3989
rect 8126 3937 8138 3989
rect 8190 3937 8196 3989
rect 8004 3924 8011 3937
rect 8045 3924 8083 3937
rect 8117 3924 8155 3937
rect 8189 3924 8196 3937
rect 8004 1568 8010 3924
rect 8190 1568 8196 3924
rect 8004 1562 8196 1568
rect 8500 4124 8692 4130
rect 8500 4072 8506 4124
rect 8558 4072 8570 4124
rect 8622 4072 8634 4124
rect 8686 4072 8692 4124
rect 8500 4059 8507 4072
rect 8541 4059 8651 4072
rect 8685 4059 8692 4072
rect 8500 4007 8506 4059
rect 8558 4007 8570 4059
rect 8622 4007 8634 4059
rect 8686 4007 8692 4059
rect 8500 3994 8507 4007
rect 8541 3994 8651 4007
rect 8685 3994 8692 4007
rect 8500 3942 8506 3994
rect 8558 3942 8570 3994
rect 8622 3942 8634 3994
rect 8686 3942 8692 3994
rect 8500 3929 8507 3942
rect 8541 3929 8651 3942
rect 8685 3929 8692 3942
rect 8500 3877 8506 3929
rect 8558 3877 8570 3929
rect 8622 3877 8634 3929
rect 8686 3877 8692 3929
rect 8500 3876 8692 3877
rect 8500 3864 8507 3876
rect 8541 3864 8651 3876
rect 8685 3864 8692 3876
rect 8500 3812 8506 3864
rect 8558 3812 8570 3864
rect 8622 3812 8634 3864
rect 8686 3812 8692 3864
rect 8500 3804 8692 3812
rect 8500 3799 8507 3804
rect 8541 3799 8651 3804
rect 8685 3799 8692 3804
rect 8500 3747 8506 3799
rect 8558 3747 8570 3799
rect 8622 3747 8634 3799
rect 8686 3747 8692 3799
rect 8500 3734 8692 3747
rect 8500 3682 8506 3734
rect 8558 3682 8570 3734
rect 8622 3682 8634 3734
rect 8686 3682 8692 3734
rect 8500 3669 8692 3682
rect 8500 3617 8506 3669
rect 8558 3617 8570 3669
rect 8622 3617 8634 3669
rect 8686 3617 8692 3669
rect 8500 3604 8692 3617
rect 8500 1568 8506 3604
rect 8686 1568 8692 3604
rect 8500 1562 8692 1568
rect 8996 4119 9188 4125
rect 8996 4067 9002 4119
rect 9054 4067 9066 4119
rect 9118 4067 9130 4119
rect 9182 4067 9188 4119
rect 8996 4064 9003 4067
rect 9037 4064 9075 4067
rect 9109 4064 9147 4067
rect 9181 4064 9188 4067
rect 8996 4054 9188 4064
rect 8996 4002 9002 4054
rect 9054 4002 9066 4054
rect 9118 4002 9130 4054
rect 9182 4002 9188 4054
rect 8996 3991 9003 4002
rect 9037 3991 9075 4002
rect 9109 3991 9147 4002
rect 9181 3991 9188 4002
rect 8996 3989 9188 3991
rect 8996 3937 9002 3989
rect 9054 3937 9066 3989
rect 9118 3937 9130 3989
rect 9182 3937 9188 3989
rect 8996 3924 9003 3937
rect 9037 3924 9075 3937
rect 9109 3924 9147 3937
rect 9181 3924 9188 3937
rect 8996 1568 9002 3924
rect 9182 1568 9188 3924
rect 8996 1562 9188 1568
rect 9492 4124 9684 4130
rect 9492 4072 9498 4124
rect 9550 4072 9562 4124
rect 9614 4072 9626 4124
rect 9678 4072 9684 4124
rect 9492 4059 9499 4072
rect 9533 4059 9643 4072
rect 9677 4059 9684 4072
rect 9492 4007 9498 4059
rect 9550 4007 9562 4059
rect 9614 4007 9626 4059
rect 9678 4007 9684 4059
rect 9492 3994 9499 4007
rect 9533 3994 9643 4007
rect 9677 3994 9684 4007
rect 9492 3942 9498 3994
rect 9550 3942 9562 3994
rect 9614 3942 9626 3994
rect 9678 3942 9684 3994
rect 9492 3929 9499 3942
rect 9533 3929 9643 3942
rect 9677 3929 9684 3942
rect 9492 3877 9498 3929
rect 9550 3877 9562 3929
rect 9614 3877 9626 3929
rect 9678 3877 9684 3929
rect 9492 3876 9684 3877
rect 9492 3864 9499 3876
rect 9533 3864 9643 3876
rect 9677 3864 9684 3876
rect 9492 3812 9498 3864
rect 9550 3812 9562 3864
rect 9614 3812 9626 3864
rect 9678 3812 9684 3864
rect 9492 3804 9684 3812
rect 9492 3799 9499 3804
rect 9533 3799 9643 3804
rect 9677 3799 9684 3804
rect 9492 3747 9498 3799
rect 9550 3747 9562 3799
rect 9614 3747 9626 3799
rect 9678 3747 9684 3799
rect 9492 3734 9684 3747
rect 9492 3682 9498 3734
rect 9550 3682 9562 3734
rect 9614 3682 9626 3734
rect 9678 3682 9684 3734
rect 9492 3669 9684 3682
rect 9492 3617 9498 3669
rect 9550 3617 9562 3669
rect 9614 3617 9626 3669
rect 9678 3617 9684 3669
rect 9492 3604 9684 3617
rect 9492 1568 9498 3604
rect 9678 1568 9684 3604
rect 9492 1562 9684 1568
rect 9988 4119 10180 4125
rect 9988 4067 9994 4119
rect 10046 4067 10058 4119
rect 10110 4067 10122 4119
rect 10174 4067 10180 4119
rect 9988 4064 9995 4067
rect 10029 4064 10067 4067
rect 10101 4064 10139 4067
rect 10173 4064 10180 4067
rect 9988 4054 10180 4064
rect 9988 4002 9994 4054
rect 10046 4002 10058 4054
rect 10110 4002 10122 4054
rect 10174 4002 10180 4054
rect 9988 3991 9995 4002
rect 10029 3991 10067 4002
rect 10101 3991 10139 4002
rect 10173 3991 10180 4002
rect 9988 3989 10180 3991
rect 9988 3937 9994 3989
rect 10046 3937 10058 3989
rect 10110 3937 10122 3989
rect 10174 3937 10180 3989
rect 9988 3924 9995 3937
rect 10029 3924 10067 3937
rect 10101 3924 10139 3937
rect 10173 3924 10180 3937
rect 9988 1568 9994 3924
rect 10174 1568 10180 3924
rect 9988 1562 10180 1568
rect 10484 4124 10676 4130
rect 10484 4072 10490 4124
rect 10542 4072 10554 4124
rect 10606 4072 10618 4124
rect 10670 4072 10676 4124
rect 10484 4059 10491 4072
rect 10525 4059 10635 4072
rect 10669 4059 10676 4072
rect 10484 4007 10490 4059
rect 10542 4007 10554 4059
rect 10606 4007 10618 4059
rect 10670 4007 10676 4059
rect 10484 3994 10491 4007
rect 10525 3994 10635 4007
rect 10669 3994 10676 4007
rect 10484 3942 10490 3994
rect 10542 3942 10554 3994
rect 10606 3942 10618 3994
rect 10670 3942 10676 3994
rect 10484 3929 10491 3942
rect 10525 3929 10635 3942
rect 10669 3929 10676 3942
rect 10484 3877 10490 3929
rect 10542 3877 10554 3929
rect 10606 3877 10618 3929
rect 10670 3877 10676 3929
rect 10484 3876 10676 3877
rect 10484 3864 10491 3876
rect 10525 3864 10635 3876
rect 10669 3864 10676 3876
rect 10484 3812 10490 3864
rect 10542 3812 10554 3864
rect 10606 3812 10618 3864
rect 10670 3812 10676 3864
rect 10484 3804 10676 3812
rect 10484 3799 10491 3804
rect 10525 3799 10635 3804
rect 10669 3799 10676 3804
rect 10484 3747 10490 3799
rect 10542 3747 10554 3799
rect 10606 3747 10618 3799
rect 10670 3747 10676 3799
rect 10484 3734 10676 3747
rect 10484 3682 10490 3734
rect 10542 3682 10554 3734
rect 10606 3682 10618 3734
rect 10670 3682 10676 3734
rect 10484 3669 10676 3682
rect 10484 3617 10490 3669
rect 10542 3617 10554 3669
rect 10606 3617 10618 3669
rect 10670 3617 10676 3669
rect 10484 3604 10676 3617
rect 10484 1568 10490 3604
rect 10670 1568 10676 3604
rect 10484 1562 10676 1568
rect 10980 4119 11172 4125
rect 10980 4067 10986 4119
rect 11038 4067 11050 4119
rect 11102 4067 11114 4119
rect 11166 4067 11172 4119
rect 10980 4064 10987 4067
rect 11021 4064 11059 4067
rect 11093 4064 11131 4067
rect 11165 4064 11172 4067
rect 10980 4054 11172 4064
rect 10980 4002 10986 4054
rect 11038 4002 11050 4054
rect 11102 4002 11114 4054
rect 11166 4002 11172 4054
rect 10980 3991 10987 4002
rect 11021 3991 11059 4002
rect 11093 3991 11131 4002
rect 11165 3991 11172 4002
rect 10980 3989 11172 3991
rect 10980 3937 10986 3989
rect 11038 3937 11050 3989
rect 11102 3937 11114 3989
rect 11166 3937 11172 3989
rect 10980 3924 10987 3937
rect 11021 3924 11059 3937
rect 11093 3924 11131 3937
rect 11165 3924 11172 3937
rect 10980 1568 10986 3924
rect 11166 1568 11172 3924
rect 10980 1562 11172 1568
rect 11476 4124 11668 4130
rect 11476 4072 11482 4124
rect 11534 4072 11546 4124
rect 11598 4072 11610 4124
rect 11662 4072 11668 4124
rect 11476 4059 11483 4072
rect 11517 4059 11627 4072
rect 11661 4059 11668 4072
rect 11476 4007 11482 4059
rect 11534 4007 11546 4059
rect 11598 4007 11610 4059
rect 11662 4007 11668 4059
rect 11476 3994 11483 4007
rect 11517 3994 11627 4007
rect 11661 3994 11668 4007
rect 11476 3942 11482 3994
rect 11534 3942 11546 3994
rect 11598 3942 11610 3994
rect 11662 3942 11668 3994
rect 11476 3929 11483 3942
rect 11517 3929 11627 3942
rect 11661 3929 11668 3942
rect 11476 3877 11482 3929
rect 11534 3877 11546 3929
rect 11598 3877 11610 3929
rect 11662 3877 11668 3929
rect 11476 3876 11668 3877
rect 11476 3864 11483 3876
rect 11517 3864 11627 3876
rect 11661 3864 11668 3876
rect 11476 3812 11482 3864
rect 11534 3812 11546 3864
rect 11598 3812 11610 3864
rect 11662 3812 11668 3864
rect 11476 3804 11668 3812
rect 11476 3799 11483 3804
rect 11517 3799 11627 3804
rect 11661 3799 11668 3804
rect 11476 3747 11482 3799
rect 11534 3747 11546 3799
rect 11598 3747 11610 3799
rect 11662 3747 11668 3799
rect 11476 3734 11668 3747
rect 11476 3682 11482 3734
rect 11534 3682 11546 3734
rect 11598 3682 11610 3734
rect 11662 3682 11668 3734
rect 11476 3669 11668 3682
rect 11476 3617 11482 3669
rect 11534 3617 11546 3669
rect 11598 3617 11610 3669
rect 11662 3617 11668 3669
rect 11476 3604 11668 3617
rect 11476 1568 11482 3604
rect 11662 1568 11668 3604
rect 11476 1562 11668 1568
rect 11972 4119 12164 4125
rect 11972 4067 11978 4119
rect 12030 4067 12042 4119
rect 12094 4067 12106 4119
rect 12158 4067 12164 4119
rect 11972 4064 11979 4067
rect 12013 4064 12051 4067
rect 12085 4064 12123 4067
rect 12157 4064 12164 4067
rect 11972 4054 12164 4064
rect 11972 4002 11978 4054
rect 12030 4002 12042 4054
rect 12094 4002 12106 4054
rect 12158 4002 12164 4054
rect 11972 3991 11979 4002
rect 12013 3991 12051 4002
rect 12085 3991 12123 4002
rect 12157 3991 12164 4002
rect 11972 3989 12164 3991
rect 11972 3937 11978 3989
rect 12030 3937 12042 3989
rect 12094 3937 12106 3989
rect 12158 3937 12164 3989
rect 11972 3924 11979 3937
rect 12013 3924 12051 3937
rect 12085 3924 12123 3937
rect 12157 3924 12164 3937
rect 11972 1568 11978 3924
rect 12158 1568 12164 3924
rect 11972 1562 12164 1568
rect 12468 4124 12660 4130
rect 12468 4072 12474 4124
rect 12526 4072 12538 4124
rect 12590 4072 12602 4124
rect 12654 4072 12660 4124
rect 12468 4059 12475 4072
rect 12509 4059 12619 4072
rect 12653 4059 12660 4072
rect 12468 4007 12474 4059
rect 12526 4007 12538 4059
rect 12590 4007 12602 4059
rect 12654 4007 12660 4059
rect 12468 3994 12475 4007
rect 12509 3994 12619 4007
rect 12653 3994 12660 4007
rect 12468 3942 12474 3994
rect 12526 3942 12538 3994
rect 12590 3942 12602 3994
rect 12654 3942 12660 3994
rect 12468 3929 12475 3942
rect 12509 3929 12619 3942
rect 12653 3929 12660 3942
rect 12468 3877 12474 3929
rect 12526 3877 12538 3929
rect 12590 3877 12602 3929
rect 12654 3877 12660 3929
rect 12468 3876 12660 3877
rect 12468 3864 12475 3876
rect 12509 3864 12619 3876
rect 12653 3864 12660 3876
rect 12468 3812 12474 3864
rect 12526 3812 12538 3864
rect 12590 3812 12602 3864
rect 12654 3812 12660 3864
rect 12468 3804 12660 3812
rect 12468 3799 12475 3804
rect 12509 3799 12619 3804
rect 12653 3799 12660 3804
rect 12468 3747 12474 3799
rect 12526 3747 12538 3799
rect 12590 3747 12602 3799
rect 12654 3747 12660 3799
rect 12468 3734 12660 3747
rect 12468 3682 12474 3734
rect 12526 3682 12538 3734
rect 12590 3682 12602 3734
rect 12654 3682 12660 3734
rect 12468 3669 12660 3682
rect 12468 3617 12474 3669
rect 12526 3617 12538 3669
rect 12590 3617 12602 3669
rect 12654 3617 12660 3669
rect 12468 3604 12660 3617
rect 12468 1568 12474 3604
rect 12654 1568 12660 3604
rect 12468 1562 12660 1568
rect 12964 4119 13156 4125
rect 12964 4067 12970 4119
rect 13022 4067 13034 4119
rect 13086 4067 13098 4119
rect 13150 4067 13156 4119
rect 12964 4064 12971 4067
rect 13005 4064 13043 4067
rect 13077 4064 13115 4067
rect 13149 4064 13156 4067
rect 12964 4054 13156 4064
rect 12964 4002 12970 4054
rect 13022 4002 13034 4054
rect 13086 4002 13098 4054
rect 13150 4002 13156 4054
rect 12964 3991 12971 4002
rect 13005 3991 13043 4002
rect 13077 3991 13115 4002
rect 13149 3991 13156 4002
rect 12964 3989 13156 3991
rect 12964 3937 12970 3989
rect 13022 3937 13034 3989
rect 13086 3937 13098 3989
rect 13150 3937 13156 3989
rect 12964 3924 12971 3937
rect 13005 3924 13043 3937
rect 13077 3924 13115 3937
rect 13149 3924 13156 3937
rect 12964 1568 12970 3924
rect 13150 1568 13156 3924
rect 12964 1562 13156 1568
rect 13460 4124 13652 4130
rect 13460 4072 13466 4124
rect 13518 4072 13530 4124
rect 13582 4072 13594 4124
rect 13646 4072 13652 4124
rect 13460 4059 13467 4072
rect 13501 4059 13611 4072
rect 13645 4059 13652 4072
rect 13460 4007 13466 4059
rect 13518 4007 13530 4059
rect 13582 4007 13594 4059
rect 13646 4007 13652 4059
rect 13460 3994 13467 4007
rect 13501 3994 13611 4007
rect 13645 3994 13652 4007
rect 13460 3942 13466 3994
rect 13518 3942 13530 3994
rect 13582 3942 13594 3994
rect 13646 3942 13652 3994
rect 13460 3929 13467 3942
rect 13501 3929 13611 3942
rect 13645 3929 13652 3942
rect 13460 3877 13466 3929
rect 13518 3877 13530 3929
rect 13582 3877 13594 3929
rect 13646 3877 13652 3929
rect 13460 3876 13652 3877
rect 13460 3864 13467 3876
rect 13501 3864 13611 3876
rect 13645 3864 13652 3876
rect 13460 3812 13466 3864
rect 13518 3812 13530 3864
rect 13582 3812 13594 3864
rect 13646 3812 13652 3864
rect 13460 3804 13652 3812
rect 13460 3799 13467 3804
rect 13501 3799 13611 3804
rect 13645 3799 13652 3804
rect 13460 3747 13466 3799
rect 13518 3747 13530 3799
rect 13582 3747 13594 3799
rect 13646 3747 13652 3799
rect 13460 3734 13652 3747
rect 13460 3682 13466 3734
rect 13518 3682 13530 3734
rect 13582 3682 13594 3734
rect 13646 3682 13652 3734
rect 13460 3669 13652 3682
rect 13460 3617 13466 3669
rect 13518 3617 13530 3669
rect 13582 3617 13594 3669
rect 13646 3617 13652 3669
rect 13460 3604 13652 3617
rect 13460 1568 13466 3604
rect 13646 1568 13652 3604
rect 13460 1562 13652 1568
rect 13990 4124 14135 4130
rect 13990 4072 13991 4124
rect 14043 4072 14083 4124
rect 13990 4064 13999 4072
rect 14033 4064 14135 4072
rect 13990 4060 14135 4064
rect 13990 4008 13991 4060
rect 14043 4008 14083 4060
rect 13990 3996 13999 4008
rect 14033 3996 14135 4008
rect 13990 3944 13991 3996
rect 14043 3944 14083 3996
rect 13990 3932 13999 3944
rect 14033 3932 14135 3944
rect 13990 3880 13991 3932
rect 14043 3880 14083 3932
rect 13990 3879 14135 3880
rect 13990 3868 13999 3879
rect 14033 3868 14135 3879
rect 13990 3816 13991 3868
rect 14043 3816 14083 3868
rect 13990 3806 14135 3816
rect 13990 3804 13999 3806
rect 14033 3804 14135 3806
rect 13990 3752 13991 3804
rect 14043 3752 14083 3804
rect 13990 3740 14135 3752
rect 13990 3688 13991 3740
rect 14043 3688 14083 3740
rect 13990 3676 14135 3688
rect 13990 3624 13991 3676
rect 14043 3624 14083 3676
rect 13990 3612 14135 3624
rect 13990 3560 13991 3612
rect 14043 3560 14083 3612
rect 13990 3553 13999 3560
rect 14033 3553 14135 3560
rect 13990 3548 14135 3553
rect 13990 3496 13991 3548
rect 14043 3496 14083 3548
rect 13990 3484 13999 3496
rect 14033 3484 14135 3496
rect 13990 3432 13991 3484
rect 14043 3432 14083 3484
rect 13990 3420 13999 3432
rect 14033 3420 14135 3432
rect 13990 3368 13991 3420
rect 14043 3368 14083 3420
rect 13990 3356 13999 3368
rect 14033 3356 14135 3368
rect 13990 3304 13991 3356
rect 14043 3304 14083 3356
rect 13990 3295 14135 3304
rect 13990 3292 13999 3295
rect 14033 3292 14135 3295
rect 13990 3240 13991 3292
rect 14043 3240 14083 3292
rect 13990 3228 14135 3240
rect 13990 3176 13991 3228
rect 14043 3176 14083 3228
rect 13990 3164 14135 3176
rect 13990 3112 13991 3164
rect 14043 3112 14083 3164
rect 13990 3100 14135 3112
rect 13990 3048 13991 3100
rect 14043 3048 14083 3100
rect 13990 3042 13999 3048
rect 14033 3042 14135 3048
rect 13990 3036 14135 3042
rect 13990 2984 13991 3036
rect 14043 2984 14083 3036
rect 13990 2972 13999 2984
rect 14033 2972 14135 2984
rect 13990 2920 13991 2972
rect 14043 2920 14083 2972
rect 13990 2908 13999 2920
rect 14033 2908 14135 2920
rect 13990 2856 13991 2908
rect 14043 2856 14083 2908
rect 13990 2844 13999 2856
rect 14033 2844 14135 2856
rect 13990 2792 13991 2844
rect 14043 2792 14083 2844
rect 13990 2784 14135 2792
rect 13990 2780 13999 2784
rect 14033 2780 14135 2784
rect 13990 2728 13991 2780
rect 14043 2728 14083 2780
rect 13990 2716 14135 2728
rect 13990 2664 13991 2716
rect 14043 2664 14083 2716
rect 13990 2652 14135 2664
rect 13990 2600 13991 2652
rect 14043 2600 14083 2652
rect 13990 2588 14135 2600
rect 13990 2536 13991 2588
rect 14043 2536 14083 2588
rect 13990 2531 13999 2536
rect 14033 2531 14135 2536
rect 13990 2524 14135 2531
rect 13990 2472 13991 2524
rect 14043 2472 14083 2524
rect 13990 2460 13999 2472
rect 14033 2460 14135 2472
rect 13990 2408 13991 2460
rect 14043 2408 14083 2460
rect 13990 2396 13999 2408
rect 14033 2396 14135 2408
rect 13990 2344 13991 2396
rect 14043 2344 14083 2396
rect 13990 2332 13999 2344
rect 14033 2332 14135 2344
rect 13990 2280 13991 2332
rect 14043 2280 14083 2332
rect 13990 2273 14135 2280
rect 13990 2268 13999 2273
rect 14033 2268 14135 2273
rect 13990 2216 13991 2268
rect 14043 2216 14083 2268
rect 13990 2204 14135 2216
rect 13990 2152 13991 2204
rect 14043 2152 14083 2204
rect 13990 2140 14135 2152
rect 13990 2088 13991 2140
rect 14043 2088 14083 2140
rect 13990 2075 14135 2088
rect 13990 2023 13991 2075
rect 14043 2023 14083 2075
rect 13990 2018 13999 2023
rect 14033 2018 14135 2023
rect 13990 2010 14135 2018
rect 13990 1958 13991 2010
rect 14043 1958 14083 2010
rect 13990 1945 13999 1958
rect 14033 1945 14135 1958
rect 13990 1893 13991 1945
rect 14043 1893 14083 1945
rect 13990 1880 13999 1893
rect 14033 1880 14135 1893
rect 13990 1828 13991 1880
rect 14043 1828 14083 1880
rect 13990 1815 13999 1828
rect 14033 1815 14135 1828
rect 13990 1763 13991 1815
rect 14043 1763 14083 1815
rect 13990 1756 14135 1763
rect 13990 1750 13999 1756
rect 14033 1750 14135 1756
rect 13990 1698 13991 1750
rect 14043 1698 14083 1750
rect 13990 1685 14135 1698
rect 13990 1633 13991 1685
rect 14043 1633 14083 1685
rect 13990 1620 14135 1633
rect 13990 1568 13991 1620
rect 14043 1568 14083 1620
rect 13990 1562 14135 1568
rect 14350 4124 14356 4140
rect 14390 4124 14428 4140
rect 14606 4124 14618 4426
rect 14402 4072 14422 4124
rect 14350 4067 14428 4072
rect 14350 4059 14356 4067
rect 14390 4059 14428 4067
rect 14606 4059 14618 4072
rect 14402 4007 14422 4059
rect 14350 3994 14428 4007
rect 14606 3994 14618 4007
rect 14402 3942 14422 3994
rect 14474 3942 14494 3960
rect 14546 3942 14566 3960
rect 14350 3929 14428 3942
rect 14462 3929 14618 3942
rect 14402 3877 14422 3929
rect 14474 3877 14494 3929
rect 14546 3877 14566 3929
rect 14350 3864 14428 3877
rect 14462 3864 14618 3877
rect 14402 3812 14422 3864
rect 14474 3812 14494 3864
rect 14546 3812 14566 3864
rect 14350 3808 14618 3812
rect 14350 3799 14428 3808
rect 14462 3799 14618 3808
rect 14402 3747 14422 3799
rect 14474 3747 14494 3799
rect 14546 3747 14566 3799
rect 14350 3741 14356 3747
rect 14390 3741 14500 3747
rect 14534 3741 14572 3747
rect 14606 3741 14618 3747
rect 14350 3736 14618 3741
rect 14350 3734 14428 3736
rect 14462 3734 14618 3736
rect 14402 3682 14422 3734
rect 14474 3682 14494 3734
rect 14546 3682 14566 3734
rect 14350 3669 14356 3682
rect 14390 3669 14500 3682
rect 14534 3669 14572 3682
rect 14606 3669 14618 3682
rect 14402 3617 14422 3669
rect 14474 3617 14494 3669
rect 14546 3617 14566 3669
rect 14350 3604 14356 3617
rect 14390 3604 14500 3617
rect 14534 3604 14572 3617
rect 14606 3604 14618 3617
rect 14402 3552 14422 3604
rect 14474 3552 14494 3604
rect 14546 3552 14566 3604
rect 14350 3540 14356 3552
rect 14390 3540 14500 3552
rect 14534 3540 14572 3552
rect 14606 3540 14618 3552
rect 14402 3488 14422 3540
rect 14474 3488 14494 3540
rect 14546 3488 14566 3540
rect 14350 3486 14428 3488
rect 14462 3486 14618 3488
rect 14350 3483 14618 3486
rect 14350 3476 14356 3483
rect 14390 3476 14500 3483
rect 14534 3476 14572 3483
rect 14606 3476 14618 3483
rect 14402 3424 14422 3476
rect 14474 3424 14494 3476
rect 14546 3424 14566 3476
rect 14350 3414 14428 3424
rect 14462 3414 14618 3424
rect 14350 3412 14618 3414
rect 14402 3360 14422 3412
rect 14474 3360 14494 3412
rect 14546 3360 14566 3412
rect 14350 3348 14428 3360
rect 14462 3348 14618 3360
rect 14402 3296 14422 3348
rect 14474 3296 14494 3348
rect 14546 3296 14566 3348
rect 14350 3284 14428 3296
rect 14462 3284 14618 3296
rect 14402 3232 14422 3284
rect 14474 3232 14494 3284
rect 14546 3232 14566 3284
rect 14350 3230 14356 3232
rect 14390 3230 14428 3232
rect 14350 3220 14428 3230
rect 14462 3230 14500 3232
rect 14534 3230 14572 3232
rect 14606 3230 14618 3232
rect 14462 3220 14618 3230
rect 14402 3168 14422 3220
rect 14474 3168 14494 3220
rect 14546 3168 14566 3220
rect 14350 3157 14356 3168
rect 14390 3160 14500 3168
rect 14390 3157 14428 3160
rect 14350 3156 14428 3157
rect 14462 3157 14500 3160
rect 14534 3157 14572 3168
rect 14606 3157 14618 3168
rect 14462 3156 14618 3157
rect 14402 3104 14422 3156
rect 14474 3104 14494 3156
rect 14546 3104 14566 3156
rect 14350 3092 14356 3104
rect 14390 3092 14500 3104
rect 14534 3092 14572 3104
rect 14606 3092 14618 3104
rect 14402 3040 14422 3092
rect 14474 3040 14494 3092
rect 14546 3040 14566 3092
rect 14350 3028 14356 3040
rect 14390 3028 14500 3040
rect 14534 3028 14572 3040
rect 14606 3028 14618 3040
rect 14402 2976 14422 3028
rect 14474 2976 14494 3028
rect 14546 2976 14566 3028
rect 14350 2972 14618 2976
rect 14350 2964 14356 2972
rect 14390 2964 14500 2972
rect 14534 2964 14572 2972
rect 14606 2964 14618 2972
rect 14402 2912 14422 2964
rect 14474 2912 14494 2964
rect 14546 2912 14566 2964
rect 14350 2910 14428 2912
rect 14462 2910 14618 2912
rect 14350 2900 14618 2910
rect 14402 2848 14422 2900
rect 14474 2848 14494 2900
rect 14546 2848 14566 2900
rect 14350 2838 14428 2848
rect 14462 2838 14618 2848
rect 14350 2836 14618 2838
rect 14402 2784 14422 2836
rect 14474 2784 14494 2836
rect 14546 2784 14566 2836
rect 14350 2772 14428 2784
rect 14462 2772 14618 2784
rect 14402 2720 14422 2772
rect 14474 2720 14494 2772
rect 14546 2720 14566 2772
rect 14350 2719 14356 2720
rect 14390 2719 14428 2720
rect 14350 2708 14428 2719
rect 14462 2719 14500 2720
rect 14534 2719 14572 2720
rect 14606 2719 14618 2720
rect 14462 2708 14618 2719
rect 14402 2656 14422 2708
rect 14474 2656 14494 2708
rect 14546 2656 14566 2708
rect 14350 2646 14356 2656
rect 14390 2646 14428 2656
rect 14350 2644 14428 2646
rect 14462 2646 14500 2656
rect 14534 2646 14572 2656
rect 14606 2646 14618 2656
rect 14462 2644 14618 2646
rect 14402 2592 14422 2644
rect 14474 2592 14494 2644
rect 14546 2592 14566 2644
rect 14350 2580 14356 2592
rect 14390 2584 14500 2592
rect 14390 2580 14428 2584
rect 14462 2580 14500 2584
rect 14534 2580 14572 2592
rect 14606 2580 14618 2592
rect 14402 2528 14422 2580
rect 14474 2528 14494 2580
rect 14546 2528 14566 2580
rect 14350 2516 14356 2528
rect 14390 2516 14500 2528
rect 14534 2516 14572 2528
rect 14606 2516 14618 2528
rect 14402 2464 14422 2516
rect 14474 2464 14494 2516
rect 14546 2464 14566 2516
rect 14350 2461 14618 2464
rect 14350 2452 14356 2461
rect 14390 2452 14500 2461
rect 14534 2452 14572 2461
rect 14606 2452 14618 2461
rect 14402 2400 14422 2452
rect 14474 2400 14494 2452
rect 14546 2400 14566 2452
rect 14350 2388 14618 2400
rect 14402 2336 14422 2388
rect 14474 2336 14494 2388
rect 14546 2336 14566 2388
rect 14350 2334 14428 2336
rect 14462 2334 14618 2336
rect 14350 2324 14618 2334
rect 14402 2272 14422 2324
rect 14474 2272 14494 2324
rect 14546 2272 14566 2324
rect 14350 2262 14428 2272
rect 14462 2262 14618 2272
rect 14350 2260 14618 2262
rect 14402 2208 14422 2260
rect 14474 2208 14494 2260
rect 14546 2208 14566 2260
rect 14350 2196 14428 2208
rect 14462 2196 14618 2208
rect 14402 2144 14422 2196
rect 14474 2144 14494 2196
rect 14546 2144 14566 2196
rect 14350 2135 14356 2144
rect 14390 2135 14428 2144
rect 14350 2132 14428 2135
rect 14462 2135 14500 2144
rect 14534 2135 14572 2144
rect 14606 2135 14618 2144
rect 14462 2132 14618 2135
rect 14402 2080 14422 2132
rect 14474 2080 14494 2132
rect 14546 2080 14566 2132
rect 14350 2068 14356 2080
rect 14390 2068 14428 2080
rect 14462 2068 14500 2080
rect 14534 2068 14572 2080
rect 14606 2068 14618 2080
rect 14402 2016 14422 2068
rect 14474 2016 14494 2068
rect 14546 2016 14566 2068
rect 14350 2004 14356 2016
rect 14390 2008 14500 2016
rect 14390 2004 14428 2008
rect 14462 2004 14500 2008
rect 14534 2004 14572 2016
rect 14606 2004 14618 2016
rect 14402 1952 14422 2004
rect 14474 1952 14494 2004
rect 14546 1952 14566 2004
rect 14350 1950 14618 1952
rect 14350 1940 14356 1950
rect 14390 1940 14500 1950
rect 14534 1940 14572 1950
rect 14606 1940 14618 1950
rect 14402 1888 14422 1940
rect 14474 1888 14494 1940
rect 14546 1888 14566 1940
rect 14350 1877 14618 1888
rect 14350 1876 14356 1877
rect 14390 1876 14500 1877
rect 14534 1876 14572 1877
rect 14606 1876 14618 1877
rect 14402 1824 14422 1876
rect 14474 1824 14494 1876
rect 14546 1824 14566 1876
rect 14350 1812 14618 1824
rect 14402 1760 14422 1812
rect 14474 1760 14494 1812
rect 14546 1760 14566 1812
rect 14350 1758 14428 1760
rect 14462 1758 14618 1760
rect 14350 1748 14618 1758
rect 14402 1696 14422 1748
rect 14474 1696 14494 1748
rect 14546 1696 14566 1748
rect 14350 1686 14428 1696
rect 14462 1686 14618 1696
rect 14350 1684 14618 1686
rect 14402 1632 14422 1684
rect 14474 1632 14494 1684
rect 14546 1632 14566 1684
rect 14350 1623 14356 1632
rect 14390 1623 14428 1632
rect 14350 1620 14428 1623
rect 14462 1624 14500 1632
rect 14534 1624 14572 1632
rect 14606 1624 14618 1632
rect 14462 1620 14618 1624
rect 14402 1568 14422 1620
rect 14474 1568 14494 1620
rect 14546 1568 14566 1620
rect 517 1530 674 1543
rect 780 1530 786 1543
rect 517 1478 518 1530
rect 570 1478 590 1530
rect 642 1478 662 1530
rect 517 1465 674 1478
rect 780 1465 786 1478
rect 517 1413 518 1465
rect 570 1413 590 1465
rect 642 1413 662 1465
rect 517 1406 529 1413
rect 563 1406 601 1413
rect 635 1406 674 1413
rect 517 1400 674 1406
rect 780 1400 786 1413
rect 517 1348 518 1400
rect 570 1348 590 1400
rect 642 1348 662 1400
rect 517 1335 529 1348
rect 563 1335 601 1348
rect 635 1335 674 1348
rect 780 1335 786 1348
rect 517 1283 518 1335
rect 570 1283 590 1335
rect 642 1283 662 1335
rect 517 1270 529 1283
rect 563 1270 601 1283
rect 635 1270 674 1283
rect 780 1270 786 1283
rect 517 1218 518 1270
rect 570 1218 590 1270
rect 642 1218 662 1270
rect 14350 1549 14356 1568
rect 14390 1549 14428 1568
rect 14350 1542 14428 1549
rect 14462 1551 14500 1568
rect 14534 1551 14572 1568
rect 14606 1551 14618 1568
rect 14462 1542 14618 1551
rect 14350 1512 14618 1542
rect 14350 1509 14500 1512
rect 14350 1475 14356 1509
rect 14390 1504 14500 1509
rect 14390 1475 14428 1504
rect 14350 1470 14428 1475
rect 14462 1478 14500 1504
rect 14534 1478 14572 1512
rect 14606 1478 14618 1512
rect 14462 1470 14618 1478
rect 14350 1439 14618 1470
rect 14350 1435 14500 1439
rect 14350 1401 14356 1435
rect 14390 1432 14500 1435
rect 14390 1401 14428 1432
rect 14350 1398 14428 1401
rect 14462 1405 14500 1432
rect 14534 1405 14572 1439
rect 14606 1405 14618 1439
rect 14462 1398 14618 1405
rect 14350 1366 14618 1398
rect 14350 1361 14500 1366
rect 14350 1327 14356 1361
rect 14390 1360 14500 1361
rect 14390 1327 14428 1360
rect 14350 1326 14428 1327
rect 14462 1332 14500 1360
rect 14534 1332 14572 1366
rect 14606 1332 14618 1366
rect 14462 1326 14618 1332
rect 14350 1293 14618 1326
rect 14350 1288 14500 1293
rect 14350 1287 14428 1288
rect 517 1205 529 1218
rect 563 1205 601 1218
rect 635 1205 674 1218
rect 780 1205 786 1218
rect 517 1153 518 1205
rect 570 1153 590 1205
rect 642 1153 662 1205
rect 517 1148 674 1153
rect 517 1140 529 1148
rect 563 1140 601 1148
rect 635 1140 674 1148
rect 780 1140 786 1153
rect 517 1088 518 1140
rect 570 1088 590 1140
rect 642 1088 662 1140
rect 912 1250 970 1262
rect 912 1216 924 1250
rect 958 1216 970 1250
rect 912 1178 970 1216
rect 912 1144 924 1178
rect 958 1144 970 1178
rect 912 1132 970 1144
rect 1306 1250 1436 1262
rect 1306 1144 1318 1250
rect 1424 1144 1436 1250
rect 1306 1132 1436 1144
rect 1868 1250 1998 1262
rect 1868 1144 1880 1250
rect 1986 1144 1998 1250
rect 1868 1132 1998 1144
rect 2298 1250 2428 1262
rect 2298 1144 2310 1250
rect 2416 1144 2428 1250
rect 2298 1132 2428 1144
rect 2860 1250 2990 1262
rect 2860 1144 2872 1250
rect 2978 1144 2990 1250
rect 2860 1132 2990 1144
rect 3290 1250 3420 1262
rect 3290 1144 3302 1250
rect 3408 1144 3420 1250
rect 3290 1132 3420 1144
rect 3852 1250 3982 1262
rect 3852 1144 3864 1250
rect 3970 1144 3982 1250
rect 3852 1132 3982 1144
rect 4282 1250 4412 1262
rect 4282 1144 4294 1250
rect 4400 1144 4412 1250
rect 4282 1132 4412 1144
rect 4844 1250 4974 1262
rect 4844 1144 4856 1250
rect 4962 1144 4974 1250
rect 4844 1132 4974 1144
rect 5274 1250 5404 1262
rect 5274 1144 5286 1250
rect 5392 1144 5404 1250
rect 5274 1132 5404 1144
rect 5836 1250 5966 1262
rect 5836 1144 5848 1250
rect 5954 1144 5966 1250
rect 5836 1132 5966 1144
rect 6266 1250 6396 1262
rect 6266 1144 6278 1250
rect 6384 1144 6396 1250
rect 6266 1132 6396 1144
rect 6828 1250 6958 1262
rect 6828 1144 6840 1250
rect 6946 1144 6958 1250
rect 6828 1132 6958 1144
rect 7258 1250 7388 1262
rect 7258 1144 7270 1250
rect 7376 1144 7388 1250
rect 7258 1132 7388 1144
rect 7820 1250 7950 1262
rect 7820 1144 7832 1250
rect 7938 1144 7950 1250
rect 7820 1132 7950 1144
rect 8250 1250 8380 1262
rect 8250 1144 8262 1250
rect 8368 1144 8380 1250
rect 8250 1132 8380 1144
rect 8812 1250 8942 1262
rect 8812 1144 8824 1250
rect 8930 1144 8942 1250
rect 8812 1132 8942 1144
rect 9242 1250 9372 1262
rect 9242 1144 9254 1250
rect 9360 1144 9372 1250
rect 9242 1132 9372 1144
rect 9804 1250 9934 1262
rect 9804 1144 9816 1250
rect 9922 1144 9934 1250
rect 9804 1132 9934 1144
rect 10234 1250 10364 1262
rect 10234 1144 10246 1250
rect 10352 1144 10364 1250
rect 10234 1132 10364 1144
rect 10796 1250 10926 1262
rect 10796 1144 10808 1250
rect 10914 1144 10926 1250
rect 10796 1132 10926 1144
rect 11226 1250 11356 1262
rect 11226 1144 11238 1250
rect 11344 1144 11356 1250
rect 11226 1132 11356 1144
rect 11788 1250 11918 1262
rect 11788 1144 11800 1250
rect 11906 1144 11918 1250
rect 11788 1132 11918 1144
rect 12218 1250 12348 1262
rect 12218 1144 12230 1250
rect 12336 1144 12348 1250
rect 12218 1132 12348 1144
rect 12780 1250 12910 1262
rect 12780 1144 12792 1250
rect 12898 1144 12910 1250
rect 12780 1132 12910 1144
rect 13210 1250 13340 1262
rect 13210 1144 13222 1250
rect 13328 1144 13340 1250
rect 13210 1132 13340 1144
rect 13772 1250 13902 1262
rect 13772 1144 13784 1250
rect 13890 1144 13902 1250
rect 13772 1132 13902 1144
rect 14130 1250 14260 1262
rect 14130 1144 14142 1250
rect 14248 1144 14260 1250
rect 14130 1132 14260 1144
rect 14350 1253 14356 1287
rect 14390 1254 14428 1287
rect 14462 1259 14500 1288
rect 14534 1259 14572 1293
rect 14606 1259 14618 1293
rect 14462 1254 14618 1259
rect 14390 1253 14618 1254
rect 14350 1220 14618 1253
rect 14350 1216 14500 1220
rect 14350 1213 14428 1216
rect 14350 1179 14356 1213
rect 14390 1182 14428 1213
rect 14462 1186 14500 1216
rect 14534 1186 14572 1220
rect 14606 1186 14618 1220
rect 14462 1182 14618 1186
rect 14390 1179 14618 1182
rect 14350 1147 14618 1179
rect 14350 1144 14500 1147
rect 14350 1139 14428 1144
rect 517 1075 674 1088
rect 780 1075 786 1088
rect 517 1023 518 1075
rect 570 1023 590 1075
rect 642 1023 662 1075
rect 14350 1105 14356 1139
rect 14390 1110 14428 1139
rect 14462 1113 14500 1144
rect 14534 1113 14572 1147
rect 14606 1113 14618 1147
rect 14462 1110 14618 1113
rect 14390 1105 14618 1110
rect 14350 1074 14618 1105
rect 14350 1072 14500 1074
rect 14350 1065 14428 1072
rect 14350 1031 14356 1065
rect 14390 1038 14428 1065
rect 14462 1040 14500 1072
rect 14534 1040 14572 1074
rect 14606 1040 14618 1074
rect 14462 1038 14618 1040
rect 14390 1031 14618 1038
tri 14349 1024 14350 1025 se
rect 14350 1024 14618 1031
rect 517 1010 674 1023
rect 780 1010 786 1023
rect 517 958 518 1010
rect 570 958 590 1010
rect 642 958 662 1010
tri 786 1001 809 1024 sw
tri 14326 1001 14349 1024 se
rect 14349 1001 14618 1024
rect 786 1000 809 1001
tri 809 1000 810 1001 sw
tri 14325 1000 14326 1001 se
rect 14326 1000 14500 1001
rect 786 991 810 1000
tri 810 991 819 1000 sw
tri 14316 991 14325 1000 se
rect 14325 991 14428 1000
rect 786 958 819 991
rect 517 945 674 958
rect 780 957 819 958
tri 819 957 853 991 sw
tri 14282 957 14316 991 se
rect 14316 957 14356 991
rect 14390 966 14428 991
rect 14462 967 14500 1000
rect 14534 967 14572 1001
rect 14606 967 14618 1001
rect 14462 966 14618 967
rect 14390 957 14618 966
rect 780 945 853 957
rect 517 893 518 945
rect 570 893 590 945
rect 642 893 662 945
rect 714 893 734 894
rect 786 928 853 945
tri 853 928 882 957 sw
tri 14253 928 14282 957 se
rect 14282 928 14618 957
rect 786 917 882 928
tri 882 917 893 928 sw
tri 14242 917 14253 928 se
rect 14253 917 14428 928
rect 786 893 893 917
rect 517 883 746 893
rect 780 883 893 893
tri 893 883 927 917 sw
tri 14208 883 14242 917 se
rect 14242 883 14356 917
rect 14390 894 14428 917
rect 14462 894 14500 928
rect 14534 894 14572 928
rect 14606 894 14618 928
rect 14390 883 14618 894
rect 39 829 269 863
rect 303 845 329 863
tri 329 845 366 882 sw
rect 517 880 927 883
rect 303 829 366 845
rect 39 820 366 829
tri 366 820 391 845 sw
rect 517 828 518 880
rect 570 828 590 880
rect 642 828 662 880
rect 714 828 734 880
rect 786 845 927 880
tri 927 845 965 883 sw
tri 14170 845 14208 883 se
rect 14208 845 14618 883
rect 14807 4420 14832 4454
rect 14866 4420 15097 4454
rect 14807 4382 15097 4420
rect 14807 4348 14832 4382
rect 14866 4348 15097 4382
rect 14807 4310 15097 4348
rect 14807 4276 14832 4310
rect 14866 4276 15097 4310
rect 14807 4238 15097 4276
rect 14807 4204 14832 4238
rect 14866 4204 15097 4238
rect 14807 4166 15097 4204
rect 14807 4132 14832 4166
rect 14866 4132 15097 4166
rect 14807 4094 15097 4132
rect 14807 4060 14832 4094
rect 14866 4060 15097 4094
rect 14807 4022 15097 4060
rect 14807 3988 14832 4022
rect 14866 3988 15097 4022
rect 14807 3950 15097 3988
rect 14807 3916 14832 3950
rect 14866 3916 15097 3950
rect 14807 3878 15097 3916
rect 14807 3844 14832 3878
rect 14866 3844 15097 3878
rect 14807 3806 15097 3844
rect 14807 3772 14832 3806
rect 14866 3772 15097 3806
rect 14807 3734 15097 3772
rect 14807 3700 14832 3734
rect 14866 3700 15097 3734
rect 14807 3662 15097 3700
rect 14807 3628 14832 3662
rect 14866 3628 15097 3662
rect 14807 3590 15097 3628
rect 14807 3556 14832 3590
rect 14866 3556 15097 3590
rect 14807 3518 15097 3556
rect 14807 3484 14832 3518
rect 14866 3484 15097 3518
rect 14807 3446 15097 3484
rect 14807 3412 14832 3446
rect 14866 3412 15097 3446
rect 14807 3374 15097 3412
rect 14807 3340 14832 3374
rect 14866 3340 15097 3374
rect 14807 3302 15097 3340
rect 14807 3268 14832 3302
rect 14866 3268 15097 3302
rect 14807 3230 15097 3268
rect 14807 3196 14832 3230
rect 14866 3196 15097 3230
rect 14807 3158 15097 3196
rect 14807 3124 14832 3158
rect 14866 3124 15097 3158
rect 14807 3086 15097 3124
rect 14807 3052 14832 3086
rect 14866 3052 15097 3086
rect 14807 3014 15097 3052
rect 14807 2980 14832 3014
rect 14866 2980 15097 3014
rect 14807 2942 15097 2980
rect 14807 2908 14832 2942
rect 14866 2908 15097 2942
rect 14807 2870 15097 2908
rect 14807 2836 14832 2870
rect 14866 2836 15097 2870
rect 14807 2798 15097 2836
rect 14807 2764 14832 2798
rect 14866 2764 15097 2798
rect 14807 2726 15097 2764
rect 14807 2692 14832 2726
rect 14866 2692 15097 2726
rect 14807 2654 15097 2692
rect 14807 2620 14832 2654
rect 14866 2620 15097 2654
rect 14807 2582 15097 2620
rect 14807 2548 14832 2582
rect 14866 2548 15097 2582
rect 14807 2510 15097 2548
rect 14807 2476 14832 2510
rect 14866 2476 15097 2510
rect 14807 2438 15097 2476
rect 14807 2404 14832 2438
rect 14866 2404 15097 2438
rect 14807 2366 15097 2404
rect 14807 2332 14832 2366
rect 14866 2332 15097 2366
rect 14807 2294 15097 2332
rect 14807 2260 14832 2294
rect 14866 2260 15097 2294
rect 14807 2222 15097 2260
rect 14807 2188 14832 2222
rect 14866 2188 15097 2222
rect 14807 2150 15097 2188
rect 14807 2116 14832 2150
rect 14866 2116 15097 2150
rect 14807 2078 15097 2116
rect 14807 2044 14832 2078
rect 14866 2044 15097 2078
rect 14807 2006 15097 2044
rect 14807 1972 14832 2006
rect 14866 1972 15097 2006
rect 14807 1934 15097 1972
rect 14807 1900 14832 1934
rect 14866 1900 15097 1934
rect 14807 1862 15097 1900
rect 14807 1828 14832 1862
rect 14866 1828 15097 1862
rect 14807 1790 15097 1828
rect 14807 1756 14832 1790
rect 14866 1756 15097 1790
rect 14807 1718 15097 1756
rect 14807 1684 14832 1718
rect 14866 1684 15097 1718
rect 14807 1646 15097 1684
rect 14807 1612 14832 1646
rect 14866 1612 15097 1646
rect 14807 1574 15097 1612
rect 14807 1540 14832 1574
rect 14866 1540 15097 1574
rect 14807 1502 15097 1540
rect 14807 1468 14832 1502
rect 14866 1468 15097 1502
rect 14807 1429 15097 1468
rect 14807 1395 14832 1429
rect 14866 1395 15097 1429
rect 14807 1356 15097 1395
rect 14807 1322 14832 1356
rect 14866 1322 15097 1356
rect 14807 1283 15097 1322
rect 14807 1249 14832 1283
rect 14866 1249 15097 1283
rect 14807 1210 15097 1249
rect 14807 1176 14832 1210
rect 14866 1176 15097 1210
rect 14807 1137 15097 1176
rect 14807 1103 14832 1137
rect 14866 1103 15097 1137
rect 14807 1064 15097 1103
rect 14807 1030 14832 1064
rect 14866 1030 15097 1064
rect 14807 991 15097 1030
rect 14807 957 14832 991
rect 14866 957 15097 991
rect 14807 918 15097 957
rect 14807 884 14832 918
rect 14866 884 15097 918
tri 14793 845 14807 859 se
rect 14807 845 15097 884
rect 786 832 965 845
tri 965 832 978 845 sw
tri 14157 832 14170 845 se
rect 14170 832 14618 845
rect 786 828 14618 832
rect 517 820 14618 828
rect 39 789 391 820
rect 39 755 269 789
rect 303 786 391 789
tri 391 786 425 820 sw
rect 517 818 709 820
tri 517 786 549 818 ne
rect 549 786 709 818
rect 743 786 782 820
rect 816 786 855 820
rect 889 786 928 820
rect 303 755 425 786
rect 39 748 425 755
tri 425 748 463 786 sw
tri 549 748 587 786 ne
rect 587 748 928 786
rect 39 715 463 748
rect 39 681 269 715
rect 303 714 463 715
tri 463 714 497 748 sw
tri 587 714 621 748 ne
rect 621 714 709 748
rect 743 714 782 748
rect 816 714 855 748
rect 889 714 928 748
rect 14426 818 14618 820
rect 14426 811 14611 818
tri 14611 811 14618 818 nw
tri 14759 811 14793 845 se
rect 14793 811 14832 845
rect 14866 811 15097 845
rect 14426 772 14572 811
tri 14572 772 14611 811 nw
tri 14720 772 14759 811 se
rect 14759 772 15097 811
rect 14426 738 14538 772
tri 14538 738 14572 772 nw
tri 14686 738 14720 772 se
rect 14720 738 14832 772
rect 14866 738 15097 772
rect 14426 714 14502 738
rect 303 702 497 714
tri 497 702 509 714 sw
tri 621 702 633 714 ne
rect 633 702 14502 714
tri 14502 702 14538 738 nw
tri 14650 702 14686 738 se
rect 14686 702 15097 738
rect 303 699 509 702
tri 509 699 512 702 sw
tri 14647 699 14650 702 se
rect 14650 699 15097 702
rect 303 681 512 699
rect 39 665 512 681
tri 512 665 546 699 sw
tri 14613 665 14647 699 se
rect 14647 665 14832 699
rect 14866 665 15097 699
rect 39 641 546 665
rect 39 607 269 641
rect 303 626 546 641
tri 546 626 585 665 sw
tri 14574 626 14613 665 se
rect 14613 626 15097 665
rect 303 607 585 626
rect 39 592 585 607
tri 585 592 619 626 sw
tri 14540 592 14574 626 se
rect 14574 592 14832 626
rect 14866 592 15097 626
rect 39 567 619 592
rect 39 533 269 567
rect 303 553 619 567
tri 619 553 658 592 sw
tri 14501 553 14540 592 se
rect 14540 553 15097 592
rect 303 533 658 553
rect 39 519 658 533
tri 658 519 692 553 sw
tri 14467 519 14501 553 se
rect 14501 519 14832 553
rect 14866 519 15097 553
rect 39 497 692 519
tri 692 497 714 519 sw
tri 14445 497 14467 519 se
rect 14467 497 15097 519
rect 39 463 343 497
rect 377 463 419 497
rect 453 463 495 497
rect 529 463 571 497
rect 605 463 648 497
rect 682 481 714 497
tri 714 481 730 497 sw
tri 14429 481 14445 497 se
rect 14445 481 15097 497
rect 682 463 730 481
tri 730 463 748 481 sw
tri 14411 463 14429 481 se
rect 14429 463 14465 481
rect 39 447 748 463
tri 748 447 764 463 sw
tri 14395 447 14411 463 se
rect 14411 447 14465 463
rect 14499 447 14539 481
rect 14573 447 14613 481
rect 14647 447 14686 481
rect 14720 447 14759 481
rect 14793 447 15097 481
rect 39 402 764 447
tri 764 402 809 447 sw
tri 14350 402 14395 447 se
rect 14395 402 15097 447
rect 39 375 15097 402
rect 39 341 361 375
rect 395 341 434 375
rect 468 341 507 375
rect 541 341 580 375
rect 614 341 653 375
rect 687 341 726 375
rect 760 341 799 375
rect 833 341 872 375
rect 906 341 945 375
rect 979 341 1018 375
rect 1052 341 1091 375
rect 1125 341 1164 375
rect 1198 341 1237 375
rect 1271 341 1310 375
rect 1344 341 1383 375
rect 1417 341 1456 375
rect 1490 341 1529 375
rect 1563 341 1602 375
rect 1636 341 1675 375
rect 1709 341 1748 375
rect 1782 341 1821 375
rect 1855 341 1894 375
rect 1928 341 1967 375
rect 2001 341 2040 375
rect 2074 341 2113 375
rect 2147 341 2186 375
rect 2220 341 2259 375
rect 2293 341 2332 375
rect 2366 341 2405 375
rect 2439 341 2478 375
rect 2512 341 2551 375
rect 2585 341 2624 375
rect 2658 341 2697 375
rect 2731 341 2770 375
rect 2804 341 2843 375
rect 2877 341 2916 375
rect 2950 341 2989 375
rect 3023 341 3062 375
rect 3096 341 3135 375
rect 3169 341 3208 375
rect 3242 341 3281 375
rect 3315 341 3354 375
rect 3388 341 3427 375
rect 3461 341 3500 375
rect 3534 341 3573 375
rect 3607 341 3646 375
rect 3680 341 3719 375
rect 3753 341 3792 375
rect 3826 341 3865 375
rect 3899 341 3938 375
rect 3972 341 4011 375
rect 4045 341 4084 375
rect 4118 341 4157 375
rect 4191 341 4229 375
rect 4263 341 4301 375
rect 4335 341 4373 375
rect 4407 341 4445 375
rect 4479 341 4517 375
rect 4551 341 4589 375
rect 4623 341 4661 375
rect 4695 341 4733 375
rect 4767 341 4805 375
rect 4839 341 4877 375
rect 4911 341 4949 375
rect 4983 341 5021 375
rect 5055 341 5093 375
rect 5127 341 5165 375
rect 5199 341 5237 375
rect 5271 341 5309 375
rect 5343 341 5381 375
rect 5415 341 5453 375
rect 5487 341 5525 375
rect 5559 341 5597 375
rect 5631 341 5669 375
rect 5703 341 5741 375
rect 5775 341 5813 375
rect 5847 341 5885 375
rect 5919 341 5957 375
rect 5991 341 6029 375
rect 6063 341 6101 375
rect 6135 341 6173 375
rect 6207 341 6245 375
rect 6279 341 6317 375
rect 6351 341 6389 375
rect 6423 341 6461 375
rect 6495 341 6533 375
rect 6567 341 6605 375
rect 6639 341 6677 375
rect 6711 341 6749 375
rect 6783 341 6821 375
rect 6855 341 6893 375
rect 6927 341 6965 375
rect 6999 341 7037 375
rect 7071 341 7109 375
rect 7143 341 7181 375
rect 7215 341 7253 375
rect 7287 341 7325 375
rect 7359 341 7397 375
rect 7431 341 7469 375
rect 7503 341 7541 375
rect 7575 341 7613 375
rect 7647 341 7685 375
rect 7719 341 7757 375
rect 7791 341 7829 375
rect 7863 341 7901 375
rect 7935 341 7973 375
rect 8007 341 8045 375
rect 8079 341 8117 375
rect 8151 341 8189 375
rect 8223 341 8261 375
rect 8295 341 8333 375
rect 8367 341 8405 375
rect 8439 341 8477 375
rect 8511 341 8549 375
rect 8583 341 8621 375
rect 8655 341 8693 375
rect 8727 341 8765 375
rect 8799 341 8837 375
rect 8871 341 8909 375
rect 8943 341 8981 375
rect 9015 341 9053 375
rect 9087 341 9125 375
rect 9159 341 9197 375
rect 9231 341 9269 375
rect 9303 341 9341 375
rect 9375 341 9413 375
rect 9447 341 9485 375
rect 9519 341 9557 375
rect 9591 341 9629 375
rect 9663 341 9701 375
rect 9735 341 9773 375
rect 9807 341 9845 375
rect 9879 341 9917 375
rect 9951 341 9989 375
rect 10023 341 10061 375
rect 10095 341 10133 375
rect 10167 341 10205 375
rect 10239 341 10277 375
rect 10311 341 10349 375
rect 10383 341 10421 375
rect 10455 341 10493 375
rect 10527 341 10565 375
rect 10599 341 10637 375
rect 10671 341 10709 375
rect 10743 341 10781 375
rect 10815 341 10853 375
rect 10887 341 10925 375
rect 10959 341 10997 375
rect 11031 341 11069 375
rect 11103 341 11141 375
rect 11175 341 11213 375
rect 11247 341 11285 375
rect 11319 341 11357 375
rect 11391 341 11429 375
rect 11463 341 11501 375
rect 11535 341 11573 375
rect 11607 341 11645 375
rect 11679 341 11717 375
rect 11751 341 11789 375
rect 11823 341 11861 375
rect 11895 341 11933 375
rect 11967 341 12005 375
rect 12039 341 12077 375
rect 12111 341 12149 375
rect 12183 341 12221 375
rect 12255 341 12293 375
rect 12327 341 12365 375
rect 12399 341 12437 375
rect 12471 341 12509 375
rect 12543 341 12581 375
rect 12615 341 12653 375
rect 12687 341 12725 375
rect 12759 341 12797 375
rect 12831 341 12869 375
rect 12903 341 12941 375
rect 12975 341 13013 375
rect 13047 341 13085 375
rect 13119 341 13157 375
rect 13191 341 13229 375
rect 13263 341 13301 375
rect 13335 341 13373 375
rect 13407 341 13445 375
rect 13479 341 13517 375
rect 13551 341 13589 375
rect 13623 341 13661 375
rect 13695 341 13733 375
rect 13767 341 13805 375
rect 13839 341 13877 375
rect 13911 341 13949 375
rect 13983 341 14021 375
rect 14055 341 14093 375
rect 14127 341 14165 375
rect 14199 341 14237 375
rect 14271 341 14309 375
rect 14343 341 14381 375
rect 14415 341 14453 375
rect 14487 341 14525 375
rect 14559 341 14597 375
rect 14631 341 14669 375
rect 14703 341 14741 375
rect 14775 341 15097 375
rect 39 314 15097 341
<< via1 >>
rect 518 4426 570 4456
rect 518 4404 529 4426
rect 529 4404 563 4426
rect 563 4404 570 4426
rect 590 4426 642 4456
rect 590 4404 601 4426
rect 601 4404 635 4426
rect 635 4404 642 4426
rect 662 4404 674 4456
rect 674 4445 708 4456
rect 708 4445 714 4456
rect 734 4445 786 4456
rect 674 4404 714 4445
rect 734 4404 780 4445
rect 780 4404 786 4445
rect 518 4351 570 4390
rect 518 4338 529 4351
rect 529 4338 563 4351
rect 563 4338 570 4351
rect 590 4351 642 4390
rect 590 4338 601 4351
rect 601 4338 635 4351
rect 635 4338 642 4351
rect 662 4338 674 4390
rect 674 4338 714 4390
rect 734 4338 780 4390
rect 780 4338 786 4390
rect 518 4317 529 4325
rect 529 4317 563 4325
rect 563 4317 570 4325
rect 518 4276 570 4317
rect 518 4273 529 4276
rect 529 4273 563 4276
rect 563 4273 570 4276
rect 590 4317 601 4325
rect 601 4317 635 4325
rect 635 4317 642 4325
rect 590 4276 642 4317
rect 590 4273 601 4276
rect 601 4273 635 4276
rect 635 4273 642 4276
rect 662 4273 674 4325
rect 674 4273 714 4325
rect 734 4273 780 4325
rect 780 4273 786 4325
rect 518 4242 529 4260
rect 529 4242 563 4260
rect 563 4242 570 4260
rect 518 4208 570 4242
rect 590 4242 601 4260
rect 601 4242 635 4260
rect 635 4242 642 4260
rect 590 4208 642 4242
rect 662 4208 674 4260
rect 674 4208 714 4260
rect 734 4208 780 4260
rect 780 4208 786 4260
rect 518 4167 529 4195
rect 529 4167 563 4195
rect 563 4167 570 4195
rect 518 4143 570 4167
rect 590 4167 601 4195
rect 601 4167 635 4195
rect 635 4167 642 4195
rect 590 4143 642 4167
rect 662 4143 674 4195
rect 674 4143 714 4195
rect 734 4143 780 4195
rect 780 4143 786 4195
rect 518 4126 570 4130
rect 518 4092 529 4126
rect 529 4092 563 4126
rect 563 4092 570 4126
rect 518 4078 570 4092
rect 590 4126 642 4130
rect 590 4092 601 4126
rect 601 4092 635 4126
rect 635 4092 642 4126
rect 590 4078 642 4092
rect 662 4078 674 4130
rect 674 4078 714 4130
rect 734 4078 780 4130
rect 780 4078 786 4130
rect 518 4052 570 4065
rect 518 4018 529 4052
rect 529 4018 563 4052
rect 563 4018 570 4052
rect 518 4013 570 4018
rect 590 4052 642 4065
rect 590 4018 601 4052
rect 601 4018 635 4052
rect 635 4018 642 4052
rect 590 4013 642 4018
rect 662 4013 674 4065
rect 674 4013 714 4065
rect 734 4013 780 4065
rect 780 4013 786 4065
rect 518 3978 570 4000
rect 518 3948 529 3978
rect 529 3948 563 3978
rect 563 3948 570 3978
rect 590 3978 642 4000
rect 590 3948 601 3978
rect 601 3948 635 3978
rect 635 3948 642 3978
rect 662 3948 674 4000
rect 674 3948 714 4000
rect 734 3948 780 4000
rect 780 3948 786 4000
rect 518 3904 570 3935
rect 518 3883 529 3904
rect 529 3883 563 3904
rect 563 3883 570 3904
rect 590 3904 642 3935
rect 590 3883 601 3904
rect 601 3883 635 3904
rect 635 3883 642 3904
rect 662 3883 674 3935
rect 674 3883 714 3935
rect 734 3883 780 3935
rect 780 3883 786 3935
rect 518 3818 570 3870
rect 590 3818 642 3870
rect 662 3818 674 3870
rect 674 3818 714 3870
rect 734 3818 780 3870
rect 780 3818 786 3870
rect 518 3794 570 3805
rect 518 3760 529 3794
rect 529 3760 563 3794
rect 563 3760 570 3794
rect 518 3753 570 3760
rect 590 3794 642 3805
rect 590 3760 601 3794
rect 601 3760 635 3794
rect 635 3760 642 3794
rect 590 3753 642 3760
rect 662 3753 674 3805
rect 674 3753 714 3805
rect 734 3753 780 3805
rect 780 3753 786 3805
rect 518 3720 570 3740
rect 518 3688 529 3720
rect 529 3688 563 3720
rect 563 3688 570 3720
rect 590 3720 642 3740
rect 590 3688 601 3720
rect 601 3688 635 3720
rect 635 3688 642 3720
rect 662 3688 674 3740
rect 674 3688 714 3740
rect 734 3688 780 3740
rect 780 3688 786 3740
rect 518 3646 570 3675
rect 518 3623 529 3646
rect 529 3623 563 3646
rect 563 3623 570 3646
rect 590 3646 642 3675
rect 590 3623 601 3646
rect 601 3623 635 3646
rect 635 3623 642 3646
rect 662 3623 674 3675
rect 674 3623 714 3675
rect 734 3623 780 3675
rect 780 3623 786 3675
rect 518 3572 570 3610
rect 518 3558 529 3572
rect 529 3558 563 3572
rect 563 3558 570 3572
rect 590 3572 642 3610
rect 590 3558 601 3572
rect 601 3558 635 3572
rect 635 3558 642 3572
rect 662 3558 674 3610
rect 674 3558 714 3610
rect 734 3558 780 3610
rect 780 3558 786 3610
rect 518 3538 529 3545
rect 529 3538 563 3545
rect 563 3538 570 3545
rect 518 3498 570 3538
rect 518 3493 529 3498
rect 529 3493 563 3498
rect 563 3493 570 3498
rect 590 3538 601 3545
rect 601 3538 635 3545
rect 635 3538 642 3545
rect 590 3498 642 3538
rect 590 3493 601 3498
rect 601 3493 635 3498
rect 635 3493 642 3498
rect 662 3493 674 3545
rect 674 3493 714 3545
rect 734 3493 780 3545
rect 780 3493 786 3545
rect 518 3464 529 3480
rect 529 3464 563 3480
rect 563 3464 570 3480
rect 518 3428 570 3464
rect 590 3464 601 3480
rect 601 3464 635 3480
rect 635 3464 642 3480
rect 590 3428 642 3464
rect 662 3428 674 3480
rect 674 3428 714 3480
rect 734 3428 780 3480
rect 780 3428 786 3480
rect 518 3390 529 3415
rect 529 3390 563 3415
rect 563 3390 570 3415
rect 518 3363 570 3390
rect 590 3390 601 3415
rect 601 3390 635 3415
rect 635 3390 642 3415
rect 590 3363 642 3390
rect 662 3363 674 3415
rect 674 3363 714 3415
rect 734 3363 780 3415
rect 780 3363 786 3415
rect 518 3316 529 3350
rect 529 3316 563 3350
rect 563 3316 570 3350
rect 518 3298 570 3316
rect 590 3316 601 3350
rect 601 3316 635 3350
rect 635 3316 642 3350
rect 590 3298 642 3316
rect 662 3298 674 3350
rect 674 3298 714 3350
rect 734 3298 780 3350
rect 780 3298 786 3350
rect 518 3276 570 3285
rect 518 3242 529 3276
rect 529 3242 563 3276
rect 563 3242 570 3276
rect 518 3233 570 3242
rect 590 3276 642 3285
rect 590 3242 601 3276
rect 601 3242 635 3276
rect 635 3242 642 3276
rect 590 3233 642 3242
rect 662 3233 674 3285
rect 674 3233 714 3285
rect 734 3233 780 3285
rect 780 3233 786 3285
rect 518 3202 570 3220
rect 518 3168 529 3202
rect 529 3168 563 3202
rect 563 3168 570 3202
rect 590 3202 642 3220
rect 590 3168 601 3202
rect 601 3168 635 3202
rect 635 3168 642 3202
rect 662 3168 674 3220
rect 674 3168 714 3220
rect 734 3168 780 3220
rect 780 3168 786 3220
rect 518 3128 570 3155
rect 518 3103 529 3128
rect 529 3103 563 3128
rect 563 3103 570 3128
rect 590 3128 642 3155
rect 590 3103 601 3128
rect 601 3103 635 3128
rect 635 3103 642 3128
rect 662 3103 674 3155
rect 674 3103 714 3155
rect 734 3103 780 3155
rect 780 3103 786 3155
rect 518 3054 570 3090
rect 518 3038 529 3054
rect 529 3038 563 3054
rect 563 3038 570 3054
rect 590 3054 642 3090
rect 590 3038 601 3054
rect 601 3038 635 3054
rect 635 3038 642 3054
rect 662 3038 674 3090
rect 674 3038 714 3090
rect 734 3038 780 3090
rect 780 3038 786 3090
rect 518 3020 529 3025
rect 529 3020 563 3025
rect 563 3020 570 3025
rect 518 2980 570 3020
rect 518 2973 529 2980
rect 529 2973 563 2980
rect 563 2973 570 2980
rect 590 3020 601 3025
rect 601 3020 635 3025
rect 635 3020 642 3025
rect 590 2980 642 3020
rect 590 2973 601 2980
rect 601 2973 635 2980
rect 635 2973 642 2980
rect 662 2973 674 3025
rect 674 2973 714 3025
rect 734 2973 780 3025
rect 780 2973 786 3025
rect 518 2946 529 2960
rect 529 2946 563 2960
rect 563 2946 570 2960
rect 518 2908 570 2946
rect 590 2946 601 2960
rect 601 2946 635 2960
rect 635 2946 642 2960
rect 590 2908 642 2946
rect 662 2908 674 2960
rect 674 2908 714 2960
rect 734 2908 780 2960
rect 780 2908 786 2960
rect 518 2872 529 2895
rect 529 2872 563 2895
rect 563 2872 570 2895
rect 518 2843 570 2872
rect 590 2872 601 2895
rect 601 2872 635 2895
rect 635 2872 642 2895
rect 590 2843 642 2872
rect 662 2843 674 2895
rect 674 2843 714 2895
rect 734 2843 780 2895
rect 780 2843 786 2895
rect 518 2798 529 2830
rect 529 2798 563 2830
rect 563 2798 570 2830
rect 518 2778 570 2798
rect 590 2798 601 2830
rect 601 2798 635 2830
rect 635 2798 642 2830
rect 590 2778 642 2798
rect 662 2778 674 2830
rect 674 2778 714 2830
rect 734 2778 780 2830
rect 780 2778 786 2830
rect 518 2758 570 2765
rect 518 2724 529 2758
rect 529 2724 563 2758
rect 563 2724 570 2758
rect 518 2713 570 2724
rect 590 2758 642 2765
rect 590 2724 601 2758
rect 601 2724 635 2758
rect 635 2724 642 2758
rect 590 2713 642 2724
rect 662 2713 674 2765
rect 674 2713 714 2765
rect 734 2713 780 2765
rect 780 2713 786 2765
rect 518 2684 570 2700
rect 518 2650 529 2684
rect 529 2650 563 2684
rect 563 2650 570 2684
rect 518 2648 570 2650
rect 590 2684 642 2700
rect 590 2650 601 2684
rect 601 2650 635 2684
rect 635 2650 642 2684
rect 590 2648 642 2650
rect 662 2648 674 2700
rect 674 2648 714 2700
rect 734 2648 780 2700
rect 780 2648 786 2700
rect 518 2610 570 2635
rect 518 2583 529 2610
rect 529 2583 563 2610
rect 563 2583 570 2610
rect 590 2610 642 2635
rect 590 2583 601 2610
rect 601 2583 635 2610
rect 635 2583 642 2610
rect 662 2583 674 2635
rect 674 2583 714 2635
rect 734 2583 780 2635
rect 780 2583 786 2635
rect 518 2536 570 2570
rect 518 2518 529 2536
rect 529 2518 563 2536
rect 563 2518 570 2536
rect 590 2536 642 2570
rect 590 2518 601 2536
rect 601 2518 635 2536
rect 635 2518 642 2536
rect 662 2518 674 2570
rect 674 2518 714 2570
rect 734 2518 780 2570
rect 780 2518 786 2570
rect 518 2502 529 2505
rect 529 2502 563 2505
rect 563 2502 570 2505
rect 518 2462 570 2502
rect 518 2453 529 2462
rect 529 2453 563 2462
rect 563 2453 570 2462
rect 590 2502 601 2505
rect 601 2502 635 2505
rect 635 2502 642 2505
rect 590 2462 642 2502
rect 590 2453 601 2462
rect 601 2453 635 2462
rect 635 2453 642 2462
rect 662 2453 674 2505
rect 674 2453 714 2505
rect 734 2453 780 2505
rect 780 2453 786 2505
rect 518 2428 529 2440
rect 529 2428 563 2440
rect 563 2428 570 2440
rect 518 2389 570 2428
rect 518 2388 529 2389
rect 529 2388 563 2389
rect 563 2388 570 2389
rect 590 2428 601 2440
rect 601 2428 635 2440
rect 635 2428 642 2440
rect 590 2389 642 2428
rect 590 2388 601 2389
rect 601 2388 635 2389
rect 635 2388 642 2389
rect 662 2388 674 2440
rect 674 2388 714 2440
rect 734 2388 780 2440
rect 780 2388 786 2440
rect 518 2355 529 2375
rect 529 2355 563 2375
rect 563 2355 570 2375
rect 518 2323 570 2355
rect 590 2355 601 2375
rect 601 2355 635 2375
rect 635 2355 642 2375
rect 590 2323 642 2355
rect 662 2323 674 2375
rect 674 2323 714 2375
rect 734 2323 780 2375
rect 780 2323 786 2375
rect 518 2282 529 2310
rect 529 2282 563 2310
rect 563 2282 570 2310
rect 518 2258 570 2282
rect 590 2282 601 2310
rect 601 2282 635 2310
rect 635 2282 642 2310
rect 590 2258 642 2282
rect 662 2258 674 2310
rect 674 2258 714 2310
rect 734 2258 780 2310
rect 780 2258 786 2310
rect 518 2243 570 2245
rect 518 2209 529 2243
rect 529 2209 563 2243
rect 563 2209 570 2243
rect 518 2193 570 2209
rect 590 2243 642 2245
rect 590 2209 601 2243
rect 601 2209 635 2243
rect 635 2209 642 2243
rect 590 2193 642 2209
rect 662 2193 674 2245
rect 674 2193 714 2245
rect 734 2193 780 2245
rect 780 2193 786 2245
rect 518 2170 570 2180
rect 518 2136 529 2170
rect 529 2136 563 2170
rect 563 2136 570 2170
rect 518 2128 570 2136
rect 590 2170 642 2180
rect 590 2136 601 2170
rect 601 2136 635 2170
rect 635 2136 642 2170
rect 590 2128 642 2136
rect 662 2128 674 2180
rect 674 2128 714 2180
rect 734 2128 780 2180
rect 780 2128 786 2180
rect 518 2097 570 2115
rect 518 2063 529 2097
rect 529 2063 563 2097
rect 563 2063 570 2097
rect 590 2097 642 2115
rect 590 2063 601 2097
rect 601 2063 635 2097
rect 635 2063 642 2097
rect 662 2063 674 2115
rect 674 2063 714 2115
rect 734 2063 780 2115
rect 780 2063 786 2115
rect 518 2024 570 2050
rect 518 1998 529 2024
rect 529 1998 563 2024
rect 563 1998 570 2024
rect 590 2024 642 2050
rect 590 1998 601 2024
rect 601 1998 635 2024
rect 635 1998 642 2024
rect 662 1998 674 2050
rect 674 1998 714 2050
rect 734 1998 780 2050
rect 780 1998 786 2050
rect 518 1951 570 1985
rect 518 1933 529 1951
rect 529 1933 563 1951
rect 563 1933 570 1951
rect 590 1951 642 1985
rect 590 1933 601 1951
rect 601 1933 635 1951
rect 635 1933 642 1951
rect 662 1933 674 1985
rect 674 1933 714 1985
rect 734 1933 780 1985
rect 780 1933 786 1985
rect 518 1917 529 1920
rect 529 1917 563 1920
rect 563 1917 570 1920
rect 518 1878 570 1917
rect 518 1868 529 1878
rect 529 1868 563 1878
rect 563 1868 570 1878
rect 590 1917 601 1920
rect 601 1917 635 1920
rect 635 1917 642 1920
rect 590 1878 642 1917
rect 590 1868 601 1878
rect 601 1868 635 1878
rect 635 1868 642 1878
rect 662 1868 674 1920
rect 674 1868 714 1920
rect 734 1868 780 1920
rect 780 1868 786 1920
rect 518 1844 529 1855
rect 529 1844 563 1855
rect 563 1844 570 1855
rect 518 1805 570 1844
rect 518 1803 529 1805
rect 529 1803 563 1805
rect 563 1803 570 1805
rect 590 1844 601 1855
rect 601 1844 635 1855
rect 635 1844 642 1855
rect 590 1805 642 1844
rect 590 1803 601 1805
rect 601 1803 635 1805
rect 635 1803 642 1805
rect 662 1803 674 1855
rect 674 1803 714 1855
rect 734 1803 780 1855
rect 780 1803 786 1855
rect 518 1771 529 1790
rect 529 1771 563 1790
rect 563 1771 570 1790
rect 518 1738 570 1771
rect 590 1771 601 1790
rect 601 1771 635 1790
rect 635 1771 642 1790
rect 590 1738 642 1771
rect 662 1738 674 1790
rect 674 1738 714 1790
rect 734 1738 780 1790
rect 780 1738 786 1790
rect 518 1698 529 1725
rect 529 1698 563 1725
rect 563 1698 570 1725
rect 518 1673 570 1698
rect 590 1698 601 1725
rect 601 1698 635 1725
rect 635 1698 642 1725
rect 590 1673 642 1698
rect 662 1673 674 1725
rect 674 1673 714 1725
rect 734 1673 780 1725
rect 780 1673 786 1725
rect 518 1659 570 1660
rect 518 1625 529 1659
rect 529 1625 563 1659
rect 563 1625 570 1659
rect 518 1608 570 1625
rect 590 1659 642 1660
rect 590 1625 601 1659
rect 601 1625 635 1659
rect 635 1625 642 1659
rect 590 1608 642 1625
rect 662 1608 674 1660
rect 674 1608 714 1660
rect 734 1608 780 1660
rect 780 1608 786 1660
rect 518 1586 570 1595
rect 518 1552 529 1586
rect 529 1552 563 1586
rect 563 1552 570 1586
rect 518 1543 570 1552
rect 590 1586 642 1595
rect 590 1552 601 1586
rect 601 1552 635 1586
rect 635 1552 642 1586
rect 590 1543 642 1552
rect 662 1543 674 1595
rect 674 1543 714 1595
rect 734 1543 780 1595
rect 780 1543 786 1595
rect 1066 4098 1118 4119
rect 1066 4067 1067 4098
rect 1067 4067 1101 4098
rect 1101 4067 1118 4098
rect 1130 4098 1182 4119
rect 1130 4067 1139 4098
rect 1139 4067 1173 4098
rect 1173 4067 1182 4098
rect 1194 4098 1246 4119
rect 1194 4067 1211 4098
rect 1211 4067 1245 4098
rect 1245 4067 1246 4098
rect 1066 4025 1118 4054
rect 1066 4002 1067 4025
rect 1067 4002 1101 4025
rect 1101 4002 1118 4025
rect 1130 4025 1182 4054
rect 1130 4002 1139 4025
rect 1139 4002 1173 4025
rect 1173 4002 1182 4025
rect 1194 4025 1246 4054
rect 1194 4002 1211 4025
rect 1211 4002 1245 4025
rect 1245 4002 1246 4025
rect 1066 3952 1118 3989
rect 1066 3937 1067 3952
rect 1067 3937 1101 3952
rect 1101 3937 1118 3952
rect 1130 3952 1182 3989
rect 1130 3937 1139 3952
rect 1139 3937 1173 3952
rect 1173 3937 1182 3952
rect 1194 3952 1246 3989
rect 1194 3937 1211 3952
rect 1211 3937 1245 3952
rect 1245 3937 1246 3952
rect 1066 3918 1067 3924
rect 1067 3918 1101 3924
rect 1101 3918 1139 3924
rect 1139 3918 1173 3924
rect 1173 3918 1211 3924
rect 1211 3918 1245 3924
rect 1245 3918 1246 3924
rect 1066 3879 1246 3918
rect 1066 3845 1067 3879
rect 1067 3845 1101 3879
rect 1101 3845 1139 3879
rect 1139 3845 1173 3879
rect 1173 3845 1211 3879
rect 1211 3845 1245 3879
rect 1245 3845 1246 3879
rect 1066 3806 1246 3845
rect 1066 3772 1067 3806
rect 1067 3772 1101 3806
rect 1101 3772 1139 3806
rect 1139 3772 1173 3806
rect 1173 3772 1211 3806
rect 1211 3772 1245 3806
rect 1245 3772 1246 3806
rect 1066 3733 1246 3772
rect 1066 3699 1067 3733
rect 1067 3699 1101 3733
rect 1101 3699 1139 3733
rect 1139 3699 1173 3733
rect 1173 3699 1211 3733
rect 1211 3699 1245 3733
rect 1245 3699 1246 3733
rect 1066 3660 1246 3699
rect 1066 3626 1067 3660
rect 1067 3626 1101 3660
rect 1101 3626 1139 3660
rect 1139 3626 1173 3660
rect 1173 3626 1211 3660
rect 1211 3626 1245 3660
rect 1245 3626 1246 3660
rect 1066 3587 1246 3626
rect 1066 3553 1067 3587
rect 1067 3553 1101 3587
rect 1101 3553 1139 3587
rect 1139 3553 1173 3587
rect 1173 3553 1211 3587
rect 1211 3553 1245 3587
rect 1245 3553 1246 3587
rect 1066 3514 1246 3553
rect 1066 3480 1067 3514
rect 1067 3480 1101 3514
rect 1101 3480 1139 3514
rect 1139 3480 1173 3514
rect 1173 3480 1211 3514
rect 1211 3480 1245 3514
rect 1245 3480 1246 3514
rect 1066 3441 1246 3480
rect 1066 3407 1067 3441
rect 1067 3407 1101 3441
rect 1101 3407 1139 3441
rect 1139 3407 1173 3441
rect 1173 3407 1211 3441
rect 1211 3407 1245 3441
rect 1245 3407 1246 3441
rect 1066 3368 1246 3407
rect 1066 3334 1067 3368
rect 1067 3334 1101 3368
rect 1101 3334 1139 3368
rect 1139 3334 1173 3368
rect 1173 3334 1211 3368
rect 1211 3334 1245 3368
rect 1245 3334 1246 3368
rect 1066 3295 1246 3334
rect 1066 3261 1067 3295
rect 1067 3261 1101 3295
rect 1101 3261 1139 3295
rect 1139 3261 1173 3295
rect 1173 3261 1211 3295
rect 1211 3261 1245 3295
rect 1245 3261 1246 3295
rect 1066 3222 1246 3261
rect 1066 3188 1067 3222
rect 1067 3188 1101 3222
rect 1101 3188 1139 3222
rect 1139 3188 1173 3222
rect 1173 3188 1211 3222
rect 1211 3188 1245 3222
rect 1245 3188 1246 3222
rect 1066 3149 1246 3188
rect 1066 3115 1067 3149
rect 1067 3115 1101 3149
rect 1101 3115 1139 3149
rect 1139 3115 1173 3149
rect 1173 3115 1211 3149
rect 1211 3115 1245 3149
rect 1245 3115 1246 3149
rect 1066 3076 1246 3115
rect 1066 3042 1067 3076
rect 1067 3042 1101 3076
rect 1101 3042 1139 3076
rect 1139 3042 1173 3076
rect 1173 3042 1211 3076
rect 1211 3042 1245 3076
rect 1245 3042 1246 3076
rect 1066 3003 1246 3042
rect 1066 2969 1067 3003
rect 1067 2969 1101 3003
rect 1101 2969 1139 3003
rect 1139 2969 1173 3003
rect 1173 2969 1211 3003
rect 1211 2969 1245 3003
rect 1245 2969 1246 3003
rect 1066 2930 1246 2969
rect 1066 2896 1067 2930
rect 1067 2896 1101 2930
rect 1101 2896 1139 2930
rect 1139 2896 1173 2930
rect 1173 2896 1211 2930
rect 1211 2896 1245 2930
rect 1245 2896 1246 2930
rect 1066 2857 1246 2896
rect 1066 2823 1067 2857
rect 1067 2823 1101 2857
rect 1101 2823 1139 2857
rect 1139 2823 1173 2857
rect 1173 2823 1211 2857
rect 1211 2823 1245 2857
rect 1245 2823 1246 2857
rect 1066 2784 1246 2823
rect 1066 2750 1067 2784
rect 1067 2750 1101 2784
rect 1101 2750 1139 2784
rect 1139 2750 1173 2784
rect 1173 2750 1211 2784
rect 1211 2750 1245 2784
rect 1245 2750 1246 2784
rect 1066 2711 1246 2750
rect 1066 2677 1067 2711
rect 1067 2677 1101 2711
rect 1101 2677 1139 2711
rect 1139 2677 1173 2711
rect 1173 2677 1211 2711
rect 1211 2677 1245 2711
rect 1245 2677 1246 2711
rect 1066 2638 1246 2677
rect 1066 2604 1067 2638
rect 1067 2604 1101 2638
rect 1101 2604 1139 2638
rect 1139 2604 1173 2638
rect 1173 2604 1211 2638
rect 1211 2604 1245 2638
rect 1245 2604 1246 2638
rect 1066 2565 1246 2604
rect 1066 2531 1067 2565
rect 1067 2531 1101 2565
rect 1101 2531 1139 2565
rect 1139 2531 1173 2565
rect 1173 2531 1211 2565
rect 1211 2531 1245 2565
rect 1245 2531 1246 2565
rect 1066 2492 1246 2531
rect 1066 2458 1067 2492
rect 1067 2458 1101 2492
rect 1101 2458 1139 2492
rect 1139 2458 1173 2492
rect 1173 2458 1211 2492
rect 1211 2458 1245 2492
rect 1245 2458 1246 2492
rect 1066 2419 1246 2458
rect 1066 2385 1067 2419
rect 1067 2385 1101 2419
rect 1101 2385 1139 2419
rect 1139 2385 1173 2419
rect 1173 2385 1211 2419
rect 1211 2385 1245 2419
rect 1245 2385 1246 2419
rect 1066 2346 1246 2385
rect 1066 2312 1067 2346
rect 1067 2312 1101 2346
rect 1101 2312 1139 2346
rect 1139 2312 1173 2346
rect 1173 2312 1211 2346
rect 1211 2312 1245 2346
rect 1245 2312 1246 2346
rect 1066 2273 1246 2312
rect 1066 2239 1067 2273
rect 1067 2239 1101 2273
rect 1101 2239 1139 2273
rect 1139 2239 1173 2273
rect 1173 2239 1211 2273
rect 1211 2239 1245 2273
rect 1245 2239 1246 2273
rect 1066 2200 1246 2239
rect 1066 2166 1067 2200
rect 1067 2166 1101 2200
rect 1101 2166 1139 2200
rect 1139 2166 1173 2200
rect 1173 2166 1211 2200
rect 1211 2166 1245 2200
rect 1245 2166 1246 2200
rect 1066 2126 1246 2166
rect 1066 2092 1067 2126
rect 1067 2092 1101 2126
rect 1101 2092 1139 2126
rect 1139 2092 1173 2126
rect 1173 2092 1211 2126
rect 1211 2092 1245 2126
rect 1245 2092 1246 2126
rect 1066 2052 1246 2092
rect 1066 2018 1067 2052
rect 1067 2018 1101 2052
rect 1101 2018 1139 2052
rect 1139 2018 1173 2052
rect 1173 2018 1211 2052
rect 1211 2018 1245 2052
rect 1245 2018 1246 2052
rect 1066 1978 1246 2018
rect 1066 1944 1067 1978
rect 1067 1944 1101 1978
rect 1101 1944 1139 1978
rect 1139 1944 1173 1978
rect 1173 1944 1211 1978
rect 1211 1944 1245 1978
rect 1245 1944 1246 1978
rect 1066 1904 1246 1944
rect 1066 1870 1067 1904
rect 1067 1870 1101 1904
rect 1101 1870 1139 1904
rect 1139 1870 1173 1904
rect 1173 1870 1211 1904
rect 1211 1870 1245 1904
rect 1245 1870 1246 1904
rect 1066 1830 1246 1870
rect 1066 1796 1067 1830
rect 1067 1796 1101 1830
rect 1101 1796 1139 1830
rect 1139 1796 1173 1830
rect 1173 1796 1211 1830
rect 1211 1796 1245 1830
rect 1245 1796 1246 1830
rect 1066 1756 1246 1796
rect 1066 1722 1067 1756
rect 1067 1722 1101 1756
rect 1101 1722 1139 1756
rect 1139 1722 1173 1756
rect 1173 1722 1211 1756
rect 1211 1722 1245 1756
rect 1245 1722 1246 1756
rect 1066 1682 1246 1722
rect 1066 1648 1067 1682
rect 1067 1648 1101 1682
rect 1101 1648 1139 1682
rect 1139 1648 1173 1682
rect 1173 1648 1211 1682
rect 1211 1648 1245 1682
rect 1245 1648 1246 1682
rect 1066 1608 1246 1648
rect 1066 1574 1067 1608
rect 1067 1574 1101 1608
rect 1101 1574 1139 1608
rect 1139 1574 1173 1608
rect 1173 1574 1211 1608
rect 1211 1574 1245 1608
rect 1245 1574 1246 1608
rect 1066 1568 1246 1574
rect 1562 4092 1614 4124
rect 1562 4072 1563 4092
rect 1563 4072 1597 4092
rect 1597 4072 1614 4092
rect 1626 4072 1678 4124
rect 1690 4092 1742 4124
rect 1690 4072 1707 4092
rect 1707 4072 1741 4092
rect 1741 4072 1742 4092
rect 1562 4058 1563 4059
rect 1563 4058 1597 4059
rect 1597 4058 1614 4059
rect 1562 4020 1614 4058
rect 1562 4007 1563 4020
rect 1563 4007 1597 4020
rect 1597 4007 1614 4020
rect 1626 4007 1678 4059
rect 1690 4058 1707 4059
rect 1707 4058 1741 4059
rect 1741 4058 1742 4059
rect 1690 4020 1742 4058
rect 1690 4007 1707 4020
rect 1707 4007 1741 4020
rect 1741 4007 1742 4020
rect 1562 3986 1563 3994
rect 1563 3986 1597 3994
rect 1597 3986 1614 3994
rect 1562 3948 1614 3986
rect 1562 3942 1563 3948
rect 1563 3942 1597 3948
rect 1597 3942 1614 3948
rect 1626 3942 1678 3994
rect 1690 3986 1707 3994
rect 1707 3986 1741 3994
rect 1741 3986 1742 3994
rect 1690 3948 1742 3986
rect 1690 3942 1707 3948
rect 1707 3942 1741 3948
rect 1741 3942 1742 3948
rect 1562 3914 1563 3929
rect 1563 3914 1597 3929
rect 1597 3914 1614 3929
rect 1562 3877 1614 3914
rect 1626 3877 1678 3929
rect 1690 3914 1707 3929
rect 1707 3914 1741 3929
rect 1741 3914 1742 3929
rect 1690 3877 1742 3914
rect 1562 3842 1563 3864
rect 1563 3842 1597 3864
rect 1597 3842 1614 3864
rect 1562 3812 1614 3842
rect 1626 3812 1678 3864
rect 1690 3842 1707 3864
rect 1707 3842 1741 3864
rect 1741 3842 1742 3864
rect 1690 3812 1742 3842
rect 1562 3770 1563 3799
rect 1563 3770 1597 3799
rect 1597 3770 1614 3799
rect 1562 3747 1614 3770
rect 1626 3747 1678 3799
rect 1690 3770 1707 3799
rect 1707 3770 1741 3799
rect 1741 3770 1742 3799
rect 1690 3747 1742 3770
rect 1562 3732 1614 3734
rect 1562 3698 1563 3732
rect 1563 3698 1597 3732
rect 1597 3698 1614 3732
rect 1562 3682 1614 3698
rect 1626 3682 1678 3734
rect 1690 3732 1742 3734
rect 1690 3698 1707 3732
rect 1707 3698 1741 3732
rect 1741 3698 1742 3732
rect 1690 3682 1742 3698
rect 1562 3660 1614 3669
rect 1562 3626 1563 3660
rect 1563 3626 1597 3660
rect 1597 3626 1614 3660
rect 1562 3617 1614 3626
rect 1626 3617 1678 3669
rect 1690 3660 1742 3669
rect 1690 3626 1707 3660
rect 1707 3626 1741 3660
rect 1741 3626 1742 3660
rect 1690 3617 1742 3626
rect 1562 3588 1742 3604
rect 1562 3554 1563 3588
rect 1563 3554 1597 3588
rect 1597 3554 1707 3588
rect 1707 3554 1741 3588
rect 1741 3554 1742 3588
rect 1562 3516 1742 3554
rect 1562 3482 1563 3516
rect 1563 3482 1597 3516
rect 1597 3482 1707 3516
rect 1707 3482 1741 3516
rect 1741 3482 1742 3516
rect 1562 3444 1742 3482
rect 1562 3410 1563 3444
rect 1563 3410 1597 3444
rect 1597 3410 1707 3444
rect 1707 3410 1741 3444
rect 1741 3410 1742 3444
rect 1562 3372 1742 3410
rect 1562 3338 1563 3372
rect 1563 3338 1597 3372
rect 1597 3338 1707 3372
rect 1707 3338 1741 3372
rect 1741 3338 1742 3372
rect 1562 3300 1742 3338
rect 1562 3266 1563 3300
rect 1563 3266 1597 3300
rect 1597 3266 1707 3300
rect 1707 3266 1741 3300
rect 1741 3266 1742 3300
rect 1562 3228 1742 3266
rect 1562 3194 1563 3228
rect 1563 3194 1597 3228
rect 1597 3194 1707 3228
rect 1707 3194 1741 3228
rect 1741 3194 1742 3228
rect 1562 3108 1742 3194
rect 1562 3074 1563 3108
rect 1563 3074 1597 3108
rect 1597 3074 1635 3108
rect 1635 3074 1669 3108
rect 1669 3074 1707 3108
rect 1707 3074 1741 3108
rect 1741 3074 1742 3108
rect 1562 3028 1742 3074
rect 1562 2994 1563 3028
rect 1563 2994 1597 3028
rect 1597 2994 1635 3028
rect 1635 2994 1669 3028
rect 1669 2994 1707 3028
rect 1707 2994 1741 3028
rect 1741 2994 1742 3028
rect 1562 2948 1742 2994
rect 1562 2914 1563 2948
rect 1563 2914 1597 2948
rect 1597 2914 1635 2948
rect 1635 2914 1669 2948
rect 1669 2914 1707 2948
rect 1707 2914 1741 2948
rect 1741 2914 1742 2948
rect 1562 2868 1742 2914
rect 1562 2834 1563 2868
rect 1563 2834 1597 2868
rect 1597 2834 1635 2868
rect 1635 2834 1669 2868
rect 1669 2834 1707 2868
rect 1707 2834 1741 2868
rect 1741 2834 1742 2868
rect 1562 2788 1742 2834
rect 1562 2754 1563 2788
rect 1563 2754 1597 2788
rect 1597 2754 1635 2788
rect 1635 2754 1669 2788
rect 1669 2754 1707 2788
rect 1707 2754 1741 2788
rect 1741 2754 1742 2788
rect 1562 2708 1742 2754
rect 1562 2674 1563 2708
rect 1563 2674 1597 2708
rect 1597 2674 1635 2708
rect 1635 2674 1669 2708
rect 1669 2674 1707 2708
rect 1707 2674 1741 2708
rect 1741 2674 1742 2708
rect 1562 2628 1742 2674
rect 1562 2594 1563 2628
rect 1563 2594 1597 2628
rect 1597 2594 1635 2628
rect 1635 2594 1669 2628
rect 1669 2594 1707 2628
rect 1707 2594 1741 2628
rect 1741 2594 1742 2628
rect 1562 2518 1742 2594
rect 1562 2484 1563 2518
rect 1563 2484 1597 2518
rect 1597 2484 1707 2518
rect 1707 2484 1741 2518
rect 1741 2484 1742 2518
rect 1562 2446 1742 2484
rect 1562 2412 1563 2446
rect 1563 2412 1597 2446
rect 1597 2412 1707 2446
rect 1707 2412 1741 2446
rect 1741 2412 1742 2446
rect 1562 2374 1742 2412
rect 1562 2340 1563 2374
rect 1563 2340 1597 2374
rect 1597 2340 1707 2374
rect 1707 2340 1741 2374
rect 1741 2340 1742 2374
rect 1562 2302 1742 2340
rect 1562 2268 1563 2302
rect 1563 2268 1597 2302
rect 1597 2268 1707 2302
rect 1707 2268 1741 2302
rect 1741 2268 1742 2302
rect 1562 2230 1742 2268
rect 1562 2196 1563 2230
rect 1563 2196 1597 2230
rect 1597 2196 1707 2230
rect 1707 2196 1741 2230
rect 1741 2196 1742 2230
rect 1562 2158 1742 2196
rect 1562 2124 1563 2158
rect 1563 2124 1597 2158
rect 1597 2124 1707 2158
rect 1707 2124 1741 2158
rect 1741 2124 1742 2158
rect 1562 2086 1742 2124
rect 1562 2052 1563 2086
rect 1563 2052 1597 2086
rect 1597 2052 1707 2086
rect 1707 2052 1741 2086
rect 1741 2052 1742 2086
rect 1562 2014 1742 2052
rect 1562 1980 1563 2014
rect 1563 1980 1597 2014
rect 1597 1980 1707 2014
rect 1707 1980 1741 2014
rect 1741 1980 1742 2014
rect 1562 1942 1742 1980
rect 1562 1908 1563 1942
rect 1563 1908 1597 1942
rect 1597 1908 1707 1942
rect 1707 1908 1741 1942
rect 1741 1908 1742 1942
rect 1562 1870 1742 1908
rect 1562 1836 1563 1870
rect 1563 1836 1597 1870
rect 1597 1836 1707 1870
rect 1707 1836 1741 1870
rect 1741 1836 1742 1870
rect 1562 1798 1742 1836
rect 1562 1764 1563 1798
rect 1563 1764 1597 1798
rect 1597 1764 1707 1798
rect 1707 1764 1741 1798
rect 1741 1764 1742 1798
rect 1562 1726 1742 1764
rect 1562 1692 1563 1726
rect 1563 1692 1597 1726
rect 1597 1692 1707 1726
rect 1707 1692 1741 1726
rect 1741 1692 1742 1726
rect 1562 1654 1742 1692
rect 1562 1620 1563 1654
rect 1563 1620 1597 1654
rect 1597 1620 1707 1654
rect 1707 1620 1741 1654
rect 1741 1620 1742 1654
rect 1562 1568 1742 1620
rect 2058 4098 2110 4119
rect 2058 4067 2059 4098
rect 2059 4067 2093 4098
rect 2093 4067 2110 4098
rect 2122 4098 2174 4119
rect 2122 4067 2131 4098
rect 2131 4067 2165 4098
rect 2165 4067 2174 4098
rect 2186 4098 2238 4119
rect 2186 4067 2203 4098
rect 2203 4067 2237 4098
rect 2237 4067 2238 4098
rect 2058 4025 2110 4054
rect 2058 4002 2059 4025
rect 2059 4002 2093 4025
rect 2093 4002 2110 4025
rect 2122 4025 2174 4054
rect 2122 4002 2131 4025
rect 2131 4002 2165 4025
rect 2165 4002 2174 4025
rect 2186 4025 2238 4054
rect 2186 4002 2203 4025
rect 2203 4002 2237 4025
rect 2237 4002 2238 4025
rect 2058 3952 2110 3989
rect 2058 3937 2059 3952
rect 2059 3937 2093 3952
rect 2093 3937 2110 3952
rect 2122 3952 2174 3989
rect 2122 3937 2131 3952
rect 2131 3937 2165 3952
rect 2165 3937 2174 3952
rect 2186 3952 2238 3989
rect 2186 3937 2203 3952
rect 2203 3937 2237 3952
rect 2237 3937 2238 3952
rect 2058 3918 2059 3924
rect 2059 3918 2093 3924
rect 2093 3918 2131 3924
rect 2131 3918 2165 3924
rect 2165 3918 2203 3924
rect 2203 3918 2237 3924
rect 2237 3918 2238 3924
rect 2058 3879 2238 3918
rect 2058 3845 2059 3879
rect 2059 3845 2093 3879
rect 2093 3845 2131 3879
rect 2131 3845 2165 3879
rect 2165 3845 2203 3879
rect 2203 3845 2237 3879
rect 2237 3845 2238 3879
rect 2058 3806 2238 3845
rect 2058 3772 2059 3806
rect 2059 3772 2093 3806
rect 2093 3772 2131 3806
rect 2131 3772 2165 3806
rect 2165 3772 2203 3806
rect 2203 3772 2237 3806
rect 2237 3772 2238 3806
rect 2058 3733 2238 3772
rect 2058 3699 2059 3733
rect 2059 3699 2093 3733
rect 2093 3699 2131 3733
rect 2131 3699 2165 3733
rect 2165 3699 2203 3733
rect 2203 3699 2237 3733
rect 2237 3699 2238 3733
rect 2058 3660 2238 3699
rect 2058 3626 2059 3660
rect 2059 3626 2093 3660
rect 2093 3626 2131 3660
rect 2131 3626 2165 3660
rect 2165 3626 2203 3660
rect 2203 3626 2237 3660
rect 2237 3626 2238 3660
rect 2058 3587 2238 3626
rect 2058 3553 2059 3587
rect 2059 3553 2093 3587
rect 2093 3553 2131 3587
rect 2131 3553 2165 3587
rect 2165 3553 2203 3587
rect 2203 3553 2237 3587
rect 2237 3553 2238 3587
rect 2058 3514 2238 3553
rect 2058 3480 2059 3514
rect 2059 3480 2093 3514
rect 2093 3480 2131 3514
rect 2131 3480 2165 3514
rect 2165 3480 2203 3514
rect 2203 3480 2237 3514
rect 2237 3480 2238 3514
rect 2058 3441 2238 3480
rect 2058 3407 2059 3441
rect 2059 3407 2093 3441
rect 2093 3407 2131 3441
rect 2131 3407 2165 3441
rect 2165 3407 2203 3441
rect 2203 3407 2237 3441
rect 2237 3407 2238 3441
rect 2058 3368 2238 3407
rect 2058 3334 2059 3368
rect 2059 3334 2093 3368
rect 2093 3334 2131 3368
rect 2131 3334 2165 3368
rect 2165 3334 2203 3368
rect 2203 3334 2237 3368
rect 2237 3334 2238 3368
rect 2058 3295 2238 3334
rect 2058 3261 2059 3295
rect 2059 3261 2093 3295
rect 2093 3261 2131 3295
rect 2131 3261 2165 3295
rect 2165 3261 2203 3295
rect 2203 3261 2237 3295
rect 2237 3261 2238 3295
rect 2058 3222 2238 3261
rect 2058 3188 2059 3222
rect 2059 3188 2093 3222
rect 2093 3188 2131 3222
rect 2131 3188 2165 3222
rect 2165 3188 2203 3222
rect 2203 3188 2237 3222
rect 2237 3188 2238 3222
rect 2058 3149 2238 3188
rect 2058 3115 2059 3149
rect 2059 3115 2093 3149
rect 2093 3115 2131 3149
rect 2131 3115 2165 3149
rect 2165 3115 2203 3149
rect 2203 3115 2237 3149
rect 2237 3115 2238 3149
rect 2058 3076 2238 3115
rect 2058 3042 2059 3076
rect 2059 3042 2093 3076
rect 2093 3042 2131 3076
rect 2131 3042 2165 3076
rect 2165 3042 2203 3076
rect 2203 3042 2237 3076
rect 2237 3042 2238 3076
rect 2058 3003 2238 3042
rect 2058 2969 2059 3003
rect 2059 2969 2093 3003
rect 2093 2969 2131 3003
rect 2131 2969 2165 3003
rect 2165 2969 2203 3003
rect 2203 2969 2237 3003
rect 2237 2969 2238 3003
rect 2058 2930 2238 2969
rect 2058 2896 2059 2930
rect 2059 2896 2093 2930
rect 2093 2896 2131 2930
rect 2131 2896 2165 2930
rect 2165 2896 2203 2930
rect 2203 2896 2237 2930
rect 2237 2896 2238 2930
rect 2058 2857 2238 2896
rect 2058 2823 2059 2857
rect 2059 2823 2093 2857
rect 2093 2823 2131 2857
rect 2131 2823 2165 2857
rect 2165 2823 2203 2857
rect 2203 2823 2237 2857
rect 2237 2823 2238 2857
rect 2058 2784 2238 2823
rect 2058 2750 2059 2784
rect 2059 2750 2093 2784
rect 2093 2750 2131 2784
rect 2131 2750 2165 2784
rect 2165 2750 2203 2784
rect 2203 2750 2237 2784
rect 2237 2750 2238 2784
rect 2058 2711 2238 2750
rect 2058 2677 2059 2711
rect 2059 2677 2093 2711
rect 2093 2677 2131 2711
rect 2131 2677 2165 2711
rect 2165 2677 2203 2711
rect 2203 2677 2237 2711
rect 2237 2677 2238 2711
rect 2058 2638 2238 2677
rect 2058 2604 2059 2638
rect 2059 2604 2093 2638
rect 2093 2604 2131 2638
rect 2131 2604 2165 2638
rect 2165 2604 2203 2638
rect 2203 2604 2237 2638
rect 2237 2604 2238 2638
rect 2058 2565 2238 2604
rect 2058 2531 2059 2565
rect 2059 2531 2093 2565
rect 2093 2531 2131 2565
rect 2131 2531 2165 2565
rect 2165 2531 2203 2565
rect 2203 2531 2237 2565
rect 2237 2531 2238 2565
rect 2058 2492 2238 2531
rect 2058 2458 2059 2492
rect 2059 2458 2093 2492
rect 2093 2458 2131 2492
rect 2131 2458 2165 2492
rect 2165 2458 2203 2492
rect 2203 2458 2237 2492
rect 2237 2458 2238 2492
rect 2058 2419 2238 2458
rect 2058 2385 2059 2419
rect 2059 2385 2093 2419
rect 2093 2385 2131 2419
rect 2131 2385 2165 2419
rect 2165 2385 2203 2419
rect 2203 2385 2237 2419
rect 2237 2385 2238 2419
rect 2058 2346 2238 2385
rect 2058 2312 2059 2346
rect 2059 2312 2093 2346
rect 2093 2312 2131 2346
rect 2131 2312 2165 2346
rect 2165 2312 2203 2346
rect 2203 2312 2237 2346
rect 2237 2312 2238 2346
rect 2058 2273 2238 2312
rect 2058 2239 2059 2273
rect 2059 2239 2093 2273
rect 2093 2239 2131 2273
rect 2131 2239 2165 2273
rect 2165 2239 2203 2273
rect 2203 2239 2237 2273
rect 2237 2239 2238 2273
rect 2058 2200 2238 2239
rect 2058 2166 2059 2200
rect 2059 2166 2093 2200
rect 2093 2166 2131 2200
rect 2131 2166 2165 2200
rect 2165 2166 2203 2200
rect 2203 2166 2237 2200
rect 2237 2166 2238 2200
rect 2058 2126 2238 2166
rect 2058 2092 2059 2126
rect 2059 2092 2093 2126
rect 2093 2092 2131 2126
rect 2131 2092 2165 2126
rect 2165 2092 2203 2126
rect 2203 2092 2237 2126
rect 2237 2092 2238 2126
rect 2058 2052 2238 2092
rect 2058 2018 2059 2052
rect 2059 2018 2093 2052
rect 2093 2018 2131 2052
rect 2131 2018 2165 2052
rect 2165 2018 2203 2052
rect 2203 2018 2237 2052
rect 2237 2018 2238 2052
rect 2058 1978 2238 2018
rect 2058 1944 2059 1978
rect 2059 1944 2093 1978
rect 2093 1944 2131 1978
rect 2131 1944 2165 1978
rect 2165 1944 2203 1978
rect 2203 1944 2237 1978
rect 2237 1944 2238 1978
rect 2058 1904 2238 1944
rect 2058 1870 2059 1904
rect 2059 1870 2093 1904
rect 2093 1870 2131 1904
rect 2131 1870 2165 1904
rect 2165 1870 2203 1904
rect 2203 1870 2237 1904
rect 2237 1870 2238 1904
rect 2058 1830 2238 1870
rect 2058 1796 2059 1830
rect 2059 1796 2093 1830
rect 2093 1796 2131 1830
rect 2131 1796 2165 1830
rect 2165 1796 2203 1830
rect 2203 1796 2237 1830
rect 2237 1796 2238 1830
rect 2058 1756 2238 1796
rect 2058 1722 2059 1756
rect 2059 1722 2093 1756
rect 2093 1722 2131 1756
rect 2131 1722 2165 1756
rect 2165 1722 2203 1756
rect 2203 1722 2237 1756
rect 2237 1722 2238 1756
rect 2058 1682 2238 1722
rect 2058 1648 2059 1682
rect 2059 1648 2093 1682
rect 2093 1648 2131 1682
rect 2131 1648 2165 1682
rect 2165 1648 2203 1682
rect 2203 1648 2237 1682
rect 2237 1648 2238 1682
rect 2058 1608 2238 1648
rect 2058 1574 2059 1608
rect 2059 1574 2093 1608
rect 2093 1574 2131 1608
rect 2131 1574 2165 1608
rect 2165 1574 2203 1608
rect 2203 1574 2237 1608
rect 2237 1574 2238 1608
rect 2058 1568 2238 1574
rect 2554 4092 2606 4124
rect 2554 4072 2555 4092
rect 2555 4072 2589 4092
rect 2589 4072 2606 4092
rect 2618 4072 2670 4124
rect 2682 4092 2734 4124
rect 2682 4072 2699 4092
rect 2699 4072 2733 4092
rect 2733 4072 2734 4092
rect 2554 4058 2555 4059
rect 2555 4058 2589 4059
rect 2589 4058 2606 4059
rect 2554 4020 2606 4058
rect 2554 4007 2555 4020
rect 2555 4007 2589 4020
rect 2589 4007 2606 4020
rect 2618 4007 2670 4059
rect 2682 4058 2699 4059
rect 2699 4058 2733 4059
rect 2733 4058 2734 4059
rect 2682 4020 2734 4058
rect 2682 4007 2699 4020
rect 2699 4007 2733 4020
rect 2733 4007 2734 4020
rect 2554 3986 2555 3994
rect 2555 3986 2589 3994
rect 2589 3986 2606 3994
rect 2554 3948 2606 3986
rect 2554 3942 2555 3948
rect 2555 3942 2589 3948
rect 2589 3942 2606 3948
rect 2618 3942 2670 3994
rect 2682 3986 2699 3994
rect 2699 3986 2733 3994
rect 2733 3986 2734 3994
rect 2682 3948 2734 3986
rect 2682 3942 2699 3948
rect 2699 3942 2733 3948
rect 2733 3942 2734 3948
rect 2554 3914 2555 3929
rect 2555 3914 2589 3929
rect 2589 3914 2606 3929
rect 2554 3877 2606 3914
rect 2618 3877 2670 3929
rect 2682 3914 2699 3929
rect 2699 3914 2733 3929
rect 2733 3914 2734 3929
rect 2682 3877 2734 3914
rect 2554 3842 2555 3864
rect 2555 3842 2589 3864
rect 2589 3842 2606 3864
rect 2554 3812 2606 3842
rect 2618 3812 2670 3864
rect 2682 3842 2699 3864
rect 2699 3842 2733 3864
rect 2733 3842 2734 3864
rect 2682 3812 2734 3842
rect 2554 3770 2555 3799
rect 2555 3770 2589 3799
rect 2589 3770 2606 3799
rect 2554 3747 2606 3770
rect 2618 3747 2670 3799
rect 2682 3770 2699 3799
rect 2699 3770 2733 3799
rect 2733 3770 2734 3799
rect 2682 3747 2734 3770
rect 2554 3732 2606 3734
rect 2554 3698 2555 3732
rect 2555 3698 2589 3732
rect 2589 3698 2606 3732
rect 2554 3682 2606 3698
rect 2618 3682 2670 3734
rect 2682 3732 2734 3734
rect 2682 3698 2699 3732
rect 2699 3698 2733 3732
rect 2733 3698 2734 3732
rect 2682 3682 2734 3698
rect 2554 3660 2606 3669
rect 2554 3626 2555 3660
rect 2555 3626 2589 3660
rect 2589 3626 2606 3660
rect 2554 3617 2606 3626
rect 2618 3617 2670 3669
rect 2682 3660 2734 3669
rect 2682 3626 2699 3660
rect 2699 3626 2733 3660
rect 2733 3626 2734 3660
rect 2682 3617 2734 3626
rect 2554 3588 2734 3604
rect 2554 3554 2555 3588
rect 2555 3554 2589 3588
rect 2589 3554 2699 3588
rect 2699 3554 2733 3588
rect 2733 3554 2734 3588
rect 2554 3516 2734 3554
rect 2554 3482 2555 3516
rect 2555 3482 2589 3516
rect 2589 3482 2699 3516
rect 2699 3482 2733 3516
rect 2733 3482 2734 3516
rect 2554 3444 2734 3482
rect 2554 3410 2555 3444
rect 2555 3410 2589 3444
rect 2589 3410 2699 3444
rect 2699 3410 2733 3444
rect 2733 3410 2734 3444
rect 2554 3372 2734 3410
rect 2554 3338 2555 3372
rect 2555 3338 2589 3372
rect 2589 3338 2699 3372
rect 2699 3338 2733 3372
rect 2733 3338 2734 3372
rect 2554 3300 2734 3338
rect 2554 3266 2555 3300
rect 2555 3266 2589 3300
rect 2589 3266 2699 3300
rect 2699 3266 2733 3300
rect 2733 3266 2734 3300
rect 2554 3228 2734 3266
rect 2554 3194 2555 3228
rect 2555 3194 2589 3228
rect 2589 3194 2699 3228
rect 2699 3194 2733 3228
rect 2733 3194 2734 3228
rect 2554 3108 2734 3194
rect 2554 3074 2555 3108
rect 2555 3074 2589 3108
rect 2589 3074 2627 3108
rect 2627 3074 2661 3108
rect 2661 3074 2699 3108
rect 2699 3074 2733 3108
rect 2733 3074 2734 3108
rect 2554 3028 2734 3074
rect 2554 2994 2555 3028
rect 2555 2994 2589 3028
rect 2589 2994 2627 3028
rect 2627 2994 2661 3028
rect 2661 2994 2699 3028
rect 2699 2994 2733 3028
rect 2733 2994 2734 3028
rect 2554 2948 2734 2994
rect 2554 2914 2555 2948
rect 2555 2914 2589 2948
rect 2589 2914 2627 2948
rect 2627 2914 2661 2948
rect 2661 2914 2699 2948
rect 2699 2914 2733 2948
rect 2733 2914 2734 2948
rect 2554 2868 2734 2914
rect 2554 2834 2555 2868
rect 2555 2834 2589 2868
rect 2589 2834 2627 2868
rect 2627 2834 2661 2868
rect 2661 2834 2699 2868
rect 2699 2834 2733 2868
rect 2733 2834 2734 2868
rect 2554 2788 2734 2834
rect 2554 2754 2555 2788
rect 2555 2754 2589 2788
rect 2589 2754 2627 2788
rect 2627 2754 2661 2788
rect 2661 2754 2699 2788
rect 2699 2754 2733 2788
rect 2733 2754 2734 2788
rect 2554 2708 2734 2754
rect 2554 2674 2555 2708
rect 2555 2674 2589 2708
rect 2589 2674 2627 2708
rect 2627 2674 2661 2708
rect 2661 2674 2699 2708
rect 2699 2674 2733 2708
rect 2733 2674 2734 2708
rect 2554 2628 2734 2674
rect 2554 2594 2555 2628
rect 2555 2594 2589 2628
rect 2589 2594 2627 2628
rect 2627 2594 2661 2628
rect 2661 2594 2699 2628
rect 2699 2594 2733 2628
rect 2733 2594 2734 2628
rect 2554 2518 2734 2594
rect 2554 2484 2555 2518
rect 2555 2484 2589 2518
rect 2589 2484 2699 2518
rect 2699 2484 2733 2518
rect 2733 2484 2734 2518
rect 2554 2446 2734 2484
rect 2554 2412 2555 2446
rect 2555 2412 2589 2446
rect 2589 2412 2699 2446
rect 2699 2412 2733 2446
rect 2733 2412 2734 2446
rect 2554 2374 2734 2412
rect 2554 2340 2555 2374
rect 2555 2340 2589 2374
rect 2589 2340 2699 2374
rect 2699 2340 2733 2374
rect 2733 2340 2734 2374
rect 2554 2302 2734 2340
rect 2554 2268 2555 2302
rect 2555 2268 2589 2302
rect 2589 2268 2699 2302
rect 2699 2268 2733 2302
rect 2733 2268 2734 2302
rect 2554 2230 2734 2268
rect 2554 2196 2555 2230
rect 2555 2196 2589 2230
rect 2589 2196 2699 2230
rect 2699 2196 2733 2230
rect 2733 2196 2734 2230
rect 2554 2158 2734 2196
rect 2554 2124 2555 2158
rect 2555 2124 2589 2158
rect 2589 2124 2699 2158
rect 2699 2124 2733 2158
rect 2733 2124 2734 2158
rect 2554 2086 2734 2124
rect 2554 2052 2555 2086
rect 2555 2052 2589 2086
rect 2589 2052 2699 2086
rect 2699 2052 2733 2086
rect 2733 2052 2734 2086
rect 2554 2014 2734 2052
rect 2554 1980 2555 2014
rect 2555 1980 2589 2014
rect 2589 1980 2699 2014
rect 2699 1980 2733 2014
rect 2733 1980 2734 2014
rect 2554 1942 2734 1980
rect 2554 1908 2555 1942
rect 2555 1908 2589 1942
rect 2589 1908 2699 1942
rect 2699 1908 2733 1942
rect 2733 1908 2734 1942
rect 2554 1870 2734 1908
rect 2554 1836 2555 1870
rect 2555 1836 2589 1870
rect 2589 1836 2699 1870
rect 2699 1836 2733 1870
rect 2733 1836 2734 1870
rect 2554 1798 2734 1836
rect 2554 1764 2555 1798
rect 2555 1764 2589 1798
rect 2589 1764 2699 1798
rect 2699 1764 2733 1798
rect 2733 1764 2734 1798
rect 2554 1726 2734 1764
rect 2554 1692 2555 1726
rect 2555 1692 2589 1726
rect 2589 1692 2699 1726
rect 2699 1692 2733 1726
rect 2733 1692 2734 1726
rect 2554 1654 2734 1692
rect 2554 1620 2555 1654
rect 2555 1620 2589 1654
rect 2589 1620 2699 1654
rect 2699 1620 2733 1654
rect 2733 1620 2734 1654
rect 2554 1568 2734 1620
rect 3050 4098 3102 4119
rect 3050 4067 3051 4098
rect 3051 4067 3085 4098
rect 3085 4067 3102 4098
rect 3114 4098 3166 4119
rect 3114 4067 3123 4098
rect 3123 4067 3157 4098
rect 3157 4067 3166 4098
rect 3178 4098 3230 4119
rect 3178 4067 3195 4098
rect 3195 4067 3229 4098
rect 3229 4067 3230 4098
rect 3050 4025 3102 4054
rect 3050 4002 3051 4025
rect 3051 4002 3085 4025
rect 3085 4002 3102 4025
rect 3114 4025 3166 4054
rect 3114 4002 3123 4025
rect 3123 4002 3157 4025
rect 3157 4002 3166 4025
rect 3178 4025 3230 4054
rect 3178 4002 3195 4025
rect 3195 4002 3229 4025
rect 3229 4002 3230 4025
rect 3050 3952 3102 3989
rect 3050 3937 3051 3952
rect 3051 3937 3085 3952
rect 3085 3937 3102 3952
rect 3114 3952 3166 3989
rect 3114 3937 3123 3952
rect 3123 3937 3157 3952
rect 3157 3937 3166 3952
rect 3178 3952 3230 3989
rect 3178 3937 3195 3952
rect 3195 3937 3229 3952
rect 3229 3937 3230 3952
rect 3050 3918 3051 3924
rect 3051 3918 3085 3924
rect 3085 3918 3123 3924
rect 3123 3918 3157 3924
rect 3157 3918 3195 3924
rect 3195 3918 3229 3924
rect 3229 3918 3230 3924
rect 3050 3879 3230 3918
rect 3050 3845 3051 3879
rect 3051 3845 3085 3879
rect 3085 3845 3123 3879
rect 3123 3845 3157 3879
rect 3157 3845 3195 3879
rect 3195 3845 3229 3879
rect 3229 3845 3230 3879
rect 3050 3806 3230 3845
rect 3050 3772 3051 3806
rect 3051 3772 3085 3806
rect 3085 3772 3123 3806
rect 3123 3772 3157 3806
rect 3157 3772 3195 3806
rect 3195 3772 3229 3806
rect 3229 3772 3230 3806
rect 3050 3733 3230 3772
rect 3050 3699 3051 3733
rect 3051 3699 3085 3733
rect 3085 3699 3123 3733
rect 3123 3699 3157 3733
rect 3157 3699 3195 3733
rect 3195 3699 3229 3733
rect 3229 3699 3230 3733
rect 3050 3660 3230 3699
rect 3050 3626 3051 3660
rect 3051 3626 3085 3660
rect 3085 3626 3123 3660
rect 3123 3626 3157 3660
rect 3157 3626 3195 3660
rect 3195 3626 3229 3660
rect 3229 3626 3230 3660
rect 3050 3587 3230 3626
rect 3050 3553 3051 3587
rect 3051 3553 3085 3587
rect 3085 3553 3123 3587
rect 3123 3553 3157 3587
rect 3157 3553 3195 3587
rect 3195 3553 3229 3587
rect 3229 3553 3230 3587
rect 3050 3514 3230 3553
rect 3050 3480 3051 3514
rect 3051 3480 3085 3514
rect 3085 3480 3123 3514
rect 3123 3480 3157 3514
rect 3157 3480 3195 3514
rect 3195 3480 3229 3514
rect 3229 3480 3230 3514
rect 3050 3441 3230 3480
rect 3050 3407 3051 3441
rect 3051 3407 3085 3441
rect 3085 3407 3123 3441
rect 3123 3407 3157 3441
rect 3157 3407 3195 3441
rect 3195 3407 3229 3441
rect 3229 3407 3230 3441
rect 3050 3368 3230 3407
rect 3050 3334 3051 3368
rect 3051 3334 3085 3368
rect 3085 3334 3123 3368
rect 3123 3334 3157 3368
rect 3157 3334 3195 3368
rect 3195 3334 3229 3368
rect 3229 3334 3230 3368
rect 3050 3295 3230 3334
rect 3050 3261 3051 3295
rect 3051 3261 3085 3295
rect 3085 3261 3123 3295
rect 3123 3261 3157 3295
rect 3157 3261 3195 3295
rect 3195 3261 3229 3295
rect 3229 3261 3230 3295
rect 3050 3222 3230 3261
rect 3050 3188 3051 3222
rect 3051 3188 3085 3222
rect 3085 3188 3123 3222
rect 3123 3188 3157 3222
rect 3157 3188 3195 3222
rect 3195 3188 3229 3222
rect 3229 3188 3230 3222
rect 3050 3149 3230 3188
rect 3050 3115 3051 3149
rect 3051 3115 3085 3149
rect 3085 3115 3123 3149
rect 3123 3115 3157 3149
rect 3157 3115 3195 3149
rect 3195 3115 3229 3149
rect 3229 3115 3230 3149
rect 3050 3076 3230 3115
rect 3050 3042 3051 3076
rect 3051 3042 3085 3076
rect 3085 3042 3123 3076
rect 3123 3042 3157 3076
rect 3157 3042 3195 3076
rect 3195 3042 3229 3076
rect 3229 3042 3230 3076
rect 3050 3003 3230 3042
rect 3050 2969 3051 3003
rect 3051 2969 3085 3003
rect 3085 2969 3123 3003
rect 3123 2969 3157 3003
rect 3157 2969 3195 3003
rect 3195 2969 3229 3003
rect 3229 2969 3230 3003
rect 3050 2930 3230 2969
rect 3050 2896 3051 2930
rect 3051 2896 3085 2930
rect 3085 2896 3123 2930
rect 3123 2896 3157 2930
rect 3157 2896 3195 2930
rect 3195 2896 3229 2930
rect 3229 2896 3230 2930
rect 3050 2857 3230 2896
rect 3050 2823 3051 2857
rect 3051 2823 3085 2857
rect 3085 2823 3123 2857
rect 3123 2823 3157 2857
rect 3157 2823 3195 2857
rect 3195 2823 3229 2857
rect 3229 2823 3230 2857
rect 3050 2784 3230 2823
rect 3050 2750 3051 2784
rect 3051 2750 3085 2784
rect 3085 2750 3123 2784
rect 3123 2750 3157 2784
rect 3157 2750 3195 2784
rect 3195 2750 3229 2784
rect 3229 2750 3230 2784
rect 3050 2711 3230 2750
rect 3050 2677 3051 2711
rect 3051 2677 3085 2711
rect 3085 2677 3123 2711
rect 3123 2677 3157 2711
rect 3157 2677 3195 2711
rect 3195 2677 3229 2711
rect 3229 2677 3230 2711
rect 3050 2638 3230 2677
rect 3050 2604 3051 2638
rect 3051 2604 3085 2638
rect 3085 2604 3123 2638
rect 3123 2604 3157 2638
rect 3157 2604 3195 2638
rect 3195 2604 3229 2638
rect 3229 2604 3230 2638
rect 3050 2565 3230 2604
rect 3050 2531 3051 2565
rect 3051 2531 3085 2565
rect 3085 2531 3123 2565
rect 3123 2531 3157 2565
rect 3157 2531 3195 2565
rect 3195 2531 3229 2565
rect 3229 2531 3230 2565
rect 3050 2492 3230 2531
rect 3050 2458 3051 2492
rect 3051 2458 3085 2492
rect 3085 2458 3123 2492
rect 3123 2458 3157 2492
rect 3157 2458 3195 2492
rect 3195 2458 3229 2492
rect 3229 2458 3230 2492
rect 3050 2419 3230 2458
rect 3050 2385 3051 2419
rect 3051 2385 3085 2419
rect 3085 2385 3123 2419
rect 3123 2385 3157 2419
rect 3157 2385 3195 2419
rect 3195 2385 3229 2419
rect 3229 2385 3230 2419
rect 3050 2346 3230 2385
rect 3050 2312 3051 2346
rect 3051 2312 3085 2346
rect 3085 2312 3123 2346
rect 3123 2312 3157 2346
rect 3157 2312 3195 2346
rect 3195 2312 3229 2346
rect 3229 2312 3230 2346
rect 3050 2273 3230 2312
rect 3050 2239 3051 2273
rect 3051 2239 3085 2273
rect 3085 2239 3123 2273
rect 3123 2239 3157 2273
rect 3157 2239 3195 2273
rect 3195 2239 3229 2273
rect 3229 2239 3230 2273
rect 3050 2200 3230 2239
rect 3050 2166 3051 2200
rect 3051 2166 3085 2200
rect 3085 2166 3123 2200
rect 3123 2166 3157 2200
rect 3157 2166 3195 2200
rect 3195 2166 3229 2200
rect 3229 2166 3230 2200
rect 3050 2126 3230 2166
rect 3050 2092 3051 2126
rect 3051 2092 3085 2126
rect 3085 2092 3123 2126
rect 3123 2092 3157 2126
rect 3157 2092 3195 2126
rect 3195 2092 3229 2126
rect 3229 2092 3230 2126
rect 3050 2052 3230 2092
rect 3050 2018 3051 2052
rect 3051 2018 3085 2052
rect 3085 2018 3123 2052
rect 3123 2018 3157 2052
rect 3157 2018 3195 2052
rect 3195 2018 3229 2052
rect 3229 2018 3230 2052
rect 3050 1978 3230 2018
rect 3050 1944 3051 1978
rect 3051 1944 3085 1978
rect 3085 1944 3123 1978
rect 3123 1944 3157 1978
rect 3157 1944 3195 1978
rect 3195 1944 3229 1978
rect 3229 1944 3230 1978
rect 3050 1904 3230 1944
rect 3050 1870 3051 1904
rect 3051 1870 3085 1904
rect 3085 1870 3123 1904
rect 3123 1870 3157 1904
rect 3157 1870 3195 1904
rect 3195 1870 3229 1904
rect 3229 1870 3230 1904
rect 3050 1830 3230 1870
rect 3050 1796 3051 1830
rect 3051 1796 3085 1830
rect 3085 1796 3123 1830
rect 3123 1796 3157 1830
rect 3157 1796 3195 1830
rect 3195 1796 3229 1830
rect 3229 1796 3230 1830
rect 3050 1756 3230 1796
rect 3050 1722 3051 1756
rect 3051 1722 3085 1756
rect 3085 1722 3123 1756
rect 3123 1722 3157 1756
rect 3157 1722 3195 1756
rect 3195 1722 3229 1756
rect 3229 1722 3230 1756
rect 3050 1682 3230 1722
rect 3050 1648 3051 1682
rect 3051 1648 3085 1682
rect 3085 1648 3123 1682
rect 3123 1648 3157 1682
rect 3157 1648 3195 1682
rect 3195 1648 3229 1682
rect 3229 1648 3230 1682
rect 3050 1608 3230 1648
rect 3050 1574 3051 1608
rect 3051 1574 3085 1608
rect 3085 1574 3123 1608
rect 3123 1574 3157 1608
rect 3157 1574 3195 1608
rect 3195 1574 3229 1608
rect 3229 1574 3230 1608
rect 3050 1568 3230 1574
rect 3546 4092 3598 4124
rect 3546 4072 3547 4092
rect 3547 4072 3581 4092
rect 3581 4072 3598 4092
rect 3610 4072 3662 4124
rect 3674 4092 3726 4124
rect 3674 4072 3691 4092
rect 3691 4072 3725 4092
rect 3725 4072 3726 4092
rect 3546 4058 3547 4059
rect 3547 4058 3581 4059
rect 3581 4058 3598 4059
rect 3546 4020 3598 4058
rect 3546 4007 3547 4020
rect 3547 4007 3581 4020
rect 3581 4007 3598 4020
rect 3610 4007 3662 4059
rect 3674 4058 3691 4059
rect 3691 4058 3725 4059
rect 3725 4058 3726 4059
rect 3674 4020 3726 4058
rect 3674 4007 3691 4020
rect 3691 4007 3725 4020
rect 3725 4007 3726 4020
rect 3546 3986 3547 3994
rect 3547 3986 3581 3994
rect 3581 3986 3598 3994
rect 3546 3948 3598 3986
rect 3546 3942 3547 3948
rect 3547 3942 3581 3948
rect 3581 3942 3598 3948
rect 3610 3942 3662 3994
rect 3674 3986 3691 3994
rect 3691 3986 3725 3994
rect 3725 3986 3726 3994
rect 3674 3948 3726 3986
rect 3674 3942 3691 3948
rect 3691 3942 3725 3948
rect 3725 3942 3726 3948
rect 3546 3914 3547 3929
rect 3547 3914 3581 3929
rect 3581 3914 3598 3929
rect 3546 3877 3598 3914
rect 3610 3877 3662 3929
rect 3674 3914 3691 3929
rect 3691 3914 3725 3929
rect 3725 3914 3726 3929
rect 3674 3877 3726 3914
rect 3546 3842 3547 3864
rect 3547 3842 3581 3864
rect 3581 3842 3598 3864
rect 3546 3812 3598 3842
rect 3610 3812 3662 3864
rect 3674 3842 3691 3864
rect 3691 3842 3725 3864
rect 3725 3842 3726 3864
rect 3674 3812 3726 3842
rect 3546 3770 3547 3799
rect 3547 3770 3581 3799
rect 3581 3770 3598 3799
rect 3546 3747 3598 3770
rect 3610 3747 3662 3799
rect 3674 3770 3691 3799
rect 3691 3770 3725 3799
rect 3725 3770 3726 3799
rect 3674 3747 3726 3770
rect 3546 3732 3598 3734
rect 3546 3698 3547 3732
rect 3547 3698 3581 3732
rect 3581 3698 3598 3732
rect 3546 3682 3598 3698
rect 3610 3682 3662 3734
rect 3674 3732 3726 3734
rect 3674 3698 3691 3732
rect 3691 3698 3725 3732
rect 3725 3698 3726 3732
rect 3674 3682 3726 3698
rect 3546 3660 3598 3669
rect 3546 3626 3547 3660
rect 3547 3626 3581 3660
rect 3581 3626 3598 3660
rect 3546 3617 3598 3626
rect 3610 3617 3662 3669
rect 3674 3660 3726 3669
rect 3674 3626 3691 3660
rect 3691 3626 3725 3660
rect 3725 3626 3726 3660
rect 3674 3617 3726 3626
rect 3546 3588 3726 3604
rect 3546 3554 3547 3588
rect 3547 3554 3581 3588
rect 3581 3554 3691 3588
rect 3691 3554 3725 3588
rect 3725 3554 3726 3588
rect 3546 3516 3726 3554
rect 3546 3482 3547 3516
rect 3547 3482 3581 3516
rect 3581 3482 3691 3516
rect 3691 3482 3725 3516
rect 3725 3482 3726 3516
rect 3546 3444 3726 3482
rect 3546 3410 3547 3444
rect 3547 3410 3581 3444
rect 3581 3410 3691 3444
rect 3691 3410 3725 3444
rect 3725 3410 3726 3444
rect 3546 3372 3726 3410
rect 3546 3338 3547 3372
rect 3547 3338 3581 3372
rect 3581 3338 3691 3372
rect 3691 3338 3725 3372
rect 3725 3338 3726 3372
rect 3546 3300 3726 3338
rect 3546 3266 3547 3300
rect 3547 3266 3581 3300
rect 3581 3266 3691 3300
rect 3691 3266 3725 3300
rect 3725 3266 3726 3300
rect 3546 3228 3726 3266
rect 3546 3194 3547 3228
rect 3547 3194 3581 3228
rect 3581 3194 3691 3228
rect 3691 3194 3725 3228
rect 3725 3194 3726 3228
rect 3546 3108 3726 3194
rect 3546 3074 3547 3108
rect 3547 3074 3581 3108
rect 3581 3074 3619 3108
rect 3619 3074 3653 3108
rect 3653 3074 3691 3108
rect 3691 3074 3725 3108
rect 3725 3074 3726 3108
rect 3546 3028 3726 3074
rect 3546 2994 3547 3028
rect 3547 2994 3581 3028
rect 3581 2994 3619 3028
rect 3619 2994 3653 3028
rect 3653 2994 3691 3028
rect 3691 2994 3725 3028
rect 3725 2994 3726 3028
rect 3546 2948 3726 2994
rect 3546 2914 3547 2948
rect 3547 2914 3581 2948
rect 3581 2914 3619 2948
rect 3619 2914 3653 2948
rect 3653 2914 3691 2948
rect 3691 2914 3725 2948
rect 3725 2914 3726 2948
rect 3546 2868 3726 2914
rect 3546 2834 3547 2868
rect 3547 2834 3581 2868
rect 3581 2834 3619 2868
rect 3619 2834 3653 2868
rect 3653 2834 3691 2868
rect 3691 2834 3725 2868
rect 3725 2834 3726 2868
rect 3546 2788 3726 2834
rect 3546 2754 3547 2788
rect 3547 2754 3581 2788
rect 3581 2754 3619 2788
rect 3619 2754 3653 2788
rect 3653 2754 3691 2788
rect 3691 2754 3725 2788
rect 3725 2754 3726 2788
rect 3546 2708 3726 2754
rect 3546 2674 3547 2708
rect 3547 2674 3581 2708
rect 3581 2674 3619 2708
rect 3619 2674 3653 2708
rect 3653 2674 3691 2708
rect 3691 2674 3725 2708
rect 3725 2674 3726 2708
rect 3546 2628 3726 2674
rect 3546 2594 3547 2628
rect 3547 2594 3581 2628
rect 3581 2594 3619 2628
rect 3619 2594 3653 2628
rect 3653 2594 3691 2628
rect 3691 2594 3725 2628
rect 3725 2594 3726 2628
rect 3546 2518 3726 2594
rect 3546 2484 3547 2518
rect 3547 2484 3581 2518
rect 3581 2484 3691 2518
rect 3691 2484 3725 2518
rect 3725 2484 3726 2518
rect 3546 2446 3726 2484
rect 3546 2412 3547 2446
rect 3547 2412 3581 2446
rect 3581 2412 3691 2446
rect 3691 2412 3725 2446
rect 3725 2412 3726 2446
rect 3546 2374 3726 2412
rect 3546 2340 3547 2374
rect 3547 2340 3581 2374
rect 3581 2340 3691 2374
rect 3691 2340 3725 2374
rect 3725 2340 3726 2374
rect 3546 2302 3726 2340
rect 3546 2268 3547 2302
rect 3547 2268 3581 2302
rect 3581 2268 3691 2302
rect 3691 2268 3725 2302
rect 3725 2268 3726 2302
rect 3546 2230 3726 2268
rect 3546 2196 3547 2230
rect 3547 2196 3581 2230
rect 3581 2196 3691 2230
rect 3691 2196 3725 2230
rect 3725 2196 3726 2230
rect 3546 2158 3726 2196
rect 3546 2124 3547 2158
rect 3547 2124 3581 2158
rect 3581 2124 3691 2158
rect 3691 2124 3725 2158
rect 3725 2124 3726 2158
rect 3546 2086 3726 2124
rect 3546 2052 3547 2086
rect 3547 2052 3581 2086
rect 3581 2052 3691 2086
rect 3691 2052 3725 2086
rect 3725 2052 3726 2086
rect 3546 2014 3726 2052
rect 3546 1980 3547 2014
rect 3547 1980 3581 2014
rect 3581 1980 3691 2014
rect 3691 1980 3725 2014
rect 3725 1980 3726 2014
rect 3546 1942 3726 1980
rect 3546 1908 3547 1942
rect 3547 1908 3581 1942
rect 3581 1908 3691 1942
rect 3691 1908 3725 1942
rect 3725 1908 3726 1942
rect 3546 1870 3726 1908
rect 3546 1836 3547 1870
rect 3547 1836 3581 1870
rect 3581 1836 3691 1870
rect 3691 1836 3725 1870
rect 3725 1836 3726 1870
rect 3546 1798 3726 1836
rect 3546 1764 3547 1798
rect 3547 1764 3581 1798
rect 3581 1764 3691 1798
rect 3691 1764 3725 1798
rect 3725 1764 3726 1798
rect 3546 1726 3726 1764
rect 3546 1692 3547 1726
rect 3547 1692 3581 1726
rect 3581 1692 3691 1726
rect 3691 1692 3725 1726
rect 3725 1692 3726 1726
rect 3546 1654 3726 1692
rect 3546 1620 3547 1654
rect 3547 1620 3581 1654
rect 3581 1620 3691 1654
rect 3691 1620 3725 1654
rect 3725 1620 3726 1654
rect 3546 1568 3726 1620
rect 4042 4098 4094 4119
rect 4042 4067 4043 4098
rect 4043 4067 4077 4098
rect 4077 4067 4094 4098
rect 4106 4098 4158 4119
rect 4106 4067 4115 4098
rect 4115 4067 4149 4098
rect 4149 4067 4158 4098
rect 4170 4098 4222 4119
rect 4170 4067 4187 4098
rect 4187 4067 4221 4098
rect 4221 4067 4222 4098
rect 4042 4025 4094 4054
rect 4042 4002 4043 4025
rect 4043 4002 4077 4025
rect 4077 4002 4094 4025
rect 4106 4025 4158 4054
rect 4106 4002 4115 4025
rect 4115 4002 4149 4025
rect 4149 4002 4158 4025
rect 4170 4025 4222 4054
rect 4170 4002 4187 4025
rect 4187 4002 4221 4025
rect 4221 4002 4222 4025
rect 4042 3952 4094 3989
rect 4042 3937 4043 3952
rect 4043 3937 4077 3952
rect 4077 3937 4094 3952
rect 4106 3952 4158 3989
rect 4106 3937 4115 3952
rect 4115 3937 4149 3952
rect 4149 3937 4158 3952
rect 4170 3952 4222 3989
rect 4170 3937 4187 3952
rect 4187 3937 4221 3952
rect 4221 3937 4222 3952
rect 4042 3918 4043 3924
rect 4043 3918 4077 3924
rect 4077 3918 4115 3924
rect 4115 3918 4149 3924
rect 4149 3918 4187 3924
rect 4187 3918 4221 3924
rect 4221 3918 4222 3924
rect 4042 3879 4222 3918
rect 4042 3845 4043 3879
rect 4043 3845 4077 3879
rect 4077 3845 4115 3879
rect 4115 3845 4149 3879
rect 4149 3845 4187 3879
rect 4187 3845 4221 3879
rect 4221 3845 4222 3879
rect 4042 3806 4222 3845
rect 4042 3772 4043 3806
rect 4043 3772 4077 3806
rect 4077 3772 4115 3806
rect 4115 3772 4149 3806
rect 4149 3772 4187 3806
rect 4187 3772 4221 3806
rect 4221 3772 4222 3806
rect 4042 3733 4222 3772
rect 4042 3699 4043 3733
rect 4043 3699 4077 3733
rect 4077 3699 4115 3733
rect 4115 3699 4149 3733
rect 4149 3699 4187 3733
rect 4187 3699 4221 3733
rect 4221 3699 4222 3733
rect 4042 3660 4222 3699
rect 4042 3626 4043 3660
rect 4043 3626 4077 3660
rect 4077 3626 4115 3660
rect 4115 3626 4149 3660
rect 4149 3626 4187 3660
rect 4187 3626 4221 3660
rect 4221 3626 4222 3660
rect 4042 3587 4222 3626
rect 4042 3553 4043 3587
rect 4043 3553 4077 3587
rect 4077 3553 4115 3587
rect 4115 3553 4149 3587
rect 4149 3553 4187 3587
rect 4187 3553 4221 3587
rect 4221 3553 4222 3587
rect 4042 3514 4222 3553
rect 4042 3480 4043 3514
rect 4043 3480 4077 3514
rect 4077 3480 4115 3514
rect 4115 3480 4149 3514
rect 4149 3480 4187 3514
rect 4187 3480 4221 3514
rect 4221 3480 4222 3514
rect 4042 3441 4222 3480
rect 4042 3407 4043 3441
rect 4043 3407 4077 3441
rect 4077 3407 4115 3441
rect 4115 3407 4149 3441
rect 4149 3407 4187 3441
rect 4187 3407 4221 3441
rect 4221 3407 4222 3441
rect 4042 3368 4222 3407
rect 4042 3334 4043 3368
rect 4043 3334 4077 3368
rect 4077 3334 4115 3368
rect 4115 3334 4149 3368
rect 4149 3334 4187 3368
rect 4187 3334 4221 3368
rect 4221 3334 4222 3368
rect 4042 3295 4222 3334
rect 4042 3261 4043 3295
rect 4043 3261 4077 3295
rect 4077 3261 4115 3295
rect 4115 3261 4149 3295
rect 4149 3261 4187 3295
rect 4187 3261 4221 3295
rect 4221 3261 4222 3295
rect 4042 3222 4222 3261
rect 4042 3188 4043 3222
rect 4043 3188 4077 3222
rect 4077 3188 4115 3222
rect 4115 3188 4149 3222
rect 4149 3188 4187 3222
rect 4187 3188 4221 3222
rect 4221 3188 4222 3222
rect 4042 3149 4222 3188
rect 4042 3115 4043 3149
rect 4043 3115 4077 3149
rect 4077 3115 4115 3149
rect 4115 3115 4149 3149
rect 4149 3115 4187 3149
rect 4187 3115 4221 3149
rect 4221 3115 4222 3149
rect 4042 3076 4222 3115
rect 4042 3042 4043 3076
rect 4043 3042 4077 3076
rect 4077 3042 4115 3076
rect 4115 3042 4149 3076
rect 4149 3042 4187 3076
rect 4187 3042 4221 3076
rect 4221 3042 4222 3076
rect 4042 3003 4222 3042
rect 4042 2969 4043 3003
rect 4043 2969 4077 3003
rect 4077 2969 4115 3003
rect 4115 2969 4149 3003
rect 4149 2969 4187 3003
rect 4187 2969 4221 3003
rect 4221 2969 4222 3003
rect 4042 2930 4222 2969
rect 4042 2896 4043 2930
rect 4043 2896 4077 2930
rect 4077 2896 4115 2930
rect 4115 2896 4149 2930
rect 4149 2896 4187 2930
rect 4187 2896 4221 2930
rect 4221 2896 4222 2930
rect 4042 2857 4222 2896
rect 4042 2823 4043 2857
rect 4043 2823 4077 2857
rect 4077 2823 4115 2857
rect 4115 2823 4149 2857
rect 4149 2823 4187 2857
rect 4187 2823 4221 2857
rect 4221 2823 4222 2857
rect 4042 2784 4222 2823
rect 4042 2750 4043 2784
rect 4043 2750 4077 2784
rect 4077 2750 4115 2784
rect 4115 2750 4149 2784
rect 4149 2750 4187 2784
rect 4187 2750 4221 2784
rect 4221 2750 4222 2784
rect 4042 2711 4222 2750
rect 4042 2677 4043 2711
rect 4043 2677 4077 2711
rect 4077 2677 4115 2711
rect 4115 2677 4149 2711
rect 4149 2677 4187 2711
rect 4187 2677 4221 2711
rect 4221 2677 4222 2711
rect 4042 2638 4222 2677
rect 4042 2604 4043 2638
rect 4043 2604 4077 2638
rect 4077 2604 4115 2638
rect 4115 2604 4149 2638
rect 4149 2604 4187 2638
rect 4187 2604 4221 2638
rect 4221 2604 4222 2638
rect 4042 2565 4222 2604
rect 4042 2531 4043 2565
rect 4043 2531 4077 2565
rect 4077 2531 4115 2565
rect 4115 2531 4149 2565
rect 4149 2531 4187 2565
rect 4187 2531 4221 2565
rect 4221 2531 4222 2565
rect 4042 2492 4222 2531
rect 4042 2458 4043 2492
rect 4043 2458 4077 2492
rect 4077 2458 4115 2492
rect 4115 2458 4149 2492
rect 4149 2458 4187 2492
rect 4187 2458 4221 2492
rect 4221 2458 4222 2492
rect 4042 2419 4222 2458
rect 4042 2385 4043 2419
rect 4043 2385 4077 2419
rect 4077 2385 4115 2419
rect 4115 2385 4149 2419
rect 4149 2385 4187 2419
rect 4187 2385 4221 2419
rect 4221 2385 4222 2419
rect 4042 2346 4222 2385
rect 4042 2312 4043 2346
rect 4043 2312 4077 2346
rect 4077 2312 4115 2346
rect 4115 2312 4149 2346
rect 4149 2312 4187 2346
rect 4187 2312 4221 2346
rect 4221 2312 4222 2346
rect 4042 2273 4222 2312
rect 4042 2239 4043 2273
rect 4043 2239 4077 2273
rect 4077 2239 4115 2273
rect 4115 2239 4149 2273
rect 4149 2239 4187 2273
rect 4187 2239 4221 2273
rect 4221 2239 4222 2273
rect 4042 2200 4222 2239
rect 4042 2166 4043 2200
rect 4043 2166 4077 2200
rect 4077 2166 4115 2200
rect 4115 2166 4149 2200
rect 4149 2166 4187 2200
rect 4187 2166 4221 2200
rect 4221 2166 4222 2200
rect 4042 2126 4222 2166
rect 4042 2092 4043 2126
rect 4043 2092 4077 2126
rect 4077 2092 4115 2126
rect 4115 2092 4149 2126
rect 4149 2092 4187 2126
rect 4187 2092 4221 2126
rect 4221 2092 4222 2126
rect 4042 2052 4222 2092
rect 4042 2018 4043 2052
rect 4043 2018 4077 2052
rect 4077 2018 4115 2052
rect 4115 2018 4149 2052
rect 4149 2018 4187 2052
rect 4187 2018 4221 2052
rect 4221 2018 4222 2052
rect 4042 1978 4222 2018
rect 4042 1944 4043 1978
rect 4043 1944 4077 1978
rect 4077 1944 4115 1978
rect 4115 1944 4149 1978
rect 4149 1944 4187 1978
rect 4187 1944 4221 1978
rect 4221 1944 4222 1978
rect 4042 1904 4222 1944
rect 4042 1870 4043 1904
rect 4043 1870 4077 1904
rect 4077 1870 4115 1904
rect 4115 1870 4149 1904
rect 4149 1870 4187 1904
rect 4187 1870 4221 1904
rect 4221 1870 4222 1904
rect 4042 1830 4222 1870
rect 4042 1796 4043 1830
rect 4043 1796 4077 1830
rect 4077 1796 4115 1830
rect 4115 1796 4149 1830
rect 4149 1796 4187 1830
rect 4187 1796 4221 1830
rect 4221 1796 4222 1830
rect 4042 1756 4222 1796
rect 4042 1722 4043 1756
rect 4043 1722 4077 1756
rect 4077 1722 4115 1756
rect 4115 1722 4149 1756
rect 4149 1722 4187 1756
rect 4187 1722 4221 1756
rect 4221 1722 4222 1756
rect 4042 1682 4222 1722
rect 4042 1648 4043 1682
rect 4043 1648 4077 1682
rect 4077 1648 4115 1682
rect 4115 1648 4149 1682
rect 4149 1648 4187 1682
rect 4187 1648 4221 1682
rect 4221 1648 4222 1682
rect 4042 1608 4222 1648
rect 4042 1574 4043 1608
rect 4043 1574 4077 1608
rect 4077 1574 4115 1608
rect 4115 1574 4149 1608
rect 4149 1574 4187 1608
rect 4187 1574 4221 1608
rect 4221 1574 4222 1608
rect 4042 1568 4222 1574
rect 4538 4092 4590 4124
rect 4538 4072 4539 4092
rect 4539 4072 4573 4092
rect 4573 4072 4590 4092
rect 4602 4072 4654 4124
rect 4666 4092 4718 4124
rect 4666 4072 4683 4092
rect 4683 4072 4717 4092
rect 4717 4072 4718 4092
rect 4538 4058 4539 4059
rect 4539 4058 4573 4059
rect 4573 4058 4590 4059
rect 4538 4020 4590 4058
rect 4538 4007 4539 4020
rect 4539 4007 4573 4020
rect 4573 4007 4590 4020
rect 4602 4007 4654 4059
rect 4666 4058 4683 4059
rect 4683 4058 4717 4059
rect 4717 4058 4718 4059
rect 4666 4020 4718 4058
rect 4666 4007 4683 4020
rect 4683 4007 4717 4020
rect 4717 4007 4718 4020
rect 4538 3986 4539 3994
rect 4539 3986 4573 3994
rect 4573 3986 4590 3994
rect 4538 3948 4590 3986
rect 4538 3942 4539 3948
rect 4539 3942 4573 3948
rect 4573 3942 4590 3948
rect 4602 3942 4654 3994
rect 4666 3986 4683 3994
rect 4683 3986 4717 3994
rect 4717 3986 4718 3994
rect 4666 3948 4718 3986
rect 4666 3942 4683 3948
rect 4683 3942 4717 3948
rect 4717 3942 4718 3948
rect 4538 3914 4539 3929
rect 4539 3914 4573 3929
rect 4573 3914 4590 3929
rect 4538 3877 4590 3914
rect 4602 3877 4654 3929
rect 4666 3914 4683 3929
rect 4683 3914 4717 3929
rect 4717 3914 4718 3929
rect 4666 3877 4718 3914
rect 4538 3842 4539 3864
rect 4539 3842 4573 3864
rect 4573 3842 4590 3864
rect 4538 3812 4590 3842
rect 4602 3812 4654 3864
rect 4666 3842 4683 3864
rect 4683 3842 4717 3864
rect 4717 3842 4718 3864
rect 4666 3812 4718 3842
rect 4538 3770 4539 3799
rect 4539 3770 4573 3799
rect 4573 3770 4590 3799
rect 4538 3747 4590 3770
rect 4602 3747 4654 3799
rect 4666 3770 4683 3799
rect 4683 3770 4717 3799
rect 4717 3770 4718 3799
rect 4666 3747 4718 3770
rect 4538 3732 4590 3734
rect 4538 3698 4539 3732
rect 4539 3698 4573 3732
rect 4573 3698 4590 3732
rect 4538 3682 4590 3698
rect 4602 3682 4654 3734
rect 4666 3732 4718 3734
rect 4666 3698 4683 3732
rect 4683 3698 4717 3732
rect 4717 3698 4718 3732
rect 4666 3682 4718 3698
rect 4538 3660 4590 3669
rect 4538 3626 4539 3660
rect 4539 3626 4573 3660
rect 4573 3626 4590 3660
rect 4538 3617 4590 3626
rect 4602 3617 4654 3669
rect 4666 3660 4718 3669
rect 4666 3626 4683 3660
rect 4683 3626 4717 3660
rect 4717 3626 4718 3660
rect 4666 3617 4718 3626
rect 4538 3588 4718 3604
rect 4538 3554 4539 3588
rect 4539 3554 4573 3588
rect 4573 3554 4683 3588
rect 4683 3554 4717 3588
rect 4717 3554 4718 3588
rect 4538 3516 4718 3554
rect 4538 3482 4539 3516
rect 4539 3482 4573 3516
rect 4573 3482 4683 3516
rect 4683 3482 4717 3516
rect 4717 3482 4718 3516
rect 4538 3444 4718 3482
rect 4538 3410 4539 3444
rect 4539 3410 4573 3444
rect 4573 3410 4683 3444
rect 4683 3410 4717 3444
rect 4717 3410 4718 3444
rect 4538 3372 4718 3410
rect 4538 3338 4539 3372
rect 4539 3338 4573 3372
rect 4573 3338 4683 3372
rect 4683 3338 4717 3372
rect 4717 3338 4718 3372
rect 4538 3300 4718 3338
rect 4538 3266 4539 3300
rect 4539 3266 4573 3300
rect 4573 3266 4683 3300
rect 4683 3266 4717 3300
rect 4717 3266 4718 3300
rect 4538 3228 4718 3266
rect 4538 3194 4539 3228
rect 4539 3194 4573 3228
rect 4573 3194 4683 3228
rect 4683 3194 4717 3228
rect 4717 3194 4718 3228
rect 4538 3108 4718 3194
rect 4538 3074 4539 3108
rect 4539 3074 4573 3108
rect 4573 3074 4611 3108
rect 4611 3074 4645 3108
rect 4645 3074 4683 3108
rect 4683 3074 4717 3108
rect 4717 3074 4718 3108
rect 4538 3028 4718 3074
rect 4538 2994 4539 3028
rect 4539 2994 4573 3028
rect 4573 2994 4611 3028
rect 4611 2994 4645 3028
rect 4645 2994 4683 3028
rect 4683 2994 4717 3028
rect 4717 2994 4718 3028
rect 4538 2948 4718 2994
rect 4538 2914 4539 2948
rect 4539 2914 4573 2948
rect 4573 2914 4611 2948
rect 4611 2914 4645 2948
rect 4645 2914 4683 2948
rect 4683 2914 4717 2948
rect 4717 2914 4718 2948
rect 4538 2868 4718 2914
rect 4538 2834 4539 2868
rect 4539 2834 4573 2868
rect 4573 2834 4611 2868
rect 4611 2834 4645 2868
rect 4645 2834 4683 2868
rect 4683 2834 4717 2868
rect 4717 2834 4718 2868
rect 4538 2788 4718 2834
rect 4538 2754 4539 2788
rect 4539 2754 4573 2788
rect 4573 2754 4611 2788
rect 4611 2754 4645 2788
rect 4645 2754 4683 2788
rect 4683 2754 4717 2788
rect 4717 2754 4718 2788
rect 4538 2708 4718 2754
rect 4538 2674 4539 2708
rect 4539 2674 4573 2708
rect 4573 2674 4611 2708
rect 4611 2674 4645 2708
rect 4645 2674 4683 2708
rect 4683 2674 4717 2708
rect 4717 2674 4718 2708
rect 4538 2628 4718 2674
rect 4538 2594 4539 2628
rect 4539 2594 4573 2628
rect 4573 2594 4611 2628
rect 4611 2594 4645 2628
rect 4645 2594 4683 2628
rect 4683 2594 4717 2628
rect 4717 2594 4718 2628
rect 4538 2518 4718 2594
rect 4538 2484 4539 2518
rect 4539 2484 4573 2518
rect 4573 2484 4683 2518
rect 4683 2484 4717 2518
rect 4717 2484 4718 2518
rect 4538 2446 4718 2484
rect 4538 2412 4539 2446
rect 4539 2412 4573 2446
rect 4573 2412 4683 2446
rect 4683 2412 4717 2446
rect 4717 2412 4718 2446
rect 4538 2374 4718 2412
rect 4538 2340 4539 2374
rect 4539 2340 4573 2374
rect 4573 2340 4683 2374
rect 4683 2340 4717 2374
rect 4717 2340 4718 2374
rect 4538 2302 4718 2340
rect 4538 2268 4539 2302
rect 4539 2268 4573 2302
rect 4573 2268 4683 2302
rect 4683 2268 4717 2302
rect 4717 2268 4718 2302
rect 4538 2230 4718 2268
rect 4538 2196 4539 2230
rect 4539 2196 4573 2230
rect 4573 2196 4683 2230
rect 4683 2196 4717 2230
rect 4717 2196 4718 2230
rect 4538 2158 4718 2196
rect 4538 2124 4539 2158
rect 4539 2124 4573 2158
rect 4573 2124 4683 2158
rect 4683 2124 4717 2158
rect 4717 2124 4718 2158
rect 4538 2086 4718 2124
rect 4538 2052 4539 2086
rect 4539 2052 4573 2086
rect 4573 2052 4683 2086
rect 4683 2052 4717 2086
rect 4717 2052 4718 2086
rect 4538 2014 4718 2052
rect 4538 1980 4539 2014
rect 4539 1980 4573 2014
rect 4573 1980 4683 2014
rect 4683 1980 4717 2014
rect 4717 1980 4718 2014
rect 4538 1942 4718 1980
rect 4538 1908 4539 1942
rect 4539 1908 4573 1942
rect 4573 1908 4683 1942
rect 4683 1908 4717 1942
rect 4717 1908 4718 1942
rect 4538 1870 4718 1908
rect 4538 1836 4539 1870
rect 4539 1836 4573 1870
rect 4573 1836 4683 1870
rect 4683 1836 4717 1870
rect 4717 1836 4718 1870
rect 4538 1798 4718 1836
rect 4538 1764 4539 1798
rect 4539 1764 4573 1798
rect 4573 1764 4683 1798
rect 4683 1764 4717 1798
rect 4717 1764 4718 1798
rect 4538 1726 4718 1764
rect 4538 1692 4539 1726
rect 4539 1692 4573 1726
rect 4573 1692 4683 1726
rect 4683 1692 4717 1726
rect 4717 1692 4718 1726
rect 4538 1654 4718 1692
rect 4538 1620 4539 1654
rect 4539 1620 4573 1654
rect 4573 1620 4683 1654
rect 4683 1620 4717 1654
rect 4717 1620 4718 1654
rect 4538 1568 4718 1620
rect 5034 4098 5086 4119
rect 5034 4067 5035 4098
rect 5035 4067 5069 4098
rect 5069 4067 5086 4098
rect 5098 4098 5150 4119
rect 5098 4067 5107 4098
rect 5107 4067 5141 4098
rect 5141 4067 5150 4098
rect 5162 4098 5214 4119
rect 5162 4067 5179 4098
rect 5179 4067 5213 4098
rect 5213 4067 5214 4098
rect 5034 4025 5086 4054
rect 5034 4002 5035 4025
rect 5035 4002 5069 4025
rect 5069 4002 5086 4025
rect 5098 4025 5150 4054
rect 5098 4002 5107 4025
rect 5107 4002 5141 4025
rect 5141 4002 5150 4025
rect 5162 4025 5214 4054
rect 5162 4002 5179 4025
rect 5179 4002 5213 4025
rect 5213 4002 5214 4025
rect 5034 3952 5086 3989
rect 5034 3937 5035 3952
rect 5035 3937 5069 3952
rect 5069 3937 5086 3952
rect 5098 3952 5150 3989
rect 5098 3937 5107 3952
rect 5107 3937 5141 3952
rect 5141 3937 5150 3952
rect 5162 3952 5214 3989
rect 5162 3937 5179 3952
rect 5179 3937 5213 3952
rect 5213 3937 5214 3952
rect 5034 3918 5035 3924
rect 5035 3918 5069 3924
rect 5069 3918 5107 3924
rect 5107 3918 5141 3924
rect 5141 3918 5179 3924
rect 5179 3918 5213 3924
rect 5213 3918 5214 3924
rect 5034 3879 5214 3918
rect 5034 3845 5035 3879
rect 5035 3845 5069 3879
rect 5069 3845 5107 3879
rect 5107 3845 5141 3879
rect 5141 3845 5179 3879
rect 5179 3845 5213 3879
rect 5213 3845 5214 3879
rect 5034 3806 5214 3845
rect 5034 3772 5035 3806
rect 5035 3772 5069 3806
rect 5069 3772 5107 3806
rect 5107 3772 5141 3806
rect 5141 3772 5179 3806
rect 5179 3772 5213 3806
rect 5213 3772 5214 3806
rect 5034 3733 5214 3772
rect 5034 3699 5035 3733
rect 5035 3699 5069 3733
rect 5069 3699 5107 3733
rect 5107 3699 5141 3733
rect 5141 3699 5179 3733
rect 5179 3699 5213 3733
rect 5213 3699 5214 3733
rect 5034 3660 5214 3699
rect 5034 3626 5035 3660
rect 5035 3626 5069 3660
rect 5069 3626 5107 3660
rect 5107 3626 5141 3660
rect 5141 3626 5179 3660
rect 5179 3626 5213 3660
rect 5213 3626 5214 3660
rect 5034 3587 5214 3626
rect 5034 3553 5035 3587
rect 5035 3553 5069 3587
rect 5069 3553 5107 3587
rect 5107 3553 5141 3587
rect 5141 3553 5179 3587
rect 5179 3553 5213 3587
rect 5213 3553 5214 3587
rect 5034 3514 5214 3553
rect 5034 3480 5035 3514
rect 5035 3480 5069 3514
rect 5069 3480 5107 3514
rect 5107 3480 5141 3514
rect 5141 3480 5179 3514
rect 5179 3480 5213 3514
rect 5213 3480 5214 3514
rect 5034 3441 5214 3480
rect 5034 3407 5035 3441
rect 5035 3407 5069 3441
rect 5069 3407 5107 3441
rect 5107 3407 5141 3441
rect 5141 3407 5179 3441
rect 5179 3407 5213 3441
rect 5213 3407 5214 3441
rect 5034 3368 5214 3407
rect 5034 3334 5035 3368
rect 5035 3334 5069 3368
rect 5069 3334 5107 3368
rect 5107 3334 5141 3368
rect 5141 3334 5179 3368
rect 5179 3334 5213 3368
rect 5213 3334 5214 3368
rect 5034 3295 5214 3334
rect 5034 3261 5035 3295
rect 5035 3261 5069 3295
rect 5069 3261 5107 3295
rect 5107 3261 5141 3295
rect 5141 3261 5179 3295
rect 5179 3261 5213 3295
rect 5213 3261 5214 3295
rect 5034 3222 5214 3261
rect 5034 3188 5035 3222
rect 5035 3188 5069 3222
rect 5069 3188 5107 3222
rect 5107 3188 5141 3222
rect 5141 3188 5179 3222
rect 5179 3188 5213 3222
rect 5213 3188 5214 3222
rect 5034 3149 5214 3188
rect 5034 3115 5035 3149
rect 5035 3115 5069 3149
rect 5069 3115 5107 3149
rect 5107 3115 5141 3149
rect 5141 3115 5179 3149
rect 5179 3115 5213 3149
rect 5213 3115 5214 3149
rect 5034 3076 5214 3115
rect 5034 3042 5035 3076
rect 5035 3042 5069 3076
rect 5069 3042 5107 3076
rect 5107 3042 5141 3076
rect 5141 3042 5179 3076
rect 5179 3042 5213 3076
rect 5213 3042 5214 3076
rect 5034 3003 5214 3042
rect 5034 2969 5035 3003
rect 5035 2969 5069 3003
rect 5069 2969 5107 3003
rect 5107 2969 5141 3003
rect 5141 2969 5179 3003
rect 5179 2969 5213 3003
rect 5213 2969 5214 3003
rect 5034 2930 5214 2969
rect 5034 2896 5035 2930
rect 5035 2896 5069 2930
rect 5069 2896 5107 2930
rect 5107 2896 5141 2930
rect 5141 2896 5179 2930
rect 5179 2896 5213 2930
rect 5213 2896 5214 2930
rect 5034 2857 5214 2896
rect 5034 2823 5035 2857
rect 5035 2823 5069 2857
rect 5069 2823 5107 2857
rect 5107 2823 5141 2857
rect 5141 2823 5179 2857
rect 5179 2823 5213 2857
rect 5213 2823 5214 2857
rect 5034 2784 5214 2823
rect 5034 2750 5035 2784
rect 5035 2750 5069 2784
rect 5069 2750 5107 2784
rect 5107 2750 5141 2784
rect 5141 2750 5179 2784
rect 5179 2750 5213 2784
rect 5213 2750 5214 2784
rect 5034 2711 5214 2750
rect 5034 2677 5035 2711
rect 5035 2677 5069 2711
rect 5069 2677 5107 2711
rect 5107 2677 5141 2711
rect 5141 2677 5179 2711
rect 5179 2677 5213 2711
rect 5213 2677 5214 2711
rect 5034 2638 5214 2677
rect 5034 2604 5035 2638
rect 5035 2604 5069 2638
rect 5069 2604 5107 2638
rect 5107 2604 5141 2638
rect 5141 2604 5179 2638
rect 5179 2604 5213 2638
rect 5213 2604 5214 2638
rect 5034 2565 5214 2604
rect 5034 2531 5035 2565
rect 5035 2531 5069 2565
rect 5069 2531 5107 2565
rect 5107 2531 5141 2565
rect 5141 2531 5179 2565
rect 5179 2531 5213 2565
rect 5213 2531 5214 2565
rect 5034 2492 5214 2531
rect 5034 2458 5035 2492
rect 5035 2458 5069 2492
rect 5069 2458 5107 2492
rect 5107 2458 5141 2492
rect 5141 2458 5179 2492
rect 5179 2458 5213 2492
rect 5213 2458 5214 2492
rect 5034 2419 5214 2458
rect 5034 2385 5035 2419
rect 5035 2385 5069 2419
rect 5069 2385 5107 2419
rect 5107 2385 5141 2419
rect 5141 2385 5179 2419
rect 5179 2385 5213 2419
rect 5213 2385 5214 2419
rect 5034 2346 5214 2385
rect 5034 2312 5035 2346
rect 5035 2312 5069 2346
rect 5069 2312 5107 2346
rect 5107 2312 5141 2346
rect 5141 2312 5179 2346
rect 5179 2312 5213 2346
rect 5213 2312 5214 2346
rect 5034 2273 5214 2312
rect 5034 2239 5035 2273
rect 5035 2239 5069 2273
rect 5069 2239 5107 2273
rect 5107 2239 5141 2273
rect 5141 2239 5179 2273
rect 5179 2239 5213 2273
rect 5213 2239 5214 2273
rect 5034 2200 5214 2239
rect 5034 2166 5035 2200
rect 5035 2166 5069 2200
rect 5069 2166 5107 2200
rect 5107 2166 5141 2200
rect 5141 2166 5179 2200
rect 5179 2166 5213 2200
rect 5213 2166 5214 2200
rect 5034 2126 5214 2166
rect 5034 2092 5035 2126
rect 5035 2092 5069 2126
rect 5069 2092 5107 2126
rect 5107 2092 5141 2126
rect 5141 2092 5179 2126
rect 5179 2092 5213 2126
rect 5213 2092 5214 2126
rect 5034 2052 5214 2092
rect 5034 2018 5035 2052
rect 5035 2018 5069 2052
rect 5069 2018 5107 2052
rect 5107 2018 5141 2052
rect 5141 2018 5179 2052
rect 5179 2018 5213 2052
rect 5213 2018 5214 2052
rect 5034 1978 5214 2018
rect 5034 1944 5035 1978
rect 5035 1944 5069 1978
rect 5069 1944 5107 1978
rect 5107 1944 5141 1978
rect 5141 1944 5179 1978
rect 5179 1944 5213 1978
rect 5213 1944 5214 1978
rect 5034 1904 5214 1944
rect 5034 1870 5035 1904
rect 5035 1870 5069 1904
rect 5069 1870 5107 1904
rect 5107 1870 5141 1904
rect 5141 1870 5179 1904
rect 5179 1870 5213 1904
rect 5213 1870 5214 1904
rect 5034 1830 5214 1870
rect 5034 1796 5035 1830
rect 5035 1796 5069 1830
rect 5069 1796 5107 1830
rect 5107 1796 5141 1830
rect 5141 1796 5179 1830
rect 5179 1796 5213 1830
rect 5213 1796 5214 1830
rect 5034 1756 5214 1796
rect 5034 1722 5035 1756
rect 5035 1722 5069 1756
rect 5069 1722 5107 1756
rect 5107 1722 5141 1756
rect 5141 1722 5179 1756
rect 5179 1722 5213 1756
rect 5213 1722 5214 1756
rect 5034 1682 5214 1722
rect 5034 1648 5035 1682
rect 5035 1648 5069 1682
rect 5069 1648 5107 1682
rect 5107 1648 5141 1682
rect 5141 1648 5179 1682
rect 5179 1648 5213 1682
rect 5213 1648 5214 1682
rect 5034 1608 5214 1648
rect 5034 1574 5035 1608
rect 5035 1574 5069 1608
rect 5069 1574 5107 1608
rect 5107 1574 5141 1608
rect 5141 1574 5179 1608
rect 5179 1574 5213 1608
rect 5213 1574 5214 1608
rect 5034 1568 5214 1574
rect 5530 4092 5582 4124
rect 5530 4072 5531 4092
rect 5531 4072 5565 4092
rect 5565 4072 5582 4092
rect 5594 4072 5646 4124
rect 5658 4092 5710 4124
rect 5658 4072 5675 4092
rect 5675 4072 5709 4092
rect 5709 4072 5710 4092
rect 5530 4058 5531 4059
rect 5531 4058 5565 4059
rect 5565 4058 5582 4059
rect 5530 4020 5582 4058
rect 5530 4007 5531 4020
rect 5531 4007 5565 4020
rect 5565 4007 5582 4020
rect 5594 4007 5646 4059
rect 5658 4058 5675 4059
rect 5675 4058 5709 4059
rect 5709 4058 5710 4059
rect 5658 4020 5710 4058
rect 5658 4007 5675 4020
rect 5675 4007 5709 4020
rect 5709 4007 5710 4020
rect 5530 3986 5531 3994
rect 5531 3986 5565 3994
rect 5565 3986 5582 3994
rect 5530 3948 5582 3986
rect 5530 3942 5531 3948
rect 5531 3942 5565 3948
rect 5565 3942 5582 3948
rect 5594 3942 5646 3994
rect 5658 3986 5675 3994
rect 5675 3986 5709 3994
rect 5709 3986 5710 3994
rect 5658 3948 5710 3986
rect 5658 3942 5675 3948
rect 5675 3942 5709 3948
rect 5709 3942 5710 3948
rect 5530 3914 5531 3929
rect 5531 3914 5565 3929
rect 5565 3914 5582 3929
rect 5530 3877 5582 3914
rect 5594 3877 5646 3929
rect 5658 3914 5675 3929
rect 5675 3914 5709 3929
rect 5709 3914 5710 3929
rect 5658 3877 5710 3914
rect 5530 3842 5531 3864
rect 5531 3842 5565 3864
rect 5565 3842 5582 3864
rect 5530 3812 5582 3842
rect 5594 3812 5646 3864
rect 5658 3842 5675 3864
rect 5675 3842 5709 3864
rect 5709 3842 5710 3864
rect 5658 3812 5710 3842
rect 5530 3770 5531 3799
rect 5531 3770 5565 3799
rect 5565 3770 5582 3799
rect 5530 3747 5582 3770
rect 5594 3747 5646 3799
rect 5658 3770 5675 3799
rect 5675 3770 5709 3799
rect 5709 3770 5710 3799
rect 5658 3747 5710 3770
rect 5530 3732 5582 3734
rect 5530 3698 5531 3732
rect 5531 3698 5565 3732
rect 5565 3698 5582 3732
rect 5530 3682 5582 3698
rect 5594 3682 5646 3734
rect 5658 3732 5710 3734
rect 5658 3698 5675 3732
rect 5675 3698 5709 3732
rect 5709 3698 5710 3732
rect 5658 3682 5710 3698
rect 5530 3660 5582 3669
rect 5530 3626 5531 3660
rect 5531 3626 5565 3660
rect 5565 3626 5582 3660
rect 5530 3617 5582 3626
rect 5594 3617 5646 3669
rect 5658 3660 5710 3669
rect 5658 3626 5675 3660
rect 5675 3626 5709 3660
rect 5709 3626 5710 3660
rect 5658 3617 5710 3626
rect 5530 3588 5710 3604
rect 5530 3554 5531 3588
rect 5531 3554 5565 3588
rect 5565 3554 5675 3588
rect 5675 3554 5709 3588
rect 5709 3554 5710 3588
rect 5530 3516 5710 3554
rect 5530 3482 5531 3516
rect 5531 3482 5565 3516
rect 5565 3482 5675 3516
rect 5675 3482 5709 3516
rect 5709 3482 5710 3516
rect 5530 3444 5710 3482
rect 5530 3410 5531 3444
rect 5531 3410 5565 3444
rect 5565 3410 5675 3444
rect 5675 3410 5709 3444
rect 5709 3410 5710 3444
rect 5530 3372 5710 3410
rect 5530 3338 5531 3372
rect 5531 3338 5565 3372
rect 5565 3338 5675 3372
rect 5675 3338 5709 3372
rect 5709 3338 5710 3372
rect 5530 3300 5710 3338
rect 5530 3266 5531 3300
rect 5531 3266 5565 3300
rect 5565 3266 5675 3300
rect 5675 3266 5709 3300
rect 5709 3266 5710 3300
rect 5530 3228 5710 3266
rect 5530 3194 5531 3228
rect 5531 3194 5565 3228
rect 5565 3194 5675 3228
rect 5675 3194 5709 3228
rect 5709 3194 5710 3228
rect 5530 3108 5710 3194
rect 5530 3074 5531 3108
rect 5531 3074 5565 3108
rect 5565 3074 5603 3108
rect 5603 3074 5637 3108
rect 5637 3074 5675 3108
rect 5675 3074 5709 3108
rect 5709 3074 5710 3108
rect 5530 3028 5710 3074
rect 5530 2994 5531 3028
rect 5531 2994 5565 3028
rect 5565 2994 5603 3028
rect 5603 2994 5637 3028
rect 5637 2994 5675 3028
rect 5675 2994 5709 3028
rect 5709 2994 5710 3028
rect 5530 2948 5710 2994
rect 5530 2914 5531 2948
rect 5531 2914 5565 2948
rect 5565 2914 5603 2948
rect 5603 2914 5637 2948
rect 5637 2914 5675 2948
rect 5675 2914 5709 2948
rect 5709 2914 5710 2948
rect 5530 2868 5710 2914
rect 5530 2834 5531 2868
rect 5531 2834 5565 2868
rect 5565 2834 5603 2868
rect 5603 2834 5637 2868
rect 5637 2834 5675 2868
rect 5675 2834 5709 2868
rect 5709 2834 5710 2868
rect 5530 2788 5710 2834
rect 5530 2754 5531 2788
rect 5531 2754 5565 2788
rect 5565 2754 5603 2788
rect 5603 2754 5637 2788
rect 5637 2754 5675 2788
rect 5675 2754 5709 2788
rect 5709 2754 5710 2788
rect 5530 2708 5710 2754
rect 5530 2674 5531 2708
rect 5531 2674 5565 2708
rect 5565 2674 5603 2708
rect 5603 2674 5637 2708
rect 5637 2674 5675 2708
rect 5675 2674 5709 2708
rect 5709 2674 5710 2708
rect 5530 2628 5710 2674
rect 5530 2594 5531 2628
rect 5531 2594 5565 2628
rect 5565 2594 5603 2628
rect 5603 2594 5637 2628
rect 5637 2594 5675 2628
rect 5675 2594 5709 2628
rect 5709 2594 5710 2628
rect 5530 2518 5710 2594
rect 5530 2484 5531 2518
rect 5531 2484 5565 2518
rect 5565 2484 5675 2518
rect 5675 2484 5709 2518
rect 5709 2484 5710 2518
rect 5530 2446 5710 2484
rect 5530 2412 5531 2446
rect 5531 2412 5565 2446
rect 5565 2412 5675 2446
rect 5675 2412 5709 2446
rect 5709 2412 5710 2446
rect 5530 2374 5710 2412
rect 5530 2340 5531 2374
rect 5531 2340 5565 2374
rect 5565 2340 5675 2374
rect 5675 2340 5709 2374
rect 5709 2340 5710 2374
rect 5530 2302 5710 2340
rect 5530 2268 5531 2302
rect 5531 2268 5565 2302
rect 5565 2268 5675 2302
rect 5675 2268 5709 2302
rect 5709 2268 5710 2302
rect 5530 2230 5710 2268
rect 5530 2196 5531 2230
rect 5531 2196 5565 2230
rect 5565 2196 5675 2230
rect 5675 2196 5709 2230
rect 5709 2196 5710 2230
rect 5530 2158 5710 2196
rect 5530 2124 5531 2158
rect 5531 2124 5565 2158
rect 5565 2124 5675 2158
rect 5675 2124 5709 2158
rect 5709 2124 5710 2158
rect 5530 2086 5710 2124
rect 5530 2052 5531 2086
rect 5531 2052 5565 2086
rect 5565 2052 5675 2086
rect 5675 2052 5709 2086
rect 5709 2052 5710 2086
rect 5530 2014 5710 2052
rect 5530 1980 5531 2014
rect 5531 1980 5565 2014
rect 5565 1980 5675 2014
rect 5675 1980 5709 2014
rect 5709 1980 5710 2014
rect 5530 1942 5710 1980
rect 5530 1908 5531 1942
rect 5531 1908 5565 1942
rect 5565 1908 5675 1942
rect 5675 1908 5709 1942
rect 5709 1908 5710 1942
rect 5530 1870 5710 1908
rect 5530 1836 5531 1870
rect 5531 1836 5565 1870
rect 5565 1836 5675 1870
rect 5675 1836 5709 1870
rect 5709 1836 5710 1870
rect 5530 1798 5710 1836
rect 5530 1764 5531 1798
rect 5531 1764 5565 1798
rect 5565 1764 5675 1798
rect 5675 1764 5709 1798
rect 5709 1764 5710 1798
rect 5530 1726 5710 1764
rect 5530 1692 5531 1726
rect 5531 1692 5565 1726
rect 5565 1692 5675 1726
rect 5675 1692 5709 1726
rect 5709 1692 5710 1726
rect 5530 1654 5710 1692
rect 5530 1620 5531 1654
rect 5531 1620 5565 1654
rect 5565 1620 5675 1654
rect 5675 1620 5709 1654
rect 5709 1620 5710 1654
rect 5530 1568 5710 1620
rect 6026 4098 6078 4119
rect 6026 4067 6027 4098
rect 6027 4067 6061 4098
rect 6061 4067 6078 4098
rect 6090 4098 6142 4119
rect 6090 4067 6099 4098
rect 6099 4067 6133 4098
rect 6133 4067 6142 4098
rect 6154 4098 6206 4119
rect 6154 4067 6171 4098
rect 6171 4067 6205 4098
rect 6205 4067 6206 4098
rect 6026 4025 6078 4054
rect 6026 4002 6027 4025
rect 6027 4002 6061 4025
rect 6061 4002 6078 4025
rect 6090 4025 6142 4054
rect 6090 4002 6099 4025
rect 6099 4002 6133 4025
rect 6133 4002 6142 4025
rect 6154 4025 6206 4054
rect 6154 4002 6171 4025
rect 6171 4002 6205 4025
rect 6205 4002 6206 4025
rect 6026 3952 6078 3989
rect 6026 3937 6027 3952
rect 6027 3937 6061 3952
rect 6061 3937 6078 3952
rect 6090 3952 6142 3989
rect 6090 3937 6099 3952
rect 6099 3937 6133 3952
rect 6133 3937 6142 3952
rect 6154 3952 6206 3989
rect 6154 3937 6171 3952
rect 6171 3937 6205 3952
rect 6205 3937 6206 3952
rect 6026 3918 6027 3924
rect 6027 3918 6061 3924
rect 6061 3918 6099 3924
rect 6099 3918 6133 3924
rect 6133 3918 6171 3924
rect 6171 3918 6205 3924
rect 6205 3918 6206 3924
rect 6026 3879 6206 3918
rect 6026 3845 6027 3879
rect 6027 3845 6061 3879
rect 6061 3845 6099 3879
rect 6099 3845 6133 3879
rect 6133 3845 6171 3879
rect 6171 3845 6205 3879
rect 6205 3845 6206 3879
rect 6026 3806 6206 3845
rect 6026 3772 6027 3806
rect 6027 3772 6061 3806
rect 6061 3772 6099 3806
rect 6099 3772 6133 3806
rect 6133 3772 6171 3806
rect 6171 3772 6205 3806
rect 6205 3772 6206 3806
rect 6026 3733 6206 3772
rect 6026 3699 6027 3733
rect 6027 3699 6061 3733
rect 6061 3699 6099 3733
rect 6099 3699 6133 3733
rect 6133 3699 6171 3733
rect 6171 3699 6205 3733
rect 6205 3699 6206 3733
rect 6026 3660 6206 3699
rect 6026 3626 6027 3660
rect 6027 3626 6061 3660
rect 6061 3626 6099 3660
rect 6099 3626 6133 3660
rect 6133 3626 6171 3660
rect 6171 3626 6205 3660
rect 6205 3626 6206 3660
rect 6026 3587 6206 3626
rect 6026 3553 6027 3587
rect 6027 3553 6061 3587
rect 6061 3553 6099 3587
rect 6099 3553 6133 3587
rect 6133 3553 6171 3587
rect 6171 3553 6205 3587
rect 6205 3553 6206 3587
rect 6026 3514 6206 3553
rect 6026 3480 6027 3514
rect 6027 3480 6061 3514
rect 6061 3480 6099 3514
rect 6099 3480 6133 3514
rect 6133 3480 6171 3514
rect 6171 3480 6205 3514
rect 6205 3480 6206 3514
rect 6026 3441 6206 3480
rect 6026 3407 6027 3441
rect 6027 3407 6061 3441
rect 6061 3407 6099 3441
rect 6099 3407 6133 3441
rect 6133 3407 6171 3441
rect 6171 3407 6205 3441
rect 6205 3407 6206 3441
rect 6026 3368 6206 3407
rect 6026 3334 6027 3368
rect 6027 3334 6061 3368
rect 6061 3334 6099 3368
rect 6099 3334 6133 3368
rect 6133 3334 6171 3368
rect 6171 3334 6205 3368
rect 6205 3334 6206 3368
rect 6026 3295 6206 3334
rect 6026 3261 6027 3295
rect 6027 3261 6061 3295
rect 6061 3261 6099 3295
rect 6099 3261 6133 3295
rect 6133 3261 6171 3295
rect 6171 3261 6205 3295
rect 6205 3261 6206 3295
rect 6026 3222 6206 3261
rect 6026 3188 6027 3222
rect 6027 3188 6061 3222
rect 6061 3188 6099 3222
rect 6099 3188 6133 3222
rect 6133 3188 6171 3222
rect 6171 3188 6205 3222
rect 6205 3188 6206 3222
rect 6026 3149 6206 3188
rect 6026 3115 6027 3149
rect 6027 3115 6061 3149
rect 6061 3115 6099 3149
rect 6099 3115 6133 3149
rect 6133 3115 6171 3149
rect 6171 3115 6205 3149
rect 6205 3115 6206 3149
rect 6026 3076 6206 3115
rect 6026 3042 6027 3076
rect 6027 3042 6061 3076
rect 6061 3042 6099 3076
rect 6099 3042 6133 3076
rect 6133 3042 6171 3076
rect 6171 3042 6205 3076
rect 6205 3042 6206 3076
rect 6026 3003 6206 3042
rect 6026 2969 6027 3003
rect 6027 2969 6061 3003
rect 6061 2969 6099 3003
rect 6099 2969 6133 3003
rect 6133 2969 6171 3003
rect 6171 2969 6205 3003
rect 6205 2969 6206 3003
rect 6026 2930 6206 2969
rect 6026 2896 6027 2930
rect 6027 2896 6061 2930
rect 6061 2896 6099 2930
rect 6099 2896 6133 2930
rect 6133 2896 6171 2930
rect 6171 2896 6205 2930
rect 6205 2896 6206 2930
rect 6026 2857 6206 2896
rect 6026 2823 6027 2857
rect 6027 2823 6061 2857
rect 6061 2823 6099 2857
rect 6099 2823 6133 2857
rect 6133 2823 6171 2857
rect 6171 2823 6205 2857
rect 6205 2823 6206 2857
rect 6026 2784 6206 2823
rect 6026 2750 6027 2784
rect 6027 2750 6061 2784
rect 6061 2750 6099 2784
rect 6099 2750 6133 2784
rect 6133 2750 6171 2784
rect 6171 2750 6205 2784
rect 6205 2750 6206 2784
rect 6026 2711 6206 2750
rect 6026 2677 6027 2711
rect 6027 2677 6061 2711
rect 6061 2677 6099 2711
rect 6099 2677 6133 2711
rect 6133 2677 6171 2711
rect 6171 2677 6205 2711
rect 6205 2677 6206 2711
rect 6026 2638 6206 2677
rect 6026 2604 6027 2638
rect 6027 2604 6061 2638
rect 6061 2604 6099 2638
rect 6099 2604 6133 2638
rect 6133 2604 6171 2638
rect 6171 2604 6205 2638
rect 6205 2604 6206 2638
rect 6026 2565 6206 2604
rect 6026 2531 6027 2565
rect 6027 2531 6061 2565
rect 6061 2531 6099 2565
rect 6099 2531 6133 2565
rect 6133 2531 6171 2565
rect 6171 2531 6205 2565
rect 6205 2531 6206 2565
rect 6026 2492 6206 2531
rect 6026 2458 6027 2492
rect 6027 2458 6061 2492
rect 6061 2458 6099 2492
rect 6099 2458 6133 2492
rect 6133 2458 6171 2492
rect 6171 2458 6205 2492
rect 6205 2458 6206 2492
rect 6026 2419 6206 2458
rect 6026 2385 6027 2419
rect 6027 2385 6061 2419
rect 6061 2385 6099 2419
rect 6099 2385 6133 2419
rect 6133 2385 6171 2419
rect 6171 2385 6205 2419
rect 6205 2385 6206 2419
rect 6026 2346 6206 2385
rect 6026 2312 6027 2346
rect 6027 2312 6061 2346
rect 6061 2312 6099 2346
rect 6099 2312 6133 2346
rect 6133 2312 6171 2346
rect 6171 2312 6205 2346
rect 6205 2312 6206 2346
rect 6026 2273 6206 2312
rect 6026 2239 6027 2273
rect 6027 2239 6061 2273
rect 6061 2239 6099 2273
rect 6099 2239 6133 2273
rect 6133 2239 6171 2273
rect 6171 2239 6205 2273
rect 6205 2239 6206 2273
rect 6026 2200 6206 2239
rect 6026 2166 6027 2200
rect 6027 2166 6061 2200
rect 6061 2166 6099 2200
rect 6099 2166 6133 2200
rect 6133 2166 6171 2200
rect 6171 2166 6205 2200
rect 6205 2166 6206 2200
rect 6026 2126 6206 2166
rect 6026 2092 6027 2126
rect 6027 2092 6061 2126
rect 6061 2092 6099 2126
rect 6099 2092 6133 2126
rect 6133 2092 6171 2126
rect 6171 2092 6205 2126
rect 6205 2092 6206 2126
rect 6026 2052 6206 2092
rect 6026 2018 6027 2052
rect 6027 2018 6061 2052
rect 6061 2018 6099 2052
rect 6099 2018 6133 2052
rect 6133 2018 6171 2052
rect 6171 2018 6205 2052
rect 6205 2018 6206 2052
rect 6026 1978 6206 2018
rect 6026 1944 6027 1978
rect 6027 1944 6061 1978
rect 6061 1944 6099 1978
rect 6099 1944 6133 1978
rect 6133 1944 6171 1978
rect 6171 1944 6205 1978
rect 6205 1944 6206 1978
rect 6026 1904 6206 1944
rect 6026 1870 6027 1904
rect 6027 1870 6061 1904
rect 6061 1870 6099 1904
rect 6099 1870 6133 1904
rect 6133 1870 6171 1904
rect 6171 1870 6205 1904
rect 6205 1870 6206 1904
rect 6026 1830 6206 1870
rect 6026 1796 6027 1830
rect 6027 1796 6061 1830
rect 6061 1796 6099 1830
rect 6099 1796 6133 1830
rect 6133 1796 6171 1830
rect 6171 1796 6205 1830
rect 6205 1796 6206 1830
rect 6026 1756 6206 1796
rect 6026 1722 6027 1756
rect 6027 1722 6061 1756
rect 6061 1722 6099 1756
rect 6099 1722 6133 1756
rect 6133 1722 6171 1756
rect 6171 1722 6205 1756
rect 6205 1722 6206 1756
rect 6026 1682 6206 1722
rect 6026 1648 6027 1682
rect 6027 1648 6061 1682
rect 6061 1648 6099 1682
rect 6099 1648 6133 1682
rect 6133 1648 6171 1682
rect 6171 1648 6205 1682
rect 6205 1648 6206 1682
rect 6026 1608 6206 1648
rect 6026 1574 6027 1608
rect 6027 1574 6061 1608
rect 6061 1574 6099 1608
rect 6099 1574 6133 1608
rect 6133 1574 6171 1608
rect 6171 1574 6205 1608
rect 6205 1574 6206 1608
rect 6026 1568 6206 1574
rect 6522 4092 6574 4124
rect 6522 4072 6523 4092
rect 6523 4072 6557 4092
rect 6557 4072 6574 4092
rect 6586 4072 6638 4124
rect 6650 4092 6702 4124
rect 6650 4072 6667 4092
rect 6667 4072 6701 4092
rect 6701 4072 6702 4092
rect 6522 4058 6523 4059
rect 6523 4058 6557 4059
rect 6557 4058 6574 4059
rect 6522 4020 6574 4058
rect 6522 4007 6523 4020
rect 6523 4007 6557 4020
rect 6557 4007 6574 4020
rect 6586 4007 6638 4059
rect 6650 4058 6667 4059
rect 6667 4058 6701 4059
rect 6701 4058 6702 4059
rect 6650 4020 6702 4058
rect 6650 4007 6667 4020
rect 6667 4007 6701 4020
rect 6701 4007 6702 4020
rect 6522 3986 6523 3994
rect 6523 3986 6557 3994
rect 6557 3986 6574 3994
rect 6522 3948 6574 3986
rect 6522 3942 6523 3948
rect 6523 3942 6557 3948
rect 6557 3942 6574 3948
rect 6586 3942 6638 3994
rect 6650 3986 6667 3994
rect 6667 3986 6701 3994
rect 6701 3986 6702 3994
rect 6650 3948 6702 3986
rect 6650 3942 6667 3948
rect 6667 3942 6701 3948
rect 6701 3942 6702 3948
rect 6522 3914 6523 3929
rect 6523 3914 6557 3929
rect 6557 3914 6574 3929
rect 6522 3877 6574 3914
rect 6586 3877 6638 3929
rect 6650 3914 6667 3929
rect 6667 3914 6701 3929
rect 6701 3914 6702 3929
rect 6650 3877 6702 3914
rect 6522 3842 6523 3864
rect 6523 3842 6557 3864
rect 6557 3842 6574 3864
rect 6522 3812 6574 3842
rect 6586 3812 6638 3864
rect 6650 3842 6667 3864
rect 6667 3842 6701 3864
rect 6701 3842 6702 3864
rect 6650 3812 6702 3842
rect 6522 3770 6523 3799
rect 6523 3770 6557 3799
rect 6557 3770 6574 3799
rect 6522 3747 6574 3770
rect 6586 3747 6638 3799
rect 6650 3770 6667 3799
rect 6667 3770 6701 3799
rect 6701 3770 6702 3799
rect 6650 3747 6702 3770
rect 6522 3732 6574 3734
rect 6522 3698 6523 3732
rect 6523 3698 6557 3732
rect 6557 3698 6574 3732
rect 6522 3682 6574 3698
rect 6586 3682 6638 3734
rect 6650 3732 6702 3734
rect 6650 3698 6667 3732
rect 6667 3698 6701 3732
rect 6701 3698 6702 3732
rect 6650 3682 6702 3698
rect 6522 3660 6574 3669
rect 6522 3626 6523 3660
rect 6523 3626 6557 3660
rect 6557 3626 6574 3660
rect 6522 3617 6574 3626
rect 6586 3617 6638 3669
rect 6650 3660 6702 3669
rect 6650 3626 6667 3660
rect 6667 3626 6701 3660
rect 6701 3626 6702 3660
rect 6650 3617 6702 3626
rect 6522 3588 6702 3604
rect 6522 3554 6523 3588
rect 6523 3554 6557 3588
rect 6557 3554 6667 3588
rect 6667 3554 6701 3588
rect 6701 3554 6702 3588
rect 6522 3516 6702 3554
rect 6522 3482 6523 3516
rect 6523 3482 6557 3516
rect 6557 3482 6667 3516
rect 6667 3482 6701 3516
rect 6701 3482 6702 3516
rect 6522 3444 6702 3482
rect 6522 3410 6523 3444
rect 6523 3410 6557 3444
rect 6557 3410 6667 3444
rect 6667 3410 6701 3444
rect 6701 3410 6702 3444
rect 6522 3372 6702 3410
rect 6522 3338 6523 3372
rect 6523 3338 6557 3372
rect 6557 3338 6667 3372
rect 6667 3338 6701 3372
rect 6701 3338 6702 3372
rect 6522 3300 6702 3338
rect 6522 3266 6523 3300
rect 6523 3266 6557 3300
rect 6557 3266 6667 3300
rect 6667 3266 6701 3300
rect 6701 3266 6702 3300
rect 6522 3228 6702 3266
rect 6522 3194 6523 3228
rect 6523 3194 6557 3228
rect 6557 3194 6667 3228
rect 6667 3194 6701 3228
rect 6701 3194 6702 3228
rect 6522 3108 6702 3194
rect 6522 3074 6523 3108
rect 6523 3074 6557 3108
rect 6557 3074 6595 3108
rect 6595 3074 6629 3108
rect 6629 3074 6667 3108
rect 6667 3074 6701 3108
rect 6701 3074 6702 3108
rect 6522 3028 6702 3074
rect 6522 2994 6523 3028
rect 6523 2994 6557 3028
rect 6557 2994 6595 3028
rect 6595 2994 6629 3028
rect 6629 2994 6667 3028
rect 6667 2994 6701 3028
rect 6701 2994 6702 3028
rect 6522 2948 6702 2994
rect 6522 2914 6523 2948
rect 6523 2914 6557 2948
rect 6557 2914 6595 2948
rect 6595 2914 6629 2948
rect 6629 2914 6667 2948
rect 6667 2914 6701 2948
rect 6701 2914 6702 2948
rect 6522 2868 6702 2914
rect 6522 2834 6523 2868
rect 6523 2834 6557 2868
rect 6557 2834 6595 2868
rect 6595 2834 6629 2868
rect 6629 2834 6667 2868
rect 6667 2834 6701 2868
rect 6701 2834 6702 2868
rect 6522 2788 6702 2834
rect 6522 2754 6523 2788
rect 6523 2754 6557 2788
rect 6557 2754 6595 2788
rect 6595 2754 6629 2788
rect 6629 2754 6667 2788
rect 6667 2754 6701 2788
rect 6701 2754 6702 2788
rect 6522 2708 6702 2754
rect 6522 2674 6523 2708
rect 6523 2674 6557 2708
rect 6557 2674 6595 2708
rect 6595 2674 6629 2708
rect 6629 2674 6667 2708
rect 6667 2674 6701 2708
rect 6701 2674 6702 2708
rect 6522 2628 6702 2674
rect 6522 2594 6523 2628
rect 6523 2594 6557 2628
rect 6557 2594 6595 2628
rect 6595 2594 6629 2628
rect 6629 2594 6667 2628
rect 6667 2594 6701 2628
rect 6701 2594 6702 2628
rect 6522 2518 6702 2594
rect 6522 2484 6523 2518
rect 6523 2484 6557 2518
rect 6557 2484 6667 2518
rect 6667 2484 6701 2518
rect 6701 2484 6702 2518
rect 6522 2446 6702 2484
rect 6522 2412 6523 2446
rect 6523 2412 6557 2446
rect 6557 2412 6667 2446
rect 6667 2412 6701 2446
rect 6701 2412 6702 2446
rect 6522 2374 6702 2412
rect 6522 2340 6523 2374
rect 6523 2340 6557 2374
rect 6557 2340 6667 2374
rect 6667 2340 6701 2374
rect 6701 2340 6702 2374
rect 6522 2302 6702 2340
rect 6522 2268 6523 2302
rect 6523 2268 6557 2302
rect 6557 2268 6667 2302
rect 6667 2268 6701 2302
rect 6701 2268 6702 2302
rect 6522 2230 6702 2268
rect 6522 2196 6523 2230
rect 6523 2196 6557 2230
rect 6557 2196 6667 2230
rect 6667 2196 6701 2230
rect 6701 2196 6702 2230
rect 6522 2158 6702 2196
rect 6522 2124 6523 2158
rect 6523 2124 6557 2158
rect 6557 2124 6667 2158
rect 6667 2124 6701 2158
rect 6701 2124 6702 2158
rect 6522 2086 6702 2124
rect 6522 2052 6523 2086
rect 6523 2052 6557 2086
rect 6557 2052 6667 2086
rect 6667 2052 6701 2086
rect 6701 2052 6702 2086
rect 6522 2014 6702 2052
rect 6522 1980 6523 2014
rect 6523 1980 6557 2014
rect 6557 1980 6667 2014
rect 6667 1980 6701 2014
rect 6701 1980 6702 2014
rect 6522 1942 6702 1980
rect 6522 1908 6523 1942
rect 6523 1908 6557 1942
rect 6557 1908 6667 1942
rect 6667 1908 6701 1942
rect 6701 1908 6702 1942
rect 6522 1870 6702 1908
rect 6522 1836 6523 1870
rect 6523 1836 6557 1870
rect 6557 1836 6667 1870
rect 6667 1836 6701 1870
rect 6701 1836 6702 1870
rect 6522 1798 6702 1836
rect 6522 1764 6523 1798
rect 6523 1764 6557 1798
rect 6557 1764 6667 1798
rect 6667 1764 6701 1798
rect 6701 1764 6702 1798
rect 6522 1726 6702 1764
rect 6522 1692 6523 1726
rect 6523 1692 6557 1726
rect 6557 1692 6667 1726
rect 6667 1692 6701 1726
rect 6701 1692 6702 1726
rect 6522 1654 6702 1692
rect 6522 1620 6523 1654
rect 6523 1620 6557 1654
rect 6557 1620 6667 1654
rect 6667 1620 6701 1654
rect 6701 1620 6702 1654
rect 6522 1568 6702 1620
rect 7018 4098 7070 4119
rect 7018 4067 7019 4098
rect 7019 4067 7053 4098
rect 7053 4067 7070 4098
rect 7082 4098 7134 4119
rect 7082 4067 7091 4098
rect 7091 4067 7125 4098
rect 7125 4067 7134 4098
rect 7146 4098 7198 4119
rect 7146 4067 7163 4098
rect 7163 4067 7197 4098
rect 7197 4067 7198 4098
rect 7018 4025 7070 4054
rect 7018 4002 7019 4025
rect 7019 4002 7053 4025
rect 7053 4002 7070 4025
rect 7082 4025 7134 4054
rect 7082 4002 7091 4025
rect 7091 4002 7125 4025
rect 7125 4002 7134 4025
rect 7146 4025 7198 4054
rect 7146 4002 7163 4025
rect 7163 4002 7197 4025
rect 7197 4002 7198 4025
rect 7018 3952 7070 3989
rect 7018 3937 7019 3952
rect 7019 3937 7053 3952
rect 7053 3937 7070 3952
rect 7082 3952 7134 3989
rect 7082 3937 7091 3952
rect 7091 3937 7125 3952
rect 7125 3937 7134 3952
rect 7146 3952 7198 3989
rect 7146 3937 7163 3952
rect 7163 3937 7197 3952
rect 7197 3937 7198 3952
rect 7018 3918 7019 3924
rect 7019 3918 7053 3924
rect 7053 3918 7091 3924
rect 7091 3918 7125 3924
rect 7125 3918 7163 3924
rect 7163 3918 7197 3924
rect 7197 3918 7198 3924
rect 7018 3879 7198 3918
rect 7018 3845 7019 3879
rect 7019 3845 7053 3879
rect 7053 3845 7091 3879
rect 7091 3845 7125 3879
rect 7125 3845 7163 3879
rect 7163 3845 7197 3879
rect 7197 3845 7198 3879
rect 7018 3806 7198 3845
rect 7018 3772 7019 3806
rect 7019 3772 7053 3806
rect 7053 3772 7091 3806
rect 7091 3772 7125 3806
rect 7125 3772 7163 3806
rect 7163 3772 7197 3806
rect 7197 3772 7198 3806
rect 7018 3733 7198 3772
rect 7018 3699 7019 3733
rect 7019 3699 7053 3733
rect 7053 3699 7091 3733
rect 7091 3699 7125 3733
rect 7125 3699 7163 3733
rect 7163 3699 7197 3733
rect 7197 3699 7198 3733
rect 7018 3660 7198 3699
rect 7018 3626 7019 3660
rect 7019 3626 7053 3660
rect 7053 3626 7091 3660
rect 7091 3626 7125 3660
rect 7125 3626 7163 3660
rect 7163 3626 7197 3660
rect 7197 3626 7198 3660
rect 7018 3587 7198 3626
rect 7018 3553 7019 3587
rect 7019 3553 7053 3587
rect 7053 3553 7091 3587
rect 7091 3553 7125 3587
rect 7125 3553 7163 3587
rect 7163 3553 7197 3587
rect 7197 3553 7198 3587
rect 7018 3514 7198 3553
rect 7018 3480 7019 3514
rect 7019 3480 7053 3514
rect 7053 3480 7091 3514
rect 7091 3480 7125 3514
rect 7125 3480 7163 3514
rect 7163 3480 7197 3514
rect 7197 3480 7198 3514
rect 7018 3441 7198 3480
rect 7018 3407 7019 3441
rect 7019 3407 7053 3441
rect 7053 3407 7091 3441
rect 7091 3407 7125 3441
rect 7125 3407 7163 3441
rect 7163 3407 7197 3441
rect 7197 3407 7198 3441
rect 7018 3368 7198 3407
rect 7018 3334 7019 3368
rect 7019 3334 7053 3368
rect 7053 3334 7091 3368
rect 7091 3334 7125 3368
rect 7125 3334 7163 3368
rect 7163 3334 7197 3368
rect 7197 3334 7198 3368
rect 7018 3295 7198 3334
rect 7018 3261 7019 3295
rect 7019 3261 7053 3295
rect 7053 3261 7091 3295
rect 7091 3261 7125 3295
rect 7125 3261 7163 3295
rect 7163 3261 7197 3295
rect 7197 3261 7198 3295
rect 7018 3222 7198 3261
rect 7018 3188 7019 3222
rect 7019 3188 7053 3222
rect 7053 3188 7091 3222
rect 7091 3188 7125 3222
rect 7125 3188 7163 3222
rect 7163 3188 7197 3222
rect 7197 3188 7198 3222
rect 7018 3149 7198 3188
rect 7018 3115 7019 3149
rect 7019 3115 7053 3149
rect 7053 3115 7091 3149
rect 7091 3115 7125 3149
rect 7125 3115 7163 3149
rect 7163 3115 7197 3149
rect 7197 3115 7198 3149
rect 7018 3076 7198 3115
rect 7018 3042 7019 3076
rect 7019 3042 7053 3076
rect 7053 3042 7091 3076
rect 7091 3042 7125 3076
rect 7125 3042 7163 3076
rect 7163 3042 7197 3076
rect 7197 3042 7198 3076
rect 7018 3003 7198 3042
rect 7018 2969 7019 3003
rect 7019 2969 7053 3003
rect 7053 2969 7091 3003
rect 7091 2969 7125 3003
rect 7125 2969 7163 3003
rect 7163 2969 7197 3003
rect 7197 2969 7198 3003
rect 7018 2930 7198 2969
rect 7018 2896 7019 2930
rect 7019 2896 7053 2930
rect 7053 2896 7091 2930
rect 7091 2896 7125 2930
rect 7125 2896 7163 2930
rect 7163 2896 7197 2930
rect 7197 2896 7198 2930
rect 7018 2857 7198 2896
rect 7018 2823 7019 2857
rect 7019 2823 7053 2857
rect 7053 2823 7091 2857
rect 7091 2823 7125 2857
rect 7125 2823 7163 2857
rect 7163 2823 7197 2857
rect 7197 2823 7198 2857
rect 7018 2784 7198 2823
rect 7018 2750 7019 2784
rect 7019 2750 7053 2784
rect 7053 2750 7091 2784
rect 7091 2750 7125 2784
rect 7125 2750 7163 2784
rect 7163 2750 7197 2784
rect 7197 2750 7198 2784
rect 7018 2711 7198 2750
rect 7018 2677 7019 2711
rect 7019 2677 7053 2711
rect 7053 2677 7091 2711
rect 7091 2677 7125 2711
rect 7125 2677 7163 2711
rect 7163 2677 7197 2711
rect 7197 2677 7198 2711
rect 7018 2638 7198 2677
rect 7018 2604 7019 2638
rect 7019 2604 7053 2638
rect 7053 2604 7091 2638
rect 7091 2604 7125 2638
rect 7125 2604 7163 2638
rect 7163 2604 7197 2638
rect 7197 2604 7198 2638
rect 7018 2565 7198 2604
rect 7018 2531 7019 2565
rect 7019 2531 7053 2565
rect 7053 2531 7091 2565
rect 7091 2531 7125 2565
rect 7125 2531 7163 2565
rect 7163 2531 7197 2565
rect 7197 2531 7198 2565
rect 7018 2492 7198 2531
rect 7018 2458 7019 2492
rect 7019 2458 7053 2492
rect 7053 2458 7091 2492
rect 7091 2458 7125 2492
rect 7125 2458 7163 2492
rect 7163 2458 7197 2492
rect 7197 2458 7198 2492
rect 7018 2419 7198 2458
rect 7018 2385 7019 2419
rect 7019 2385 7053 2419
rect 7053 2385 7091 2419
rect 7091 2385 7125 2419
rect 7125 2385 7163 2419
rect 7163 2385 7197 2419
rect 7197 2385 7198 2419
rect 7018 2346 7198 2385
rect 7018 2312 7019 2346
rect 7019 2312 7053 2346
rect 7053 2312 7091 2346
rect 7091 2312 7125 2346
rect 7125 2312 7163 2346
rect 7163 2312 7197 2346
rect 7197 2312 7198 2346
rect 7018 2273 7198 2312
rect 7018 2239 7019 2273
rect 7019 2239 7053 2273
rect 7053 2239 7091 2273
rect 7091 2239 7125 2273
rect 7125 2239 7163 2273
rect 7163 2239 7197 2273
rect 7197 2239 7198 2273
rect 7018 2200 7198 2239
rect 7018 2166 7019 2200
rect 7019 2166 7053 2200
rect 7053 2166 7091 2200
rect 7091 2166 7125 2200
rect 7125 2166 7163 2200
rect 7163 2166 7197 2200
rect 7197 2166 7198 2200
rect 7018 2126 7198 2166
rect 7018 2092 7019 2126
rect 7019 2092 7053 2126
rect 7053 2092 7091 2126
rect 7091 2092 7125 2126
rect 7125 2092 7163 2126
rect 7163 2092 7197 2126
rect 7197 2092 7198 2126
rect 7018 2052 7198 2092
rect 7018 2018 7019 2052
rect 7019 2018 7053 2052
rect 7053 2018 7091 2052
rect 7091 2018 7125 2052
rect 7125 2018 7163 2052
rect 7163 2018 7197 2052
rect 7197 2018 7198 2052
rect 7018 1978 7198 2018
rect 7018 1944 7019 1978
rect 7019 1944 7053 1978
rect 7053 1944 7091 1978
rect 7091 1944 7125 1978
rect 7125 1944 7163 1978
rect 7163 1944 7197 1978
rect 7197 1944 7198 1978
rect 7018 1904 7198 1944
rect 7018 1870 7019 1904
rect 7019 1870 7053 1904
rect 7053 1870 7091 1904
rect 7091 1870 7125 1904
rect 7125 1870 7163 1904
rect 7163 1870 7197 1904
rect 7197 1870 7198 1904
rect 7018 1830 7198 1870
rect 7018 1796 7019 1830
rect 7019 1796 7053 1830
rect 7053 1796 7091 1830
rect 7091 1796 7125 1830
rect 7125 1796 7163 1830
rect 7163 1796 7197 1830
rect 7197 1796 7198 1830
rect 7018 1756 7198 1796
rect 7018 1722 7019 1756
rect 7019 1722 7053 1756
rect 7053 1722 7091 1756
rect 7091 1722 7125 1756
rect 7125 1722 7163 1756
rect 7163 1722 7197 1756
rect 7197 1722 7198 1756
rect 7018 1682 7198 1722
rect 7018 1648 7019 1682
rect 7019 1648 7053 1682
rect 7053 1648 7091 1682
rect 7091 1648 7125 1682
rect 7125 1648 7163 1682
rect 7163 1648 7197 1682
rect 7197 1648 7198 1682
rect 7018 1608 7198 1648
rect 7018 1574 7019 1608
rect 7019 1574 7053 1608
rect 7053 1574 7091 1608
rect 7091 1574 7125 1608
rect 7125 1574 7163 1608
rect 7163 1574 7197 1608
rect 7197 1574 7198 1608
rect 7018 1568 7198 1574
rect 7514 4092 7566 4124
rect 7514 4072 7515 4092
rect 7515 4072 7549 4092
rect 7549 4072 7566 4092
rect 7578 4072 7630 4124
rect 7642 4092 7694 4124
rect 7642 4072 7659 4092
rect 7659 4072 7693 4092
rect 7693 4072 7694 4092
rect 7514 4058 7515 4059
rect 7515 4058 7549 4059
rect 7549 4058 7566 4059
rect 7514 4020 7566 4058
rect 7514 4007 7515 4020
rect 7515 4007 7549 4020
rect 7549 4007 7566 4020
rect 7578 4007 7630 4059
rect 7642 4058 7659 4059
rect 7659 4058 7693 4059
rect 7693 4058 7694 4059
rect 7642 4020 7694 4058
rect 7642 4007 7659 4020
rect 7659 4007 7693 4020
rect 7693 4007 7694 4020
rect 7514 3986 7515 3994
rect 7515 3986 7549 3994
rect 7549 3986 7566 3994
rect 7514 3948 7566 3986
rect 7514 3942 7515 3948
rect 7515 3942 7549 3948
rect 7549 3942 7566 3948
rect 7578 3942 7630 3994
rect 7642 3986 7659 3994
rect 7659 3986 7693 3994
rect 7693 3986 7694 3994
rect 7642 3948 7694 3986
rect 7642 3942 7659 3948
rect 7659 3942 7693 3948
rect 7693 3942 7694 3948
rect 7514 3914 7515 3929
rect 7515 3914 7549 3929
rect 7549 3914 7566 3929
rect 7514 3877 7566 3914
rect 7578 3877 7630 3929
rect 7642 3914 7659 3929
rect 7659 3914 7693 3929
rect 7693 3914 7694 3929
rect 7642 3877 7694 3914
rect 7514 3842 7515 3864
rect 7515 3842 7549 3864
rect 7549 3842 7566 3864
rect 7514 3812 7566 3842
rect 7578 3812 7630 3864
rect 7642 3842 7659 3864
rect 7659 3842 7693 3864
rect 7693 3842 7694 3864
rect 7642 3812 7694 3842
rect 7514 3770 7515 3799
rect 7515 3770 7549 3799
rect 7549 3770 7566 3799
rect 7514 3747 7566 3770
rect 7578 3747 7630 3799
rect 7642 3770 7659 3799
rect 7659 3770 7693 3799
rect 7693 3770 7694 3799
rect 7642 3747 7694 3770
rect 7514 3732 7566 3734
rect 7514 3698 7515 3732
rect 7515 3698 7549 3732
rect 7549 3698 7566 3732
rect 7514 3682 7566 3698
rect 7578 3682 7630 3734
rect 7642 3732 7694 3734
rect 7642 3698 7659 3732
rect 7659 3698 7693 3732
rect 7693 3698 7694 3732
rect 7642 3682 7694 3698
rect 7514 3660 7566 3669
rect 7514 3626 7515 3660
rect 7515 3626 7549 3660
rect 7549 3626 7566 3660
rect 7514 3617 7566 3626
rect 7578 3617 7630 3669
rect 7642 3660 7694 3669
rect 7642 3626 7659 3660
rect 7659 3626 7693 3660
rect 7693 3626 7694 3660
rect 7642 3617 7694 3626
rect 7514 3588 7694 3604
rect 7514 3554 7515 3588
rect 7515 3554 7549 3588
rect 7549 3554 7659 3588
rect 7659 3554 7693 3588
rect 7693 3554 7694 3588
rect 7514 3516 7694 3554
rect 7514 3482 7515 3516
rect 7515 3482 7549 3516
rect 7549 3482 7659 3516
rect 7659 3482 7693 3516
rect 7693 3482 7694 3516
rect 7514 3444 7694 3482
rect 7514 3410 7515 3444
rect 7515 3410 7549 3444
rect 7549 3410 7659 3444
rect 7659 3410 7693 3444
rect 7693 3410 7694 3444
rect 7514 3372 7694 3410
rect 7514 3338 7515 3372
rect 7515 3338 7549 3372
rect 7549 3338 7659 3372
rect 7659 3338 7693 3372
rect 7693 3338 7694 3372
rect 7514 3300 7694 3338
rect 7514 3266 7515 3300
rect 7515 3266 7549 3300
rect 7549 3266 7659 3300
rect 7659 3266 7693 3300
rect 7693 3266 7694 3300
rect 7514 3228 7694 3266
rect 7514 3194 7515 3228
rect 7515 3194 7549 3228
rect 7549 3194 7659 3228
rect 7659 3194 7693 3228
rect 7693 3194 7694 3228
rect 7514 3108 7694 3194
rect 7514 3074 7515 3108
rect 7515 3074 7549 3108
rect 7549 3074 7587 3108
rect 7587 3074 7621 3108
rect 7621 3074 7659 3108
rect 7659 3074 7693 3108
rect 7693 3074 7694 3108
rect 7514 3028 7694 3074
rect 7514 2994 7515 3028
rect 7515 2994 7549 3028
rect 7549 2994 7587 3028
rect 7587 2994 7621 3028
rect 7621 2994 7659 3028
rect 7659 2994 7693 3028
rect 7693 2994 7694 3028
rect 7514 2948 7694 2994
rect 7514 2914 7515 2948
rect 7515 2914 7549 2948
rect 7549 2914 7587 2948
rect 7587 2914 7621 2948
rect 7621 2914 7659 2948
rect 7659 2914 7693 2948
rect 7693 2914 7694 2948
rect 7514 2868 7694 2914
rect 7514 2834 7515 2868
rect 7515 2834 7549 2868
rect 7549 2834 7587 2868
rect 7587 2834 7621 2868
rect 7621 2834 7659 2868
rect 7659 2834 7693 2868
rect 7693 2834 7694 2868
rect 7514 2788 7694 2834
rect 7514 2754 7515 2788
rect 7515 2754 7549 2788
rect 7549 2754 7587 2788
rect 7587 2754 7621 2788
rect 7621 2754 7659 2788
rect 7659 2754 7693 2788
rect 7693 2754 7694 2788
rect 7514 2708 7694 2754
rect 7514 2674 7515 2708
rect 7515 2674 7549 2708
rect 7549 2674 7587 2708
rect 7587 2674 7621 2708
rect 7621 2674 7659 2708
rect 7659 2674 7693 2708
rect 7693 2674 7694 2708
rect 7514 2628 7694 2674
rect 7514 2594 7515 2628
rect 7515 2594 7549 2628
rect 7549 2594 7587 2628
rect 7587 2594 7621 2628
rect 7621 2594 7659 2628
rect 7659 2594 7693 2628
rect 7693 2594 7694 2628
rect 7514 2518 7694 2594
rect 7514 2484 7515 2518
rect 7515 2484 7549 2518
rect 7549 2484 7659 2518
rect 7659 2484 7693 2518
rect 7693 2484 7694 2518
rect 7514 2446 7694 2484
rect 7514 2412 7515 2446
rect 7515 2412 7549 2446
rect 7549 2412 7659 2446
rect 7659 2412 7693 2446
rect 7693 2412 7694 2446
rect 7514 2374 7694 2412
rect 7514 2340 7515 2374
rect 7515 2340 7549 2374
rect 7549 2340 7659 2374
rect 7659 2340 7693 2374
rect 7693 2340 7694 2374
rect 7514 2302 7694 2340
rect 7514 2268 7515 2302
rect 7515 2268 7549 2302
rect 7549 2268 7659 2302
rect 7659 2268 7693 2302
rect 7693 2268 7694 2302
rect 7514 2230 7694 2268
rect 7514 2196 7515 2230
rect 7515 2196 7549 2230
rect 7549 2196 7659 2230
rect 7659 2196 7693 2230
rect 7693 2196 7694 2230
rect 7514 2158 7694 2196
rect 7514 2124 7515 2158
rect 7515 2124 7549 2158
rect 7549 2124 7659 2158
rect 7659 2124 7693 2158
rect 7693 2124 7694 2158
rect 7514 2086 7694 2124
rect 7514 2052 7515 2086
rect 7515 2052 7549 2086
rect 7549 2052 7659 2086
rect 7659 2052 7693 2086
rect 7693 2052 7694 2086
rect 7514 2014 7694 2052
rect 7514 1980 7515 2014
rect 7515 1980 7549 2014
rect 7549 1980 7659 2014
rect 7659 1980 7693 2014
rect 7693 1980 7694 2014
rect 7514 1942 7694 1980
rect 7514 1908 7515 1942
rect 7515 1908 7549 1942
rect 7549 1908 7659 1942
rect 7659 1908 7693 1942
rect 7693 1908 7694 1942
rect 7514 1870 7694 1908
rect 7514 1836 7515 1870
rect 7515 1836 7549 1870
rect 7549 1836 7659 1870
rect 7659 1836 7693 1870
rect 7693 1836 7694 1870
rect 7514 1798 7694 1836
rect 7514 1764 7515 1798
rect 7515 1764 7549 1798
rect 7549 1764 7659 1798
rect 7659 1764 7693 1798
rect 7693 1764 7694 1798
rect 7514 1726 7694 1764
rect 7514 1692 7515 1726
rect 7515 1692 7549 1726
rect 7549 1692 7659 1726
rect 7659 1692 7693 1726
rect 7693 1692 7694 1726
rect 7514 1654 7694 1692
rect 7514 1620 7515 1654
rect 7515 1620 7549 1654
rect 7549 1620 7659 1654
rect 7659 1620 7693 1654
rect 7693 1620 7694 1654
rect 7514 1568 7694 1620
rect 8010 4098 8062 4119
rect 8010 4067 8011 4098
rect 8011 4067 8045 4098
rect 8045 4067 8062 4098
rect 8074 4098 8126 4119
rect 8074 4067 8083 4098
rect 8083 4067 8117 4098
rect 8117 4067 8126 4098
rect 8138 4098 8190 4119
rect 8138 4067 8155 4098
rect 8155 4067 8189 4098
rect 8189 4067 8190 4098
rect 8010 4025 8062 4054
rect 8010 4002 8011 4025
rect 8011 4002 8045 4025
rect 8045 4002 8062 4025
rect 8074 4025 8126 4054
rect 8074 4002 8083 4025
rect 8083 4002 8117 4025
rect 8117 4002 8126 4025
rect 8138 4025 8190 4054
rect 8138 4002 8155 4025
rect 8155 4002 8189 4025
rect 8189 4002 8190 4025
rect 8010 3952 8062 3989
rect 8010 3937 8011 3952
rect 8011 3937 8045 3952
rect 8045 3937 8062 3952
rect 8074 3952 8126 3989
rect 8074 3937 8083 3952
rect 8083 3937 8117 3952
rect 8117 3937 8126 3952
rect 8138 3952 8190 3989
rect 8138 3937 8155 3952
rect 8155 3937 8189 3952
rect 8189 3937 8190 3952
rect 8010 3918 8011 3924
rect 8011 3918 8045 3924
rect 8045 3918 8083 3924
rect 8083 3918 8117 3924
rect 8117 3918 8155 3924
rect 8155 3918 8189 3924
rect 8189 3918 8190 3924
rect 8010 3879 8190 3918
rect 8010 3845 8011 3879
rect 8011 3845 8045 3879
rect 8045 3845 8083 3879
rect 8083 3845 8117 3879
rect 8117 3845 8155 3879
rect 8155 3845 8189 3879
rect 8189 3845 8190 3879
rect 8010 3806 8190 3845
rect 8010 3772 8011 3806
rect 8011 3772 8045 3806
rect 8045 3772 8083 3806
rect 8083 3772 8117 3806
rect 8117 3772 8155 3806
rect 8155 3772 8189 3806
rect 8189 3772 8190 3806
rect 8010 3733 8190 3772
rect 8010 3699 8011 3733
rect 8011 3699 8045 3733
rect 8045 3699 8083 3733
rect 8083 3699 8117 3733
rect 8117 3699 8155 3733
rect 8155 3699 8189 3733
rect 8189 3699 8190 3733
rect 8010 3660 8190 3699
rect 8010 3626 8011 3660
rect 8011 3626 8045 3660
rect 8045 3626 8083 3660
rect 8083 3626 8117 3660
rect 8117 3626 8155 3660
rect 8155 3626 8189 3660
rect 8189 3626 8190 3660
rect 8010 3587 8190 3626
rect 8010 3553 8011 3587
rect 8011 3553 8045 3587
rect 8045 3553 8083 3587
rect 8083 3553 8117 3587
rect 8117 3553 8155 3587
rect 8155 3553 8189 3587
rect 8189 3553 8190 3587
rect 8010 3514 8190 3553
rect 8010 3480 8011 3514
rect 8011 3480 8045 3514
rect 8045 3480 8083 3514
rect 8083 3480 8117 3514
rect 8117 3480 8155 3514
rect 8155 3480 8189 3514
rect 8189 3480 8190 3514
rect 8010 3441 8190 3480
rect 8010 3407 8011 3441
rect 8011 3407 8045 3441
rect 8045 3407 8083 3441
rect 8083 3407 8117 3441
rect 8117 3407 8155 3441
rect 8155 3407 8189 3441
rect 8189 3407 8190 3441
rect 8010 3368 8190 3407
rect 8010 3334 8011 3368
rect 8011 3334 8045 3368
rect 8045 3334 8083 3368
rect 8083 3334 8117 3368
rect 8117 3334 8155 3368
rect 8155 3334 8189 3368
rect 8189 3334 8190 3368
rect 8010 3295 8190 3334
rect 8010 3261 8011 3295
rect 8011 3261 8045 3295
rect 8045 3261 8083 3295
rect 8083 3261 8117 3295
rect 8117 3261 8155 3295
rect 8155 3261 8189 3295
rect 8189 3261 8190 3295
rect 8010 3222 8190 3261
rect 8010 3188 8011 3222
rect 8011 3188 8045 3222
rect 8045 3188 8083 3222
rect 8083 3188 8117 3222
rect 8117 3188 8155 3222
rect 8155 3188 8189 3222
rect 8189 3188 8190 3222
rect 8010 3149 8190 3188
rect 8010 3115 8011 3149
rect 8011 3115 8045 3149
rect 8045 3115 8083 3149
rect 8083 3115 8117 3149
rect 8117 3115 8155 3149
rect 8155 3115 8189 3149
rect 8189 3115 8190 3149
rect 8010 3076 8190 3115
rect 8010 3042 8011 3076
rect 8011 3042 8045 3076
rect 8045 3042 8083 3076
rect 8083 3042 8117 3076
rect 8117 3042 8155 3076
rect 8155 3042 8189 3076
rect 8189 3042 8190 3076
rect 8010 3003 8190 3042
rect 8010 2969 8011 3003
rect 8011 2969 8045 3003
rect 8045 2969 8083 3003
rect 8083 2969 8117 3003
rect 8117 2969 8155 3003
rect 8155 2969 8189 3003
rect 8189 2969 8190 3003
rect 8010 2930 8190 2969
rect 8010 2896 8011 2930
rect 8011 2896 8045 2930
rect 8045 2896 8083 2930
rect 8083 2896 8117 2930
rect 8117 2896 8155 2930
rect 8155 2896 8189 2930
rect 8189 2896 8190 2930
rect 8010 2857 8190 2896
rect 8010 2823 8011 2857
rect 8011 2823 8045 2857
rect 8045 2823 8083 2857
rect 8083 2823 8117 2857
rect 8117 2823 8155 2857
rect 8155 2823 8189 2857
rect 8189 2823 8190 2857
rect 8010 2784 8190 2823
rect 8010 2750 8011 2784
rect 8011 2750 8045 2784
rect 8045 2750 8083 2784
rect 8083 2750 8117 2784
rect 8117 2750 8155 2784
rect 8155 2750 8189 2784
rect 8189 2750 8190 2784
rect 8010 2711 8190 2750
rect 8010 2677 8011 2711
rect 8011 2677 8045 2711
rect 8045 2677 8083 2711
rect 8083 2677 8117 2711
rect 8117 2677 8155 2711
rect 8155 2677 8189 2711
rect 8189 2677 8190 2711
rect 8010 2638 8190 2677
rect 8010 2604 8011 2638
rect 8011 2604 8045 2638
rect 8045 2604 8083 2638
rect 8083 2604 8117 2638
rect 8117 2604 8155 2638
rect 8155 2604 8189 2638
rect 8189 2604 8190 2638
rect 8010 2565 8190 2604
rect 8010 2531 8011 2565
rect 8011 2531 8045 2565
rect 8045 2531 8083 2565
rect 8083 2531 8117 2565
rect 8117 2531 8155 2565
rect 8155 2531 8189 2565
rect 8189 2531 8190 2565
rect 8010 2492 8190 2531
rect 8010 2458 8011 2492
rect 8011 2458 8045 2492
rect 8045 2458 8083 2492
rect 8083 2458 8117 2492
rect 8117 2458 8155 2492
rect 8155 2458 8189 2492
rect 8189 2458 8190 2492
rect 8010 2419 8190 2458
rect 8010 2385 8011 2419
rect 8011 2385 8045 2419
rect 8045 2385 8083 2419
rect 8083 2385 8117 2419
rect 8117 2385 8155 2419
rect 8155 2385 8189 2419
rect 8189 2385 8190 2419
rect 8010 2346 8190 2385
rect 8010 2312 8011 2346
rect 8011 2312 8045 2346
rect 8045 2312 8083 2346
rect 8083 2312 8117 2346
rect 8117 2312 8155 2346
rect 8155 2312 8189 2346
rect 8189 2312 8190 2346
rect 8010 2273 8190 2312
rect 8010 2239 8011 2273
rect 8011 2239 8045 2273
rect 8045 2239 8083 2273
rect 8083 2239 8117 2273
rect 8117 2239 8155 2273
rect 8155 2239 8189 2273
rect 8189 2239 8190 2273
rect 8010 2200 8190 2239
rect 8010 2166 8011 2200
rect 8011 2166 8045 2200
rect 8045 2166 8083 2200
rect 8083 2166 8117 2200
rect 8117 2166 8155 2200
rect 8155 2166 8189 2200
rect 8189 2166 8190 2200
rect 8010 2126 8190 2166
rect 8010 2092 8011 2126
rect 8011 2092 8045 2126
rect 8045 2092 8083 2126
rect 8083 2092 8117 2126
rect 8117 2092 8155 2126
rect 8155 2092 8189 2126
rect 8189 2092 8190 2126
rect 8010 2052 8190 2092
rect 8010 2018 8011 2052
rect 8011 2018 8045 2052
rect 8045 2018 8083 2052
rect 8083 2018 8117 2052
rect 8117 2018 8155 2052
rect 8155 2018 8189 2052
rect 8189 2018 8190 2052
rect 8010 1978 8190 2018
rect 8010 1944 8011 1978
rect 8011 1944 8045 1978
rect 8045 1944 8083 1978
rect 8083 1944 8117 1978
rect 8117 1944 8155 1978
rect 8155 1944 8189 1978
rect 8189 1944 8190 1978
rect 8010 1904 8190 1944
rect 8010 1870 8011 1904
rect 8011 1870 8045 1904
rect 8045 1870 8083 1904
rect 8083 1870 8117 1904
rect 8117 1870 8155 1904
rect 8155 1870 8189 1904
rect 8189 1870 8190 1904
rect 8010 1830 8190 1870
rect 8010 1796 8011 1830
rect 8011 1796 8045 1830
rect 8045 1796 8083 1830
rect 8083 1796 8117 1830
rect 8117 1796 8155 1830
rect 8155 1796 8189 1830
rect 8189 1796 8190 1830
rect 8010 1756 8190 1796
rect 8010 1722 8011 1756
rect 8011 1722 8045 1756
rect 8045 1722 8083 1756
rect 8083 1722 8117 1756
rect 8117 1722 8155 1756
rect 8155 1722 8189 1756
rect 8189 1722 8190 1756
rect 8010 1682 8190 1722
rect 8010 1648 8011 1682
rect 8011 1648 8045 1682
rect 8045 1648 8083 1682
rect 8083 1648 8117 1682
rect 8117 1648 8155 1682
rect 8155 1648 8189 1682
rect 8189 1648 8190 1682
rect 8010 1608 8190 1648
rect 8010 1574 8011 1608
rect 8011 1574 8045 1608
rect 8045 1574 8083 1608
rect 8083 1574 8117 1608
rect 8117 1574 8155 1608
rect 8155 1574 8189 1608
rect 8189 1574 8190 1608
rect 8010 1568 8190 1574
rect 8506 4092 8558 4124
rect 8506 4072 8507 4092
rect 8507 4072 8541 4092
rect 8541 4072 8558 4092
rect 8570 4072 8622 4124
rect 8634 4092 8686 4124
rect 8634 4072 8651 4092
rect 8651 4072 8685 4092
rect 8685 4072 8686 4092
rect 8506 4058 8507 4059
rect 8507 4058 8541 4059
rect 8541 4058 8558 4059
rect 8506 4020 8558 4058
rect 8506 4007 8507 4020
rect 8507 4007 8541 4020
rect 8541 4007 8558 4020
rect 8570 4007 8622 4059
rect 8634 4058 8651 4059
rect 8651 4058 8685 4059
rect 8685 4058 8686 4059
rect 8634 4020 8686 4058
rect 8634 4007 8651 4020
rect 8651 4007 8685 4020
rect 8685 4007 8686 4020
rect 8506 3986 8507 3994
rect 8507 3986 8541 3994
rect 8541 3986 8558 3994
rect 8506 3948 8558 3986
rect 8506 3942 8507 3948
rect 8507 3942 8541 3948
rect 8541 3942 8558 3948
rect 8570 3942 8622 3994
rect 8634 3986 8651 3994
rect 8651 3986 8685 3994
rect 8685 3986 8686 3994
rect 8634 3948 8686 3986
rect 8634 3942 8651 3948
rect 8651 3942 8685 3948
rect 8685 3942 8686 3948
rect 8506 3914 8507 3929
rect 8507 3914 8541 3929
rect 8541 3914 8558 3929
rect 8506 3877 8558 3914
rect 8570 3877 8622 3929
rect 8634 3914 8651 3929
rect 8651 3914 8685 3929
rect 8685 3914 8686 3929
rect 8634 3877 8686 3914
rect 8506 3842 8507 3864
rect 8507 3842 8541 3864
rect 8541 3842 8558 3864
rect 8506 3812 8558 3842
rect 8570 3812 8622 3864
rect 8634 3842 8651 3864
rect 8651 3842 8685 3864
rect 8685 3842 8686 3864
rect 8634 3812 8686 3842
rect 8506 3770 8507 3799
rect 8507 3770 8541 3799
rect 8541 3770 8558 3799
rect 8506 3747 8558 3770
rect 8570 3747 8622 3799
rect 8634 3770 8651 3799
rect 8651 3770 8685 3799
rect 8685 3770 8686 3799
rect 8634 3747 8686 3770
rect 8506 3732 8558 3734
rect 8506 3698 8507 3732
rect 8507 3698 8541 3732
rect 8541 3698 8558 3732
rect 8506 3682 8558 3698
rect 8570 3682 8622 3734
rect 8634 3732 8686 3734
rect 8634 3698 8651 3732
rect 8651 3698 8685 3732
rect 8685 3698 8686 3732
rect 8634 3682 8686 3698
rect 8506 3660 8558 3669
rect 8506 3626 8507 3660
rect 8507 3626 8541 3660
rect 8541 3626 8558 3660
rect 8506 3617 8558 3626
rect 8570 3617 8622 3669
rect 8634 3660 8686 3669
rect 8634 3626 8651 3660
rect 8651 3626 8685 3660
rect 8685 3626 8686 3660
rect 8634 3617 8686 3626
rect 8506 3588 8686 3604
rect 8506 3554 8507 3588
rect 8507 3554 8541 3588
rect 8541 3554 8651 3588
rect 8651 3554 8685 3588
rect 8685 3554 8686 3588
rect 8506 3516 8686 3554
rect 8506 3482 8507 3516
rect 8507 3482 8541 3516
rect 8541 3482 8651 3516
rect 8651 3482 8685 3516
rect 8685 3482 8686 3516
rect 8506 3444 8686 3482
rect 8506 3410 8507 3444
rect 8507 3410 8541 3444
rect 8541 3410 8651 3444
rect 8651 3410 8685 3444
rect 8685 3410 8686 3444
rect 8506 3372 8686 3410
rect 8506 3338 8507 3372
rect 8507 3338 8541 3372
rect 8541 3338 8651 3372
rect 8651 3338 8685 3372
rect 8685 3338 8686 3372
rect 8506 3300 8686 3338
rect 8506 3266 8507 3300
rect 8507 3266 8541 3300
rect 8541 3266 8651 3300
rect 8651 3266 8685 3300
rect 8685 3266 8686 3300
rect 8506 3228 8686 3266
rect 8506 3194 8507 3228
rect 8507 3194 8541 3228
rect 8541 3194 8651 3228
rect 8651 3194 8685 3228
rect 8685 3194 8686 3228
rect 8506 3108 8686 3194
rect 8506 3074 8507 3108
rect 8507 3074 8541 3108
rect 8541 3074 8579 3108
rect 8579 3074 8613 3108
rect 8613 3074 8651 3108
rect 8651 3074 8685 3108
rect 8685 3074 8686 3108
rect 8506 3028 8686 3074
rect 8506 2994 8507 3028
rect 8507 2994 8541 3028
rect 8541 2994 8579 3028
rect 8579 2994 8613 3028
rect 8613 2994 8651 3028
rect 8651 2994 8685 3028
rect 8685 2994 8686 3028
rect 8506 2948 8686 2994
rect 8506 2914 8507 2948
rect 8507 2914 8541 2948
rect 8541 2914 8579 2948
rect 8579 2914 8613 2948
rect 8613 2914 8651 2948
rect 8651 2914 8685 2948
rect 8685 2914 8686 2948
rect 8506 2868 8686 2914
rect 8506 2834 8507 2868
rect 8507 2834 8541 2868
rect 8541 2834 8579 2868
rect 8579 2834 8613 2868
rect 8613 2834 8651 2868
rect 8651 2834 8685 2868
rect 8685 2834 8686 2868
rect 8506 2788 8686 2834
rect 8506 2754 8507 2788
rect 8507 2754 8541 2788
rect 8541 2754 8579 2788
rect 8579 2754 8613 2788
rect 8613 2754 8651 2788
rect 8651 2754 8685 2788
rect 8685 2754 8686 2788
rect 8506 2708 8686 2754
rect 8506 2674 8507 2708
rect 8507 2674 8541 2708
rect 8541 2674 8579 2708
rect 8579 2674 8613 2708
rect 8613 2674 8651 2708
rect 8651 2674 8685 2708
rect 8685 2674 8686 2708
rect 8506 2628 8686 2674
rect 8506 2594 8507 2628
rect 8507 2594 8541 2628
rect 8541 2594 8579 2628
rect 8579 2594 8613 2628
rect 8613 2594 8651 2628
rect 8651 2594 8685 2628
rect 8685 2594 8686 2628
rect 8506 2518 8686 2594
rect 8506 2484 8507 2518
rect 8507 2484 8541 2518
rect 8541 2484 8651 2518
rect 8651 2484 8685 2518
rect 8685 2484 8686 2518
rect 8506 2446 8686 2484
rect 8506 2412 8507 2446
rect 8507 2412 8541 2446
rect 8541 2412 8651 2446
rect 8651 2412 8685 2446
rect 8685 2412 8686 2446
rect 8506 2374 8686 2412
rect 8506 2340 8507 2374
rect 8507 2340 8541 2374
rect 8541 2340 8651 2374
rect 8651 2340 8685 2374
rect 8685 2340 8686 2374
rect 8506 2302 8686 2340
rect 8506 2268 8507 2302
rect 8507 2268 8541 2302
rect 8541 2268 8651 2302
rect 8651 2268 8685 2302
rect 8685 2268 8686 2302
rect 8506 2230 8686 2268
rect 8506 2196 8507 2230
rect 8507 2196 8541 2230
rect 8541 2196 8651 2230
rect 8651 2196 8685 2230
rect 8685 2196 8686 2230
rect 8506 2158 8686 2196
rect 8506 2124 8507 2158
rect 8507 2124 8541 2158
rect 8541 2124 8651 2158
rect 8651 2124 8685 2158
rect 8685 2124 8686 2158
rect 8506 2086 8686 2124
rect 8506 2052 8507 2086
rect 8507 2052 8541 2086
rect 8541 2052 8651 2086
rect 8651 2052 8685 2086
rect 8685 2052 8686 2086
rect 8506 2014 8686 2052
rect 8506 1980 8507 2014
rect 8507 1980 8541 2014
rect 8541 1980 8651 2014
rect 8651 1980 8685 2014
rect 8685 1980 8686 2014
rect 8506 1942 8686 1980
rect 8506 1908 8507 1942
rect 8507 1908 8541 1942
rect 8541 1908 8651 1942
rect 8651 1908 8685 1942
rect 8685 1908 8686 1942
rect 8506 1870 8686 1908
rect 8506 1836 8507 1870
rect 8507 1836 8541 1870
rect 8541 1836 8651 1870
rect 8651 1836 8685 1870
rect 8685 1836 8686 1870
rect 8506 1798 8686 1836
rect 8506 1764 8507 1798
rect 8507 1764 8541 1798
rect 8541 1764 8651 1798
rect 8651 1764 8685 1798
rect 8685 1764 8686 1798
rect 8506 1726 8686 1764
rect 8506 1692 8507 1726
rect 8507 1692 8541 1726
rect 8541 1692 8651 1726
rect 8651 1692 8685 1726
rect 8685 1692 8686 1726
rect 8506 1654 8686 1692
rect 8506 1620 8507 1654
rect 8507 1620 8541 1654
rect 8541 1620 8651 1654
rect 8651 1620 8685 1654
rect 8685 1620 8686 1654
rect 8506 1568 8686 1620
rect 9002 4098 9054 4119
rect 9002 4067 9003 4098
rect 9003 4067 9037 4098
rect 9037 4067 9054 4098
rect 9066 4098 9118 4119
rect 9066 4067 9075 4098
rect 9075 4067 9109 4098
rect 9109 4067 9118 4098
rect 9130 4098 9182 4119
rect 9130 4067 9147 4098
rect 9147 4067 9181 4098
rect 9181 4067 9182 4098
rect 9002 4025 9054 4054
rect 9002 4002 9003 4025
rect 9003 4002 9037 4025
rect 9037 4002 9054 4025
rect 9066 4025 9118 4054
rect 9066 4002 9075 4025
rect 9075 4002 9109 4025
rect 9109 4002 9118 4025
rect 9130 4025 9182 4054
rect 9130 4002 9147 4025
rect 9147 4002 9181 4025
rect 9181 4002 9182 4025
rect 9002 3952 9054 3989
rect 9002 3937 9003 3952
rect 9003 3937 9037 3952
rect 9037 3937 9054 3952
rect 9066 3952 9118 3989
rect 9066 3937 9075 3952
rect 9075 3937 9109 3952
rect 9109 3937 9118 3952
rect 9130 3952 9182 3989
rect 9130 3937 9147 3952
rect 9147 3937 9181 3952
rect 9181 3937 9182 3952
rect 9002 3918 9003 3924
rect 9003 3918 9037 3924
rect 9037 3918 9075 3924
rect 9075 3918 9109 3924
rect 9109 3918 9147 3924
rect 9147 3918 9181 3924
rect 9181 3918 9182 3924
rect 9002 3879 9182 3918
rect 9002 3845 9003 3879
rect 9003 3845 9037 3879
rect 9037 3845 9075 3879
rect 9075 3845 9109 3879
rect 9109 3845 9147 3879
rect 9147 3845 9181 3879
rect 9181 3845 9182 3879
rect 9002 3806 9182 3845
rect 9002 3772 9003 3806
rect 9003 3772 9037 3806
rect 9037 3772 9075 3806
rect 9075 3772 9109 3806
rect 9109 3772 9147 3806
rect 9147 3772 9181 3806
rect 9181 3772 9182 3806
rect 9002 3733 9182 3772
rect 9002 3699 9003 3733
rect 9003 3699 9037 3733
rect 9037 3699 9075 3733
rect 9075 3699 9109 3733
rect 9109 3699 9147 3733
rect 9147 3699 9181 3733
rect 9181 3699 9182 3733
rect 9002 3660 9182 3699
rect 9002 3626 9003 3660
rect 9003 3626 9037 3660
rect 9037 3626 9075 3660
rect 9075 3626 9109 3660
rect 9109 3626 9147 3660
rect 9147 3626 9181 3660
rect 9181 3626 9182 3660
rect 9002 3587 9182 3626
rect 9002 3553 9003 3587
rect 9003 3553 9037 3587
rect 9037 3553 9075 3587
rect 9075 3553 9109 3587
rect 9109 3553 9147 3587
rect 9147 3553 9181 3587
rect 9181 3553 9182 3587
rect 9002 3514 9182 3553
rect 9002 3480 9003 3514
rect 9003 3480 9037 3514
rect 9037 3480 9075 3514
rect 9075 3480 9109 3514
rect 9109 3480 9147 3514
rect 9147 3480 9181 3514
rect 9181 3480 9182 3514
rect 9002 3441 9182 3480
rect 9002 3407 9003 3441
rect 9003 3407 9037 3441
rect 9037 3407 9075 3441
rect 9075 3407 9109 3441
rect 9109 3407 9147 3441
rect 9147 3407 9181 3441
rect 9181 3407 9182 3441
rect 9002 3368 9182 3407
rect 9002 3334 9003 3368
rect 9003 3334 9037 3368
rect 9037 3334 9075 3368
rect 9075 3334 9109 3368
rect 9109 3334 9147 3368
rect 9147 3334 9181 3368
rect 9181 3334 9182 3368
rect 9002 3295 9182 3334
rect 9002 3261 9003 3295
rect 9003 3261 9037 3295
rect 9037 3261 9075 3295
rect 9075 3261 9109 3295
rect 9109 3261 9147 3295
rect 9147 3261 9181 3295
rect 9181 3261 9182 3295
rect 9002 3222 9182 3261
rect 9002 3188 9003 3222
rect 9003 3188 9037 3222
rect 9037 3188 9075 3222
rect 9075 3188 9109 3222
rect 9109 3188 9147 3222
rect 9147 3188 9181 3222
rect 9181 3188 9182 3222
rect 9002 3149 9182 3188
rect 9002 3115 9003 3149
rect 9003 3115 9037 3149
rect 9037 3115 9075 3149
rect 9075 3115 9109 3149
rect 9109 3115 9147 3149
rect 9147 3115 9181 3149
rect 9181 3115 9182 3149
rect 9002 3076 9182 3115
rect 9002 3042 9003 3076
rect 9003 3042 9037 3076
rect 9037 3042 9075 3076
rect 9075 3042 9109 3076
rect 9109 3042 9147 3076
rect 9147 3042 9181 3076
rect 9181 3042 9182 3076
rect 9002 3003 9182 3042
rect 9002 2969 9003 3003
rect 9003 2969 9037 3003
rect 9037 2969 9075 3003
rect 9075 2969 9109 3003
rect 9109 2969 9147 3003
rect 9147 2969 9181 3003
rect 9181 2969 9182 3003
rect 9002 2930 9182 2969
rect 9002 2896 9003 2930
rect 9003 2896 9037 2930
rect 9037 2896 9075 2930
rect 9075 2896 9109 2930
rect 9109 2896 9147 2930
rect 9147 2896 9181 2930
rect 9181 2896 9182 2930
rect 9002 2857 9182 2896
rect 9002 2823 9003 2857
rect 9003 2823 9037 2857
rect 9037 2823 9075 2857
rect 9075 2823 9109 2857
rect 9109 2823 9147 2857
rect 9147 2823 9181 2857
rect 9181 2823 9182 2857
rect 9002 2784 9182 2823
rect 9002 2750 9003 2784
rect 9003 2750 9037 2784
rect 9037 2750 9075 2784
rect 9075 2750 9109 2784
rect 9109 2750 9147 2784
rect 9147 2750 9181 2784
rect 9181 2750 9182 2784
rect 9002 2711 9182 2750
rect 9002 2677 9003 2711
rect 9003 2677 9037 2711
rect 9037 2677 9075 2711
rect 9075 2677 9109 2711
rect 9109 2677 9147 2711
rect 9147 2677 9181 2711
rect 9181 2677 9182 2711
rect 9002 2638 9182 2677
rect 9002 2604 9003 2638
rect 9003 2604 9037 2638
rect 9037 2604 9075 2638
rect 9075 2604 9109 2638
rect 9109 2604 9147 2638
rect 9147 2604 9181 2638
rect 9181 2604 9182 2638
rect 9002 2565 9182 2604
rect 9002 2531 9003 2565
rect 9003 2531 9037 2565
rect 9037 2531 9075 2565
rect 9075 2531 9109 2565
rect 9109 2531 9147 2565
rect 9147 2531 9181 2565
rect 9181 2531 9182 2565
rect 9002 2492 9182 2531
rect 9002 2458 9003 2492
rect 9003 2458 9037 2492
rect 9037 2458 9075 2492
rect 9075 2458 9109 2492
rect 9109 2458 9147 2492
rect 9147 2458 9181 2492
rect 9181 2458 9182 2492
rect 9002 2419 9182 2458
rect 9002 2385 9003 2419
rect 9003 2385 9037 2419
rect 9037 2385 9075 2419
rect 9075 2385 9109 2419
rect 9109 2385 9147 2419
rect 9147 2385 9181 2419
rect 9181 2385 9182 2419
rect 9002 2346 9182 2385
rect 9002 2312 9003 2346
rect 9003 2312 9037 2346
rect 9037 2312 9075 2346
rect 9075 2312 9109 2346
rect 9109 2312 9147 2346
rect 9147 2312 9181 2346
rect 9181 2312 9182 2346
rect 9002 2273 9182 2312
rect 9002 2239 9003 2273
rect 9003 2239 9037 2273
rect 9037 2239 9075 2273
rect 9075 2239 9109 2273
rect 9109 2239 9147 2273
rect 9147 2239 9181 2273
rect 9181 2239 9182 2273
rect 9002 2200 9182 2239
rect 9002 2166 9003 2200
rect 9003 2166 9037 2200
rect 9037 2166 9075 2200
rect 9075 2166 9109 2200
rect 9109 2166 9147 2200
rect 9147 2166 9181 2200
rect 9181 2166 9182 2200
rect 9002 2126 9182 2166
rect 9002 2092 9003 2126
rect 9003 2092 9037 2126
rect 9037 2092 9075 2126
rect 9075 2092 9109 2126
rect 9109 2092 9147 2126
rect 9147 2092 9181 2126
rect 9181 2092 9182 2126
rect 9002 2052 9182 2092
rect 9002 2018 9003 2052
rect 9003 2018 9037 2052
rect 9037 2018 9075 2052
rect 9075 2018 9109 2052
rect 9109 2018 9147 2052
rect 9147 2018 9181 2052
rect 9181 2018 9182 2052
rect 9002 1978 9182 2018
rect 9002 1944 9003 1978
rect 9003 1944 9037 1978
rect 9037 1944 9075 1978
rect 9075 1944 9109 1978
rect 9109 1944 9147 1978
rect 9147 1944 9181 1978
rect 9181 1944 9182 1978
rect 9002 1904 9182 1944
rect 9002 1870 9003 1904
rect 9003 1870 9037 1904
rect 9037 1870 9075 1904
rect 9075 1870 9109 1904
rect 9109 1870 9147 1904
rect 9147 1870 9181 1904
rect 9181 1870 9182 1904
rect 9002 1830 9182 1870
rect 9002 1796 9003 1830
rect 9003 1796 9037 1830
rect 9037 1796 9075 1830
rect 9075 1796 9109 1830
rect 9109 1796 9147 1830
rect 9147 1796 9181 1830
rect 9181 1796 9182 1830
rect 9002 1756 9182 1796
rect 9002 1722 9003 1756
rect 9003 1722 9037 1756
rect 9037 1722 9075 1756
rect 9075 1722 9109 1756
rect 9109 1722 9147 1756
rect 9147 1722 9181 1756
rect 9181 1722 9182 1756
rect 9002 1682 9182 1722
rect 9002 1648 9003 1682
rect 9003 1648 9037 1682
rect 9037 1648 9075 1682
rect 9075 1648 9109 1682
rect 9109 1648 9147 1682
rect 9147 1648 9181 1682
rect 9181 1648 9182 1682
rect 9002 1608 9182 1648
rect 9002 1574 9003 1608
rect 9003 1574 9037 1608
rect 9037 1574 9075 1608
rect 9075 1574 9109 1608
rect 9109 1574 9147 1608
rect 9147 1574 9181 1608
rect 9181 1574 9182 1608
rect 9002 1568 9182 1574
rect 9498 4092 9550 4124
rect 9498 4072 9499 4092
rect 9499 4072 9533 4092
rect 9533 4072 9550 4092
rect 9562 4072 9614 4124
rect 9626 4092 9678 4124
rect 9626 4072 9643 4092
rect 9643 4072 9677 4092
rect 9677 4072 9678 4092
rect 9498 4058 9499 4059
rect 9499 4058 9533 4059
rect 9533 4058 9550 4059
rect 9498 4020 9550 4058
rect 9498 4007 9499 4020
rect 9499 4007 9533 4020
rect 9533 4007 9550 4020
rect 9562 4007 9614 4059
rect 9626 4058 9643 4059
rect 9643 4058 9677 4059
rect 9677 4058 9678 4059
rect 9626 4020 9678 4058
rect 9626 4007 9643 4020
rect 9643 4007 9677 4020
rect 9677 4007 9678 4020
rect 9498 3986 9499 3994
rect 9499 3986 9533 3994
rect 9533 3986 9550 3994
rect 9498 3948 9550 3986
rect 9498 3942 9499 3948
rect 9499 3942 9533 3948
rect 9533 3942 9550 3948
rect 9562 3942 9614 3994
rect 9626 3986 9643 3994
rect 9643 3986 9677 3994
rect 9677 3986 9678 3994
rect 9626 3948 9678 3986
rect 9626 3942 9643 3948
rect 9643 3942 9677 3948
rect 9677 3942 9678 3948
rect 9498 3914 9499 3929
rect 9499 3914 9533 3929
rect 9533 3914 9550 3929
rect 9498 3877 9550 3914
rect 9562 3877 9614 3929
rect 9626 3914 9643 3929
rect 9643 3914 9677 3929
rect 9677 3914 9678 3929
rect 9626 3877 9678 3914
rect 9498 3842 9499 3864
rect 9499 3842 9533 3864
rect 9533 3842 9550 3864
rect 9498 3812 9550 3842
rect 9562 3812 9614 3864
rect 9626 3842 9643 3864
rect 9643 3842 9677 3864
rect 9677 3842 9678 3864
rect 9626 3812 9678 3842
rect 9498 3770 9499 3799
rect 9499 3770 9533 3799
rect 9533 3770 9550 3799
rect 9498 3747 9550 3770
rect 9562 3747 9614 3799
rect 9626 3770 9643 3799
rect 9643 3770 9677 3799
rect 9677 3770 9678 3799
rect 9626 3747 9678 3770
rect 9498 3732 9550 3734
rect 9498 3698 9499 3732
rect 9499 3698 9533 3732
rect 9533 3698 9550 3732
rect 9498 3682 9550 3698
rect 9562 3682 9614 3734
rect 9626 3732 9678 3734
rect 9626 3698 9643 3732
rect 9643 3698 9677 3732
rect 9677 3698 9678 3732
rect 9626 3682 9678 3698
rect 9498 3660 9550 3669
rect 9498 3626 9499 3660
rect 9499 3626 9533 3660
rect 9533 3626 9550 3660
rect 9498 3617 9550 3626
rect 9562 3617 9614 3669
rect 9626 3660 9678 3669
rect 9626 3626 9643 3660
rect 9643 3626 9677 3660
rect 9677 3626 9678 3660
rect 9626 3617 9678 3626
rect 9498 3588 9678 3604
rect 9498 3554 9499 3588
rect 9499 3554 9533 3588
rect 9533 3554 9643 3588
rect 9643 3554 9677 3588
rect 9677 3554 9678 3588
rect 9498 3516 9678 3554
rect 9498 3482 9499 3516
rect 9499 3482 9533 3516
rect 9533 3482 9643 3516
rect 9643 3482 9677 3516
rect 9677 3482 9678 3516
rect 9498 3444 9678 3482
rect 9498 3410 9499 3444
rect 9499 3410 9533 3444
rect 9533 3410 9643 3444
rect 9643 3410 9677 3444
rect 9677 3410 9678 3444
rect 9498 3372 9678 3410
rect 9498 3338 9499 3372
rect 9499 3338 9533 3372
rect 9533 3338 9643 3372
rect 9643 3338 9677 3372
rect 9677 3338 9678 3372
rect 9498 3300 9678 3338
rect 9498 3266 9499 3300
rect 9499 3266 9533 3300
rect 9533 3266 9643 3300
rect 9643 3266 9677 3300
rect 9677 3266 9678 3300
rect 9498 3228 9678 3266
rect 9498 3194 9499 3228
rect 9499 3194 9533 3228
rect 9533 3194 9643 3228
rect 9643 3194 9677 3228
rect 9677 3194 9678 3228
rect 9498 3108 9678 3194
rect 9498 3074 9499 3108
rect 9499 3074 9533 3108
rect 9533 3074 9571 3108
rect 9571 3074 9605 3108
rect 9605 3074 9643 3108
rect 9643 3074 9677 3108
rect 9677 3074 9678 3108
rect 9498 3028 9678 3074
rect 9498 2994 9499 3028
rect 9499 2994 9533 3028
rect 9533 2994 9571 3028
rect 9571 2994 9605 3028
rect 9605 2994 9643 3028
rect 9643 2994 9677 3028
rect 9677 2994 9678 3028
rect 9498 2948 9678 2994
rect 9498 2914 9499 2948
rect 9499 2914 9533 2948
rect 9533 2914 9571 2948
rect 9571 2914 9605 2948
rect 9605 2914 9643 2948
rect 9643 2914 9677 2948
rect 9677 2914 9678 2948
rect 9498 2868 9678 2914
rect 9498 2834 9499 2868
rect 9499 2834 9533 2868
rect 9533 2834 9571 2868
rect 9571 2834 9605 2868
rect 9605 2834 9643 2868
rect 9643 2834 9677 2868
rect 9677 2834 9678 2868
rect 9498 2788 9678 2834
rect 9498 2754 9499 2788
rect 9499 2754 9533 2788
rect 9533 2754 9571 2788
rect 9571 2754 9605 2788
rect 9605 2754 9643 2788
rect 9643 2754 9677 2788
rect 9677 2754 9678 2788
rect 9498 2708 9678 2754
rect 9498 2674 9499 2708
rect 9499 2674 9533 2708
rect 9533 2674 9571 2708
rect 9571 2674 9605 2708
rect 9605 2674 9643 2708
rect 9643 2674 9677 2708
rect 9677 2674 9678 2708
rect 9498 2628 9678 2674
rect 9498 2594 9499 2628
rect 9499 2594 9533 2628
rect 9533 2594 9571 2628
rect 9571 2594 9605 2628
rect 9605 2594 9643 2628
rect 9643 2594 9677 2628
rect 9677 2594 9678 2628
rect 9498 2518 9678 2594
rect 9498 2484 9499 2518
rect 9499 2484 9533 2518
rect 9533 2484 9643 2518
rect 9643 2484 9677 2518
rect 9677 2484 9678 2518
rect 9498 2446 9678 2484
rect 9498 2412 9499 2446
rect 9499 2412 9533 2446
rect 9533 2412 9643 2446
rect 9643 2412 9677 2446
rect 9677 2412 9678 2446
rect 9498 2374 9678 2412
rect 9498 2340 9499 2374
rect 9499 2340 9533 2374
rect 9533 2340 9643 2374
rect 9643 2340 9677 2374
rect 9677 2340 9678 2374
rect 9498 2302 9678 2340
rect 9498 2268 9499 2302
rect 9499 2268 9533 2302
rect 9533 2268 9643 2302
rect 9643 2268 9677 2302
rect 9677 2268 9678 2302
rect 9498 2230 9678 2268
rect 9498 2196 9499 2230
rect 9499 2196 9533 2230
rect 9533 2196 9643 2230
rect 9643 2196 9677 2230
rect 9677 2196 9678 2230
rect 9498 2158 9678 2196
rect 9498 2124 9499 2158
rect 9499 2124 9533 2158
rect 9533 2124 9643 2158
rect 9643 2124 9677 2158
rect 9677 2124 9678 2158
rect 9498 2086 9678 2124
rect 9498 2052 9499 2086
rect 9499 2052 9533 2086
rect 9533 2052 9643 2086
rect 9643 2052 9677 2086
rect 9677 2052 9678 2086
rect 9498 2014 9678 2052
rect 9498 1980 9499 2014
rect 9499 1980 9533 2014
rect 9533 1980 9643 2014
rect 9643 1980 9677 2014
rect 9677 1980 9678 2014
rect 9498 1942 9678 1980
rect 9498 1908 9499 1942
rect 9499 1908 9533 1942
rect 9533 1908 9643 1942
rect 9643 1908 9677 1942
rect 9677 1908 9678 1942
rect 9498 1870 9678 1908
rect 9498 1836 9499 1870
rect 9499 1836 9533 1870
rect 9533 1836 9643 1870
rect 9643 1836 9677 1870
rect 9677 1836 9678 1870
rect 9498 1798 9678 1836
rect 9498 1764 9499 1798
rect 9499 1764 9533 1798
rect 9533 1764 9643 1798
rect 9643 1764 9677 1798
rect 9677 1764 9678 1798
rect 9498 1726 9678 1764
rect 9498 1692 9499 1726
rect 9499 1692 9533 1726
rect 9533 1692 9643 1726
rect 9643 1692 9677 1726
rect 9677 1692 9678 1726
rect 9498 1654 9678 1692
rect 9498 1620 9499 1654
rect 9499 1620 9533 1654
rect 9533 1620 9643 1654
rect 9643 1620 9677 1654
rect 9677 1620 9678 1654
rect 9498 1568 9678 1620
rect 9994 4098 10046 4119
rect 9994 4067 9995 4098
rect 9995 4067 10029 4098
rect 10029 4067 10046 4098
rect 10058 4098 10110 4119
rect 10058 4067 10067 4098
rect 10067 4067 10101 4098
rect 10101 4067 10110 4098
rect 10122 4098 10174 4119
rect 10122 4067 10139 4098
rect 10139 4067 10173 4098
rect 10173 4067 10174 4098
rect 9994 4025 10046 4054
rect 9994 4002 9995 4025
rect 9995 4002 10029 4025
rect 10029 4002 10046 4025
rect 10058 4025 10110 4054
rect 10058 4002 10067 4025
rect 10067 4002 10101 4025
rect 10101 4002 10110 4025
rect 10122 4025 10174 4054
rect 10122 4002 10139 4025
rect 10139 4002 10173 4025
rect 10173 4002 10174 4025
rect 9994 3952 10046 3989
rect 9994 3937 9995 3952
rect 9995 3937 10029 3952
rect 10029 3937 10046 3952
rect 10058 3952 10110 3989
rect 10058 3937 10067 3952
rect 10067 3937 10101 3952
rect 10101 3937 10110 3952
rect 10122 3952 10174 3989
rect 10122 3937 10139 3952
rect 10139 3937 10173 3952
rect 10173 3937 10174 3952
rect 9994 3918 9995 3924
rect 9995 3918 10029 3924
rect 10029 3918 10067 3924
rect 10067 3918 10101 3924
rect 10101 3918 10139 3924
rect 10139 3918 10173 3924
rect 10173 3918 10174 3924
rect 9994 3879 10174 3918
rect 9994 3845 9995 3879
rect 9995 3845 10029 3879
rect 10029 3845 10067 3879
rect 10067 3845 10101 3879
rect 10101 3845 10139 3879
rect 10139 3845 10173 3879
rect 10173 3845 10174 3879
rect 9994 3806 10174 3845
rect 9994 3772 9995 3806
rect 9995 3772 10029 3806
rect 10029 3772 10067 3806
rect 10067 3772 10101 3806
rect 10101 3772 10139 3806
rect 10139 3772 10173 3806
rect 10173 3772 10174 3806
rect 9994 3733 10174 3772
rect 9994 3699 9995 3733
rect 9995 3699 10029 3733
rect 10029 3699 10067 3733
rect 10067 3699 10101 3733
rect 10101 3699 10139 3733
rect 10139 3699 10173 3733
rect 10173 3699 10174 3733
rect 9994 3660 10174 3699
rect 9994 3626 9995 3660
rect 9995 3626 10029 3660
rect 10029 3626 10067 3660
rect 10067 3626 10101 3660
rect 10101 3626 10139 3660
rect 10139 3626 10173 3660
rect 10173 3626 10174 3660
rect 9994 3587 10174 3626
rect 9994 3553 9995 3587
rect 9995 3553 10029 3587
rect 10029 3553 10067 3587
rect 10067 3553 10101 3587
rect 10101 3553 10139 3587
rect 10139 3553 10173 3587
rect 10173 3553 10174 3587
rect 9994 3514 10174 3553
rect 9994 3480 9995 3514
rect 9995 3480 10029 3514
rect 10029 3480 10067 3514
rect 10067 3480 10101 3514
rect 10101 3480 10139 3514
rect 10139 3480 10173 3514
rect 10173 3480 10174 3514
rect 9994 3441 10174 3480
rect 9994 3407 9995 3441
rect 9995 3407 10029 3441
rect 10029 3407 10067 3441
rect 10067 3407 10101 3441
rect 10101 3407 10139 3441
rect 10139 3407 10173 3441
rect 10173 3407 10174 3441
rect 9994 3368 10174 3407
rect 9994 3334 9995 3368
rect 9995 3334 10029 3368
rect 10029 3334 10067 3368
rect 10067 3334 10101 3368
rect 10101 3334 10139 3368
rect 10139 3334 10173 3368
rect 10173 3334 10174 3368
rect 9994 3295 10174 3334
rect 9994 3261 9995 3295
rect 9995 3261 10029 3295
rect 10029 3261 10067 3295
rect 10067 3261 10101 3295
rect 10101 3261 10139 3295
rect 10139 3261 10173 3295
rect 10173 3261 10174 3295
rect 9994 3222 10174 3261
rect 9994 3188 9995 3222
rect 9995 3188 10029 3222
rect 10029 3188 10067 3222
rect 10067 3188 10101 3222
rect 10101 3188 10139 3222
rect 10139 3188 10173 3222
rect 10173 3188 10174 3222
rect 9994 3149 10174 3188
rect 9994 3115 9995 3149
rect 9995 3115 10029 3149
rect 10029 3115 10067 3149
rect 10067 3115 10101 3149
rect 10101 3115 10139 3149
rect 10139 3115 10173 3149
rect 10173 3115 10174 3149
rect 9994 3076 10174 3115
rect 9994 3042 9995 3076
rect 9995 3042 10029 3076
rect 10029 3042 10067 3076
rect 10067 3042 10101 3076
rect 10101 3042 10139 3076
rect 10139 3042 10173 3076
rect 10173 3042 10174 3076
rect 9994 3003 10174 3042
rect 9994 2969 9995 3003
rect 9995 2969 10029 3003
rect 10029 2969 10067 3003
rect 10067 2969 10101 3003
rect 10101 2969 10139 3003
rect 10139 2969 10173 3003
rect 10173 2969 10174 3003
rect 9994 2930 10174 2969
rect 9994 2896 9995 2930
rect 9995 2896 10029 2930
rect 10029 2896 10067 2930
rect 10067 2896 10101 2930
rect 10101 2896 10139 2930
rect 10139 2896 10173 2930
rect 10173 2896 10174 2930
rect 9994 2857 10174 2896
rect 9994 2823 9995 2857
rect 9995 2823 10029 2857
rect 10029 2823 10067 2857
rect 10067 2823 10101 2857
rect 10101 2823 10139 2857
rect 10139 2823 10173 2857
rect 10173 2823 10174 2857
rect 9994 2784 10174 2823
rect 9994 2750 9995 2784
rect 9995 2750 10029 2784
rect 10029 2750 10067 2784
rect 10067 2750 10101 2784
rect 10101 2750 10139 2784
rect 10139 2750 10173 2784
rect 10173 2750 10174 2784
rect 9994 2711 10174 2750
rect 9994 2677 9995 2711
rect 9995 2677 10029 2711
rect 10029 2677 10067 2711
rect 10067 2677 10101 2711
rect 10101 2677 10139 2711
rect 10139 2677 10173 2711
rect 10173 2677 10174 2711
rect 9994 2638 10174 2677
rect 9994 2604 9995 2638
rect 9995 2604 10029 2638
rect 10029 2604 10067 2638
rect 10067 2604 10101 2638
rect 10101 2604 10139 2638
rect 10139 2604 10173 2638
rect 10173 2604 10174 2638
rect 9994 2565 10174 2604
rect 9994 2531 9995 2565
rect 9995 2531 10029 2565
rect 10029 2531 10067 2565
rect 10067 2531 10101 2565
rect 10101 2531 10139 2565
rect 10139 2531 10173 2565
rect 10173 2531 10174 2565
rect 9994 2492 10174 2531
rect 9994 2458 9995 2492
rect 9995 2458 10029 2492
rect 10029 2458 10067 2492
rect 10067 2458 10101 2492
rect 10101 2458 10139 2492
rect 10139 2458 10173 2492
rect 10173 2458 10174 2492
rect 9994 2419 10174 2458
rect 9994 2385 9995 2419
rect 9995 2385 10029 2419
rect 10029 2385 10067 2419
rect 10067 2385 10101 2419
rect 10101 2385 10139 2419
rect 10139 2385 10173 2419
rect 10173 2385 10174 2419
rect 9994 2346 10174 2385
rect 9994 2312 9995 2346
rect 9995 2312 10029 2346
rect 10029 2312 10067 2346
rect 10067 2312 10101 2346
rect 10101 2312 10139 2346
rect 10139 2312 10173 2346
rect 10173 2312 10174 2346
rect 9994 2273 10174 2312
rect 9994 2239 9995 2273
rect 9995 2239 10029 2273
rect 10029 2239 10067 2273
rect 10067 2239 10101 2273
rect 10101 2239 10139 2273
rect 10139 2239 10173 2273
rect 10173 2239 10174 2273
rect 9994 2200 10174 2239
rect 9994 2166 9995 2200
rect 9995 2166 10029 2200
rect 10029 2166 10067 2200
rect 10067 2166 10101 2200
rect 10101 2166 10139 2200
rect 10139 2166 10173 2200
rect 10173 2166 10174 2200
rect 9994 2126 10174 2166
rect 9994 2092 9995 2126
rect 9995 2092 10029 2126
rect 10029 2092 10067 2126
rect 10067 2092 10101 2126
rect 10101 2092 10139 2126
rect 10139 2092 10173 2126
rect 10173 2092 10174 2126
rect 9994 2052 10174 2092
rect 9994 2018 9995 2052
rect 9995 2018 10029 2052
rect 10029 2018 10067 2052
rect 10067 2018 10101 2052
rect 10101 2018 10139 2052
rect 10139 2018 10173 2052
rect 10173 2018 10174 2052
rect 9994 1978 10174 2018
rect 9994 1944 9995 1978
rect 9995 1944 10029 1978
rect 10029 1944 10067 1978
rect 10067 1944 10101 1978
rect 10101 1944 10139 1978
rect 10139 1944 10173 1978
rect 10173 1944 10174 1978
rect 9994 1904 10174 1944
rect 9994 1870 9995 1904
rect 9995 1870 10029 1904
rect 10029 1870 10067 1904
rect 10067 1870 10101 1904
rect 10101 1870 10139 1904
rect 10139 1870 10173 1904
rect 10173 1870 10174 1904
rect 9994 1830 10174 1870
rect 9994 1796 9995 1830
rect 9995 1796 10029 1830
rect 10029 1796 10067 1830
rect 10067 1796 10101 1830
rect 10101 1796 10139 1830
rect 10139 1796 10173 1830
rect 10173 1796 10174 1830
rect 9994 1756 10174 1796
rect 9994 1722 9995 1756
rect 9995 1722 10029 1756
rect 10029 1722 10067 1756
rect 10067 1722 10101 1756
rect 10101 1722 10139 1756
rect 10139 1722 10173 1756
rect 10173 1722 10174 1756
rect 9994 1682 10174 1722
rect 9994 1648 9995 1682
rect 9995 1648 10029 1682
rect 10029 1648 10067 1682
rect 10067 1648 10101 1682
rect 10101 1648 10139 1682
rect 10139 1648 10173 1682
rect 10173 1648 10174 1682
rect 9994 1608 10174 1648
rect 9994 1574 9995 1608
rect 9995 1574 10029 1608
rect 10029 1574 10067 1608
rect 10067 1574 10101 1608
rect 10101 1574 10139 1608
rect 10139 1574 10173 1608
rect 10173 1574 10174 1608
rect 9994 1568 10174 1574
rect 10490 4092 10542 4124
rect 10490 4072 10491 4092
rect 10491 4072 10525 4092
rect 10525 4072 10542 4092
rect 10554 4072 10606 4124
rect 10618 4092 10670 4124
rect 10618 4072 10635 4092
rect 10635 4072 10669 4092
rect 10669 4072 10670 4092
rect 10490 4058 10491 4059
rect 10491 4058 10525 4059
rect 10525 4058 10542 4059
rect 10490 4020 10542 4058
rect 10490 4007 10491 4020
rect 10491 4007 10525 4020
rect 10525 4007 10542 4020
rect 10554 4007 10606 4059
rect 10618 4058 10635 4059
rect 10635 4058 10669 4059
rect 10669 4058 10670 4059
rect 10618 4020 10670 4058
rect 10618 4007 10635 4020
rect 10635 4007 10669 4020
rect 10669 4007 10670 4020
rect 10490 3986 10491 3994
rect 10491 3986 10525 3994
rect 10525 3986 10542 3994
rect 10490 3948 10542 3986
rect 10490 3942 10491 3948
rect 10491 3942 10525 3948
rect 10525 3942 10542 3948
rect 10554 3942 10606 3994
rect 10618 3986 10635 3994
rect 10635 3986 10669 3994
rect 10669 3986 10670 3994
rect 10618 3948 10670 3986
rect 10618 3942 10635 3948
rect 10635 3942 10669 3948
rect 10669 3942 10670 3948
rect 10490 3914 10491 3929
rect 10491 3914 10525 3929
rect 10525 3914 10542 3929
rect 10490 3877 10542 3914
rect 10554 3877 10606 3929
rect 10618 3914 10635 3929
rect 10635 3914 10669 3929
rect 10669 3914 10670 3929
rect 10618 3877 10670 3914
rect 10490 3842 10491 3864
rect 10491 3842 10525 3864
rect 10525 3842 10542 3864
rect 10490 3812 10542 3842
rect 10554 3812 10606 3864
rect 10618 3842 10635 3864
rect 10635 3842 10669 3864
rect 10669 3842 10670 3864
rect 10618 3812 10670 3842
rect 10490 3770 10491 3799
rect 10491 3770 10525 3799
rect 10525 3770 10542 3799
rect 10490 3747 10542 3770
rect 10554 3747 10606 3799
rect 10618 3770 10635 3799
rect 10635 3770 10669 3799
rect 10669 3770 10670 3799
rect 10618 3747 10670 3770
rect 10490 3732 10542 3734
rect 10490 3698 10491 3732
rect 10491 3698 10525 3732
rect 10525 3698 10542 3732
rect 10490 3682 10542 3698
rect 10554 3682 10606 3734
rect 10618 3732 10670 3734
rect 10618 3698 10635 3732
rect 10635 3698 10669 3732
rect 10669 3698 10670 3732
rect 10618 3682 10670 3698
rect 10490 3660 10542 3669
rect 10490 3626 10491 3660
rect 10491 3626 10525 3660
rect 10525 3626 10542 3660
rect 10490 3617 10542 3626
rect 10554 3617 10606 3669
rect 10618 3660 10670 3669
rect 10618 3626 10635 3660
rect 10635 3626 10669 3660
rect 10669 3626 10670 3660
rect 10618 3617 10670 3626
rect 10490 3588 10670 3604
rect 10490 3554 10491 3588
rect 10491 3554 10525 3588
rect 10525 3554 10635 3588
rect 10635 3554 10669 3588
rect 10669 3554 10670 3588
rect 10490 3516 10670 3554
rect 10490 3482 10491 3516
rect 10491 3482 10525 3516
rect 10525 3482 10635 3516
rect 10635 3482 10669 3516
rect 10669 3482 10670 3516
rect 10490 3444 10670 3482
rect 10490 3410 10491 3444
rect 10491 3410 10525 3444
rect 10525 3410 10635 3444
rect 10635 3410 10669 3444
rect 10669 3410 10670 3444
rect 10490 3372 10670 3410
rect 10490 3338 10491 3372
rect 10491 3338 10525 3372
rect 10525 3338 10635 3372
rect 10635 3338 10669 3372
rect 10669 3338 10670 3372
rect 10490 3300 10670 3338
rect 10490 3266 10491 3300
rect 10491 3266 10525 3300
rect 10525 3266 10635 3300
rect 10635 3266 10669 3300
rect 10669 3266 10670 3300
rect 10490 3228 10670 3266
rect 10490 3194 10491 3228
rect 10491 3194 10525 3228
rect 10525 3194 10635 3228
rect 10635 3194 10669 3228
rect 10669 3194 10670 3228
rect 10490 3108 10670 3194
rect 10490 3074 10491 3108
rect 10491 3074 10525 3108
rect 10525 3074 10563 3108
rect 10563 3074 10597 3108
rect 10597 3074 10635 3108
rect 10635 3074 10669 3108
rect 10669 3074 10670 3108
rect 10490 3028 10670 3074
rect 10490 2994 10491 3028
rect 10491 2994 10525 3028
rect 10525 2994 10563 3028
rect 10563 2994 10597 3028
rect 10597 2994 10635 3028
rect 10635 2994 10669 3028
rect 10669 2994 10670 3028
rect 10490 2948 10670 2994
rect 10490 2914 10491 2948
rect 10491 2914 10525 2948
rect 10525 2914 10563 2948
rect 10563 2914 10597 2948
rect 10597 2914 10635 2948
rect 10635 2914 10669 2948
rect 10669 2914 10670 2948
rect 10490 2868 10670 2914
rect 10490 2834 10491 2868
rect 10491 2834 10525 2868
rect 10525 2834 10563 2868
rect 10563 2834 10597 2868
rect 10597 2834 10635 2868
rect 10635 2834 10669 2868
rect 10669 2834 10670 2868
rect 10490 2788 10670 2834
rect 10490 2754 10491 2788
rect 10491 2754 10525 2788
rect 10525 2754 10563 2788
rect 10563 2754 10597 2788
rect 10597 2754 10635 2788
rect 10635 2754 10669 2788
rect 10669 2754 10670 2788
rect 10490 2708 10670 2754
rect 10490 2674 10491 2708
rect 10491 2674 10525 2708
rect 10525 2674 10563 2708
rect 10563 2674 10597 2708
rect 10597 2674 10635 2708
rect 10635 2674 10669 2708
rect 10669 2674 10670 2708
rect 10490 2628 10670 2674
rect 10490 2594 10491 2628
rect 10491 2594 10525 2628
rect 10525 2594 10563 2628
rect 10563 2594 10597 2628
rect 10597 2594 10635 2628
rect 10635 2594 10669 2628
rect 10669 2594 10670 2628
rect 10490 2518 10670 2594
rect 10490 2484 10491 2518
rect 10491 2484 10525 2518
rect 10525 2484 10635 2518
rect 10635 2484 10669 2518
rect 10669 2484 10670 2518
rect 10490 2446 10670 2484
rect 10490 2412 10491 2446
rect 10491 2412 10525 2446
rect 10525 2412 10635 2446
rect 10635 2412 10669 2446
rect 10669 2412 10670 2446
rect 10490 2374 10670 2412
rect 10490 2340 10491 2374
rect 10491 2340 10525 2374
rect 10525 2340 10635 2374
rect 10635 2340 10669 2374
rect 10669 2340 10670 2374
rect 10490 2302 10670 2340
rect 10490 2268 10491 2302
rect 10491 2268 10525 2302
rect 10525 2268 10635 2302
rect 10635 2268 10669 2302
rect 10669 2268 10670 2302
rect 10490 2230 10670 2268
rect 10490 2196 10491 2230
rect 10491 2196 10525 2230
rect 10525 2196 10635 2230
rect 10635 2196 10669 2230
rect 10669 2196 10670 2230
rect 10490 2158 10670 2196
rect 10490 2124 10491 2158
rect 10491 2124 10525 2158
rect 10525 2124 10635 2158
rect 10635 2124 10669 2158
rect 10669 2124 10670 2158
rect 10490 2086 10670 2124
rect 10490 2052 10491 2086
rect 10491 2052 10525 2086
rect 10525 2052 10635 2086
rect 10635 2052 10669 2086
rect 10669 2052 10670 2086
rect 10490 2014 10670 2052
rect 10490 1980 10491 2014
rect 10491 1980 10525 2014
rect 10525 1980 10635 2014
rect 10635 1980 10669 2014
rect 10669 1980 10670 2014
rect 10490 1942 10670 1980
rect 10490 1908 10491 1942
rect 10491 1908 10525 1942
rect 10525 1908 10635 1942
rect 10635 1908 10669 1942
rect 10669 1908 10670 1942
rect 10490 1870 10670 1908
rect 10490 1836 10491 1870
rect 10491 1836 10525 1870
rect 10525 1836 10635 1870
rect 10635 1836 10669 1870
rect 10669 1836 10670 1870
rect 10490 1798 10670 1836
rect 10490 1764 10491 1798
rect 10491 1764 10525 1798
rect 10525 1764 10635 1798
rect 10635 1764 10669 1798
rect 10669 1764 10670 1798
rect 10490 1726 10670 1764
rect 10490 1692 10491 1726
rect 10491 1692 10525 1726
rect 10525 1692 10635 1726
rect 10635 1692 10669 1726
rect 10669 1692 10670 1726
rect 10490 1654 10670 1692
rect 10490 1620 10491 1654
rect 10491 1620 10525 1654
rect 10525 1620 10635 1654
rect 10635 1620 10669 1654
rect 10669 1620 10670 1654
rect 10490 1568 10670 1620
rect 10986 4098 11038 4119
rect 10986 4067 10987 4098
rect 10987 4067 11021 4098
rect 11021 4067 11038 4098
rect 11050 4098 11102 4119
rect 11050 4067 11059 4098
rect 11059 4067 11093 4098
rect 11093 4067 11102 4098
rect 11114 4098 11166 4119
rect 11114 4067 11131 4098
rect 11131 4067 11165 4098
rect 11165 4067 11166 4098
rect 10986 4025 11038 4054
rect 10986 4002 10987 4025
rect 10987 4002 11021 4025
rect 11021 4002 11038 4025
rect 11050 4025 11102 4054
rect 11050 4002 11059 4025
rect 11059 4002 11093 4025
rect 11093 4002 11102 4025
rect 11114 4025 11166 4054
rect 11114 4002 11131 4025
rect 11131 4002 11165 4025
rect 11165 4002 11166 4025
rect 10986 3952 11038 3989
rect 10986 3937 10987 3952
rect 10987 3937 11021 3952
rect 11021 3937 11038 3952
rect 11050 3952 11102 3989
rect 11050 3937 11059 3952
rect 11059 3937 11093 3952
rect 11093 3937 11102 3952
rect 11114 3952 11166 3989
rect 11114 3937 11131 3952
rect 11131 3937 11165 3952
rect 11165 3937 11166 3952
rect 10986 3918 10987 3924
rect 10987 3918 11021 3924
rect 11021 3918 11059 3924
rect 11059 3918 11093 3924
rect 11093 3918 11131 3924
rect 11131 3918 11165 3924
rect 11165 3918 11166 3924
rect 10986 3879 11166 3918
rect 10986 3845 10987 3879
rect 10987 3845 11021 3879
rect 11021 3845 11059 3879
rect 11059 3845 11093 3879
rect 11093 3845 11131 3879
rect 11131 3845 11165 3879
rect 11165 3845 11166 3879
rect 10986 3806 11166 3845
rect 10986 3772 10987 3806
rect 10987 3772 11021 3806
rect 11021 3772 11059 3806
rect 11059 3772 11093 3806
rect 11093 3772 11131 3806
rect 11131 3772 11165 3806
rect 11165 3772 11166 3806
rect 10986 3733 11166 3772
rect 10986 3699 10987 3733
rect 10987 3699 11021 3733
rect 11021 3699 11059 3733
rect 11059 3699 11093 3733
rect 11093 3699 11131 3733
rect 11131 3699 11165 3733
rect 11165 3699 11166 3733
rect 10986 3660 11166 3699
rect 10986 3626 10987 3660
rect 10987 3626 11021 3660
rect 11021 3626 11059 3660
rect 11059 3626 11093 3660
rect 11093 3626 11131 3660
rect 11131 3626 11165 3660
rect 11165 3626 11166 3660
rect 10986 3587 11166 3626
rect 10986 3553 10987 3587
rect 10987 3553 11021 3587
rect 11021 3553 11059 3587
rect 11059 3553 11093 3587
rect 11093 3553 11131 3587
rect 11131 3553 11165 3587
rect 11165 3553 11166 3587
rect 10986 3514 11166 3553
rect 10986 3480 10987 3514
rect 10987 3480 11021 3514
rect 11021 3480 11059 3514
rect 11059 3480 11093 3514
rect 11093 3480 11131 3514
rect 11131 3480 11165 3514
rect 11165 3480 11166 3514
rect 10986 3441 11166 3480
rect 10986 3407 10987 3441
rect 10987 3407 11021 3441
rect 11021 3407 11059 3441
rect 11059 3407 11093 3441
rect 11093 3407 11131 3441
rect 11131 3407 11165 3441
rect 11165 3407 11166 3441
rect 10986 3368 11166 3407
rect 10986 3334 10987 3368
rect 10987 3334 11021 3368
rect 11021 3334 11059 3368
rect 11059 3334 11093 3368
rect 11093 3334 11131 3368
rect 11131 3334 11165 3368
rect 11165 3334 11166 3368
rect 10986 3295 11166 3334
rect 10986 3261 10987 3295
rect 10987 3261 11021 3295
rect 11021 3261 11059 3295
rect 11059 3261 11093 3295
rect 11093 3261 11131 3295
rect 11131 3261 11165 3295
rect 11165 3261 11166 3295
rect 10986 3222 11166 3261
rect 10986 3188 10987 3222
rect 10987 3188 11021 3222
rect 11021 3188 11059 3222
rect 11059 3188 11093 3222
rect 11093 3188 11131 3222
rect 11131 3188 11165 3222
rect 11165 3188 11166 3222
rect 10986 3149 11166 3188
rect 10986 3115 10987 3149
rect 10987 3115 11021 3149
rect 11021 3115 11059 3149
rect 11059 3115 11093 3149
rect 11093 3115 11131 3149
rect 11131 3115 11165 3149
rect 11165 3115 11166 3149
rect 10986 3076 11166 3115
rect 10986 3042 10987 3076
rect 10987 3042 11021 3076
rect 11021 3042 11059 3076
rect 11059 3042 11093 3076
rect 11093 3042 11131 3076
rect 11131 3042 11165 3076
rect 11165 3042 11166 3076
rect 10986 3003 11166 3042
rect 10986 2969 10987 3003
rect 10987 2969 11021 3003
rect 11021 2969 11059 3003
rect 11059 2969 11093 3003
rect 11093 2969 11131 3003
rect 11131 2969 11165 3003
rect 11165 2969 11166 3003
rect 10986 2930 11166 2969
rect 10986 2896 10987 2930
rect 10987 2896 11021 2930
rect 11021 2896 11059 2930
rect 11059 2896 11093 2930
rect 11093 2896 11131 2930
rect 11131 2896 11165 2930
rect 11165 2896 11166 2930
rect 10986 2857 11166 2896
rect 10986 2823 10987 2857
rect 10987 2823 11021 2857
rect 11021 2823 11059 2857
rect 11059 2823 11093 2857
rect 11093 2823 11131 2857
rect 11131 2823 11165 2857
rect 11165 2823 11166 2857
rect 10986 2784 11166 2823
rect 10986 2750 10987 2784
rect 10987 2750 11021 2784
rect 11021 2750 11059 2784
rect 11059 2750 11093 2784
rect 11093 2750 11131 2784
rect 11131 2750 11165 2784
rect 11165 2750 11166 2784
rect 10986 2711 11166 2750
rect 10986 2677 10987 2711
rect 10987 2677 11021 2711
rect 11021 2677 11059 2711
rect 11059 2677 11093 2711
rect 11093 2677 11131 2711
rect 11131 2677 11165 2711
rect 11165 2677 11166 2711
rect 10986 2638 11166 2677
rect 10986 2604 10987 2638
rect 10987 2604 11021 2638
rect 11021 2604 11059 2638
rect 11059 2604 11093 2638
rect 11093 2604 11131 2638
rect 11131 2604 11165 2638
rect 11165 2604 11166 2638
rect 10986 2565 11166 2604
rect 10986 2531 10987 2565
rect 10987 2531 11021 2565
rect 11021 2531 11059 2565
rect 11059 2531 11093 2565
rect 11093 2531 11131 2565
rect 11131 2531 11165 2565
rect 11165 2531 11166 2565
rect 10986 2492 11166 2531
rect 10986 2458 10987 2492
rect 10987 2458 11021 2492
rect 11021 2458 11059 2492
rect 11059 2458 11093 2492
rect 11093 2458 11131 2492
rect 11131 2458 11165 2492
rect 11165 2458 11166 2492
rect 10986 2419 11166 2458
rect 10986 2385 10987 2419
rect 10987 2385 11021 2419
rect 11021 2385 11059 2419
rect 11059 2385 11093 2419
rect 11093 2385 11131 2419
rect 11131 2385 11165 2419
rect 11165 2385 11166 2419
rect 10986 2346 11166 2385
rect 10986 2312 10987 2346
rect 10987 2312 11021 2346
rect 11021 2312 11059 2346
rect 11059 2312 11093 2346
rect 11093 2312 11131 2346
rect 11131 2312 11165 2346
rect 11165 2312 11166 2346
rect 10986 2273 11166 2312
rect 10986 2239 10987 2273
rect 10987 2239 11021 2273
rect 11021 2239 11059 2273
rect 11059 2239 11093 2273
rect 11093 2239 11131 2273
rect 11131 2239 11165 2273
rect 11165 2239 11166 2273
rect 10986 2200 11166 2239
rect 10986 2166 10987 2200
rect 10987 2166 11021 2200
rect 11021 2166 11059 2200
rect 11059 2166 11093 2200
rect 11093 2166 11131 2200
rect 11131 2166 11165 2200
rect 11165 2166 11166 2200
rect 10986 2126 11166 2166
rect 10986 2092 10987 2126
rect 10987 2092 11021 2126
rect 11021 2092 11059 2126
rect 11059 2092 11093 2126
rect 11093 2092 11131 2126
rect 11131 2092 11165 2126
rect 11165 2092 11166 2126
rect 10986 2052 11166 2092
rect 10986 2018 10987 2052
rect 10987 2018 11021 2052
rect 11021 2018 11059 2052
rect 11059 2018 11093 2052
rect 11093 2018 11131 2052
rect 11131 2018 11165 2052
rect 11165 2018 11166 2052
rect 10986 1978 11166 2018
rect 10986 1944 10987 1978
rect 10987 1944 11021 1978
rect 11021 1944 11059 1978
rect 11059 1944 11093 1978
rect 11093 1944 11131 1978
rect 11131 1944 11165 1978
rect 11165 1944 11166 1978
rect 10986 1904 11166 1944
rect 10986 1870 10987 1904
rect 10987 1870 11021 1904
rect 11021 1870 11059 1904
rect 11059 1870 11093 1904
rect 11093 1870 11131 1904
rect 11131 1870 11165 1904
rect 11165 1870 11166 1904
rect 10986 1830 11166 1870
rect 10986 1796 10987 1830
rect 10987 1796 11021 1830
rect 11021 1796 11059 1830
rect 11059 1796 11093 1830
rect 11093 1796 11131 1830
rect 11131 1796 11165 1830
rect 11165 1796 11166 1830
rect 10986 1756 11166 1796
rect 10986 1722 10987 1756
rect 10987 1722 11021 1756
rect 11021 1722 11059 1756
rect 11059 1722 11093 1756
rect 11093 1722 11131 1756
rect 11131 1722 11165 1756
rect 11165 1722 11166 1756
rect 10986 1682 11166 1722
rect 10986 1648 10987 1682
rect 10987 1648 11021 1682
rect 11021 1648 11059 1682
rect 11059 1648 11093 1682
rect 11093 1648 11131 1682
rect 11131 1648 11165 1682
rect 11165 1648 11166 1682
rect 10986 1608 11166 1648
rect 10986 1574 10987 1608
rect 10987 1574 11021 1608
rect 11021 1574 11059 1608
rect 11059 1574 11093 1608
rect 11093 1574 11131 1608
rect 11131 1574 11165 1608
rect 11165 1574 11166 1608
rect 10986 1568 11166 1574
rect 11482 4092 11534 4124
rect 11482 4072 11483 4092
rect 11483 4072 11517 4092
rect 11517 4072 11534 4092
rect 11546 4072 11598 4124
rect 11610 4092 11662 4124
rect 11610 4072 11627 4092
rect 11627 4072 11661 4092
rect 11661 4072 11662 4092
rect 11482 4058 11483 4059
rect 11483 4058 11517 4059
rect 11517 4058 11534 4059
rect 11482 4020 11534 4058
rect 11482 4007 11483 4020
rect 11483 4007 11517 4020
rect 11517 4007 11534 4020
rect 11546 4007 11598 4059
rect 11610 4058 11627 4059
rect 11627 4058 11661 4059
rect 11661 4058 11662 4059
rect 11610 4020 11662 4058
rect 11610 4007 11627 4020
rect 11627 4007 11661 4020
rect 11661 4007 11662 4020
rect 11482 3986 11483 3994
rect 11483 3986 11517 3994
rect 11517 3986 11534 3994
rect 11482 3948 11534 3986
rect 11482 3942 11483 3948
rect 11483 3942 11517 3948
rect 11517 3942 11534 3948
rect 11546 3942 11598 3994
rect 11610 3986 11627 3994
rect 11627 3986 11661 3994
rect 11661 3986 11662 3994
rect 11610 3948 11662 3986
rect 11610 3942 11627 3948
rect 11627 3942 11661 3948
rect 11661 3942 11662 3948
rect 11482 3914 11483 3929
rect 11483 3914 11517 3929
rect 11517 3914 11534 3929
rect 11482 3877 11534 3914
rect 11546 3877 11598 3929
rect 11610 3914 11627 3929
rect 11627 3914 11661 3929
rect 11661 3914 11662 3929
rect 11610 3877 11662 3914
rect 11482 3842 11483 3864
rect 11483 3842 11517 3864
rect 11517 3842 11534 3864
rect 11482 3812 11534 3842
rect 11546 3812 11598 3864
rect 11610 3842 11627 3864
rect 11627 3842 11661 3864
rect 11661 3842 11662 3864
rect 11610 3812 11662 3842
rect 11482 3770 11483 3799
rect 11483 3770 11517 3799
rect 11517 3770 11534 3799
rect 11482 3747 11534 3770
rect 11546 3747 11598 3799
rect 11610 3770 11627 3799
rect 11627 3770 11661 3799
rect 11661 3770 11662 3799
rect 11610 3747 11662 3770
rect 11482 3732 11534 3734
rect 11482 3698 11483 3732
rect 11483 3698 11517 3732
rect 11517 3698 11534 3732
rect 11482 3682 11534 3698
rect 11546 3682 11598 3734
rect 11610 3732 11662 3734
rect 11610 3698 11627 3732
rect 11627 3698 11661 3732
rect 11661 3698 11662 3732
rect 11610 3682 11662 3698
rect 11482 3660 11534 3669
rect 11482 3626 11483 3660
rect 11483 3626 11517 3660
rect 11517 3626 11534 3660
rect 11482 3617 11534 3626
rect 11546 3617 11598 3669
rect 11610 3660 11662 3669
rect 11610 3626 11627 3660
rect 11627 3626 11661 3660
rect 11661 3626 11662 3660
rect 11610 3617 11662 3626
rect 11482 3588 11662 3604
rect 11482 3554 11483 3588
rect 11483 3554 11517 3588
rect 11517 3554 11627 3588
rect 11627 3554 11661 3588
rect 11661 3554 11662 3588
rect 11482 3516 11662 3554
rect 11482 3482 11483 3516
rect 11483 3482 11517 3516
rect 11517 3482 11627 3516
rect 11627 3482 11661 3516
rect 11661 3482 11662 3516
rect 11482 3444 11662 3482
rect 11482 3410 11483 3444
rect 11483 3410 11517 3444
rect 11517 3410 11627 3444
rect 11627 3410 11661 3444
rect 11661 3410 11662 3444
rect 11482 3372 11662 3410
rect 11482 3338 11483 3372
rect 11483 3338 11517 3372
rect 11517 3338 11627 3372
rect 11627 3338 11661 3372
rect 11661 3338 11662 3372
rect 11482 3300 11662 3338
rect 11482 3266 11483 3300
rect 11483 3266 11517 3300
rect 11517 3266 11627 3300
rect 11627 3266 11661 3300
rect 11661 3266 11662 3300
rect 11482 3228 11662 3266
rect 11482 3194 11483 3228
rect 11483 3194 11517 3228
rect 11517 3194 11627 3228
rect 11627 3194 11661 3228
rect 11661 3194 11662 3228
rect 11482 3108 11662 3194
rect 11482 3074 11483 3108
rect 11483 3074 11517 3108
rect 11517 3074 11555 3108
rect 11555 3074 11589 3108
rect 11589 3074 11627 3108
rect 11627 3074 11661 3108
rect 11661 3074 11662 3108
rect 11482 3028 11662 3074
rect 11482 2994 11483 3028
rect 11483 2994 11517 3028
rect 11517 2994 11555 3028
rect 11555 2994 11589 3028
rect 11589 2994 11627 3028
rect 11627 2994 11661 3028
rect 11661 2994 11662 3028
rect 11482 2948 11662 2994
rect 11482 2914 11483 2948
rect 11483 2914 11517 2948
rect 11517 2914 11555 2948
rect 11555 2914 11589 2948
rect 11589 2914 11627 2948
rect 11627 2914 11661 2948
rect 11661 2914 11662 2948
rect 11482 2868 11662 2914
rect 11482 2834 11483 2868
rect 11483 2834 11517 2868
rect 11517 2834 11555 2868
rect 11555 2834 11589 2868
rect 11589 2834 11627 2868
rect 11627 2834 11661 2868
rect 11661 2834 11662 2868
rect 11482 2788 11662 2834
rect 11482 2754 11483 2788
rect 11483 2754 11517 2788
rect 11517 2754 11555 2788
rect 11555 2754 11589 2788
rect 11589 2754 11627 2788
rect 11627 2754 11661 2788
rect 11661 2754 11662 2788
rect 11482 2708 11662 2754
rect 11482 2674 11483 2708
rect 11483 2674 11517 2708
rect 11517 2674 11555 2708
rect 11555 2674 11589 2708
rect 11589 2674 11627 2708
rect 11627 2674 11661 2708
rect 11661 2674 11662 2708
rect 11482 2628 11662 2674
rect 11482 2594 11483 2628
rect 11483 2594 11517 2628
rect 11517 2594 11555 2628
rect 11555 2594 11589 2628
rect 11589 2594 11627 2628
rect 11627 2594 11661 2628
rect 11661 2594 11662 2628
rect 11482 2518 11662 2594
rect 11482 2484 11483 2518
rect 11483 2484 11517 2518
rect 11517 2484 11627 2518
rect 11627 2484 11661 2518
rect 11661 2484 11662 2518
rect 11482 2446 11662 2484
rect 11482 2412 11483 2446
rect 11483 2412 11517 2446
rect 11517 2412 11627 2446
rect 11627 2412 11661 2446
rect 11661 2412 11662 2446
rect 11482 2374 11662 2412
rect 11482 2340 11483 2374
rect 11483 2340 11517 2374
rect 11517 2340 11627 2374
rect 11627 2340 11661 2374
rect 11661 2340 11662 2374
rect 11482 2302 11662 2340
rect 11482 2268 11483 2302
rect 11483 2268 11517 2302
rect 11517 2268 11627 2302
rect 11627 2268 11661 2302
rect 11661 2268 11662 2302
rect 11482 2230 11662 2268
rect 11482 2196 11483 2230
rect 11483 2196 11517 2230
rect 11517 2196 11627 2230
rect 11627 2196 11661 2230
rect 11661 2196 11662 2230
rect 11482 2158 11662 2196
rect 11482 2124 11483 2158
rect 11483 2124 11517 2158
rect 11517 2124 11627 2158
rect 11627 2124 11661 2158
rect 11661 2124 11662 2158
rect 11482 2086 11662 2124
rect 11482 2052 11483 2086
rect 11483 2052 11517 2086
rect 11517 2052 11627 2086
rect 11627 2052 11661 2086
rect 11661 2052 11662 2086
rect 11482 2014 11662 2052
rect 11482 1980 11483 2014
rect 11483 1980 11517 2014
rect 11517 1980 11627 2014
rect 11627 1980 11661 2014
rect 11661 1980 11662 2014
rect 11482 1942 11662 1980
rect 11482 1908 11483 1942
rect 11483 1908 11517 1942
rect 11517 1908 11627 1942
rect 11627 1908 11661 1942
rect 11661 1908 11662 1942
rect 11482 1870 11662 1908
rect 11482 1836 11483 1870
rect 11483 1836 11517 1870
rect 11517 1836 11627 1870
rect 11627 1836 11661 1870
rect 11661 1836 11662 1870
rect 11482 1798 11662 1836
rect 11482 1764 11483 1798
rect 11483 1764 11517 1798
rect 11517 1764 11627 1798
rect 11627 1764 11661 1798
rect 11661 1764 11662 1798
rect 11482 1726 11662 1764
rect 11482 1692 11483 1726
rect 11483 1692 11517 1726
rect 11517 1692 11627 1726
rect 11627 1692 11661 1726
rect 11661 1692 11662 1726
rect 11482 1654 11662 1692
rect 11482 1620 11483 1654
rect 11483 1620 11517 1654
rect 11517 1620 11627 1654
rect 11627 1620 11661 1654
rect 11661 1620 11662 1654
rect 11482 1568 11662 1620
rect 11978 4098 12030 4119
rect 11978 4067 11979 4098
rect 11979 4067 12013 4098
rect 12013 4067 12030 4098
rect 12042 4098 12094 4119
rect 12042 4067 12051 4098
rect 12051 4067 12085 4098
rect 12085 4067 12094 4098
rect 12106 4098 12158 4119
rect 12106 4067 12123 4098
rect 12123 4067 12157 4098
rect 12157 4067 12158 4098
rect 11978 4025 12030 4054
rect 11978 4002 11979 4025
rect 11979 4002 12013 4025
rect 12013 4002 12030 4025
rect 12042 4025 12094 4054
rect 12042 4002 12051 4025
rect 12051 4002 12085 4025
rect 12085 4002 12094 4025
rect 12106 4025 12158 4054
rect 12106 4002 12123 4025
rect 12123 4002 12157 4025
rect 12157 4002 12158 4025
rect 11978 3952 12030 3989
rect 11978 3937 11979 3952
rect 11979 3937 12013 3952
rect 12013 3937 12030 3952
rect 12042 3952 12094 3989
rect 12042 3937 12051 3952
rect 12051 3937 12085 3952
rect 12085 3937 12094 3952
rect 12106 3952 12158 3989
rect 12106 3937 12123 3952
rect 12123 3937 12157 3952
rect 12157 3937 12158 3952
rect 11978 3918 11979 3924
rect 11979 3918 12013 3924
rect 12013 3918 12051 3924
rect 12051 3918 12085 3924
rect 12085 3918 12123 3924
rect 12123 3918 12157 3924
rect 12157 3918 12158 3924
rect 11978 3879 12158 3918
rect 11978 3845 11979 3879
rect 11979 3845 12013 3879
rect 12013 3845 12051 3879
rect 12051 3845 12085 3879
rect 12085 3845 12123 3879
rect 12123 3845 12157 3879
rect 12157 3845 12158 3879
rect 11978 3806 12158 3845
rect 11978 3772 11979 3806
rect 11979 3772 12013 3806
rect 12013 3772 12051 3806
rect 12051 3772 12085 3806
rect 12085 3772 12123 3806
rect 12123 3772 12157 3806
rect 12157 3772 12158 3806
rect 11978 3733 12158 3772
rect 11978 3699 11979 3733
rect 11979 3699 12013 3733
rect 12013 3699 12051 3733
rect 12051 3699 12085 3733
rect 12085 3699 12123 3733
rect 12123 3699 12157 3733
rect 12157 3699 12158 3733
rect 11978 3660 12158 3699
rect 11978 3626 11979 3660
rect 11979 3626 12013 3660
rect 12013 3626 12051 3660
rect 12051 3626 12085 3660
rect 12085 3626 12123 3660
rect 12123 3626 12157 3660
rect 12157 3626 12158 3660
rect 11978 3587 12158 3626
rect 11978 3553 11979 3587
rect 11979 3553 12013 3587
rect 12013 3553 12051 3587
rect 12051 3553 12085 3587
rect 12085 3553 12123 3587
rect 12123 3553 12157 3587
rect 12157 3553 12158 3587
rect 11978 3514 12158 3553
rect 11978 3480 11979 3514
rect 11979 3480 12013 3514
rect 12013 3480 12051 3514
rect 12051 3480 12085 3514
rect 12085 3480 12123 3514
rect 12123 3480 12157 3514
rect 12157 3480 12158 3514
rect 11978 3441 12158 3480
rect 11978 3407 11979 3441
rect 11979 3407 12013 3441
rect 12013 3407 12051 3441
rect 12051 3407 12085 3441
rect 12085 3407 12123 3441
rect 12123 3407 12157 3441
rect 12157 3407 12158 3441
rect 11978 3368 12158 3407
rect 11978 3334 11979 3368
rect 11979 3334 12013 3368
rect 12013 3334 12051 3368
rect 12051 3334 12085 3368
rect 12085 3334 12123 3368
rect 12123 3334 12157 3368
rect 12157 3334 12158 3368
rect 11978 3295 12158 3334
rect 11978 3261 11979 3295
rect 11979 3261 12013 3295
rect 12013 3261 12051 3295
rect 12051 3261 12085 3295
rect 12085 3261 12123 3295
rect 12123 3261 12157 3295
rect 12157 3261 12158 3295
rect 11978 3222 12158 3261
rect 11978 3188 11979 3222
rect 11979 3188 12013 3222
rect 12013 3188 12051 3222
rect 12051 3188 12085 3222
rect 12085 3188 12123 3222
rect 12123 3188 12157 3222
rect 12157 3188 12158 3222
rect 11978 3149 12158 3188
rect 11978 3115 11979 3149
rect 11979 3115 12013 3149
rect 12013 3115 12051 3149
rect 12051 3115 12085 3149
rect 12085 3115 12123 3149
rect 12123 3115 12157 3149
rect 12157 3115 12158 3149
rect 11978 3076 12158 3115
rect 11978 3042 11979 3076
rect 11979 3042 12013 3076
rect 12013 3042 12051 3076
rect 12051 3042 12085 3076
rect 12085 3042 12123 3076
rect 12123 3042 12157 3076
rect 12157 3042 12158 3076
rect 11978 3003 12158 3042
rect 11978 2969 11979 3003
rect 11979 2969 12013 3003
rect 12013 2969 12051 3003
rect 12051 2969 12085 3003
rect 12085 2969 12123 3003
rect 12123 2969 12157 3003
rect 12157 2969 12158 3003
rect 11978 2930 12158 2969
rect 11978 2896 11979 2930
rect 11979 2896 12013 2930
rect 12013 2896 12051 2930
rect 12051 2896 12085 2930
rect 12085 2896 12123 2930
rect 12123 2896 12157 2930
rect 12157 2896 12158 2930
rect 11978 2857 12158 2896
rect 11978 2823 11979 2857
rect 11979 2823 12013 2857
rect 12013 2823 12051 2857
rect 12051 2823 12085 2857
rect 12085 2823 12123 2857
rect 12123 2823 12157 2857
rect 12157 2823 12158 2857
rect 11978 2784 12158 2823
rect 11978 2750 11979 2784
rect 11979 2750 12013 2784
rect 12013 2750 12051 2784
rect 12051 2750 12085 2784
rect 12085 2750 12123 2784
rect 12123 2750 12157 2784
rect 12157 2750 12158 2784
rect 11978 2711 12158 2750
rect 11978 2677 11979 2711
rect 11979 2677 12013 2711
rect 12013 2677 12051 2711
rect 12051 2677 12085 2711
rect 12085 2677 12123 2711
rect 12123 2677 12157 2711
rect 12157 2677 12158 2711
rect 11978 2638 12158 2677
rect 11978 2604 11979 2638
rect 11979 2604 12013 2638
rect 12013 2604 12051 2638
rect 12051 2604 12085 2638
rect 12085 2604 12123 2638
rect 12123 2604 12157 2638
rect 12157 2604 12158 2638
rect 11978 2565 12158 2604
rect 11978 2531 11979 2565
rect 11979 2531 12013 2565
rect 12013 2531 12051 2565
rect 12051 2531 12085 2565
rect 12085 2531 12123 2565
rect 12123 2531 12157 2565
rect 12157 2531 12158 2565
rect 11978 2492 12158 2531
rect 11978 2458 11979 2492
rect 11979 2458 12013 2492
rect 12013 2458 12051 2492
rect 12051 2458 12085 2492
rect 12085 2458 12123 2492
rect 12123 2458 12157 2492
rect 12157 2458 12158 2492
rect 11978 2419 12158 2458
rect 11978 2385 11979 2419
rect 11979 2385 12013 2419
rect 12013 2385 12051 2419
rect 12051 2385 12085 2419
rect 12085 2385 12123 2419
rect 12123 2385 12157 2419
rect 12157 2385 12158 2419
rect 11978 2346 12158 2385
rect 11978 2312 11979 2346
rect 11979 2312 12013 2346
rect 12013 2312 12051 2346
rect 12051 2312 12085 2346
rect 12085 2312 12123 2346
rect 12123 2312 12157 2346
rect 12157 2312 12158 2346
rect 11978 2273 12158 2312
rect 11978 2239 11979 2273
rect 11979 2239 12013 2273
rect 12013 2239 12051 2273
rect 12051 2239 12085 2273
rect 12085 2239 12123 2273
rect 12123 2239 12157 2273
rect 12157 2239 12158 2273
rect 11978 2200 12158 2239
rect 11978 2166 11979 2200
rect 11979 2166 12013 2200
rect 12013 2166 12051 2200
rect 12051 2166 12085 2200
rect 12085 2166 12123 2200
rect 12123 2166 12157 2200
rect 12157 2166 12158 2200
rect 11978 2126 12158 2166
rect 11978 2092 11979 2126
rect 11979 2092 12013 2126
rect 12013 2092 12051 2126
rect 12051 2092 12085 2126
rect 12085 2092 12123 2126
rect 12123 2092 12157 2126
rect 12157 2092 12158 2126
rect 11978 2052 12158 2092
rect 11978 2018 11979 2052
rect 11979 2018 12013 2052
rect 12013 2018 12051 2052
rect 12051 2018 12085 2052
rect 12085 2018 12123 2052
rect 12123 2018 12157 2052
rect 12157 2018 12158 2052
rect 11978 1978 12158 2018
rect 11978 1944 11979 1978
rect 11979 1944 12013 1978
rect 12013 1944 12051 1978
rect 12051 1944 12085 1978
rect 12085 1944 12123 1978
rect 12123 1944 12157 1978
rect 12157 1944 12158 1978
rect 11978 1904 12158 1944
rect 11978 1870 11979 1904
rect 11979 1870 12013 1904
rect 12013 1870 12051 1904
rect 12051 1870 12085 1904
rect 12085 1870 12123 1904
rect 12123 1870 12157 1904
rect 12157 1870 12158 1904
rect 11978 1830 12158 1870
rect 11978 1796 11979 1830
rect 11979 1796 12013 1830
rect 12013 1796 12051 1830
rect 12051 1796 12085 1830
rect 12085 1796 12123 1830
rect 12123 1796 12157 1830
rect 12157 1796 12158 1830
rect 11978 1756 12158 1796
rect 11978 1722 11979 1756
rect 11979 1722 12013 1756
rect 12013 1722 12051 1756
rect 12051 1722 12085 1756
rect 12085 1722 12123 1756
rect 12123 1722 12157 1756
rect 12157 1722 12158 1756
rect 11978 1682 12158 1722
rect 11978 1648 11979 1682
rect 11979 1648 12013 1682
rect 12013 1648 12051 1682
rect 12051 1648 12085 1682
rect 12085 1648 12123 1682
rect 12123 1648 12157 1682
rect 12157 1648 12158 1682
rect 11978 1608 12158 1648
rect 11978 1574 11979 1608
rect 11979 1574 12013 1608
rect 12013 1574 12051 1608
rect 12051 1574 12085 1608
rect 12085 1574 12123 1608
rect 12123 1574 12157 1608
rect 12157 1574 12158 1608
rect 11978 1568 12158 1574
rect 12474 4092 12526 4124
rect 12474 4072 12475 4092
rect 12475 4072 12509 4092
rect 12509 4072 12526 4092
rect 12538 4072 12590 4124
rect 12602 4092 12654 4124
rect 12602 4072 12619 4092
rect 12619 4072 12653 4092
rect 12653 4072 12654 4092
rect 12474 4058 12475 4059
rect 12475 4058 12509 4059
rect 12509 4058 12526 4059
rect 12474 4020 12526 4058
rect 12474 4007 12475 4020
rect 12475 4007 12509 4020
rect 12509 4007 12526 4020
rect 12538 4007 12590 4059
rect 12602 4058 12619 4059
rect 12619 4058 12653 4059
rect 12653 4058 12654 4059
rect 12602 4020 12654 4058
rect 12602 4007 12619 4020
rect 12619 4007 12653 4020
rect 12653 4007 12654 4020
rect 12474 3986 12475 3994
rect 12475 3986 12509 3994
rect 12509 3986 12526 3994
rect 12474 3948 12526 3986
rect 12474 3942 12475 3948
rect 12475 3942 12509 3948
rect 12509 3942 12526 3948
rect 12538 3942 12590 3994
rect 12602 3986 12619 3994
rect 12619 3986 12653 3994
rect 12653 3986 12654 3994
rect 12602 3948 12654 3986
rect 12602 3942 12619 3948
rect 12619 3942 12653 3948
rect 12653 3942 12654 3948
rect 12474 3914 12475 3929
rect 12475 3914 12509 3929
rect 12509 3914 12526 3929
rect 12474 3877 12526 3914
rect 12538 3877 12590 3929
rect 12602 3914 12619 3929
rect 12619 3914 12653 3929
rect 12653 3914 12654 3929
rect 12602 3877 12654 3914
rect 12474 3842 12475 3864
rect 12475 3842 12509 3864
rect 12509 3842 12526 3864
rect 12474 3812 12526 3842
rect 12538 3812 12590 3864
rect 12602 3842 12619 3864
rect 12619 3842 12653 3864
rect 12653 3842 12654 3864
rect 12602 3812 12654 3842
rect 12474 3770 12475 3799
rect 12475 3770 12509 3799
rect 12509 3770 12526 3799
rect 12474 3747 12526 3770
rect 12538 3747 12590 3799
rect 12602 3770 12619 3799
rect 12619 3770 12653 3799
rect 12653 3770 12654 3799
rect 12602 3747 12654 3770
rect 12474 3732 12526 3734
rect 12474 3698 12475 3732
rect 12475 3698 12509 3732
rect 12509 3698 12526 3732
rect 12474 3682 12526 3698
rect 12538 3682 12590 3734
rect 12602 3732 12654 3734
rect 12602 3698 12619 3732
rect 12619 3698 12653 3732
rect 12653 3698 12654 3732
rect 12602 3682 12654 3698
rect 12474 3660 12526 3669
rect 12474 3626 12475 3660
rect 12475 3626 12509 3660
rect 12509 3626 12526 3660
rect 12474 3617 12526 3626
rect 12538 3617 12590 3669
rect 12602 3660 12654 3669
rect 12602 3626 12619 3660
rect 12619 3626 12653 3660
rect 12653 3626 12654 3660
rect 12602 3617 12654 3626
rect 12474 3588 12654 3604
rect 12474 3554 12475 3588
rect 12475 3554 12509 3588
rect 12509 3554 12619 3588
rect 12619 3554 12653 3588
rect 12653 3554 12654 3588
rect 12474 3516 12654 3554
rect 12474 3482 12475 3516
rect 12475 3482 12509 3516
rect 12509 3482 12619 3516
rect 12619 3482 12653 3516
rect 12653 3482 12654 3516
rect 12474 3444 12654 3482
rect 12474 3410 12475 3444
rect 12475 3410 12509 3444
rect 12509 3410 12619 3444
rect 12619 3410 12653 3444
rect 12653 3410 12654 3444
rect 12474 3372 12654 3410
rect 12474 3338 12475 3372
rect 12475 3338 12509 3372
rect 12509 3338 12619 3372
rect 12619 3338 12653 3372
rect 12653 3338 12654 3372
rect 12474 3300 12654 3338
rect 12474 3266 12475 3300
rect 12475 3266 12509 3300
rect 12509 3266 12619 3300
rect 12619 3266 12653 3300
rect 12653 3266 12654 3300
rect 12474 3228 12654 3266
rect 12474 3194 12475 3228
rect 12475 3194 12509 3228
rect 12509 3194 12619 3228
rect 12619 3194 12653 3228
rect 12653 3194 12654 3228
rect 12474 3108 12654 3194
rect 12474 3074 12475 3108
rect 12475 3074 12509 3108
rect 12509 3074 12547 3108
rect 12547 3074 12581 3108
rect 12581 3074 12619 3108
rect 12619 3074 12653 3108
rect 12653 3074 12654 3108
rect 12474 3028 12654 3074
rect 12474 2994 12475 3028
rect 12475 2994 12509 3028
rect 12509 2994 12547 3028
rect 12547 2994 12581 3028
rect 12581 2994 12619 3028
rect 12619 2994 12653 3028
rect 12653 2994 12654 3028
rect 12474 2948 12654 2994
rect 12474 2914 12475 2948
rect 12475 2914 12509 2948
rect 12509 2914 12547 2948
rect 12547 2914 12581 2948
rect 12581 2914 12619 2948
rect 12619 2914 12653 2948
rect 12653 2914 12654 2948
rect 12474 2868 12654 2914
rect 12474 2834 12475 2868
rect 12475 2834 12509 2868
rect 12509 2834 12547 2868
rect 12547 2834 12581 2868
rect 12581 2834 12619 2868
rect 12619 2834 12653 2868
rect 12653 2834 12654 2868
rect 12474 2788 12654 2834
rect 12474 2754 12475 2788
rect 12475 2754 12509 2788
rect 12509 2754 12547 2788
rect 12547 2754 12581 2788
rect 12581 2754 12619 2788
rect 12619 2754 12653 2788
rect 12653 2754 12654 2788
rect 12474 2708 12654 2754
rect 12474 2674 12475 2708
rect 12475 2674 12509 2708
rect 12509 2674 12547 2708
rect 12547 2674 12581 2708
rect 12581 2674 12619 2708
rect 12619 2674 12653 2708
rect 12653 2674 12654 2708
rect 12474 2628 12654 2674
rect 12474 2594 12475 2628
rect 12475 2594 12509 2628
rect 12509 2594 12547 2628
rect 12547 2594 12581 2628
rect 12581 2594 12619 2628
rect 12619 2594 12653 2628
rect 12653 2594 12654 2628
rect 12474 2518 12654 2594
rect 12474 2484 12475 2518
rect 12475 2484 12509 2518
rect 12509 2484 12619 2518
rect 12619 2484 12653 2518
rect 12653 2484 12654 2518
rect 12474 2446 12654 2484
rect 12474 2412 12475 2446
rect 12475 2412 12509 2446
rect 12509 2412 12619 2446
rect 12619 2412 12653 2446
rect 12653 2412 12654 2446
rect 12474 2374 12654 2412
rect 12474 2340 12475 2374
rect 12475 2340 12509 2374
rect 12509 2340 12619 2374
rect 12619 2340 12653 2374
rect 12653 2340 12654 2374
rect 12474 2302 12654 2340
rect 12474 2268 12475 2302
rect 12475 2268 12509 2302
rect 12509 2268 12619 2302
rect 12619 2268 12653 2302
rect 12653 2268 12654 2302
rect 12474 2230 12654 2268
rect 12474 2196 12475 2230
rect 12475 2196 12509 2230
rect 12509 2196 12619 2230
rect 12619 2196 12653 2230
rect 12653 2196 12654 2230
rect 12474 2158 12654 2196
rect 12474 2124 12475 2158
rect 12475 2124 12509 2158
rect 12509 2124 12619 2158
rect 12619 2124 12653 2158
rect 12653 2124 12654 2158
rect 12474 2086 12654 2124
rect 12474 2052 12475 2086
rect 12475 2052 12509 2086
rect 12509 2052 12619 2086
rect 12619 2052 12653 2086
rect 12653 2052 12654 2086
rect 12474 2014 12654 2052
rect 12474 1980 12475 2014
rect 12475 1980 12509 2014
rect 12509 1980 12619 2014
rect 12619 1980 12653 2014
rect 12653 1980 12654 2014
rect 12474 1942 12654 1980
rect 12474 1908 12475 1942
rect 12475 1908 12509 1942
rect 12509 1908 12619 1942
rect 12619 1908 12653 1942
rect 12653 1908 12654 1942
rect 12474 1870 12654 1908
rect 12474 1836 12475 1870
rect 12475 1836 12509 1870
rect 12509 1836 12619 1870
rect 12619 1836 12653 1870
rect 12653 1836 12654 1870
rect 12474 1798 12654 1836
rect 12474 1764 12475 1798
rect 12475 1764 12509 1798
rect 12509 1764 12619 1798
rect 12619 1764 12653 1798
rect 12653 1764 12654 1798
rect 12474 1726 12654 1764
rect 12474 1692 12475 1726
rect 12475 1692 12509 1726
rect 12509 1692 12619 1726
rect 12619 1692 12653 1726
rect 12653 1692 12654 1726
rect 12474 1654 12654 1692
rect 12474 1620 12475 1654
rect 12475 1620 12509 1654
rect 12509 1620 12619 1654
rect 12619 1620 12653 1654
rect 12653 1620 12654 1654
rect 12474 1568 12654 1620
rect 12970 4098 13022 4119
rect 12970 4067 12971 4098
rect 12971 4067 13005 4098
rect 13005 4067 13022 4098
rect 13034 4098 13086 4119
rect 13034 4067 13043 4098
rect 13043 4067 13077 4098
rect 13077 4067 13086 4098
rect 13098 4098 13150 4119
rect 13098 4067 13115 4098
rect 13115 4067 13149 4098
rect 13149 4067 13150 4098
rect 12970 4025 13022 4054
rect 12970 4002 12971 4025
rect 12971 4002 13005 4025
rect 13005 4002 13022 4025
rect 13034 4025 13086 4054
rect 13034 4002 13043 4025
rect 13043 4002 13077 4025
rect 13077 4002 13086 4025
rect 13098 4025 13150 4054
rect 13098 4002 13115 4025
rect 13115 4002 13149 4025
rect 13149 4002 13150 4025
rect 12970 3952 13022 3989
rect 12970 3937 12971 3952
rect 12971 3937 13005 3952
rect 13005 3937 13022 3952
rect 13034 3952 13086 3989
rect 13034 3937 13043 3952
rect 13043 3937 13077 3952
rect 13077 3937 13086 3952
rect 13098 3952 13150 3989
rect 13098 3937 13115 3952
rect 13115 3937 13149 3952
rect 13149 3937 13150 3952
rect 12970 3918 12971 3924
rect 12971 3918 13005 3924
rect 13005 3918 13043 3924
rect 13043 3918 13077 3924
rect 13077 3918 13115 3924
rect 13115 3918 13149 3924
rect 13149 3918 13150 3924
rect 12970 3879 13150 3918
rect 12970 3845 12971 3879
rect 12971 3845 13005 3879
rect 13005 3845 13043 3879
rect 13043 3845 13077 3879
rect 13077 3845 13115 3879
rect 13115 3845 13149 3879
rect 13149 3845 13150 3879
rect 12970 3806 13150 3845
rect 12970 3772 12971 3806
rect 12971 3772 13005 3806
rect 13005 3772 13043 3806
rect 13043 3772 13077 3806
rect 13077 3772 13115 3806
rect 13115 3772 13149 3806
rect 13149 3772 13150 3806
rect 12970 3733 13150 3772
rect 12970 3699 12971 3733
rect 12971 3699 13005 3733
rect 13005 3699 13043 3733
rect 13043 3699 13077 3733
rect 13077 3699 13115 3733
rect 13115 3699 13149 3733
rect 13149 3699 13150 3733
rect 12970 3660 13150 3699
rect 12970 3626 12971 3660
rect 12971 3626 13005 3660
rect 13005 3626 13043 3660
rect 13043 3626 13077 3660
rect 13077 3626 13115 3660
rect 13115 3626 13149 3660
rect 13149 3626 13150 3660
rect 12970 3587 13150 3626
rect 12970 3553 12971 3587
rect 12971 3553 13005 3587
rect 13005 3553 13043 3587
rect 13043 3553 13077 3587
rect 13077 3553 13115 3587
rect 13115 3553 13149 3587
rect 13149 3553 13150 3587
rect 12970 3514 13150 3553
rect 12970 3480 12971 3514
rect 12971 3480 13005 3514
rect 13005 3480 13043 3514
rect 13043 3480 13077 3514
rect 13077 3480 13115 3514
rect 13115 3480 13149 3514
rect 13149 3480 13150 3514
rect 12970 3441 13150 3480
rect 12970 3407 12971 3441
rect 12971 3407 13005 3441
rect 13005 3407 13043 3441
rect 13043 3407 13077 3441
rect 13077 3407 13115 3441
rect 13115 3407 13149 3441
rect 13149 3407 13150 3441
rect 12970 3368 13150 3407
rect 12970 3334 12971 3368
rect 12971 3334 13005 3368
rect 13005 3334 13043 3368
rect 13043 3334 13077 3368
rect 13077 3334 13115 3368
rect 13115 3334 13149 3368
rect 13149 3334 13150 3368
rect 12970 3295 13150 3334
rect 12970 3261 12971 3295
rect 12971 3261 13005 3295
rect 13005 3261 13043 3295
rect 13043 3261 13077 3295
rect 13077 3261 13115 3295
rect 13115 3261 13149 3295
rect 13149 3261 13150 3295
rect 12970 3222 13150 3261
rect 12970 3188 12971 3222
rect 12971 3188 13005 3222
rect 13005 3188 13043 3222
rect 13043 3188 13077 3222
rect 13077 3188 13115 3222
rect 13115 3188 13149 3222
rect 13149 3188 13150 3222
rect 12970 3149 13150 3188
rect 12970 3115 12971 3149
rect 12971 3115 13005 3149
rect 13005 3115 13043 3149
rect 13043 3115 13077 3149
rect 13077 3115 13115 3149
rect 13115 3115 13149 3149
rect 13149 3115 13150 3149
rect 12970 3076 13150 3115
rect 12970 3042 12971 3076
rect 12971 3042 13005 3076
rect 13005 3042 13043 3076
rect 13043 3042 13077 3076
rect 13077 3042 13115 3076
rect 13115 3042 13149 3076
rect 13149 3042 13150 3076
rect 12970 3003 13150 3042
rect 12970 2969 12971 3003
rect 12971 2969 13005 3003
rect 13005 2969 13043 3003
rect 13043 2969 13077 3003
rect 13077 2969 13115 3003
rect 13115 2969 13149 3003
rect 13149 2969 13150 3003
rect 12970 2930 13150 2969
rect 12970 2896 12971 2930
rect 12971 2896 13005 2930
rect 13005 2896 13043 2930
rect 13043 2896 13077 2930
rect 13077 2896 13115 2930
rect 13115 2896 13149 2930
rect 13149 2896 13150 2930
rect 12970 2857 13150 2896
rect 12970 2823 12971 2857
rect 12971 2823 13005 2857
rect 13005 2823 13043 2857
rect 13043 2823 13077 2857
rect 13077 2823 13115 2857
rect 13115 2823 13149 2857
rect 13149 2823 13150 2857
rect 12970 2784 13150 2823
rect 12970 2750 12971 2784
rect 12971 2750 13005 2784
rect 13005 2750 13043 2784
rect 13043 2750 13077 2784
rect 13077 2750 13115 2784
rect 13115 2750 13149 2784
rect 13149 2750 13150 2784
rect 12970 2711 13150 2750
rect 12970 2677 12971 2711
rect 12971 2677 13005 2711
rect 13005 2677 13043 2711
rect 13043 2677 13077 2711
rect 13077 2677 13115 2711
rect 13115 2677 13149 2711
rect 13149 2677 13150 2711
rect 12970 2638 13150 2677
rect 12970 2604 12971 2638
rect 12971 2604 13005 2638
rect 13005 2604 13043 2638
rect 13043 2604 13077 2638
rect 13077 2604 13115 2638
rect 13115 2604 13149 2638
rect 13149 2604 13150 2638
rect 12970 2565 13150 2604
rect 12970 2531 12971 2565
rect 12971 2531 13005 2565
rect 13005 2531 13043 2565
rect 13043 2531 13077 2565
rect 13077 2531 13115 2565
rect 13115 2531 13149 2565
rect 13149 2531 13150 2565
rect 12970 2492 13150 2531
rect 12970 2458 12971 2492
rect 12971 2458 13005 2492
rect 13005 2458 13043 2492
rect 13043 2458 13077 2492
rect 13077 2458 13115 2492
rect 13115 2458 13149 2492
rect 13149 2458 13150 2492
rect 12970 2419 13150 2458
rect 12970 2385 12971 2419
rect 12971 2385 13005 2419
rect 13005 2385 13043 2419
rect 13043 2385 13077 2419
rect 13077 2385 13115 2419
rect 13115 2385 13149 2419
rect 13149 2385 13150 2419
rect 12970 2346 13150 2385
rect 12970 2312 12971 2346
rect 12971 2312 13005 2346
rect 13005 2312 13043 2346
rect 13043 2312 13077 2346
rect 13077 2312 13115 2346
rect 13115 2312 13149 2346
rect 13149 2312 13150 2346
rect 12970 2273 13150 2312
rect 12970 2239 12971 2273
rect 12971 2239 13005 2273
rect 13005 2239 13043 2273
rect 13043 2239 13077 2273
rect 13077 2239 13115 2273
rect 13115 2239 13149 2273
rect 13149 2239 13150 2273
rect 12970 2200 13150 2239
rect 12970 2166 12971 2200
rect 12971 2166 13005 2200
rect 13005 2166 13043 2200
rect 13043 2166 13077 2200
rect 13077 2166 13115 2200
rect 13115 2166 13149 2200
rect 13149 2166 13150 2200
rect 12970 2126 13150 2166
rect 12970 2092 12971 2126
rect 12971 2092 13005 2126
rect 13005 2092 13043 2126
rect 13043 2092 13077 2126
rect 13077 2092 13115 2126
rect 13115 2092 13149 2126
rect 13149 2092 13150 2126
rect 12970 2052 13150 2092
rect 12970 2018 12971 2052
rect 12971 2018 13005 2052
rect 13005 2018 13043 2052
rect 13043 2018 13077 2052
rect 13077 2018 13115 2052
rect 13115 2018 13149 2052
rect 13149 2018 13150 2052
rect 12970 1978 13150 2018
rect 12970 1944 12971 1978
rect 12971 1944 13005 1978
rect 13005 1944 13043 1978
rect 13043 1944 13077 1978
rect 13077 1944 13115 1978
rect 13115 1944 13149 1978
rect 13149 1944 13150 1978
rect 12970 1904 13150 1944
rect 12970 1870 12971 1904
rect 12971 1870 13005 1904
rect 13005 1870 13043 1904
rect 13043 1870 13077 1904
rect 13077 1870 13115 1904
rect 13115 1870 13149 1904
rect 13149 1870 13150 1904
rect 12970 1830 13150 1870
rect 12970 1796 12971 1830
rect 12971 1796 13005 1830
rect 13005 1796 13043 1830
rect 13043 1796 13077 1830
rect 13077 1796 13115 1830
rect 13115 1796 13149 1830
rect 13149 1796 13150 1830
rect 12970 1756 13150 1796
rect 12970 1722 12971 1756
rect 12971 1722 13005 1756
rect 13005 1722 13043 1756
rect 13043 1722 13077 1756
rect 13077 1722 13115 1756
rect 13115 1722 13149 1756
rect 13149 1722 13150 1756
rect 12970 1682 13150 1722
rect 12970 1648 12971 1682
rect 12971 1648 13005 1682
rect 13005 1648 13043 1682
rect 13043 1648 13077 1682
rect 13077 1648 13115 1682
rect 13115 1648 13149 1682
rect 13149 1648 13150 1682
rect 12970 1608 13150 1648
rect 12970 1574 12971 1608
rect 12971 1574 13005 1608
rect 13005 1574 13043 1608
rect 13043 1574 13077 1608
rect 13077 1574 13115 1608
rect 13115 1574 13149 1608
rect 13149 1574 13150 1608
rect 12970 1568 13150 1574
rect 13466 4092 13518 4124
rect 13466 4072 13467 4092
rect 13467 4072 13501 4092
rect 13501 4072 13518 4092
rect 13530 4072 13582 4124
rect 13594 4092 13646 4124
rect 13594 4072 13611 4092
rect 13611 4072 13645 4092
rect 13645 4072 13646 4092
rect 13466 4058 13467 4059
rect 13467 4058 13501 4059
rect 13501 4058 13518 4059
rect 13466 4020 13518 4058
rect 13466 4007 13467 4020
rect 13467 4007 13501 4020
rect 13501 4007 13518 4020
rect 13530 4007 13582 4059
rect 13594 4058 13611 4059
rect 13611 4058 13645 4059
rect 13645 4058 13646 4059
rect 13594 4020 13646 4058
rect 13594 4007 13611 4020
rect 13611 4007 13645 4020
rect 13645 4007 13646 4020
rect 13466 3986 13467 3994
rect 13467 3986 13501 3994
rect 13501 3986 13518 3994
rect 13466 3948 13518 3986
rect 13466 3942 13467 3948
rect 13467 3942 13501 3948
rect 13501 3942 13518 3948
rect 13530 3942 13582 3994
rect 13594 3986 13611 3994
rect 13611 3986 13645 3994
rect 13645 3986 13646 3994
rect 13594 3948 13646 3986
rect 13594 3942 13611 3948
rect 13611 3942 13645 3948
rect 13645 3942 13646 3948
rect 13466 3914 13467 3929
rect 13467 3914 13501 3929
rect 13501 3914 13518 3929
rect 13466 3877 13518 3914
rect 13530 3877 13582 3929
rect 13594 3914 13611 3929
rect 13611 3914 13645 3929
rect 13645 3914 13646 3929
rect 13594 3877 13646 3914
rect 13466 3842 13467 3864
rect 13467 3842 13501 3864
rect 13501 3842 13518 3864
rect 13466 3812 13518 3842
rect 13530 3812 13582 3864
rect 13594 3842 13611 3864
rect 13611 3842 13645 3864
rect 13645 3842 13646 3864
rect 13594 3812 13646 3842
rect 13466 3770 13467 3799
rect 13467 3770 13501 3799
rect 13501 3770 13518 3799
rect 13466 3747 13518 3770
rect 13530 3747 13582 3799
rect 13594 3770 13611 3799
rect 13611 3770 13645 3799
rect 13645 3770 13646 3799
rect 13594 3747 13646 3770
rect 13466 3732 13518 3734
rect 13466 3698 13467 3732
rect 13467 3698 13501 3732
rect 13501 3698 13518 3732
rect 13466 3682 13518 3698
rect 13530 3682 13582 3734
rect 13594 3732 13646 3734
rect 13594 3698 13611 3732
rect 13611 3698 13645 3732
rect 13645 3698 13646 3732
rect 13594 3682 13646 3698
rect 13466 3660 13518 3669
rect 13466 3626 13467 3660
rect 13467 3626 13501 3660
rect 13501 3626 13518 3660
rect 13466 3617 13518 3626
rect 13530 3617 13582 3669
rect 13594 3660 13646 3669
rect 13594 3626 13611 3660
rect 13611 3626 13645 3660
rect 13645 3626 13646 3660
rect 13594 3617 13646 3626
rect 13466 3588 13646 3604
rect 13466 3554 13467 3588
rect 13467 3554 13501 3588
rect 13501 3554 13611 3588
rect 13611 3554 13645 3588
rect 13645 3554 13646 3588
rect 13466 3516 13646 3554
rect 13466 3482 13467 3516
rect 13467 3482 13501 3516
rect 13501 3482 13611 3516
rect 13611 3482 13645 3516
rect 13645 3482 13646 3516
rect 13466 3444 13646 3482
rect 13466 3410 13467 3444
rect 13467 3410 13501 3444
rect 13501 3410 13611 3444
rect 13611 3410 13645 3444
rect 13645 3410 13646 3444
rect 13466 3372 13646 3410
rect 13466 3338 13467 3372
rect 13467 3338 13501 3372
rect 13501 3338 13611 3372
rect 13611 3338 13645 3372
rect 13645 3338 13646 3372
rect 13466 3300 13646 3338
rect 13466 3266 13467 3300
rect 13467 3266 13501 3300
rect 13501 3266 13611 3300
rect 13611 3266 13645 3300
rect 13645 3266 13646 3300
rect 13466 3228 13646 3266
rect 13466 3194 13467 3228
rect 13467 3194 13501 3228
rect 13501 3194 13611 3228
rect 13611 3194 13645 3228
rect 13645 3194 13646 3228
rect 13466 3108 13646 3194
rect 13466 3074 13467 3108
rect 13467 3074 13501 3108
rect 13501 3074 13539 3108
rect 13539 3074 13573 3108
rect 13573 3074 13611 3108
rect 13611 3074 13645 3108
rect 13645 3074 13646 3108
rect 13466 3028 13646 3074
rect 13466 2994 13467 3028
rect 13467 2994 13501 3028
rect 13501 2994 13539 3028
rect 13539 2994 13573 3028
rect 13573 2994 13611 3028
rect 13611 2994 13645 3028
rect 13645 2994 13646 3028
rect 13466 2948 13646 2994
rect 13466 2914 13467 2948
rect 13467 2914 13501 2948
rect 13501 2914 13539 2948
rect 13539 2914 13573 2948
rect 13573 2914 13611 2948
rect 13611 2914 13645 2948
rect 13645 2914 13646 2948
rect 13466 2868 13646 2914
rect 13466 2834 13467 2868
rect 13467 2834 13501 2868
rect 13501 2834 13539 2868
rect 13539 2834 13573 2868
rect 13573 2834 13611 2868
rect 13611 2834 13645 2868
rect 13645 2834 13646 2868
rect 13466 2788 13646 2834
rect 13466 2754 13467 2788
rect 13467 2754 13501 2788
rect 13501 2754 13539 2788
rect 13539 2754 13573 2788
rect 13573 2754 13611 2788
rect 13611 2754 13645 2788
rect 13645 2754 13646 2788
rect 13466 2708 13646 2754
rect 13466 2674 13467 2708
rect 13467 2674 13501 2708
rect 13501 2674 13539 2708
rect 13539 2674 13573 2708
rect 13573 2674 13611 2708
rect 13611 2674 13645 2708
rect 13645 2674 13646 2708
rect 13466 2628 13646 2674
rect 13466 2594 13467 2628
rect 13467 2594 13501 2628
rect 13501 2594 13539 2628
rect 13539 2594 13573 2628
rect 13573 2594 13611 2628
rect 13611 2594 13645 2628
rect 13645 2594 13646 2628
rect 13466 2518 13646 2594
rect 13466 2484 13467 2518
rect 13467 2484 13501 2518
rect 13501 2484 13611 2518
rect 13611 2484 13645 2518
rect 13645 2484 13646 2518
rect 13466 2446 13646 2484
rect 13466 2412 13467 2446
rect 13467 2412 13501 2446
rect 13501 2412 13611 2446
rect 13611 2412 13645 2446
rect 13645 2412 13646 2446
rect 13466 2374 13646 2412
rect 13466 2340 13467 2374
rect 13467 2340 13501 2374
rect 13501 2340 13611 2374
rect 13611 2340 13645 2374
rect 13645 2340 13646 2374
rect 13466 2302 13646 2340
rect 13466 2268 13467 2302
rect 13467 2268 13501 2302
rect 13501 2268 13611 2302
rect 13611 2268 13645 2302
rect 13645 2268 13646 2302
rect 13466 2230 13646 2268
rect 13466 2196 13467 2230
rect 13467 2196 13501 2230
rect 13501 2196 13611 2230
rect 13611 2196 13645 2230
rect 13645 2196 13646 2230
rect 13466 2158 13646 2196
rect 13466 2124 13467 2158
rect 13467 2124 13501 2158
rect 13501 2124 13611 2158
rect 13611 2124 13645 2158
rect 13645 2124 13646 2158
rect 13466 2086 13646 2124
rect 13466 2052 13467 2086
rect 13467 2052 13501 2086
rect 13501 2052 13611 2086
rect 13611 2052 13645 2086
rect 13645 2052 13646 2086
rect 13466 2014 13646 2052
rect 13466 1980 13467 2014
rect 13467 1980 13501 2014
rect 13501 1980 13611 2014
rect 13611 1980 13645 2014
rect 13645 1980 13646 2014
rect 13466 1942 13646 1980
rect 13466 1908 13467 1942
rect 13467 1908 13501 1942
rect 13501 1908 13611 1942
rect 13611 1908 13645 1942
rect 13645 1908 13646 1942
rect 13466 1870 13646 1908
rect 13466 1836 13467 1870
rect 13467 1836 13501 1870
rect 13501 1836 13611 1870
rect 13611 1836 13645 1870
rect 13645 1836 13646 1870
rect 13466 1798 13646 1836
rect 13466 1764 13467 1798
rect 13467 1764 13501 1798
rect 13501 1764 13611 1798
rect 13611 1764 13645 1798
rect 13645 1764 13646 1798
rect 13466 1726 13646 1764
rect 13466 1692 13467 1726
rect 13467 1692 13501 1726
rect 13501 1692 13611 1726
rect 13611 1692 13645 1726
rect 13645 1692 13646 1726
rect 13466 1654 13646 1692
rect 13466 1620 13467 1654
rect 13467 1620 13501 1654
rect 13501 1620 13611 1654
rect 13611 1620 13645 1654
rect 13645 1620 13646 1654
rect 13466 1568 13646 1620
rect 13991 4098 14043 4124
rect 13991 4072 13999 4098
rect 13999 4072 14033 4098
rect 14033 4072 14043 4098
rect 14083 4072 14135 4124
rect 13991 4025 14043 4060
rect 13991 4008 13999 4025
rect 13999 4008 14033 4025
rect 14033 4008 14043 4025
rect 14083 4008 14135 4060
rect 13991 3991 13999 3996
rect 13999 3991 14033 3996
rect 14033 3991 14043 3996
rect 13991 3952 14043 3991
rect 13991 3944 13999 3952
rect 13999 3944 14033 3952
rect 14033 3944 14043 3952
rect 14083 3944 14135 3996
rect 13991 3918 13999 3932
rect 13999 3918 14033 3932
rect 14033 3918 14043 3932
rect 13991 3880 14043 3918
rect 14083 3880 14135 3932
rect 13991 3845 13999 3868
rect 13999 3845 14033 3868
rect 14033 3845 14043 3868
rect 13991 3816 14043 3845
rect 14083 3816 14135 3868
rect 13991 3772 13999 3804
rect 13999 3772 14033 3804
rect 14033 3772 14043 3804
rect 13991 3752 14043 3772
rect 14083 3752 14135 3804
rect 13991 3733 14043 3740
rect 13991 3699 13999 3733
rect 13999 3699 14033 3733
rect 14033 3699 14043 3733
rect 13991 3688 14043 3699
rect 14083 3688 14135 3740
rect 13991 3660 14043 3676
rect 13991 3626 13999 3660
rect 13999 3626 14033 3660
rect 14033 3626 14043 3660
rect 13991 3624 14043 3626
rect 14083 3624 14135 3676
rect 13991 3587 14043 3612
rect 13991 3560 13999 3587
rect 13999 3560 14033 3587
rect 14033 3560 14043 3587
rect 14083 3560 14135 3612
rect 13991 3514 14043 3548
rect 13991 3496 13999 3514
rect 13999 3496 14033 3514
rect 14033 3496 14043 3514
rect 14083 3496 14135 3548
rect 13991 3480 13999 3484
rect 13999 3480 14033 3484
rect 14033 3480 14043 3484
rect 13991 3441 14043 3480
rect 13991 3432 13999 3441
rect 13999 3432 14033 3441
rect 14033 3432 14043 3441
rect 14083 3432 14135 3484
rect 13991 3407 13999 3420
rect 13999 3407 14033 3420
rect 14033 3407 14043 3420
rect 13991 3368 14043 3407
rect 14083 3368 14135 3420
rect 13991 3334 13999 3356
rect 13999 3334 14033 3356
rect 14033 3334 14043 3356
rect 13991 3304 14043 3334
rect 14083 3304 14135 3356
rect 13991 3261 13999 3292
rect 13999 3261 14033 3292
rect 14033 3261 14043 3292
rect 13991 3240 14043 3261
rect 14083 3240 14135 3292
rect 13991 3222 14043 3228
rect 13991 3188 13999 3222
rect 13999 3188 14033 3222
rect 14033 3188 14043 3222
rect 13991 3176 14043 3188
rect 14083 3176 14135 3228
rect 13991 3149 14043 3164
rect 13991 3115 13999 3149
rect 13999 3115 14033 3149
rect 14033 3115 14043 3149
rect 13991 3112 14043 3115
rect 14083 3112 14135 3164
rect 13991 3076 14043 3100
rect 13991 3048 13999 3076
rect 13999 3048 14033 3076
rect 14033 3048 14043 3076
rect 14083 3048 14135 3100
rect 13991 3003 14043 3036
rect 13991 2984 13999 3003
rect 13999 2984 14033 3003
rect 14033 2984 14043 3003
rect 14083 2984 14135 3036
rect 13991 2969 13999 2972
rect 13999 2969 14033 2972
rect 14033 2969 14043 2972
rect 13991 2930 14043 2969
rect 13991 2920 13999 2930
rect 13999 2920 14033 2930
rect 14033 2920 14043 2930
rect 14083 2920 14135 2972
rect 13991 2896 13999 2908
rect 13999 2896 14033 2908
rect 14033 2896 14043 2908
rect 13991 2857 14043 2896
rect 13991 2856 13999 2857
rect 13999 2856 14033 2857
rect 14033 2856 14043 2857
rect 14083 2856 14135 2908
rect 13991 2823 13999 2844
rect 13999 2823 14033 2844
rect 14033 2823 14043 2844
rect 13991 2792 14043 2823
rect 14083 2792 14135 2844
rect 13991 2750 13999 2780
rect 13999 2750 14033 2780
rect 14033 2750 14043 2780
rect 13991 2728 14043 2750
rect 14083 2728 14135 2780
rect 13991 2711 14043 2716
rect 13991 2677 13999 2711
rect 13999 2677 14033 2711
rect 14033 2677 14043 2711
rect 13991 2664 14043 2677
rect 14083 2664 14135 2716
rect 13991 2638 14043 2652
rect 13991 2604 13999 2638
rect 13999 2604 14033 2638
rect 14033 2604 14043 2638
rect 13991 2600 14043 2604
rect 14083 2600 14135 2652
rect 13991 2565 14043 2588
rect 13991 2536 13999 2565
rect 13999 2536 14033 2565
rect 14033 2536 14043 2565
rect 14083 2536 14135 2588
rect 13991 2492 14043 2524
rect 13991 2472 13999 2492
rect 13999 2472 14033 2492
rect 14033 2472 14043 2492
rect 14083 2472 14135 2524
rect 13991 2458 13999 2460
rect 13999 2458 14033 2460
rect 14033 2458 14043 2460
rect 13991 2419 14043 2458
rect 13991 2408 13999 2419
rect 13999 2408 14033 2419
rect 14033 2408 14043 2419
rect 14083 2408 14135 2460
rect 13991 2385 13999 2396
rect 13999 2385 14033 2396
rect 14033 2385 14043 2396
rect 13991 2346 14043 2385
rect 13991 2344 13999 2346
rect 13999 2344 14033 2346
rect 14033 2344 14043 2346
rect 14083 2344 14135 2396
rect 13991 2312 13999 2332
rect 13999 2312 14033 2332
rect 14033 2312 14043 2332
rect 13991 2280 14043 2312
rect 14083 2280 14135 2332
rect 13991 2239 13999 2268
rect 13999 2239 14033 2268
rect 14033 2239 14043 2268
rect 13991 2216 14043 2239
rect 14083 2216 14135 2268
rect 13991 2200 14043 2204
rect 13991 2166 13999 2200
rect 13999 2166 14033 2200
rect 14033 2166 14043 2200
rect 13991 2152 14043 2166
rect 14083 2152 14135 2204
rect 13991 2126 14043 2140
rect 13991 2092 13999 2126
rect 13999 2092 14033 2126
rect 14033 2092 14043 2126
rect 13991 2088 14043 2092
rect 14083 2088 14135 2140
rect 13991 2052 14043 2075
rect 13991 2023 13999 2052
rect 13999 2023 14033 2052
rect 14033 2023 14043 2052
rect 14083 2023 14135 2075
rect 13991 1978 14043 2010
rect 13991 1958 13999 1978
rect 13999 1958 14033 1978
rect 14033 1958 14043 1978
rect 14083 1958 14135 2010
rect 13991 1944 13999 1945
rect 13999 1944 14033 1945
rect 14033 1944 14043 1945
rect 13991 1904 14043 1944
rect 13991 1893 13999 1904
rect 13999 1893 14033 1904
rect 14033 1893 14043 1904
rect 14083 1893 14135 1945
rect 13991 1870 13999 1880
rect 13999 1870 14033 1880
rect 14033 1870 14043 1880
rect 13991 1830 14043 1870
rect 13991 1828 13999 1830
rect 13999 1828 14033 1830
rect 14033 1828 14043 1830
rect 14083 1828 14135 1880
rect 13991 1796 13999 1815
rect 13999 1796 14033 1815
rect 14033 1796 14043 1815
rect 13991 1763 14043 1796
rect 14083 1763 14135 1815
rect 13991 1722 13999 1750
rect 13999 1722 14033 1750
rect 14033 1722 14043 1750
rect 13991 1698 14043 1722
rect 14083 1698 14135 1750
rect 13991 1682 14043 1685
rect 13991 1648 13999 1682
rect 13999 1648 14033 1682
rect 14033 1648 14043 1682
rect 13991 1633 14043 1648
rect 14083 1633 14135 1685
rect 13991 1608 14043 1620
rect 13991 1574 13999 1608
rect 13999 1574 14033 1608
rect 14033 1574 14043 1608
rect 13991 1568 14043 1574
rect 14083 1568 14135 1620
rect 14350 4106 14356 4124
rect 14356 4106 14390 4124
rect 14390 4106 14402 4124
rect 14350 4072 14402 4106
rect 14422 4072 14428 4124
rect 14428 4072 14474 4124
rect 14494 4072 14546 4124
rect 14566 4072 14606 4124
rect 14606 4072 14618 4124
rect 14350 4033 14356 4059
rect 14356 4033 14390 4059
rect 14390 4033 14402 4059
rect 14350 4007 14402 4033
rect 14422 4007 14428 4059
rect 14428 4007 14474 4059
rect 14494 4007 14546 4059
rect 14566 4007 14606 4059
rect 14606 4007 14618 4059
rect 14350 3960 14356 3994
rect 14356 3960 14390 3994
rect 14390 3960 14402 3994
rect 14350 3942 14402 3960
rect 14422 3960 14428 3994
rect 14428 3960 14474 3994
rect 14494 3960 14546 3994
rect 14566 3960 14606 3994
rect 14606 3960 14618 3994
rect 14422 3952 14474 3960
rect 14422 3942 14428 3952
rect 14428 3942 14462 3952
rect 14462 3942 14474 3952
rect 14494 3942 14546 3960
rect 14566 3942 14618 3960
rect 14350 3921 14402 3929
rect 14350 3887 14356 3921
rect 14356 3887 14390 3921
rect 14390 3887 14402 3921
rect 14350 3877 14402 3887
rect 14422 3918 14428 3929
rect 14428 3918 14462 3929
rect 14462 3918 14474 3929
rect 14422 3880 14474 3918
rect 14422 3877 14428 3880
rect 14428 3877 14462 3880
rect 14462 3877 14474 3880
rect 14494 3921 14546 3929
rect 14494 3887 14500 3921
rect 14500 3887 14534 3921
rect 14534 3887 14546 3921
rect 14494 3877 14546 3887
rect 14566 3921 14618 3929
rect 14566 3887 14572 3921
rect 14572 3887 14606 3921
rect 14606 3887 14618 3921
rect 14566 3877 14618 3887
rect 14350 3848 14402 3864
rect 14350 3814 14356 3848
rect 14356 3814 14390 3848
rect 14390 3814 14402 3848
rect 14350 3812 14402 3814
rect 14422 3846 14428 3864
rect 14428 3846 14462 3864
rect 14462 3846 14474 3864
rect 14422 3812 14474 3846
rect 14494 3848 14546 3864
rect 14494 3814 14500 3848
rect 14500 3814 14534 3848
rect 14534 3814 14546 3848
rect 14494 3812 14546 3814
rect 14566 3848 14618 3864
rect 14566 3814 14572 3848
rect 14572 3814 14606 3848
rect 14606 3814 14618 3848
rect 14566 3812 14618 3814
rect 14350 3775 14402 3799
rect 14350 3747 14356 3775
rect 14356 3747 14390 3775
rect 14390 3747 14402 3775
rect 14422 3774 14428 3799
rect 14428 3774 14462 3799
rect 14462 3774 14474 3799
rect 14422 3747 14474 3774
rect 14494 3775 14546 3799
rect 14494 3747 14500 3775
rect 14500 3747 14534 3775
rect 14534 3747 14546 3775
rect 14566 3775 14618 3799
rect 14566 3747 14572 3775
rect 14572 3747 14606 3775
rect 14606 3747 14618 3775
rect 14350 3702 14402 3734
rect 14350 3682 14356 3702
rect 14356 3682 14390 3702
rect 14390 3682 14402 3702
rect 14422 3702 14428 3734
rect 14428 3702 14462 3734
rect 14462 3702 14474 3734
rect 14422 3682 14474 3702
rect 14494 3702 14546 3734
rect 14494 3682 14500 3702
rect 14500 3682 14534 3702
rect 14534 3682 14546 3702
rect 14566 3702 14618 3734
rect 14566 3682 14572 3702
rect 14572 3682 14606 3702
rect 14606 3682 14618 3702
rect 14350 3668 14356 3669
rect 14356 3668 14390 3669
rect 14390 3668 14402 3669
rect 14350 3629 14402 3668
rect 14350 3617 14356 3629
rect 14356 3617 14390 3629
rect 14390 3617 14402 3629
rect 14422 3664 14474 3669
rect 14422 3630 14428 3664
rect 14428 3630 14462 3664
rect 14462 3630 14474 3664
rect 14422 3617 14474 3630
rect 14494 3668 14500 3669
rect 14500 3668 14534 3669
rect 14534 3668 14546 3669
rect 14494 3629 14546 3668
rect 14494 3617 14500 3629
rect 14500 3617 14534 3629
rect 14534 3617 14546 3629
rect 14566 3668 14572 3669
rect 14572 3668 14606 3669
rect 14606 3668 14618 3669
rect 14566 3629 14618 3668
rect 14566 3617 14572 3629
rect 14572 3617 14606 3629
rect 14606 3617 14618 3629
rect 14350 3595 14356 3604
rect 14356 3595 14390 3604
rect 14390 3595 14402 3604
rect 14350 3556 14402 3595
rect 14350 3552 14356 3556
rect 14356 3552 14390 3556
rect 14390 3552 14402 3556
rect 14422 3592 14474 3604
rect 14422 3558 14428 3592
rect 14428 3558 14462 3592
rect 14462 3558 14474 3592
rect 14422 3552 14474 3558
rect 14494 3595 14500 3604
rect 14500 3595 14534 3604
rect 14534 3595 14546 3604
rect 14494 3556 14546 3595
rect 14494 3552 14500 3556
rect 14500 3552 14534 3556
rect 14534 3552 14546 3556
rect 14566 3595 14572 3604
rect 14572 3595 14606 3604
rect 14606 3595 14618 3604
rect 14566 3556 14618 3595
rect 14566 3552 14572 3556
rect 14572 3552 14606 3556
rect 14606 3552 14618 3556
rect 14350 3522 14356 3540
rect 14356 3522 14390 3540
rect 14390 3522 14402 3540
rect 14350 3488 14402 3522
rect 14422 3520 14474 3540
rect 14422 3488 14428 3520
rect 14428 3488 14462 3520
rect 14462 3488 14474 3520
rect 14494 3522 14500 3540
rect 14500 3522 14534 3540
rect 14534 3522 14546 3540
rect 14494 3488 14546 3522
rect 14566 3522 14572 3540
rect 14572 3522 14606 3540
rect 14606 3522 14618 3540
rect 14566 3488 14618 3522
rect 14350 3449 14356 3476
rect 14356 3449 14390 3476
rect 14390 3449 14402 3476
rect 14350 3424 14402 3449
rect 14422 3448 14474 3476
rect 14422 3424 14428 3448
rect 14428 3424 14462 3448
rect 14462 3424 14474 3448
rect 14494 3449 14500 3476
rect 14500 3449 14534 3476
rect 14534 3449 14546 3476
rect 14494 3424 14546 3449
rect 14566 3449 14572 3476
rect 14572 3449 14606 3476
rect 14606 3449 14618 3476
rect 14566 3424 14618 3449
rect 14350 3410 14402 3412
rect 14350 3376 14356 3410
rect 14356 3376 14390 3410
rect 14390 3376 14402 3410
rect 14350 3360 14402 3376
rect 14422 3376 14474 3412
rect 14422 3360 14428 3376
rect 14428 3360 14462 3376
rect 14462 3360 14474 3376
rect 14494 3410 14546 3412
rect 14494 3376 14500 3410
rect 14500 3376 14534 3410
rect 14534 3376 14546 3410
rect 14494 3360 14546 3376
rect 14566 3410 14618 3412
rect 14566 3376 14572 3410
rect 14572 3376 14606 3410
rect 14606 3376 14618 3410
rect 14566 3360 14618 3376
rect 14350 3337 14402 3348
rect 14350 3303 14356 3337
rect 14356 3303 14390 3337
rect 14390 3303 14402 3337
rect 14350 3296 14402 3303
rect 14422 3342 14428 3348
rect 14428 3342 14462 3348
rect 14462 3342 14474 3348
rect 14422 3304 14474 3342
rect 14422 3296 14428 3304
rect 14428 3296 14462 3304
rect 14462 3296 14474 3304
rect 14494 3337 14546 3348
rect 14494 3303 14500 3337
rect 14500 3303 14534 3337
rect 14534 3303 14546 3337
rect 14494 3296 14546 3303
rect 14566 3337 14618 3348
rect 14566 3303 14572 3337
rect 14572 3303 14606 3337
rect 14606 3303 14618 3337
rect 14566 3296 14618 3303
rect 14350 3264 14402 3284
rect 14350 3232 14356 3264
rect 14356 3232 14390 3264
rect 14390 3232 14402 3264
rect 14422 3270 14428 3284
rect 14428 3270 14462 3284
rect 14462 3270 14474 3284
rect 14422 3232 14474 3270
rect 14494 3264 14546 3284
rect 14494 3232 14500 3264
rect 14500 3232 14534 3264
rect 14534 3232 14546 3264
rect 14566 3264 14618 3284
rect 14566 3232 14572 3264
rect 14572 3232 14606 3264
rect 14606 3232 14618 3264
rect 14350 3191 14402 3220
rect 14350 3168 14356 3191
rect 14356 3168 14390 3191
rect 14390 3168 14402 3191
rect 14422 3198 14428 3220
rect 14428 3198 14462 3220
rect 14462 3198 14474 3220
rect 14422 3168 14474 3198
rect 14494 3191 14546 3220
rect 14494 3168 14500 3191
rect 14500 3168 14534 3191
rect 14534 3168 14546 3191
rect 14566 3191 14618 3220
rect 14566 3168 14572 3191
rect 14572 3168 14606 3191
rect 14606 3168 14618 3191
rect 14350 3118 14402 3156
rect 14350 3104 14356 3118
rect 14356 3104 14390 3118
rect 14390 3104 14402 3118
rect 14422 3126 14428 3156
rect 14428 3126 14462 3156
rect 14462 3126 14474 3156
rect 14422 3104 14474 3126
rect 14494 3118 14546 3156
rect 14494 3104 14500 3118
rect 14500 3104 14534 3118
rect 14534 3104 14546 3118
rect 14566 3118 14618 3156
rect 14566 3104 14572 3118
rect 14572 3104 14606 3118
rect 14606 3104 14618 3118
rect 14350 3084 14356 3092
rect 14356 3084 14390 3092
rect 14390 3084 14402 3092
rect 14350 3045 14402 3084
rect 14350 3040 14356 3045
rect 14356 3040 14390 3045
rect 14390 3040 14402 3045
rect 14422 3088 14474 3092
rect 14422 3054 14428 3088
rect 14428 3054 14462 3088
rect 14462 3054 14474 3088
rect 14422 3040 14474 3054
rect 14494 3084 14500 3092
rect 14500 3084 14534 3092
rect 14534 3084 14546 3092
rect 14494 3045 14546 3084
rect 14494 3040 14500 3045
rect 14500 3040 14534 3045
rect 14534 3040 14546 3045
rect 14566 3084 14572 3092
rect 14572 3084 14606 3092
rect 14606 3084 14618 3092
rect 14566 3045 14618 3084
rect 14566 3040 14572 3045
rect 14572 3040 14606 3045
rect 14606 3040 14618 3045
rect 14350 3011 14356 3028
rect 14356 3011 14390 3028
rect 14390 3011 14402 3028
rect 14350 2976 14402 3011
rect 14422 3016 14474 3028
rect 14422 2982 14428 3016
rect 14428 2982 14462 3016
rect 14462 2982 14474 3016
rect 14422 2976 14474 2982
rect 14494 3011 14500 3028
rect 14500 3011 14534 3028
rect 14534 3011 14546 3028
rect 14494 2976 14546 3011
rect 14566 3011 14572 3028
rect 14572 3011 14606 3028
rect 14606 3011 14618 3028
rect 14566 2976 14618 3011
rect 14350 2938 14356 2964
rect 14356 2938 14390 2964
rect 14390 2938 14402 2964
rect 14350 2912 14402 2938
rect 14422 2944 14474 2964
rect 14422 2912 14428 2944
rect 14428 2912 14462 2944
rect 14462 2912 14474 2944
rect 14494 2938 14500 2964
rect 14500 2938 14534 2964
rect 14534 2938 14546 2964
rect 14494 2912 14546 2938
rect 14566 2938 14572 2964
rect 14572 2938 14606 2964
rect 14606 2938 14618 2964
rect 14566 2912 14618 2938
rect 14350 2899 14402 2900
rect 14350 2865 14356 2899
rect 14356 2865 14390 2899
rect 14390 2865 14402 2899
rect 14350 2848 14402 2865
rect 14422 2872 14474 2900
rect 14422 2848 14428 2872
rect 14428 2848 14462 2872
rect 14462 2848 14474 2872
rect 14494 2899 14546 2900
rect 14494 2865 14500 2899
rect 14500 2865 14534 2899
rect 14534 2865 14546 2899
rect 14494 2848 14546 2865
rect 14566 2899 14618 2900
rect 14566 2865 14572 2899
rect 14572 2865 14606 2899
rect 14606 2865 14618 2899
rect 14566 2848 14618 2865
rect 14350 2826 14402 2836
rect 14350 2792 14356 2826
rect 14356 2792 14390 2826
rect 14390 2792 14402 2826
rect 14350 2784 14402 2792
rect 14422 2800 14474 2836
rect 14422 2784 14428 2800
rect 14428 2784 14462 2800
rect 14462 2784 14474 2800
rect 14494 2826 14546 2836
rect 14494 2792 14500 2826
rect 14500 2792 14534 2826
rect 14534 2792 14546 2826
rect 14494 2784 14546 2792
rect 14566 2826 14618 2836
rect 14566 2792 14572 2826
rect 14572 2792 14606 2826
rect 14606 2792 14618 2826
rect 14566 2784 14618 2792
rect 14350 2753 14402 2772
rect 14350 2720 14356 2753
rect 14356 2720 14390 2753
rect 14390 2720 14402 2753
rect 14422 2766 14428 2772
rect 14428 2766 14462 2772
rect 14462 2766 14474 2772
rect 14422 2728 14474 2766
rect 14422 2720 14428 2728
rect 14428 2720 14462 2728
rect 14462 2720 14474 2728
rect 14494 2753 14546 2772
rect 14494 2720 14500 2753
rect 14500 2720 14534 2753
rect 14534 2720 14546 2753
rect 14566 2753 14618 2772
rect 14566 2720 14572 2753
rect 14572 2720 14606 2753
rect 14606 2720 14618 2753
rect 14350 2680 14402 2708
rect 14350 2656 14356 2680
rect 14356 2656 14390 2680
rect 14390 2656 14402 2680
rect 14422 2694 14428 2708
rect 14428 2694 14462 2708
rect 14462 2694 14474 2708
rect 14422 2656 14474 2694
rect 14494 2680 14546 2708
rect 14494 2656 14500 2680
rect 14500 2656 14534 2680
rect 14534 2656 14546 2680
rect 14566 2680 14618 2708
rect 14566 2656 14572 2680
rect 14572 2656 14606 2680
rect 14606 2656 14618 2680
rect 14350 2607 14402 2644
rect 14350 2592 14356 2607
rect 14356 2592 14390 2607
rect 14390 2592 14402 2607
rect 14422 2622 14428 2644
rect 14428 2622 14462 2644
rect 14462 2622 14474 2644
rect 14422 2592 14474 2622
rect 14494 2607 14546 2644
rect 14494 2592 14500 2607
rect 14500 2592 14534 2607
rect 14534 2592 14546 2607
rect 14566 2607 14618 2644
rect 14566 2592 14572 2607
rect 14572 2592 14606 2607
rect 14606 2592 14618 2607
rect 14350 2573 14356 2580
rect 14356 2573 14390 2580
rect 14390 2573 14402 2580
rect 14350 2534 14402 2573
rect 14350 2528 14356 2534
rect 14356 2528 14390 2534
rect 14390 2528 14402 2534
rect 14422 2550 14428 2580
rect 14428 2550 14462 2580
rect 14462 2550 14474 2580
rect 14422 2528 14474 2550
rect 14494 2573 14500 2580
rect 14500 2573 14534 2580
rect 14534 2573 14546 2580
rect 14494 2534 14546 2573
rect 14494 2528 14500 2534
rect 14500 2528 14534 2534
rect 14534 2528 14546 2534
rect 14566 2573 14572 2580
rect 14572 2573 14606 2580
rect 14606 2573 14618 2580
rect 14566 2534 14618 2573
rect 14566 2528 14572 2534
rect 14572 2528 14606 2534
rect 14606 2528 14618 2534
rect 14350 2500 14356 2516
rect 14356 2500 14390 2516
rect 14390 2500 14402 2516
rect 14350 2464 14402 2500
rect 14422 2512 14474 2516
rect 14422 2478 14428 2512
rect 14428 2478 14462 2512
rect 14462 2478 14474 2512
rect 14422 2464 14474 2478
rect 14494 2500 14500 2516
rect 14500 2500 14534 2516
rect 14534 2500 14546 2516
rect 14494 2464 14546 2500
rect 14566 2500 14572 2516
rect 14572 2500 14606 2516
rect 14606 2500 14618 2516
rect 14566 2464 14618 2500
rect 14350 2427 14356 2452
rect 14356 2427 14390 2452
rect 14390 2427 14402 2452
rect 14350 2400 14402 2427
rect 14422 2440 14474 2452
rect 14422 2406 14428 2440
rect 14428 2406 14462 2440
rect 14462 2406 14474 2440
rect 14422 2400 14474 2406
rect 14494 2427 14500 2452
rect 14500 2427 14534 2452
rect 14534 2427 14546 2452
rect 14494 2400 14546 2427
rect 14566 2427 14572 2452
rect 14572 2427 14606 2452
rect 14606 2427 14618 2452
rect 14566 2400 14618 2427
rect 14350 2354 14356 2388
rect 14356 2354 14390 2388
rect 14390 2354 14402 2388
rect 14350 2336 14402 2354
rect 14422 2368 14474 2388
rect 14422 2336 14428 2368
rect 14428 2336 14462 2368
rect 14462 2336 14474 2368
rect 14494 2354 14500 2388
rect 14500 2354 14534 2388
rect 14534 2354 14546 2388
rect 14494 2336 14546 2354
rect 14566 2354 14572 2388
rect 14572 2354 14606 2388
rect 14606 2354 14618 2388
rect 14566 2336 14618 2354
rect 14350 2315 14402 2324
rect 14350 2281 14356 2315
rect 14356 2281 14390 2315
rect 14390 2281 14402 2315
rect 14350 2272 14402 2281
rect 14422 2296 14474 2324
rect 14422 2272 14428 2296
rect 14428 2272 14462 2296
rect 14462 2272 14474 2296
rect 14494 2315 14546 2324
rect 14494 2281 14500 2315
rect 14500 2281 14534 2315
rect 14534 2281 14546 2315
rect 14494 2272 14546 2281
rect 14566 2315 14618 2324
rect 14566 2281 14572 2315
rect 14572 2281 14606 2315
rect 14606 2281 14618 2315
rect 14566 2272 14618 2281
rect 14350 2242 14402 2260
rect 14350 2208 14356 2242
rect 14356 2208 14390 2242
rect 14390 2208 14402 2242
rect 14422 2224 14474 2260
rect 14422 2208 14428 2224
rect 14428 2208 14462 2224
rect 14462 2208 14474 2224
rect 14494 2242 14546 2260
rect 14494 2208 14500 2242
rect 14500 2208 14534 2242
rect 14534 2208 14546 2242
rect 14566 2242 14618 2260
rect 14566 2208 14572 2242
rect 14572 2208 14606 2242
rect 14606 2208 14618 2242
rect 14350 2169 14402 2196
rect 14350 2144 14356 2169
rect 14356 2144 14390 2169
rect 14390 2144 14402 2169
rect 14422 2190 14428 2196
rect 14428 2190 14462 2196
rect 14462 2190 14474 2196
rect 14422 2152 14474 2190
rect 14422 2144 14428 2152
rect 14428 2144 14462 2152
rect 14462 2144 14474 2152
rect 14494 2169 14546 2196
rect 14494 2144 14500 2169
rect 14500 2144 14534 2169
rect 14534 2144 14546 2169
rect 14566 2169 14618 2196
rect 14566 2144 14572 2169
rect 14572 2144 14606 2169
rect 14606 2144 14618 2169
rect 14350 2096 14402 2132
rect 14350 2080 14356 2096
rect 14356 2080 14390 2096
rect 14390 2080 14402 2096
rect 14422 2118 14428 2132
rect 14428 2118 14462 2132
rect 14462 2118 14474 2132
rect 14422 2080 14474 2118
rect 14494 2096 14546 2132
rect 14494 2080 14500 2096
rect 14500 2080 14534 2096
rect 14534 2080 14546 2096
rect 14566 2096 14618 2132
rect 14566 2080 14572 2096
rect 14572 2080 14606 2096
rect 14606 2080 14618 2096
rect 14350 2062 14356 2068
rect 14356 2062 14390 2068
rect 14390 2062 14402 2068
rect 14350 2023 14402 2062
rect 14350 2016 14356 2023
rect 14356 2016 14390 2023
rect 14390 2016 14402 2023
rect 14422 2046 14428 2068
rect 14428 2046 14462 2068
rect 14462 2046 14474 2068
rect 14422 2016 14474 2046
rect 14494 2062 14500 2068
rect 14500 2062 14534 2068
rect 14534 2062 14546 2068
rect 14494 2023 14546 2062
rect 14494 2016 14500 2023
rect 14500 2016 14534 2023
rect 14534 2016 14546 2023
rect 14566 2062 14572 2068
rect 14572 2062 14606 2068
rect 14606 2062 14618 2068
rect 14566 2023 14618 2062
rect 14566 2016 14572 2023
rect 14572 2016 14606 2023
rect 14606 2016 14618 2023
rect 14350 1989 14356 2004
rect 14356 1989 14390 2004
rect 14390 1989 14402 2004
rect 14350 1952 14402 1989
rect 14422 1974 14428 2004
rect 14428 1974 14462 2004
rect 14462 1974 14474 2004
rect 14422 1952 14474 1974
rect 14494 1989 14500 2004
rect 14500 1989 14534 2004
rect 14534 1989 14546 2004
rect 14494 1952 14546 1989
rect 14566 1989 14572 2004
rect 14572 1989 14606 2004
rect 14606 1989 14618 2004
rect 14566 1952 14618 1989
rect 14350 1916 14356 1940
rect 14356 1916 14390 1940
rect 14390 1916 14402 1940
rect 14350 1888 14402 1916
rect 14422 1936 14474 1940
rect 14422 1902 14428 1936
rect 14428 1902 14462 1936
rect 14462 1902 14474 1936
rect 14422 1888 14474 1902
rect 14494 1916 14500 1940
rect 14500 1916 14534 1940
rect 14534 1916 14546 1940
rect 14494 1888 14546 1916
rect 14566 1916 14572 1940
rect 14572 1916 14606 1940
rect 14606 1916 14618 1940
rect 14566 1888 14618 1916
rect 14350 1843 14356 1876
rect 14356 1843 14390 1876
rect 14390 1843 14402 1876
rect 14350 1824 14402 1843
rect 14422 1864 14474 1876
rect 14422 1830 14428 1864
rect 14428 1830 14462 1864
rect 14462 1830 14474 1864
rect 14422 1824 14474 1830
rect 14494 1843 14500 1876
rect 14500 1843 14534 1876
rect 14534 1843 14546 1876
rect 14494 1824 14546 1843
rect 14566 1843 14572 1876
rect 14572 1843 14606 1876
rect 14606 1843 14618 1876
rect 14566 1824 14618 1843
rect 14350 1804 14402 1812
rect 14350 1770 14356 1804
rect 14356 1770 14390 1804
rect 14390 1770 14402 1804
rect 14350 1760 14402 1770
rect 14422 1792 14474 1812
rect 14422 1760 14428 1792
rect 14428 1760 14462 1792
rect 14462 1760 14474 1792
rect 14494 1804 14546 1812
rect 14494 1770 14500 1804
rect 14500 1770 14534 1804
rect 14534 1770 14546 1804
rect 14494 1760 14546 1770
rect 14566 1804 14618 1812
rect 14566 1770 14572 1804
rect 14572 1770 14606 1804
rect 14606 1770 14618 1804
rect 14566 1760 14618 1770
rect 14350 1731 14402 1748
rect 14350 1697 14356 1731
rect 14356 1697 14390 1731
rect 14390 1697 14402 1731
rect 14350 1696 14402 1697
rect 14422 1720 14474 1748
rect 14422 1696 14428 1720
rect 14428 1696 14462 1720
rect 14462 1696 14474 1720
rect 14494 1731 14546 1748
rect 14494 1697 14500 1731
rect 14500 1697 14534 1731
rect 14534 1697 14546 1731
rect 14494 1696 14546 1697
rect 14566 1731 14618 1748
rect 14566 1697 14572 1731
rect 14572 1697 14606 1731
rect 14606 1697 14618 1731
rect 14566 1696 14618 1697
rect 14350 1657 14402 1684
rect 14350 1632 14356 1657
rect 14356 1632 14390 1657
rect 14390 1632 14402 1657
rect 14422 1648 14474 1684
rect 14422 1632 14428 1648
rect 14428 1632 14462 1648
rect 14462 1632 14474 1648
rect 14494 1658 14546 1684
rect 14494 1632 14500 1658
rect 14500 1632 14534 1658
rect 14534 1632 14546 1658
rect 14566 1658 14618 1684
rect 14566 1632 14572 1658
rect 14572 1632 14606 1658
rect 14606 1632 14618 1658
rect 14350 1583 14402 1620
rect 14350 1568 14356 1583
rect 14356 1568 14390 1583
rect 14390 1568 14402 1583
rect 14422 1614 14428 1620
rect 14428 1614 14462 1620
rect 14462 1614 14474 1620
rect 14422 1576 14474 1614
rect 14422 1568 14428 1576
rect 14428 1568 14462 1576
rect 14462 1568 14474 1576
rect 14494 1585 14546 1620
rect 14494 1568 14500 1585
rect 14500 1568 14534 1585
rect 14534 1568 14546 1585
rect 14566 1585 14618 1620
rect 14566 1568 14572 1585
rect 14572 1568 14606 1585
rect 14606 1568 14618 1585
rect 518 1513 570 1530
rect 518 1479 529 1513
rect 529 1479 563 1513
rect 563 1479 570 1513
rect 518 1478 570 1479
rect 590 1513 642 1530
rect 590 1479 601 1513
rect 601 1479 635 1513
rect 635 1479 642 1513
rect 590 1478 642 1479
rect 662 1478 674 1530
rect 674 1478 714 1530
rect 734 1478 780 1530
rect 780 1478 786 1530
rect 518 1440 570 1465
rect 518 1413 529 1440
rect 529 1413 563 1440
rect 563 1413 570 1440
rect 590 1440 642 1465
rect 590 1413 601 1440
rect 601 1413 635 1440
rect 635 1413 642 1440
rect 662 1413 674 1465
rect 674 1413 714 1465
rect 734 1413 780 1465
rect 780 1413 786 1465
rect 518 1367 570 1400
rect 518 1348 529 1367
rect 529 1348 563 1367
rect 563 1348 570 1367
rect 590 1367 642 1400
rect 590 1348 601 1367
rect 601 1348 635 1367
rect 635 1348 642 1367
rect 662 1348 674 1400
rect 674 1348 714 1400
rect 734 1348 780 1400
rect 780 1348 786 1400
rect 518 1333 529 1335
rect 529 1333 563 1335
rect 563 1333 570 1335
rect 518 1294 570 1333
rect 518 1283 529 1294
rect 529 1283 563 1294
rect 563 1283 570 1294
rect 590 1333 601 1335
rect 601 1333 635 1335
rect 635 1333 642 1335
rect 590 1294 642 1333
rect 590 1283 601 1294
rect 601 1283 635 1294
rect 635 1283 642 1294
rect 662 1283 674 1335
rect 674 1283 714 1335
rect 734 1283 780 1335
rect 780 1283 786 1335
rect 518 1260 529 1270
rect 529 1260 563 1270
rect 563 1260 570 1270
rect 518 1221 570 1260
rect 518 1218 529 1221
rect 529 1218 563 1221
rect 563 1218 570 1221
rect 590 1260 601 1270
rect 601 1260 635 1270
rect 635 1260 642 1270
rect 590 1221 642 1260
rect 590 1218 601 1221
rect 601 1218 635 1221
rect 635 1218 642 1221
rect 662 1218 674 1270
rect 674 1218 714 1270
rect 734 1218 780 1270
rect 780 1218 786 1270
rect 518 1187 529 1205
rect 529 1187 563 1205
rect 563 1187 570 1205
rect 518 1153 570 1187
rect 590 1187 601 1205
rect 601 1187 635 1205
rect 635 1187 642 1205
rect 590 1153 642 1187
rect 662 1153 674 1205
rect 674 1153 714 1205
rect 734 1153 780 1205
rect 780 1153 786 1205
rect 518 1114 529 1140
rect 529 1114 563 1140
rect 563 1114 570 1140
rect 518 1088 570 1114
rect 590 1114 601 1140
rect 601 1114 635 1140
rect 635 1114 642 1140
rect 590 1088 642 1114
rect 662 1088 674 1140
rect 674 1088 714 1140
rect 734 1088 780 1140
rect 780 1088 786 1140
rect 518 1041 529 1075
rect 529 1041 563 1075
rect 563 1041 570 1075
rect 518 1023 570 1041
rect 590 1041 601 1075
rect 601 1041 635 1075
rect 635 1041 642 1075
rect 590 1023 642 1041
rect 662 1023 674 1075
rect 674 1023 714 1075
rect 734 1023 780 1075
rect 780 1023 786 1075
rect 518 1002 570 1010
rect 518 968 529 1002
rect 529 968 563 1002
rect 563 968 570 1002
rect 518 958 570 968
rect 590 1002 642 1010
rect 590 968 601 1002
rect 601 968 635 1002
rect 635 968 642 1002
rect 590 958 642 968
rect 662 958 674 1010
rect 674 958 714 1010
rect 734 958 780 1010
rect 780 958 786 1010
rect 518 929 570 945
rect 518 895 529 929
rect 529 895 563 929
rect 563 895 570 929
rect 518 893 570 895
rect 590 929 642 945
rect 590 895 601 929
rect 601 895 635 929
rect 635 895 642 929
rect 590 893 642 895
rect 662 894 674 945
rect 674 894 714 945
rect 734 894 780 945
rect 662 893 714 894
rect 734 893 746 894
rect 746 893 780 894
rect 780 893 786 945
rect 518 828 570 880
rect 590 828 642 880
rect 662 828 714 880
rect 734 828 786 880
<< metal2 >>
rect 518 4456 786 4462
rect 570 4404 590 4456
rect 642 4404 662 4456
rect 714 4404 734 4456
rect 518 4390 786 4404
rect 570 4338 590 4390
rect 642 4338 662 4390
rect 714 4338 734 4390
rect 518 4325 786 4338
rect 570 4273 590 4325
rect 642 4273 662 4325
rect 714 4273 734 4325
rect 518 4260 786 4273
rect 570 4208 590 4260
rect 642 4208 662 4260
rect 714 4208 734 4260
rect 518 4195 786 4208
rect 570 4143 590 4195
rect 642 4143 662 4195
rect 714 4143 734 4195
rect 518 4130 786 4143
rect 570 4078 590 4130
rect 642 4078 662 4130
rect 714 4078 734 4130
rect 518 4065 786 4078
rect 570 4013 590 4065
rect 642 4013 662 4065
rect 714 4013 734 4065
rect 518 4000 786 4013
rect 570 3948 590 4000
rect 642 3948 662 4000
rect 714 3948 734 4000
rect 518 3935 786 3948
rect 570 3883 590 3935
rect 642 3883 662 3935
rect 714 3883 734 3935
rect 518 3870 786 3883
rect 570 3818 590 3870
rect 642 3818 662 3870
rect 714 3818 734 3870
rect 518 3805 786 3818
rect 570 3753 590 3805
rect 642 3753 662 3805
rect 714 3753 734 3805
rect 518 3740 786 3753
rect 570 3688 590 3740
rect 642 3688 662 3740
rect 714 3688 734 3740
rect 518 3675 786 3688
rect 570 3623 590 3675
rect 642 3623 662 3675
rect 714 3623 734 3675
rect 518 3610 786 3623
rect 570 3558 590 3610
rect 642 3558 662 3610
rect 714 3558 734 3610
rect 518 3545 786 3558
rect 570 3493 590 3545
rect 642 3493 662 3545
rect 714 3493 734 3545
rect 518 3480 786 3493
rect 570 3428 590 3480
rect 642 3428 662 3480
rect 714 3428 734 3480
rect 518 3415 786 3428
rect 570 3363 590 3415
rect 642 3363 662 3415
rect 714 3363 734 3415
rect 518 3350 786 3363
rect 570 3298 590 3350
rect 642 3298 662 3350
rect 714 3298 734 3350
rect 518 3285 786 3298
rect 570 3233 590 3285
rect 642 3233 662 3285
rect 714 3233 734 3285
rect 518 3220 786 3233
rect 570 3168 590 3220
rect 642 3168 662 3220
rect 714 3168 734 3220
rect 518 3155 786 3168
rect 570 3103 590 3155
rect 642 3103 662 3155
rect 714 3103 734 3155
rect 518 3090 786 3103
rect 570 3038 590 3090
rect 642 3038 662 3090
rect 714 3038 734 3090
rect 518 3025 786 3038
rect 570 2973 590 3025
rect 642 2973 662 3025
rect 714 2973 734 3025
rect 518 2960 786 2973
rect 570 2908 590 2960
rect 642 2908 662 2960
rect 714 2908 734 2960
rect 518 2895 786 2908
rect 570 2843 590 2895
rect 642 2843 662 2895
rect 714 2843 734 2895
rect 518 2830 786 2843
rect 570 2778 590 2830
rect 642 2778 662 2830
rect 714 2778 734 2830
rect 518 2765 786 2778
rect 570 2713 590 2765
rect 642 2713 662 2765
rect 714 2713 734 2765
rect 518 2700 786 2713
rect 570 2648 590 2700
rect 642 2648 662 2700
rect 714 2648 734 2700
rect 518 2635 786 2648
rect 570 2583 590 2635
rect 642 2583 662 2635
rect 714 2583 734 2635
rect 518 2570 786 2583
rect 570 2518 590 2570
rect 642 2518 662 2570
rect 714 2518 734 2570
rect 518 2505 786 2518
rect 570 2453 590 2505
rect 642 2453 662 2505
rect 714 2453 734 2505
rect 518 2440 786 2453
rect 570 2388 590 2440
rect 642 2388 662 2440
rect 714 2388 734 2440
rect 518 2375 786 2388
rect 570 2323 590 2375
rect 642 2323 662 2375
rect 714 2323 734 2375
rect 518 2310 786 2323
rect 570 2258 590 2310
rect 642 2258 662 2310
rect 714 2258 734 2310
rect 518 2245 786 2258
rect 570 2193 590 2245
rect 642 2193 662 2245
rect 714 2193 734 2245
rect 518 2180 786 2193
rect 570 2128 590 2180
rect 642 2128 662 2180
rect 714 2128 734 2180
rect 518 2115 786 2128
rect 570 2063 590 2115
rect 642 2063 662 2115
rect 714 2063 734 2115
rect 518 2050 786 2063
rect 570 1998 590 2050
rect 642 1998 662 2050
rect 714 1998 734 2050
rect 518 1985 786 1998
rect 570 1933 590 1985
rect 642 1933 662 1985
rect 714 1933 734 1985
rect 518 1920 786 1933
rect 570 1868 590 1920
rect 642 1868 662 1920
rect 714 1868 734 1920
rect 518 1855 786 1868
rect 570 1803 590 1855
rect 642 1803 662 1855
rect 714 1803 734 1855
rect 518 1790 786 1803
rect 570 1738 590 1790
rect 642 1738 662 1790
rect 714 1738 734 1790
rect 518 1725 786 1738
rect 570 1673 590 1725
rect 642 1673 662 1725
rect 714 1673 734 1725
rect 518 1660 786 1673
rect 570 1608 590 1660
rect 642 1608 662 1660
rect 714 1608 734 1660
rect 518 1595 786 1608
rect 570 1543 590 1595
rect 642 1543 662 1595
rect 714 1543 734 1595
rect 1061 4119 1251 4125
rect 1061 4067 1066 4119
rect 1118 4067 1130 4119
rect 1182 4067 1194 4119
rect 1246 4067 1251 4119
rect 1061 4054 1251 4067
rect 1061 4002 1066 4054
rect 1118 4002 1130 4054
rect 1182 4002 1194 4054
rect 1246 4002 1251 4054
rect 1061 3989 1251 4002
rect 1061 3937 1066 3989
rect 1118 3937 1130 3989
rect 1182 3937 1194 3989
rect 1246 3937 1251 3989
rect 1061 3924 1251 3937
rect 1061 1568 1066 3924
rect 1246 1568 1251 3924
rect 1061 1562 1251 1568
rect 1557 4124 1747 4130
rect 1557 4072 1562 4124
rect 1614 4072 1626 4124
rect 1678 4072 1690 4124
rect 1742 4072 1747 4124
rect 1557 4059 1747 4072
rect 1557 4007 1562 4059
rect 1614 4007 1626 4059
rect 1678 4007 1690 4059
rect 1742 4007 1747 4059
rect 1557 3994 1747 4007
rect 1557 3942 1562 3994
rect 1614 3942 1626 3994
rect 1678 3942 1690 3994
rect 1742 3942 1747 3994
rect 1557 3929 1747 3942
rect 1557 3877 1562 3929
rect 1614 3877 1626 3929
rect 1678 3877 1690 3929
rect 1742 3877 1747 3929
rect 1557 3864 1747 3877
rect 1557 3812 1562 3864
rect 1614 3812 1626 3864
rect 1678 3812 1690 3864
rect 1742 3812 1747 3864
rect 1557 3799 1747 3812
rect 1557 3747 1562 3799
rect 1614 3747 1626 3799
rect 1678 3747 1690 3799
rect 1742 3747 1747 3799
rect 1557 3734 1747 3747
rect 1557 3682 1562 3734
rect 1614 3682 1626 3734
rect 1678 3682 1690 3734
rect 1742 3682 1747 3734
rect 1557 3669 1747 3682
rect 1557 3617 1562 3669
rect 1614 3617 1626 3669
rect 1678 3617 1690 3669
rect 1742 3617 1747 3669
rect 1557 3604 1747 3617
rect 1557 1568 1562 3604
rect 1742 1568 1747 3604
rect 1557 1562 1747 1568
rect 2053 4119 2243 4125
rect 2053 4067 2058 4119
rect 2110 4067 2122 4119
rect 2174 4067 2186 4119
rect 2238 4067 2243 4119
rect 2053 4054 2243 4067
rect 2053 4002 2058 4054
rect 2110 4002 2122 4054
rect 2174 4002 2186 4054
rect 2238 4002 2243 4054
rect 2053 3989 2243 4002
rect 2053 3937 2058 3989
rect 2110 3937 2122 3989
rect 2174 3937 2186 3989
rect 2238 3937 2243 3989
rect 2053 3924 2243 3937
rect 2053 1568 2058 3924
rect 2238 1568 2243 3924
rect 2053 1562 2243 1568
rect 2549 4124 2739 4130
rect 2549 4072 2554 4124
rect 2606 4072 2618 4124
rect 2670 4072 2682 4124
rect 2734 4072 2739 4124
rect 2549 4059 2739 4072
rect 2549 4007 2554 4059
rect 2606 4007 2618 4059
rect 2670 4007 2682 4059
rect 2734 4007 2739 4059
rect 2549 3994 2739 4007
rect 2549 3942 2554 3994
rect 2606 3942 2618 3994
rect 2670 3942 2682 3994
rect 2734 3942 2739 3994
rect 2549 3929 2739 3942
rect 2549 3877 2554 3929
rect 2606 3877 2618 3929
rect 2670 3877 2682 3929
rect 2734 3877 2739 3929
rect 2549 3864 2739 3877
rect 2549 3812 2554 3864
rect 2606 3812 2618 3864
rect 2670 3812 2682 3864
rect 2734 3812 2739 3864
rect 2549 3799 2739 3812
rect 2549 3747 2554 3799
rect 2606 3747 2618 3799
rect 2670 3747 2682 3799
rect 2734 3747 2739 3799
rect 2549 3734 2739 3747
rect 2549 3682 2554 3734
rect 2606 3682 2618 3734
rect 2670 3682 2682 3734
rect 2734 3682 2739 3734
rect 2549 3669 2739 3682
rect 2549 3617 2554 3669
rect 2606 3617 2618 3669
rect 2670 3617 2682 3669
rect 2734 3617 2739 3669
rect 2549 3604 2739 3617
rect 2549 1568 2554 3604
rect 2734 1568 2739 3604
rect 2549 1562 2739 1568
rect 3045 4119 3235 4125
rect 3045 4067 3050 4119
rect 3102 4067 3114 4119
rect 3166 4067 3178 4119
rect 3230 4067 3235 4119
rect 3045 4054 3235 4067
rect 3045 4002 3050 4054
rect 3102 4002 3114 4054
rect 3166 4002 3178 4054
rect 3230 4002 3235 4054
rect 3045 3989 3235 4002
rect 3045 3937 3050 3989
rect 3102 3937 3114 3989
rect 3166 3937 3178 3989
rect 3230 3937 3235 3989
rect 3045 3924 3235 3937
rect 3045 1568 3050 3924
rect 3230 1568 3235 3924
rect 3045 1562 3235 1568
rect 3541 4124 3731 4130
rect 3541 4072 3546 4124
rect 3598 4072 3610 4124
rect 3662 4072 3674 4124
rect 3726 4072 3731 4124
rect 3541 4059 3731 4072
rect 3541 4007 3546 4059
rect 3598 4007 3610 4059
rect 3662 4007 3674 4059
rect 3726 4007 3731 4059
rect 3541 3994 3731 4007
rect 3541 3942 3546 3994
rect 3598 3942 3610 3994
rect 3662 3942 3674 3994
rect 3726 3942 3731 3994
rect 3541 3929 3731 3942
rect 3541 3877 3546 3929
rect 3598 3877 3610 3929
rect 3662 3877 3674 3929
rect 3726 3877 3731 3929
rect 3541 3864 3731 3877
rect 3541 3812 3546 3864
rect 3598 3812 3610 3864
rect 3662 3812 3674 3864
rect 3726 3812 3731 3864
rect 3541 3799 3731 3812
rect 3541 3747 3546 3799
rect 3598 3747 3610 3799
rect 3662 3747 3674 3799
rect 3726 3747 3731 3799
rect 3541 3734 3731 3747
rect 3541 3682 3546 3734
rect 3598 3682 3610 3734
rect 3662 3682 3674 3734
rect 3726 3682 3731 3734
rect 3541 3669 3731 3682
rect 3541 3617 3546 3669
rect 3598 3617 3610 3669
rect 3662 3617 3674 3669
rect 3726 3617 3731 3669
rect 3541 3604 3731 3617
rect 3541 1568 3546 3604
rect 3726 1568 3731 3604
rect 3541 1562 3731 1568
rect 4037 4119 4227 4125
rect 4037 4067 4042 4119
rect 4094 4067 4106 4119
rect 4158 4067 4170 4119
rect 4222 4067 4227 4119
rect 4037 4054 4227 4067
rect 4037 4002 4042 4054
rect 4094 4002 4106 4054
rect 4158 4002 4170 4054
rect 4222 4002 4227 4054
rect 4037 3989 4227 4002
rect 4037 3937 4042 3989
rect 4094 3937 4106 3989
rect 4158 3937 4170 3989
rect 4222 3937 4227 3989
rect 4037 3924 4227 3937
rect 4037 1568 4042 3924
rect 4222 1568 4227 3924
rect 4037 1562 4227 1568
rect 4533 4124 4723 4130
rect 4533 4072 4538 4124
rect 4590 4072 4602 4124
rect 4654 4072 4666 4124
rect 4718 4072 4723 4124
rect 4533 4059 4723 4072
rect 4533 4007 4538 4059
rect 4590 4007 4602 4059
rect 4654 4007 4666 4059
rect 4718 4007 4723 4059
rect 4533 3994 4723 4007
rect 4533 3942 4538 3994
rect 4590 3942 4602 3994
rect 4654 3942 4666 3994
rect 4718 3942 4723 3994
rect 4533 3929 4723 3942
rect 4533 3877 4538 3929
rect 4590 3877 4602 3929
rect 4654 3877 4666 3929
rect 4718 3877 4723 3929
rect 4533 3864 4723 3877
rect 4533 3812 4538 3864
rect 4590 3812 4602 3864
rect 4654 3812 4666 3864
rect 4718 3812 4723 3864
rect 4533 3799 4723 3812
rect 4533 3747 4538 3799
rect 4590 3747 4602 3799
rect 4654 3747 4666 3799
rect 4718 3747 4723 3799
rect 4533 3734 4723 3747
rect 4533 3682 4538 3734
rect 4590 3682 4602 3734
rect 4654 3682 4666 3734
rect 4718 3682 4723 3734
rect 4533 3669 4723 3682
rect 4533 3617 4538 3669
rect 4590 3617 4602 3669
rect 4654 3617 4666 3669
rect 4718 3617 4723 3669
rect 4533 3604 4723 3617
rect 4533 1568 4538 3604
rect 4718 1568 4723 3604
rect 4533 1562 4723 1568
rect 5029 4119 5219 4125
rect 5029 4067 5034 4119
rect 5086 4067 5098 4119
rect 5150 4067 5162 4119
rect 5214 4067 5219 4119
rect 5029 4054 5219 4067
rect 5029 4002 5034 4054
rect 5086 4002 5098 4054
rect 5150 4002 5162 4054
rect 5214 4002 5219 4054
rect 5029 3989 5219 4002
rect 5029 3937 5034 3989
rect 5086 3937 5098 3989
rect 5150 3937 5162 3989
rect 5214 3937 5219 3989
rect 5029 3924 5219 3937
rect 5029 1568 5034 3924
rect 5214 1568 5219 3924
rect 5029 1562 5219 1568
rect 5525 4124 5715 4130
rect 5525 4072 5530 4124
rect 5582 4072 5594 4124
rect 5646 4072 5658 4124
rect 5710 4072 5715 4124
rect 5525 4059 5715 4072
rect 5525 4007 5530 4059
rect 5582 4007 5594 4059
rect 5646 4007 5658 4059
rect 5710 4007 5715 4059
rect 5525 3994 5715 4007
rect 5525 3942 5530 3994
rect 5582 3942 5594 3994
rect 5646 3942 5658 3994
rect 5710 3942 5715 3994
rect 5525 3929 5715 3942
rect 5525 3877 5530 3929
rect 5582 3877 5594 3929
rect 5646 3877 5658 3929
rect 5710 3877 5715 3929
rect 5525 3864 5715 3877
rect 5525 3812 5530 3864
rect 5582 3812 5594 3864
rect 5646 3812 5658 3864
rect 5710 3812 5715 3864
rect 5525 3799 5715 3812
rect 5525 3747 5530 3799
rect 5582 3747 5594 3799
rect 5646 3747 5658 3799
rect 5710 3747 5715 3799
rect 5525 3734 5715 3747
rect 5525 3682 5530 3734
rect 5582 3682 5594 3734
rect 5646 3682 5658 3734
rect 5710 3682 5715 3734
rect 5525 3669 5715 3682
rect 5525 3617 5530 3669
rect 5582 3617 5594 3669
rect 5646 3617 5658 3669
rect 5710 3617 5715 3669
rect 5525 3604 5715 3617
rect 5525 1568 5530 3604
rect 5710 1568 5715 3604
rect 5525 1562 5715 1568
rect 6021 4119 6211 4125
rect 6021 4067 6026 4119
rect 6078 4067 6090 4119
rect 6142 4067 6154 4119
rect 6206 4067 6211 4119
rect 6021 4054 6211 4067
rect 6021 4002 6026 4054
rect 6078 4002 6090 4054
rect 6142 4002 6154 4054
rect 6206 4002 6211 4054
rect 6021 3989 6211 4002
rect 6021 3937 6026 3989
rect 6078 3937 6090 3989
rect 6142 3937 6154 3989
rect 6206 3937 6211 3989
rect 6021 3924 6211 3937
rect 6021 1568 6026 3924
rect 6206 1568 6211 3924
rect 6021 1562 6211 1568
rect 6517 4124 6707 4130
rect 6517 4072 6522 4124
rect 6574 4072 6586 4124
rect 6638 4072 6650 4124
rect 6702 4072 6707 4124
rect 6517 4059 6707 4072
rect 6517 4007 6522 4059
rect 6574 4007 6586 4059
rect 6638 4007 6650 4059
rect 6702 4007 6707 4059
rect 6517 3994 6707 4007
rect 6517 3942 6522 3994
rect 6574 3942 6586 3994
rect 6638 3942 6650 3994
rect 6702 3942 6707 3994
rect 6517 3929 6707 3942
rect 6517 3877 6522 3929
rect 6574 3877 6586 3929
rect 6638 3877 6650 3929
rect 6702 3877 6707 3929
rect 6517 3864 6707 3877
rect 6517 3812 6522 3864
rect 6574 3812 6586 3864
rect 6638 3812 6650 3864
rect 6702 3812 6707 3864
rect 6517 3799 6707 3812
rect 6517 3747 6522 3799
rect 6574 3747 6586 3799
rect 6638 3747 6650 3799
rect 6702 3747 6707 3799
rect 6517 3734 6707 3747
rect 6517 3682 6522 3734
rect 6574 3682 6586 3734
rect 6638 3682 6650 3734
rect 6702 3682 6707 3734
rect 6517 3669 6707 3682
rect 6517 3617 6522 3669
rect 6574 3617 6586 3669
rect 6638 3617 6650 3669
rect 6702 3617 6707 3669
rect 6517 3604 6707 3617
rect 6517 1568 6522 3604
rect 6702 1568 6707 3604
rect 6517 1562 6707 1568
rect 7013 4119 7203 4125
rect 7013 4067 7018 4119
rect 7070 4067 7082 4119
rect 7134 4067 7146 4119
rect 7198 4067 7203 4119
rect 7013 4054 7203 4067
rect 7013 4002 7018 4054
rect 7070 4002 7082 4054
rect 7134 4002 7146 4054
rect 7198 4002 7203 4054
rect 7013 3989 7203 4002
rect 7013 3937 7018 3989
rect 7070 3937 7082 3989
rect 7134 3937 7146 3989
rect 7198 3937 7203 3989
rect 7013 3924 7203 3937
rect 7013 1568 7018 3924
rect 7198 1568 7203 3924
rect 7013 1562 7203 1568
rect 7509 4124 7699 4130
rect 7509 4072 7514 4124
rect 7566 4072 7578 4124
rect 7630 4072 7642 4124
rect 7694 4072 7699 4124
rect 7509 4059 7699 4072
rect 7509 4007 7514 4059
rect 7566 4007 7578 4059
rect 7630 4007 7642 4059
rect 7694 4007 7699 4059
rect 7509 3994 7699 4007
rect 7509 3942 7514 3994
rect 7566 3942 7578 3994
rect 7630 3942 7642 3994
rect 7694 3942 7699 3994
rect 7509 3929 7699 3942
rect 7509 3877 7514 3929
rect 7566 3877 7578 3929
rect 7630 3877 7642 3929
rect 7694 3877 7699 3929
rect 7509 3864 7699 3877
rect 7509 3812 7514 3864
rect 7566 3812 7578 3864
rect 7630 3812 7642 3864
rect 7694 3812 7699 3864
rect 7509 3799 7699 3812
rect 7509 3747 7514 3799
rect 7566 3747 7578 3799
rect 7630 3747 7642 3799
rect 7694 3747 7699 3799
rect 7509 3734 7699 3747
rect 7509 3682 7514 3734
rect 7566 3682 7578 3734
rect 7630 3682 7642 3734
rect 7694 3682 7699 3734
rect 7509 3669 7699 3682
rect 7509 3617 7514 3669
rect 7566 3617 7578 3669
rect 7630 3617 7642 3669
rect 7694 3617 7699 3669
rect 7509 3604 7699 3617
rect 7509 1568 7514 3604
rect 7694 1568 7699 3604
rect 7509 1562 7699 1568
rect 8005 4119 8195 4125
rect 8005 4067 8010 4119
rect 8062 4067 8074 4119
rect 8126 4067 8138 4119
rect 8190 4067 8195 4119
rect 8005 4054 8195 4067
rect 8005 4002 8010 4054
rect 8062 4002 8074 4054
rect 8126 4002 8138 4054
rect 8190 4002 8195 4054
rect 8005 3989 8195 4002
rect 8005 3937 8010 3989
rect 8062 3937 8074 3989
rect 8126 3937 8138 3989
rect 8190 3937 8195 3989
rect 8005 3924 8195 3937
rect 8005 1568 8010 3924
rect 8190 1568 8195 3924
rect 8005 1562 8195 1568
rect 8501 4124 8691 4130
rect 8501 4072 8506 4124
rect 8558 4072 8570 4124
rect 8622 4072 8634 4124
rect 8686 4072 8691 4124
rect 8501 4059 8691 4072
rect 8501 4007 8506 4059
rect 8558 4007 8570 4059
rect 8622 4007 8634 4059
rect 8686 4007 8691 4059
rect 8501 3994 8691 4007
rect 8501 3942 8506 3994
rect 8558 3942 8570 3994
rect 8622 3942 8634 3994
rect 8686 3942 8691 3994
rect 8501 3929 8691 3942
rect 8501 3877 8506 3929
rect 8558 3877 8570 3929
rect 8622 3877 8634 3929
rect 8686 3877 8691 3929
rect 8501 3864 8691 3877
rect 8501 3812 8506 3864
rect 8558 3812 8570 3864
rect 8622 3812 8634 3864
rect 8686 3812 8691 3864
rect 8501 3799 8691 3812
rect 8501 3747 8506 3799
rect 8558 3747 8570 3799
rect 8622 3747 8634 3799
rect 8686 3747 8691 3799
rect 8501 3734 8691 3747
rect 8501 3682 8506 3734
rect 8558 3682 8570 3734
rect 8622 3682 8634 3734
rect 8686 3682 8691 3734
rect 8501 3669 8691 3682
rect 8501 3617 8506 3669
rect 8558 3617 8570 3669
rect 8622 3617 8634 3669
rect 8686 3617 8691 3669
rect 8501 3604 8691 3617
rect 8501 1568 8506 3604
rect 8686 1568 8691 3604
rect 8501 1562 8691 1568
rect 8997 4119 9187 4125
rect 8997 4067 9002 4119
rect 9054 4067 9066 4119
rect 9118 4067 9130 4119
rect 9182 4067 9187 4119
rect 8997 4054 9187 4067
rect 8997 4002 9002 4054
rect 9054 4002 9066 4054
rect 9118 4002 9130 4054
rect 9182 4002 9187 4054
rect 8997 3989 9187 4002
rect 8997 3937 9002 3989
rect 9054 3937 9066 3989
rect 9118 3937 9130 3989
rect 9182 3937 9187 3989
rect 8997 3924 9187 3937
rect 8997 1568 9002 3924
rect 9182 1568 9187 3924
rect 8997 1562 9187 1568
rect 9493 4124 9683 4130
rect 9493 4072 9498 4124
rect 9550 4072 9562 4124
rect 9614 4072 9626 4124
rect 9678 4072 9683 4124
rect 9493 4059 9683 4072
rect 9493 4007 9498 4059
rect 9550 4007 9562 4059
rect 9614 4007 9626 4059
rect 9678 4007 9683 4059
rect 9493 3994 9683 4007
rect 9493 3942 9498 3994
rect 9550 3942 9562 3994
rect 9614 3942 9626 3994
rect 9678 3942 9683 3994
rect 9493 3929 9683 3942
rect 9493 3877 9498 3929
rect 9550 3877 9562 3929
rect 9614 3877 9626 3929
rect 9678 3877 9683 3929
rect 9493 3864 9683 3877
rect 9493 3812 9498 3864
rect 9550 3812 9562 3864
rect 9614 3812 9626 3864
rect 9678 3812 9683 3864
rect 9493 3799 9683 3812
rect 9493 3747 9498 3799
rect 9550 3747 9562 3799
rect 9614 3747 9626 3799
rect 9678 3747 9683 3799
rect 9493 3734 9683 3747
rect 9493 3682 9498 3734
rect 9550 3682 9562 3734
rect 9614 3682 9626 3734
rect 9678 3682 9683 3734
rect 9493 3669 9683 3682
rect 9493 3617 9498 3669
rect 9550 3617 9562 3669
rect 9614 3617 9626 3669
rect 9678 3617 9683 3669
rect 9493 3604 9683 3617
rect 9493 1568 9498 3604
rect 9678 1568 9683 3604
rect 9493 1562 9683 1568
rect 9989 4119 10179 4125
rect 9989 4067 9994 4119
rect 10046 4067 10058 4119
rect 10110 4067 10122 4119
rect 10174 4067 10179 4119
rect 9989 4054 10179 4067
rect 9989 4002 9994 4054
rect 10046 4002 10058 4054
rect 10110 4002 10122 4054
rect 10174 4002 10179 4054
rect 9989 3989 10179 4002
rect 9989 3937 9994 3989
rect 10046 3937 10058 3989
rect 10110 3937 10122 3989
rect 10174 3937 10179 3989
rect 9989 3924 10179 3937
rect 9989 1568 9994 3924
rect 10174 1568 10179 3924
rect 9989 1562 10179 1568
rect 10485 4124 10675 4130
rect 10485 4072 10490 4124
rect 10542 4072 10554 4124
rect 10606 4072 10618 4124
rect 10670 4072 10675 4124
rect 10485 4059 10675 4072
rect 10485 4007 10490 4059
rect 10542 4007 10554 4059
rect 10606 4007 10618 4059
rect 10670 4007 10675 4059
rect 10485 3994 10675 4007
rect 10485 3942 10490 3994
rect 10542 3942 10554 3994
rect 10606 3942 10618 3994
rect 10670 3942 10675 3994
rect 10485 3929 10675 3942
rect 10485 3877 10490 3929
rect 10542 3877 10554 3929
rect 10606 3877 10618 3929
rect 10670 3877 10675 3929
rect 10485 3864 10675 3877
rect 10485 3812 10490 3864
rect 10542 3812 10554 3864
rect 10606 3812 10618 3864
rect 10670 3812 10675 3864
rect 10485 3799 10675 3812
rect 10485 3747 10490 3799
rect 10542 3747 10554 3799
rect 10606 3747 10618 3799
rect 10670 3747 10675 3799
rect 10485 3734 10675 3747
rect 10485 3682 10490 3734
rect 10542 3682 10554 3734
rect 10606 3682 10618 3734
rect 10670 3682 10675 3734
rect 10485 3669 10675 3682
rect 10485 3617 10490 3669
rect 10542 3617 10554 3669
rect 10606 3617 10618 3669
rect 10670 3617 10675 3669
rect 10485 3604 10675 3617
rect 10485 1568 10490 3604
rect 10670 1568 10675 3604
rect 10485 1562 10675 1568
rect 10981 4119 11171 4125
rect 10981 4067 10986 4119
rect 11038 4067 11050 4119
rect 11102 4067 11114 4119
rect 11166 4067 11171 4119
rect 10981 4054 11171 4067
rect 10981 4002 10986 4054
rect 11038 4002 11050 4054
rect 11102 4002 11114 4054
rect 11166 4002 11171 4054
rect 10981 3989 11171 4002
rect 10981 3937 10986 3989
rect 11038 3937 11050 3989
rect 11102 3937 11114 3989
rect 11166 3937 11171 3989
rect 10981 3924 11171 3937
rect 10981 1568 10986 3924
rect 11166 1568 11171 3924
rect 10981 1562 11171 1568
rect 11477 4124 11667 4130
rect 11477 4072 11482 4124
rect 11534 4072 11546 4124
rect 11598 4072 11610 4124
rect 11662 4072 11667 4124
rect 11477 4059 11667 4072
rect 11477 4007 11482 4059
rect 11534 4007 11546 4059
rect 11598 4007 11610 4059
rect 11662 4007 11667 4059
rect 11477 3994 11667 4007
rect 11477 3942 11482 3994
rect 11534 3942 11546 3994
rect 11598 3942 11610 3994
rect 11662 3942 11667 3994
rect 11477 3929 11667 3942
rect 11477 3877 11482 3929
rect 11534 3877 11546 3929
rect 11598 3877 11610 3929
rect 11662 3877 11667 3929
rect 11477 3864 11667 3877
rect 11477 3812 11482 3864
rect 11534 3812 11546 3864
rect 11598 3812 11610 3864
rect 11662 3812 11667 3864
rect 11477 3799 11667 3812
rect 11477 3747 11482 3799
rect 11534 3747 11546 3799
rect 11598 3747 11610 3799
rect 11662 3747 11667 3799
rect 11477 3734 11667 3747
rect 11477 3682 11482 3734
rect 11534 3682 11546 3734
rect 11598 3682 11610 3734
rect 11662 3682 11667 3734
rect 11477 3669 11667 3682
rect 11477 3617 11482 3669
rect 11534 3617 11546 3669
rect 11598 3617 11610 3669
rect 11662 3617 11667 3669
rect 11477 3604 11667 3617
rect 11477 1568 11482 3604
rect 11662 1568 11667 3604
rect 11477 1562 11667 1568
rect 11973 4119 12163 4125
rect 11973 4067 11978 4119
rect 12030 4067 12042 4119
rect 12094 4067 12106 4119
rect 12158 4067 12163 4119
rect 11973 4054 12163 4067
rect 11973 4002 11978 4054
rect 12030 4002 12042 4054
rect 12094 4002 12106 4054
rect 12158 4002 12163 4054
rect 11973 3989 12163 4002
rect 11973 3937 11978 3989
rect 12030 3937 12042 3989
rect 12094 3937 12106 3989
rect 12158 3937 12163 3989
rect 11973 3924 12163 3937
rect 11973 1568 11978 3924
rect 12158 1568 12163 3924
rect 11973 1562 12163 1568
rect 12469 4124 12659 4130
rect 12469 4072 12474 4124
rect 12526 4072 12538 4124
rect 12590 4072 12602 4124
rect 12654 4072 12659 4124
rect 12469 4059 12659 4072
rect 12469 4007 12474 4059
rect 12526 4007 12538 4059
rect 12590 4007 12602 4059
rect 12654 4007 12659 4059
rect 12469 3994 12659 4007
rect 12469 3942 12474 3994
rect 12526 3942 12538 3994
rect 12590 3942 12602 3994
rect 12654 3942 12659 3994
rect 12469 3929 12659 3942
rect 12469 3877 12474 3929
rect 12526 3877 12538 3929
rect 12590 3877 12602 3929
rect 12654 3877 12659 3929
rect 12469 3864 12659 3877
rect 12469 3812 12474 3864
rect 12526 3812 12538 3864
rect 12590 3812 12602 3864
rect 12654 3812 12659 3864
rect 12469 3799 12659 3812
rect 12469 3747 12474 3799
rect 12526 3747 12538 3799
rect 12590 3747 12602 3799
rect 12654 3747 12659 3799
rect 12469 3734 12659 3747
rect 12469 3682 12474 3734
rect 12526 3682 12538 3734
rect 12590 3682 12602 3734
rect 12654 3682 12659 3734
rect 12469 3669 12659 3682
rect 12469 3617 12474 3669
rect 12526 3617 12538 3669
rect 12590 3617 12602 3669
rect 12654 3617 12659 3669
rect 12469 3604 12659 3617
rect 12469 1568 12474 3604
rect 12654 1568 12659 3604
rect 12469 1562 12659 1568
rect 12965 4119 13155 4125
rect 12965 4067 12970 4119
rect 13022 4067 13034 4119
rect 13086 4067 13098 4119
rect 13150 4067 13155 4119
rect 12965 4054 13155 4067
rect 12965 4002 12970 4054
rect 13022 4002 13034 4054
rect 13086 4002 13098 4054
rect 13150 4002 13155 4054
rect 12965 3989 13155 4002
rect 12965 3937 12970 3989
rect 13022 3937 13034 3989
rect 13086 3937 13098 3989
rect 13150 3937 13155 3989
rect 12965 3924 13155 3937
rect 12965 1568 12970 3924
rect 13150 1568 13155 3924
rect 12965 1562 13155 1568
rect 13461 4124 13651 4130
rect 13461 4072 13466 4124
rect 13518 4072 13530 4124
rect 13582 4072 13594 4124
rect 13646 4072 13651 4124
rect 13461 4059 13651 4072
rect 13461 4007 13466 4059
rect 13518 4007 13530 4059
rect 13582 4007 13594 4059
rect 13646 4007 13651 4059
rect 13461 3994 13651 4007
rect 13461 3942 13466 3994
rect 13518 3942 13530 3994
rect 13582 3942 13594 3994
rect 13646 3942 13651 3994
rect 13461 3929 13651 3942
rect 13461 3877 13466 3929
rect 13518 3877 13530 3929
rect 13582 3877 13594 3929
rect 13646 3877 13651 3929
rect 13461 3864 13651 3877
rect 13461 3812 13466 3864
rect 13518 3812 13530 3864
rect 13582 3812 13594 3864
rect 13646 3812 13651 3864
rect 13461 3799 13651 3812
rect 13461 3747 13466 3799
rect 13518 3747 13530 3799
rect 13582 3747 13594 3799
rect 13646 3747 13651 3799
rect 13461 3734 13651 3747
rect 13461 3682 13466 3734
rect 13518 3682 13530 3734
rect 13582 3682 13594 3734
rect 13646 3682 13651 3734
rect 13461 3669 13651 3682
rect 13461 3617 13466 3669
rect 13518 3617 13530 3669
rect 13582 3617 13594 3669
rect 13646 3617 13651 3669
rect 13461 3604 13651 3617
rect 13461 1568 13466 3604
rect 13646 1568 13651 3604
rect 13461 1562 13651 1568
rect 13991 4124 14135 4130
rect 14043 4072 14083 4124
rect 13991 4060 14135 4072
rect 14043 4008 14083 4060
rect 13991 3996 14135 4008
rect 14043 3944 14083 3996
rect 13991 3932 14135 3944
rect 14043 3880 14083 3932
rect 13991 3868 14135 3880
rect 14043 3816 14083 3868
rect 13991 3804 14135 3816
rect 14043 3752 14083 3804
rect 13991 3740 14135 3752
rect 14043 3688 14083 3740
rect 13991 3676 14135 3688
rect 14043 3624 14083 3676
rect 13991 3612 14135 3624
rect 14043 3560 14083 3612
rect 13991 3548 14135 3560
rect 14043 3496 14083 3548
rect 13991 3484 14135 3496
rect 14043 3432 14083 3484
rect 13991 3420 14135 3432
rect 14043 3368 14083 3420
rect 13991 3356 14135 3368
rect 14043 3304 14083 3356
rect 13991 3292 14135 3304
rect 14043 3240 14083 3292
rect 13991 3228 14135 3240
rect 14043 3176 14083 3228
rect 13991 3164 14135 3176
rect 14043 3112 14083 3164
rect 13991 3100 14135 3112
rect 14043 3048 14083 3100
rect 13991 3036 14135 3048
rect 14043 2984 14083 3036
rect 13991 2972 14135 2984
rect 14043 2920 14083 2972
rect 13991 2908 14135 2920
rect 14043 2856 14083 2908
rect 13991 2844 14135 2856
rect 14043 2792 14083 2844
rect 13991 2780 14135 2792
rect 14043 2728 14083 2780
rect 13991 2716 14135 2728
rect 14043 2664 14083 2716
rect 13991 2652 14135 2664
rect 14043 2600 14083 2652
rect 13991 2588 14135 2600
rect 14043 2536 14083 2588
rect 13991 2524 14135 2536
rect 14043 2472 14083 2524
rect 13991 2460 14135 2472
rect 14043 2408 14083 2460
rect 13991 2396 14135 2408
rect 14043 2344 14083 2396
rect 13991 2332 14135 2344
rect 14043 2280 14083 2332
rect 13991 2268 14135 2280
rect 14043 2216 14083 2268
rect 13991 2204 14135 2216
rect 14043 2152 14083 2204
rect 13991 2140 14135 2152
rect 14043 2088 14083 2140
rect 13991 2075 14135 2088
rect 14043 2023 14083 2075
rect 13991 2010 14135 2023
rect 14043 1958 14083 2010
rect 13991 1945 14135 1958
rect 14043 1893 14083 1945
rect 13991 1880 14135 1893
rect 14043 1828 14083 1880
rect 13991 1815 14135 1828
rect 14043 1763 14083 1815
rect 13991 1750 14135 1763
rect 14043 1698 14083 1750
rect 13991 1685 14135 1698
rect 14043 1633 14083 1685
rect 13991 1620 14135 1633
rect 14043 1568 14083 1620
rect 13991 1562 14135 1568
rect 14350 4124 14618 4130
rect 14402 4072 14422 4124
rect 14474 4072 14494 4124
rect 14546 4072 14566 4124
rect 14350 4059 14618 4072
rect 14402 4007 14422 4059
rect 14474 4007 14494 4059
rect 14546 4007 14566 4059
rect 14350 3994 14618 4007
rect 14402 3942 14422 3994
rect 14474 3942 14494 3994
rect 14546 3942 14566 3994
rect 14350 3929 14618 3942
rect 14402 3877 14422 3929
rect 14474 3877 14494 3929
rect 14546 3877 14566 3929
rect 14350 3864 14618 3877
rect 14402 3812 14422 3864
rect 14474 3812 14494 3864
rect 14546 3812 14566 3864
rect 14350 3799 14618 3812
rect 14402 3747 14422 3799
rect 14474 3747 14494 3799
rect 14546 3747 14566 3799
rect 14350 3734 14618 3747
rect 14402 3682 14422 3734
rect 14474 3682 14494 3734
rect 14546 3682 14566 3734
rect 14350 3669 14618 3682
rect 14402 3617 14422 3669
rect 14474 3617 14494 3669
rect 14546 3617 14566 3669
rect 14350 3604 14618 3617
rect 14402 3552 14422 3604
rect 14474 3552 14494 3604
rect 14546 3552 14566 3604
rect 14350 3540 14618 3552
rect 14402 3488 14422 3540
rect 14474 3488 14494 3540
rect 14546 3488 14566 3540
rect 14350 3476 14618 3488
rect 14402 3424 14422 3476
rect 14474 3424 14494 3476
rect 14546 3424 14566 3476
rect 14350 3412 14618 3424
rect 14402 3360 14422 3412
rect 14474 3360 14494 3412
rect 14546 3360 14566 3412
rect 14350 3348 14618 3360
rect 14402 3296 14422 3348
rect 14474 3296 14494 3348
rect 14546 3296 14566 3348
rect 14350 3284 14618 3296
rect 14402 3232 14422 3284
rect 14474 3232 14494 3284
rect 14546 3232 14566 3284
rect 14350 3220 14618 3232
rect 14402 3168 14422 3220
rect 14474 3168 14494 3220
rect 14546 3168 14566 3220
rect 14350 3156 14618 3168
rect 14402 3104 14422 3156
rect 14474 3104 14494 3156
rect 14546 3104 14566 3156
rect 14350 3092 14618 3104
rect 14402 3040 14422 3092
rect 14474 3040 14494 3092
rect 14546 3040 14566 3092
rect 14350 3028 14618 3040
rect 14402 2976 14422 3028
rect 14474 2976 14494 3028
rect 14546 2976 14566 3028
rect 14350 2964 14618 2976
rect 14402 2912 14422 2964
rect 14474 2912 14494 2964
rect 14546 2912 14566 2964
rect 14350 2900 14618 2912
rect 14402 2848 14422 2900
rect 14474 2848 14494 2900
rect 14546 2848 14566 2900
rect 14350 2836 14618 2848
rect 14402 2784 14422 2836
rect 14474 2784 14494 2836
rect 14546 2784 14566 2836
rect 14350 2772 14618 2784
rect 14402 2720 14422 2772
rect 14474 2720 14494 2772
rect 14546 2720 14566 2772
rect 14350 2708 14618 2720
rect 14402 2656 14422 2708
rect 14474 2656 14494 2708
rect 14546 2656 14566 2708
rect 14350 2644 14618 2656
rect 14402 2592 14422 2644
rect 14474 2592 14494 2644
rect 14546 2592 14566 2644
rect 14350 2580 14618 2592
rect 14402 2528 14422 2580
rect 14474 2528 14494 2580
rect 14546 2528 14566 2580
rect 14350 2516 14618 2528
rect 14402 2464 14422 2516
rect 14474 2464 14494 2516
rect 14546 2464 14566 2516
rect 14350 2452 14618 2464
rect 14402 2400 14422 2452
rect 14474 2400 14494 2452
rect 14546 2400 14566 2452
rect 14350 2388 14618 2400
rect 14402 2336 14422 2388
rect 14474 2336 14494 2388
rect 14546 2336 14566 2388
rect 14350 2324 14618 2336
rect 14402 2272 14422 2324
rect 14474 2272 14494 2324
rect 14546 2272 14566 2324
rect 14350 2260 14618 2272
rect 14402 2208 14422 2260
rect 14474 2208 14494 2260
rect 14546 2208 14566 2260
rect 14350 2196 14618 2208
rect 14402 2144 14422 2196
rect 14474 2144 14494 2196
rect 14546 2144 14566 2196
rect 14350 2132 14618 2144
rect 14402 2080 14422 2132
rect 14474 2080 14494 2132
rect 14546 2080 14566 2132
rect 14350 2068 14618 2080
rect 14402 2016 14422 2068
rect 14474 2016 14494 2068
rect 14546 2016 14566 2068
rect 14350 2004 14618 2016
rect 14402 1952 14422 2004
rect 14474 1952 14494 2004
rect 14546 1952 14566 2004
rect 14350 1940 14618 1952
rect 14402 1888 14422 1940
rect 14474 1888 14494 1940
rect 14546 1888 14566 1940
rect 14350 1876 14618 1888
rect 14402 1824 14422 1876
rect 14474 1824 14494 1876
rect 14546 1824 14566 1876
rect 14350 1812 14618 1824
rect 14402 1760 14422 1812
rect 14474 1760 14494 1812
rect 14546 1760 14566 1812
rect 14350 1748 14618 1760
rect 14402 1696 14422 1748
rect 14474 1696 14494 1748
rect 14546 1696 14566 1748
rect 14350 1684 14618 1696
rect 14402 1632 14422 1684
rect 14474 1632 14494 1684
rect 14546 1632 14566 1684
rect 14350 1620 14618 1632
rect 14402 1568 14422 1620
rect 14474 1568 14494 1620
rect 14546 1568 14566 1620
rect 14350 1562 14618 1568
rect 518 1530 786 1543
rect 570 1478 590 1530
rect 642 1478 662 1530
rect 714 1478 734 1530
rect 518 1465 786 1478
rect 570 1413 590 1465
rect 642 1413 662 1465
rect 714 1413 734 1465
rect 518 1400 786 1413
rect 570 1348 590 1400
rect 642 1348 662 1400
rect 714 1348 734 1400
rect 518 1335 786 1348
rect 570 1283 590 1335
rect 642 1283 662 1335
rect 714 1283 734 1335
rect 518 1270 786 1283
rect 570 1218 590 1270
rect 642 1218 662 1270
rect 714 1218 734 1270
rect 518 1205 786 1218
rect 570 1153 590 1205
rect 642 1153 662 1205
rect 714 1153 734 1205
rect 518 1140 786 1153
rect 570 1088 590 1140
rect 642 1088 662 1140
rect 714 1088 734 1140
rect 518 1075 786 1088
rect 570 1023 590 1075
rect 642 1023 662 1075
rect 714 1023 734 1075
rect 518 1010 786 1023
rect 570 958 590 1010
rect 642 958 662 1010
rect 714 958 734 1010
rect 518 945 786 958
rect 570 893 590 945
rect 642 893 662 945
rect 714 893 734 945
rect 518 880 786 893
rect 570 828 590 880
rect 642 828 662 880
rect 714 828 734 880
rect 518 822 786 828
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_0
timestamp 1704896540
transform -1 0 14401 0 1 3152
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_1
timestamp 1704896540
transform -1 0 14401 0 1 1552
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_2
timestamp 1704896540
transform -1 0 8164 0 1 1552
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_3
timestamp 1704896540
transform -1 0 7172 0 1 1552
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_4
timestamp 1704896540
transform -1 0 6180 0 1 1552
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_5
timestamp 1704896540
transform -1 0 5188 0 1 1552
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_6
timestamp 1704896540
transform -1 0 4196 0 1 1552
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_7
timestamp 1704896540
transform -1 0 3204 0 1 1552
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_8
timestamp 1704896540
transform -1 0 2212 0 1 1552
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_9
timestamp 1704896540
transform -1 0 1220 0 1 1552
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_10
timestamp 1704896540
transform -1 0 9156 0 1 1552
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_11
timestamp 1704896540
transform -1 0 10148 0 1 1552
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_12
timestamp 1704896540
transform -1 0 11140 0 1 1552
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_13
timestamp 1704896540
transform -1 0 12132 0 1 1552
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_14
timestamp 1704896540
transform -1 0 13124 0 1 1552
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_15
timestamp 1704896540
transform -1 0 13124 0 1 3152
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_16
timestamp 1704896540
transform -1 0 12132 0 1 3152
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_17
timestamp 1704896540
transform -1 0 11140 0 1 3152
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_18
timestamp 1704896540
transform -1 0 10148 0 1 3152
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_19
timestamp 1704896540
transform -1 0 9156 0 1 3152
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_20
timestamp 1704896540
transform -1 0 1220 0 1 3152
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_21
timestamp 1704896540
transform -1 0 2212 0 1 3152
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_22
timestamp 1704896540
transform -1 0 3204 0 1 3152
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_23
timestamp 1704896540
transform -1 0 4196 0 1 3152
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_24
timestamp 1704896540
transform -1 0 5188 0 1 3152
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_25
timestamp 1704896540
transform -1 0 6180 0 1 3152
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_26
timestamp 1704896540
transform -1 0 7172 0 1 3152
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_27
timestamp 1704896540
transform -1 0 8164 0 1 3152
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_28
timestamp 1704896540
transform 1 0 734 0 1 3152
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_29
timestamp 1704896540
transform 1 0 13988 0 1 3152
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_30
timestamp 1704896540
transform 1 0 13988 0 1 1552
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_31
timestamp 1704896540
transform 1 0 734 0 1 1552
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_32
timestamp 1704896540
transform 1 0 8036 0 1 1552
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_33
timestamp 1704896540
transform 1 0 7044 0 1 1552
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_34
timestamp 1704896540
transform 1 0 6052 0 1 1552
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_35
timestamp 1704896540
transform 1 0 5060 0 1 1552
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_36
timestamp 1704896540
transform 1 0 1092 0 1 1552
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_37
timestamp 1704896540
transform 1 0 2084 0 1 1552
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_38
timestamp 1704896540
transform 1 0 3076 0 1 1552
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_39
timestamp 1704896540
transform 1 0 4068 0 1 1552
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_40
timestamp 1704896540
transform 1 0 9028 0 1 1552
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_41
timestamp 1704896540
transform 1 0 10020 0 1 1552
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_42
timestamp 1704896540
transform 1 0 11012 0 1 1552
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_43
timestamp 1704896540
transform 1 0 12004 0 1 1552
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_44
timestamp 1704896540
transform 1 0 12996 0 1 1552
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_45
timestamp 1704896540
transform 1 0 12996 0 1 3152
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_46
timestamp 1704896540
transform 1 0 12004 0 1 3152
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_47
timestamp 1704896540
transform 1 0 11012 0 1 3152
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_48
timestamp 1704896540
transform 1 0 10020 0 1 3152
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_49
timestamp 1704896540
transform 1 0 9028 0 1 3152
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_50
timestamp 1704896540
transform 1 0 4068 0 1 3152
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_51
timestamp 1704896540
transform 1 0 3076 0 1 3152
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_52
timestamp 1704896540
transform 1 0 2084 0 1 3152
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_53
timestamp 1704896540
transform 1 0 1092 0 1 3152
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_54
timestamp 1704896540
transform 1 0 5060 0 1 3152
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_55
timestamp 1704896540
transform 1 0 6052 0 1 3152
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_56
timestamp 1704896540
transform 1 0 7044 0 1 3152
box -36 -36 92 1036
use hvDFL1sd2_CDNS_524688791850  hvDFL1sd2_CDNS_524688791850_57
timestamp 1704896540
transform 1 0 8036 0 1 3152
box -36 -36 92 1036
use L1M1_C_CDNS_524688791851  L1M1_C_CDNS_524688791851_0
timestamp 1704896540
transform -1 0 140 0 1 348
box -101 -29 29 4709
use L1M1_C_CDNS_524688791851  L1M1_C_CDNS_524688791851_1
timestamp 1704896540
transform -1 0 14924 0 1 365
box -101 -29 29 4709
use L1M1_C_CDNS_524688791852  L1M1_C_CDNS_524688791852_0
timestamp 1704896540
transform 1 0 14195 0 1 1197
box 0 0 1 1
use L1M1_C_CDNS_524688791852  L1M1_C_CDNS_524688791852_1
timestamp 1704896540
transform 1 0 13837 0 1 1197
box 0 0 1 1
use L1M1_C_CDNS_524688791852  L1M1_C_CDNS_524688791852_2
timestamp 1704896540
transform 1 0 12845 0 1 1197
box 0 0 1 1
use L1M1_C_CDNS_524688791852  L1M1_C_CDNS_524688791852_3
timestamp 1704896540
transform 1 0 13275 0 1 1197
box 0 0 1 1
use L1M1_C_CDNS_524688791852  L1M1_C_CDNS_524688791852_4
timestamp 1704896540
transform 1 0 12283 0 1 1197
box 0 0 1 1
use L1M1_C_CDNS_524688791852  L1M1_C_CDNS_524688791852_5
timestamp 1704896540
transform 1 0 11853 0 1 1197
box 0 0 1 1
use L1M1_C_CDNS_524688791852  L1M1_C_CDNS_524688791852_6
timestamp 1704896540
transform 1 0 8315 0 1 1197
box 0 0 1 1
use L1M1_C_CDNS_524688791852  L1M1_C_CDNS_524688791852_7
timestamp 1704896540
transform 1 0 7323 0 1 1197
box 0 0 1 1
use L1M1_C_CDNS_524688791852  L1M1_C_CDNS_524688791852_8
timestamp 1704896540
transform 1 0 6331 0 1 1197
box 0 0 1 1
use L1M1_C_CDNS_524688791852  L1M1_C_CDNS_524688791852_9
timestamp 1704896540
transform 1 0 5339 0 1 1197
box 0 0 1 1
use L1M1_C_CDNS_524688791852  L1M1_C_CDNS_524688791852_10
timestamp 1704896540
transform 1 0 4347 0 1 1197
box 0 0 1 1
use L1M1_C_CDNS_524688791852  L1M1_C_CDNS_524688791852_11
timestamp 1704896540
transform 1 0 3355 0 1 1197
box 0 0 1 1
use L1M1_C_CDNS_524688791852  L1M1_C_CDNS_524688791852_12
timestamp 1704896540
transform 1 0 2363 0 1 1197
box 0 0 1 1
use L1M1_C_CDNS_524688791852  L1M1_C_CDNS_524688791852_13
timestamp 1704896540
transform 1 0 9307 0 1 1197
box 0 0 1 1
use L1M1_C_CDNS_524688791852  L1M1_C_CDNS_524688791852_14
timestamp 1704896540
transform 1 0 10299 0 1 1197
box 0 0 1 1
use L1M1_C_CDNS_524688791852  L1M1_C_CDNS_524688791852_15
timestamp 1704896540
transform 1 0 11291 0 1 1197
box 0 0 1 1
use L1M1_C_CDNS_524688791852  L1M1_C_CDNS_524688791852_16
timestamp 1704896540
transform 1 0 8877 0 1 1197
box 0 0 1 1
use L1M1_C_CDNS_524688791852  L1M1_C_CDNS_524688791852_17
timestamp 1704896540
transform 1 0 9869 0 1 1197
box 0 0 1 1
use L1M1_C_CDNS_524688791852  L1M1_C_CDNS_524688791852_18
timestamp 1704896540
transform 1 0 10861 0 1 1197
box 0 0 1 1
use L1M1_C_CDNS_524688791852  L1M1_C_CDNS_524688791852_19
timestamp 1704896540
transform 1 0 1933 0 1 1197
box 0 0 1 1
use L1M1_C_CDNS_524688791852  L1M1_C_CDNS_524688791852_20
timestamp 1704896540
transform 1 0 2925 0 1 1197
box 0 0 1 1
use L1M1_C_CDNS_524688791852  L1M1_C_CDNS_524688791852_21
timestamp 1704896540
transform 1 0 3917 0 1 1197
box 0 0 1 1
use L1M1_C_CDNS_524688791852  L1M1_C_CDNS_524688791852_22
timestamp 1704896540
transform 1 0 4909 0 1 1197
box 0 0 1 1
use L1M1_C_CDNS_524688791852  L1M1_C_CDNS_524688791852_23
timestamp 1704896540
transform 1 0 5901 0 1 1197
box 0 0 1 1
use L1M1_C_CDNS_524688791852  L1M1_C_CDNS_524688791852_24
timestamp 1704896540
transform 1 0 6893 0 1 1197
box 0 0 1 1
use L1M1_C_CDNS_524688791852  L1M1_C_CDNS_524688791852_25
timestamp 1704896540
transform 1 0 7885 0 1 1197
box 0 0 1 1
use L1M1_C_CDNS_524688791852  L1M1_C_CDNS_524688791852_26
timestamp 1704896540
transform 1 0 1371 0 1 1197
box 0 0 1 1
use L1M1_C_CDNS_524688791853  L1M1_C_CDNS_524688791853_0
timestamp 1704896540
transform 1 0 941 0 1 1197
box 0 0 1 1
use pfet_CDNS_524688791851  pfet_CDNS_524688791851_0
timestamp 1704896540
transform 1 0 14135 0 1 3152
box -116 -66 236 1066
use pfet_CDNS_524688791851  pfet_CDNS_524688791851_1
timestamp 1704896540
transform 1 0 14135 0 1 1552
box -116 -66 236 1066
use pfet_CDNS_524688791852  pfet_CDNS_524688791852_0
timestamp 1704896540
transform 1 0 881 0 -1 2552
box -116 -66 13132 1066
use pfet_CDNS_524688791852  pfet_CDNS_524688791852_1
timestamp 1704896540
transform 1 0 881 0 1 3152
box -116 -66 13132 1066
<< properties >>
string GDS_END 13650052
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 12852134
string path 326.500 103.125 326.500 39.050 
<< end >>
