magic
tech sky130A
timestamp 1704896540
<< viali >>
rect 0 0 197 161
<< metal1 >>
rect -6 161 203 164
rect -6 0 0 161
rect 197 0 203 161
rect -6 -3 203 0
<< properties >>
string GDS_END 95652916
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 95650864
<< end >>
