magic
tech sky130A
timestamp 1704896540
<< metal1 >>
rect 0 0 3 346
rect 93 0 96 346
<< via1 >>
rect 3 0 93 346
<< metal2 >>
rect 0 0 3 346
rect 93 0 96 346
<< properties >>
string GDS_END 85845108
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 85842864
<< end >>
