magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -119 -66 375 366
<< mvpmos >>
rect 0 0 100 300
rect 156 0 256 300
<< mvpdiff >>
rect -50 0 0 300
rect 256 0 306 300
<< poly >>
rect 0 300 100 326
rect 0 -26 100 0
rect 156 300 256 326
rect 156 -26 256 0
<< metal1 >>
rect -51 -16 -5 258
rect 105 -16 151 258
rect 261 -16 307 258
use hvDFM1sd2_CDNS_52468879185879  hvDFM1sd2_CDNS_52468879185879_0
timestamp 1704896540
transform 1 0 100 0 1 0
box -36 -36 92 336
use hvDFM1sd_CDNS_52468879185274  hvDFM1sd_CDNS_52468879185274_0
timestamp 1704896540
transform -1 0 0 0 1 0
box -36 -36 89 336
use hvDFM1sd_CDNS_52468879185274  hvDFM1sd_CDNS_52468879185274_1
timestamp 1704896540
transform 1 0 256 0 1 0
box -36 -36 89 336
<< labels >>
flabel comment s -28 121 -28 121 0 FreeSans 300 0 0 0 S
flabel comment s 128 121 128 121 0 FreeSans 300 0 0 0 D
flabel comment s 284 121 284 121 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 86840128
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 86838610
<< end >>
