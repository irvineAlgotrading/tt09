magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< pwell >>
rect 0 66 676 720
<< nmoslvt >>
rect 194 92 224 694
rect 280 92 310 694
rect 366 92 396 694
rect 452 92 482 694
<< ndiff >>
rect 138 682 194 694
rect 138 648 149 682
rect 183 648 194 682
rect 138 614 194 648
rect 138 580 149 614
rect 183 580 194 614
rect 138 546 194 580
rect 138 512 149 546
rect 183 512 194 546
rect 138 478 194 512
rect 138 444 149 478
rect 183 444 194 478
rect 138 410 194 444
rect 138 376 149 410
rect 183 376 194 410
rect 138 342 194 376
rect 138 308 149 342
rect 183 308 194 342
rect 138 274 194 308
rect 138 240 149 274
rect 183 240 194 274
rect 138 206 194 240
rect 138 172 149 206
rect 183 172 194 206
rect 138 138 194 172
rect 138 104 149 138
rect 183 104 194 138
rect 138 92 194 104
rect 224 682 280 694
rect 224 648 235 682
rect 269 648 280 682
rect 224 614 280 648
rect 224 580 235 614
rect 269 580 280 614
rect 224 546 280 580
rect 224 512 235 546
rect 269 512 280 546
rect 224 478 280 512
rect 224 444 235 478
rect 269 444 280 478
rect 224 410 280 444
rect 224 376 235 410
rect 269 376 280 410
rect 224 342 280 376
rect 224 308 235 342
rect 269 308 280 342
rect 224 274 280 308
rect 224 240 235 274
rect 269 240 280 274
rect 224 206 280 240
rect 224 172 235 206
rect 269 172 280 206
rect 224 138 280 172
rect 224 104 235 138
rect 269 104 280 138
rect 224 92 280 104
rect 310 682 366 694
rect 310 648 321 682
rect 355 648 366 682
rect 310 614 366 648
rect 310 580 321 614
rect 355 580 366 614
rect 310 546 366 580
rect 310 512 321 546
rect 355 512 366 546
rect 310 478 366 512
rect 310 444 321 478
rect 355 444 366 478
rect 310 410 366 444
rect 310 376 321 410
rect 355 376 366 410
rect 310 342 366 376
rect 310 308 321 342
rect 355 308 366 342
rect 310 274 366 308
rect 310 240 321 274
rect 355 240 366 274
rect 310 206 366 240
rect 310 172 321 206
rect 355 172 366 206
rect 310 138 366 172
rect 310 104 321 138
rect 355 104 366 138
rect 310 92 366 104
rect 396 682 452 694
rect 396 648 407 682
rect 441 648 452 682
rect 396 614 452 648
rect 396 580 407 614
rect 441 580 452 614
rect 396 546 452 580
rect 396 512 407 546
rect 441 512 452 546
rect 396 478 452 512
rect 396 444 407 478
rect 441 444 452 478
rect 396 410 452 444
rect 396 376 407 410
rect 441 376 452 410
rect 396 342 452 376
rect 396 308 407 342
rect 441 308 452 342
rect 396 274 452 308
rect 396 240 407 274
rect 441 240 452 274
rect 396 206 452 240
rect 396 172 407 206
rect 441 172 452 206
rect 396 138 452 172
rect 396 104 407 138
rect 441 104 452 138
rect 396 92 452 104
rect 482 682 538 694
rect 482 648 493 682
rect 527 648 538 682
rect 482 614 538 648
rect 482 580 493 614
rect 527 580 538 614
rect 482 546 538 580
rect 482 512 493 546
rect 527 512 538 546
rect 482 478 538 512
rect 482 444 493 478
rect 527 444 538 478
rect 482 410 538 444
rect 482 376 493 410
rect 527 376 538 410
rect 482 342 538 376
rect 482 308 493 342
rect 527 308 538 342
rect 482 274 538 308
rect 482 240 493 274
rect 527 240 538 274
rect 482 206 538 240
rect 482 172 493 206
rect 527 172 538 206
rect 482 138 538 172
rect 482 104 493 138
rect 527 104 538 138
rect 482 92 538 104
<< ndiffc >>
rect 149 648 183 682
rect 149 580 183 614
rect 149 512 183 546
rect 149 444 183 478
rect 149 376 183 410
rect 149 308 183 342
rect 149 240 183 274
rect 149 172 183 206
rect 149 104 183 138
rect 235 648 269 682
rect 235 580 269 614
rect 235 512 269 546
rect 235 444 269 478
rect 235 376 269 410
rect 235 308 269 342
rect 235 240 269 274
rect 235 172 269 206
rect 235 104 269 138
rect 321 648 355 682
rect 321 580 355 614
rect 321 512 355 546
rect 321 444 355 478
rect 321 376 355 410
rect 321 308 355 342
rect 321 240 355 274
rect 321 172 355 206
rect 321 104 355 138
rect 407 648 441 682
rect 407 580 441 614
rect 407 512 441 546
rect 407 444 441 478
rect 407 376 441 410
rect 407 308 441 342
rect 407 240 441 274
rect 407 172 441 206
rect 407 104 441 138
rect 493 648 527 682
rect 493 580 527 614
rect 493 512 527 546
rect 493 444 527 478
rect 493 376 527 410
rect 493 308 527 342
rect 493 240 527 274
rect 493 172 527 206
rect 493 104 527 138
<< psubdiff >>
rect 26 648 84 694
rect 26 614 38 648
rect 72 614 84 648
rect 26 580 84 614
rect 26 546 38 580
rect 72 546 84 580
rect 26 512 84 546
rect 26 478 38 512
rect 72 478 84 512
rect 26 444 84 478
rect 26 410 38 444
rect 72 410 84 444
rect 26 376 84 410
rect 26 342 38 376
rect 72 342 84 376
rect 26 308 84 342
rect 26 274 38 308
rect 72 274 84 308
rect 26 240 84 274
rect 26 206 38 240
rect 72 206 84 240
rect 26 172 84 206
rect 26 138 38 172
rect 72 138 84 172
rect 26 92 84 138
rect 592 648 650 694
rect 592 614 604 648
rect 638 614 650 648
rect 592 580 650 614
rect 592 546 604 580
rect 638 546 650 580
rect 592 512 650 546
rect 592 478 604 512
rect 638 478 650 512
rect 592 444 650 478
rect 592 410 604 444
rect 638 410 650 444
rect 592 376 650 410
rect 592 342 604 376
rect 638 342 650 376
rect 592 308 650 342
rect 592 274 604 308
rect 638 274 650 308
rect 592 240 650 274
rect 592 206 604 240
rect 638 206 650 240
rect 592 172 650 206
rect 592 138 604 172
rect 638 138 650 172
rect 592 92 650 138
<< psubdiffcont >>
rect 38 614 72 648
rect 38 546 72 580
rect 38 478 72 512
rect 38 410 72 444
rect 38 342 72 376
rect 38 274 72 308
rect 38 206 72 240
rect 38 138 72 172
rect 604 614 638 648
rect 604 546 638 580
rect 604 478 638 512
rect 604 410 638 444
rect 604 342 638 376
rect 604 274 638 308
rect 604 206 638 240
rect 604 138 638 172
<< poly >>
rect 169 766 507 786
rect 169 732 185 766
rect 219 732 253 766
rect 287 732 321 766
rect 355 732 389 766
rect 423 732 457 766
rect 491 732 507 766
rect 169 716 507 732
rect 194 694 224 716
rect 280 694 310 716
rect 366 694 396 716
rect 452 694 482 716
rect 194 70 224 92
rect 280 70 310 92
rect 366 70 396 92
rect 452 70 482 92
rect 169 54 507 70
rect 169 20 185 54
rect 219 20 253 54
rect 287 20 321 54
rect 355 20 389 54
rect 423 20 457 54
rect 491 20 507 54
rect 169 0 507 20
<< polycont >>
rect 185 732 219 766
rect 253 732 287 766
rect 321 732 355 766
rect 389 732 423 766
rect 457 732 491 766
rect 185 20 219 54
rect 253 20 287 54
rect 321 20 355 54
rect 389 20 423 54
rect 457 20 491 54
<< locali >>
rect 169 732 177 766
rect 219 732 249 766
rect 287 732 321 766
rect 355 732 389 766
rect 427 732 457 766
rect 499 732 507 766
rect 149 682 183 698
rect 38 662 72 664
rect 38 590 72 614
rect 38 518 72 546
rect 38 446 72 478
rect 38 376 72 410
rect 38 308 72 340
rect 38 240 72 268
rect 38 172 72 196
rect 38 122 72 124
rect 149 614 183 628
rect 149 546 183 556
rect 149 478 183 484
rect 149 410 183 412
rect 149 374 183 376
rect 149 302 183 308
rect 149 230 183 240
rect 149 158 183 172
rect 149 88 183 104
rect 235 682 269 698
rect 235 614 269 628
rect 235 546 269 556
rect 235 478 269 484
rect 235 410 269 412
rect 235 374 269 376
rect 235 302 269 308
rect 235 230 269 240
rect 235 158 269 172
rect 235 88 269 104
rect 321 682 355 698
rect 321 614 355 628
rect 321 546 355 556
rect 321 478 355 484
rect 321 410 355 412
rect 321 374 355 376
rect 321 302 355 308
rect 321 230 355 240
rect 321 158 355 172
rect 321 88 355 104
rect 407 682 441 698
rect 407 614 441 628
rect 407 546 441 556
rect 407 478 441 484
rect 407 410 441 412
rect 407 374 441 376
rect 407 302 441 308
rect 407 230 441 240
rect 407 158 441 172
rect 407 88 441 104
rect 493 682 527 698
rect 493 614 527 628
rect 493 546 527 556
rect 493 478 527 484
rect 493 410 527 412
rect 493 374 527 376
rect 493 302 527 308
rect 493 230 527 240
rect 493 158 527 172
rect 604 662 638 664
rect 604 590 638 614
rect 604 518 638 546
rect 604 446 638 478
rect 604 376 638 410
rect 604 308 638 340
rect 604 240 638 268
rect 604 172 638 196
rect 604 122 638 124
rect 493 88 527 104
rect 169 20 177 54
rect 219 20 249 54
rect 287 20 321 54
rect 355 20 389 54
rect 427 20 457 54
rect 499 20 507 54
<< viali >>
rect 177 732 185 766
rect 185 732 211 766
rect 249 732 253 766
rect 253 732 283 766
rect 321 732 355 766
rect 393 732 423 766
rect 423 732 427 766
rect 465 732 491 766
rect 491 732 499 766
rect 38 648 72 662
rect 38 628 72 648
rect 38 580 72 590
rect 38 556 72 580
rect 38 512 72 518
rect 38 484 72 512
rect 38 444 72 446
rect 38 412 72 444
rect 38 342 72 374
rect 38 340 72 342
rect 38 274 72 302
rect 38 268 72 274
rect 38 206 72 230
rect 38 196 72 206
rect 38 138 72 158
rect 38 124 72 138
rect 149 648 183 662
rect 149 628 183 648
rect 149 580 183 590
rect 149 556 183 580
rect 149 512 183 518
rect 149 484 183 512
rect 149 444 183 446
rect 149 412 183 444
rect 149 342 183 374
rect 149 340 183 342
rect 149 274 183 302
rect 149 268 183 274
rect 149 206 183 230
rect 149 196 183 206
rect 149 138 183 158
rect 149 124 183 138
rect 235 648 269 662
rect 235 628 269 648
rect 235 580 269 590
rect 235 556 269 580
rect 235 512 269 518
rect 235 484 269 512
rect 235 444 269 446
rect 235 412 269 444
rect 235 342 269 374
rect 235 340 269 342
rect 235 274 269 302
rect 235 268 269 274
rect 235 206 269 230
rect 235 196 269 206
rect 235 138 269 158
rect 235 124 269 138
rect 321 648 355 662
rect 321 628 355 648
rect 321 580 355 590
rect 321 556 355 580
rect 321 512 355 518
rect 321 484 355 512
rect 321 444 355 446
rect 321 412 355 444
rect 321 342 355 374
rect 321 340 355 342
rect 321 274 355 302
rect 321 268 355 274
rect 321 206 355 230
rect 321 196 355 206
rect 321 138 355 158
rect 321 124 355 138
rect 407 648 441 662
rect 407 628 441 648
rect 407 580 441 590
rect 407 556 441 580
rect 407 512 441 518
rect 407 484 441 512
rect 407 444 441 446
rect 407 412 441 444
rect 407 342 441 374
rect 407 340 441 342
rect 407 274 441 302
rect 407 268 441 274
rect 407 206 441 230
rect 407 196 441 206
rect 407 138 441 158
rect 407 124 441 138
rect 493 648 527 662
rect 493 628 527 648
rect 493 580 527 590
rect 493 556 527 580
rect 493 512 527 518
rect 493 484 527 512
rect 493 444 527 446
rect 493 412 527 444
rect 493 342 527 374
rect 493 340 527 342
rect 493 274 527 302
rect 493 268 527 274
rect 493 206 527 230
rect 493 196 527 206
rect 493 138 527 158
rect 493 124 527 138
rect 604 648 638 662
rect 604 628 638 648
rect 604 580 638 590
rect 604 556 638 580
rect 604 512 638 518
rect 604 484 638 512
rect 604 444 638 446
rect 604 412 638 444
rect 604 342 638 374
rect 604 340 638 342
rect 604 274 638 302
rect 604 268 638 274
rect 604 206 638 230
rect 604 196 638 206
rect 604 138 638 158
rect 604 124 638 138
rect 177 20 185 54
rect 185 20 211 54
rect 249 20 253 54
rect 253 20 283 54
rect 321 20 355 54
rect 393 20 423 54
rect 423 20 427 54
rect 465 20 491 54
rect 491 20 499 54
<< metal1 >>
rect 165 766 511 786
rect 165 732 177 766
rect 211 732 249 766
rect 283 732 321 766
rect 355 732 393 766
rect 427 732 465 766
rect 499 732 511 766
rect 165 720 511 732
rect 26 662 84 674
rect 26 628 38 662
rect 72 628 84 662
rect 26 590 84 628
rect 26 556 38 590
rect 72 556 84 590
rect 26 518 84 556
rect 26 484 38 518
rect 72 484 84 518
rect 26 446 84 484
rect 26 412 38 446
rect 72 412 84 446
rect 26 374 84 412
rect 26 340 38 374
rect 72 340 84 374
rect 26 302 84 340
rect 26 268 38 302
rect 72 268 84 302
rect 26 230 84 268
rect 26 196 38 230
rect 72 196 84 230
rect 26 158 84 196
rect 26 124 38 158
rect 72 124 84 158
rect 26 112 84 124
rect 140 662 192 674
rect 140 628 149 662
rect 183 628 192 662
rect 140 590 192 628
rect 140 556 149 590
rect 183 556 192 590
rect 140 518 192 556
rect 140 484 149 518
rect 183 484 192 518
rect 140 446 192 484
rect 140 412 149 446
rect 183 412 192 446
rect 140 374 192 412
rect 140 362 149 374
rect 183 362 192 374
rect 140 302 192 310
rect 140 298 149 302
rect 183 298 192 302
rect 140 234 192 246
rect 140 170 192 182
rect 140 112 192 118
rect 226 668 278 674
rect 226 604 278 616
rect 226 540 278 552
rect 226 484 235 488
rect 269 484 278 488
rect 226 476 278 484
rect 226 412 235 424
rect 269 412 278 424
rect 226 374 278 412
rect 226 340 235 374
rect 269 340 278 374
rect 226 302 278 340
rect 226 268 235 302
rect 269 268 278 302
rect 226 230 278 268
rect 226 196 235 230
rect 269 196 278 230
rect 226 158 278 196
rect 226 124 235 158
rect 269 124 278 158
rect 226 112 278 124
rect 312 662 364 674
rect 312 628 321 662
rect 355 628 364 662
rect 312 590 364 628
rect 312 556 321 590
rect 355 556 364 590
rect 312 518 364 556
rect 312 484 321 518
rect 355 484 364 518
rect 312 446 364 484
rect 312 412 321 446
rect 355 412 364 446
rect 312 374 364 412
rect 312 362 321 374
rect 355 362 364 374
rect 312 302 364 310
rect 312 298 321 302
rect 355 298 364 302
rect 312 234 364 246
rect 312 170 364 182
rect 312 112 364 118
rect 398 668 450 674
rect 398 604 450 616
rect 398 540 450 552
rect 398 484 407 488
rect 441 484 450 488
rect 398 476 450 484
rect 398 412 407 424
rect 441 412 450 424
rect 398 374 450 412
rect 398 340 407 374
rect 441 340 450 374
rect 398 302 450 340
rect 398 268 407 302
rect 441 268 450 302
rect 398 230 450 268
rect 398 196 407 230
rect 441 196 450 230
rect 398 158 450 196
rect 398 124 407 158
rect 441 124 450 158
rect 398 112 450 124
rect 484 662 536 674
rect 484 628 493 662
rect 527 628 536 662
rect 484 590 536 628
rect 484 556 493 590
rect 527 556 536 590
rect 484 518 536 556
rect 484 484 493 518
rect 527 484 536 518
rect 484 446 536 484
rect 484 412 493 446
rect 527 412 536 446
rect 484 374 536 412
rect 484 362 493 374
rect 527 362 536 374
rect 484 302 536 310
rect 484 298 493 302
rect 527 298 536 302
rect 484 234 536 246
rect 484 170 536 182
rect 484 112 536 118
rect 592 662 650 674
rect 592 628 604 662
rect 638 628 650 662
rect 592 590 650 628
rect 592 556 604 590
rect 638 556 650 590
rect 592 518 650 556
rect 592 484 604 518
rect 638 484 650 518
rect 592 446 650 484
rect 592 412 604 446
rect 638 412 650 446
rect 592 374 650 412
rect 592 340 604 374
rect 638 340 650 374
rect 592 302 650 340
rect 592 268 604 302
rect 638 268 650 302
rect 592 230 650 268
rect 592 196 604 230
rect 638 196 650 230
rect 592 158 650 196
rect 592 124 604 158
rect 638 124 650 158
rect 592 112 650 124
rect 165 54 511 66
rect 165 20 177 54
rect 211 20 249 54
rect 283 20 321 54
rect 355 20 393 54
rect 427 20 465 54
rect 499 20 511 54
rect 165 0 511 20
<< via1 >>
rect 140 340 149 362
rect 149 340 183 362
rect 183 340 192 362
rect 140 310 192 340
rect 140 268 149 298
rect 149 268 183 298
rect 183 268 192 298
rect 140 246 192 268
rect 140 230 192 234
rect 140 196 149 230
rect 149 196 183 230
rect 183 196 192 230
rect 140 182 192 196
rect 140 158 192 170
rect 140 124 149 158
rect 149 124 183 158
rect 183 124 192 158
rect 140 118 192 124
rect 226 662 278 668
rect 226 628 235 662
rect 235 628 269 662
rect 269 628 278 662
rect 226 616 278 628
rect 226 590 278 604
rect 226 556 235 590
rect 235 556 269 590
rect 269 556 278 590
rect 226 552 278 556
rect 226 518 278 540
rect 226 488 235 518
rect 235 488 269 518
rect 269 488 278 518
rect 226 446 278 476
rect 226 424 235 446
rect 235 424 269 446
rect 269 424 278 446
rect 312 340 321 362
rect 321 340 355 362
rect 355 340 364 362
rect 312 310 364 340
rect 312 268 321 298
rect 321 268 355 298
rect 355 268 364 298
rect 312 246 364 268
rect 312 230 364 234
rect 312 196 321 230
rect 321 196 355 230
rect 355 196 364 230
rect 312 182 364 196
rect 312 158 364 170
rect 312 124 321 158
rect 321 124 355 158
rect 355 124 364 158
rect 312 118 364 124
rect 398 662 450 668
rect 398 628 407 662
rect 407 628 441 662
rect 441 628 450 662
rect 398 616 450 628
rect 398 590 450 604
rect 398 556 407 590
rect 407 556 441 590
rect 441 556 450 590
rect 398 552 450 556
rect 398 518 450 540
rect 398 488 407 518
rect 407 488 441 518
rect 441 488 450 518
rect 398 446 450 476
rect 398 424 407 446
rect 407 424 441 446
rect 441 424 450 446
rect 484 340 493 362
rect 493 340 527 362
rect 527 340 536 362
rect 484 310 536 340
rect 484 268 493 298
rect 493 268 527 298
rect 527 268 536 298
rect 484 246 536 268
rect 484 230 536 234
rect 484 196 493 230
rect 493 196 527 230
rect 527 196 536 230
rect 484 182 536 196
rect 484 158 536 170
rect 484 124 493 158
rect 493 124 527 158
rect 527 124 536 158
rect 484 118 536 124
<< metal2 >>
rect 0 668 676 674
rect 0 616 226 668
rect 278 616 398 668
rect 450 616 676 668
rect 0 604 676 616
rect 0 552 226 604
rect 278 552 398 604
rect 450 552 676 604
rect 0 540 676 552
rect 0 488 226 540
rect 278 488 398 540
rect 450 488 676 540
rect 0 476 676 488
rect 0 424 226 476
rect 278 424 398 476
rect 450 424 676 476
rect 0 418 676 424
rect 0 362 676 368
rect 0 310 140 362
rect 192 310 312 362
rect 364 310 484 362
rect 536 310 676 362
rect 0 298 676 310
rect 0 246 140 298
rect 192 246 312 298
rect 364 246 484 298
rect 536 246 676 298
rect 0 234 676 246
rect 0 182 140 234
rect 192 182 312 234
rect 364 182 484 234
rect 536 182 676 234
rect 0 170 676 182
rect 0 118 140 170
rect 192 118 312 170
rect 364 118 484 170
rect 536 118 676 170
rect 0 112 676 118
<< labels >>
flabel comment s 166 393 166 393 0 FreeSans 300 0 0 0 S
flabel comment s 252 393 252 393 0 FreeSans 300 0 0 0 S
flabel comment s 338 393 338 393 0 FreeSans 300 0 0 0 S
flabel comment s 424 393 424 393 0 FreeSans 300 0 0 0 S
flabel comment s 166 393 166 393 0 FreeSans 300 0 0 0 S
flabel comment s 252 393 252 393 0 FreeSans 300 0 0 0 D
flabel comment s 338 393 338 393 0 FreeSans 300 0 0 0 S
flabel comment s 424 393 424 393 0 FreeSans 300 0 0 0 D
flabel comment s 510 393 510 393 0 FreeSans 300 0 0 0 S
flabel metal1 s 53 497 53 497 7 FreeSans 300 90 0 0 SUBSTRATE
flabel metal1 s 612 497 612 497 7 FreeSans 300 90 0 0 SUBSTRATE
flabel metal1 s 313 740 395 765 0 FreeSans 300 0 0 0 GATE
port 2 nsew
flabel metal1 s 298 24 380 49 0 FreeSans 300 0 0 0 GATE
port 2 nsew
flabel metal2 s 11 503 29 573 0 FreeSans 300 90 0 0 DRAIN
port 3 nsew
flabel metal2 s 9 203 29 267 0 FreeSans 300 90 0 0 SOURCE
port 4 nsew
<< properties >>
string GDS_END 6050910
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 6035412
<< end >>
