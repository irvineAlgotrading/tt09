magic
tech sky130B
magscale 1 2
timestamp 1704896540
use sky130_fd_pr__hvdfl1sd2__example_55959141808462  sky130_fd_pr__hvdfl1sd2__example_55959141808462_0
timestamp 1704896540
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808462  sky130_fd_pr__hvdfl1sd2__example_55959141808462_1
timestamp 1704896540
transform 1 0 256 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808278  sky130_fd_pr__hvdfl1sd__example_55959141808278_0
timestamp 1704896540
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808278  sky130_fd_pr__hvdfl1sd__example_55959141808278_1
timestamp 1704896540
transform 1 0 412 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 64328830
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 64326868
<< end >>
